magic
tech gf180mcuC
magscale 1 5
timestamp 1675382720
<< obsm1 >>
rect 120 2430 89880 57225
<< metal2 >>
rect 2968 59600 3024 60000
rect 8568 59600 8624 60000
rect 14168 59600 14224 60000
rect 19768 59600 19824 60000
rect 25368 59600 25424 60000
rect 30968 59600 31024 60000
rect 36568 59600 36624 60000
rect 42168 59600 42224 60000
rect 47768 59600 47824 60000
rect 53368 59600 53424 60000
rect 58968 59600 59024 60000
rect 64568 59600 64624 60000
rect 70168 59600 70224 60000
rect 75768 59600 75824 60000
rect 81368 59600 81424 60000
rect 86968 59600 87024 60000
rect 2576 0 2632 400
rect 7560 0 7616 400
rect 12544 0 12600 400
rect 17528 0 17584 400
rect 22512 0 22568 400
rect 27496 0 27552 400
rect 32480 0 32536 400
rect 37464 0 37520 400
rect 42448 0 42504 400
rect 47432 0 47488 400
rect 52416 0 52472 400
rect 57400 0 57456 400
rect 62384 0 62440 400
rect 67368 0 67424 400
rect 72352 0 72408 400
rect 77336 0 77392 400
rect 82320 0 82376 400
rect 87304 0 87360 400
<< obsm2 >>
rect 238 59570 2938 59600
rect 3054 59570 8538 59600
rect 8654 59570 14138 59600
rect 14254 59570 19738 59600
rect 19854 59570 25338 59600
rect 25454 59570 30938 59600
rect 31054 59570 36538 59600
rect 36654 59570 42138 59600
rect 42254 59570 47738 59600
rect 47854 59570 53338 59600
rect 53454 59570 58938 59600
rect 59054 59570 64538 59600
rect 64654 59570 70138 59600
rect 70254 59570 75738 59600
rect 75854 59570 81338 59600
rect 81454 59570 86938 59600
rect 87054 59570 89810 59600
rect 238 430 89810 59570
rect 238 350 2546 430
rect 2662 350 7530 430
rect 7646 350 12514 430
rect 12630 350 17498 430
rect 17614 350 22482 430
rect 22598 350 27466 430
rect 27582 350 32450 430
rect 32566 350 37434 430
rect 37550 350 42418 430
rect 42534 350 47402 430
rect 47518 350 52386 430
rect 52502 350 57370 430
rect 57486 350 62354 430
rect 62470 350 67338 430
rect 67454 350 72322 430
rect 72438 350 77306 430
rect 77422 350 82290 430
rect 82406 350 87274 430
rect 87390 350 89810 430
<< metal3 >>
rect 0 56000 400 56056
rect 89600 56000 90000 56056
rect 0 48552 400 48608
rect 89600 48552 90000 48608
rect 0 41104 400 41160
rect 89600 41104 90000 41160
rect 0 33656 400 33712
rect 89600 33656 90000 33712
rect 0 26208 400 26264
rect 89600 26208 90000 26264
rect 0 18760 400 18816
rect 89600 18760 90000 18816
rect 0 11312 400 11368
rect 89600 11312 90000 11368
rect 0 3864 400 3920
rect 89600 3864 90000 3920
<< obsm3 >>
rect 233 56086 89815 57209
rect 430 55970 89570 56086
rect 233 48638 89815 55970
rect 430 48522 89570 48638
rect 233 41190 89815 48522
rect 430 41074 89570 41190
rect 233 33742 89815 41074
rect 430 33626 89570 33742
rect 233 26294 89815 33626
rect 430 26178 89570 26294
rect 233 18846 89815 26178
rect 430 18730 89570 18846
rect 233 11398 89815 18730
rect 430 11282 89570 11398
rect 233 3950 89815 11282
rect 430 3834 89570 3950
rect 233 2446 89815 3834
<< metal4 >>
rect 1672 2430 1832 57225
rect 9352 2430 9512 57225
rect 17032 2430 17192 57225
rect 24712 2430 24872 57225
rect 32392 2430 32552 57225
rect 40072 2430 40232 57225
rect 47752 2430 47912 57225
rect 55432 2430 55592 57225
rect 63112 2430 63272 57225
rect 70792 2430 70952 57225
rect 78472 2430 78632 57225
rect 86152 2430 86312 57225
<< obsm4 >>
rect 3374 25993 9322 37147
rect 9542 25993 17002 37147
rect 17222 25993 24682 37147
rect 24902 25993 32362 37147
rect 32582 25993 40042 37147
rect 40262 25993 47722 37147
rect 47942 25993 55402 37147
rect 55622 25993 63082 37147
rect 63302 25993 70658 37147
<< labels >>
rlabel metal3 s 89600 3864 90000 3920 6 a[0]
port 1 nsew signal input
rlabel metal3 s 89600 11312 90000 11368 6 a[1]
port 2 nsew signal input
rlabel metal3 s 89600 18760 90000 18816 6 a[2]
port 3 nsew signal input
rlabel metal3 s 89600 26208 90000 26264 6 a[3]
port 4 nsew signal input
rlabel metal3 s 89600 33656 90000 33712 6 a[4]
port 5 nsew signal input
rlabel metal3 s 89600 41104 90000 41160 6 a[5]
port 6 nsew signal input
rlabel metal3 s 89600 48552 90000 48608 6 a[6]
port 7 nsew signal input
rlabel metal3 s 89600 56000 90000 56056 6 a[7]
port 8 nsew signal input
rlabel metal3 s 0 3864 400 3920 6 b[0]
port 9 nsew signal input
rlabel metal3 s 0 11312 400 11368 6 b[1]
port 10 nsew signal input
rlabel metal3 s 0 18760 400 18816 6 b[2]
port 11 nsew signal input
rlabel metal3 s 0 26208 400 26264 6 b[3]
port 12 nsew signal input
rlabel metal3 s 0 33656 400 33712 6 b[4]
port 13 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 b[5]
port 14 nsew signal input
rlabel metal3 s 0 48552 400 48608 6 b[6]
port 15 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 b[7]
port 16 nsew signal input
rlabel metal2 s 12544 0 12600 400 6 ci[0]
port 17 nsew signal input
rlabel metal2 s 62384 0 62440 400 6 ci[10]
port 18 nsew signal input
rlabel metal2 s 67368 0 67424 400 6 ci[11]
port 19 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 ci[12]
port 20 nsew signal input
rlabel metal2 s 77336 0 77392 400 6 ci[13]
port 21 nsew signal input
rlabel metal2 s 82320 0 82376 400 6 ci[14]
port 22 nsew signal input
rlabel metal2 s 87304 0 87360 400 6 ci[15]
port 23 nsew signal input
rlabel metal2 s 17528 0 17584 400 6 ci[1]
port 24 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 ci[2]
port 25 nsew signal input
rlabel metal2 s 27496 0 27552 400 6 ci[3]
port 26 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 ci[4]
port 27 nsew signal input
rlabel metal2 s 37464 0 37520 400 6 ci[5]
port 28 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 ci[6]
port 29 nsew signal input
rlabel metal2 s 47432 0 47488 400 6 ci[7]
port 30 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 ci[8]
port 31 nsew signal input
rlabel metal2 s 57400 0 57456 400 6 ci[9]
port 32 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 clk
port 33 nsew signal input
rlabel metal2 s 2968 59600 3024 60000 6 o[0]
port 34 nsew signal output
rlabel metal2 s 58968 59600 59024 60000 6 o[10]
port 35 nsew signal output
rlabel metal2 s 64568 59600 64624 60000 6 o[11]
port 36 nsew signal output
rlabel metal2 s 70168 59600 70224 60000 6 o[12]
port 37 nsew signal output
rlabel metal2 s 75768 59600 75824 60000 6 o[13]
port 38 nsew signal output
rlabel metal2 s 81368 59600 81424 60000 6 o[14]
port 39 nsew signal output
rlabel metal2 s 86968 59600 87024 60000 6 o[15]
port 40 nsew signal output
rlabel metal2 s 8568 59600 8624 60000 6 o[1]
port 41 nsew signal output
rlabel metal2 s 14168 59600 14224 60000 6 o[2]
port 42 nsew signal output
rlabel metal2 s 19768 59600 19824 60000 6 o[3]
port 43 nsew signal output
rlabel metal2 s 25368 59600 25424 60000 6 o[4]
port 44 nsew signal output
rlabel metal2 s 30968 59600 31024 60000 6 o[5]
port 45 nsew signal output
rlabel metal2 s 36568 59600 36624 60000 6 o[6]
port 46 nsew signal output
rlabel metal2 s 42168 59600 42224 60000 6 o[7]
port 47 nsew signal output
rlabel metal2 s 47768 59600 47824 60000 6 o[8]
port 48 nsew signal output
rlabel metal2 s 53368 59600 53424 60000 6 o[9]
port 49 nsew signal output
rlabel metal2 s 7560 0 7616 400 6 rst
port 50 nsew signal input
rlabel metal4 s 1672 2430 1832 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 17032 2430 17192 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 32392 2430 32552 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 47752 2430 47912 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 63112 2430 63272 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 78472 2430 78632 57225 6 vdd
port 51 nsew power bidirectional
rlabel metal4 s 9352 2430 9512 57225 6 vss
port 52 nsew ground bidirectional
rlabel metal4 s 24712 2430 24872 57225 6 vss
port 52 nsew ground bidirectional
rlabel metal4 s 40072 2430 40232 57225 6 vss
port 52 nsew ground bidirectional
rlabel metal4 s 55432 2430 55592 57225 6 vss
port 52 nsew ground bidirectional
rlabel metal4 s 70792 2430 70952 57225 6 vss
port 52 nsew ground bidirectional
rlabel metal4 s 86152 2430 86312 57225 6 vss
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5203668
string GDS_FILE /home/brettcm/caravel/main/osu180cells/openlane/ffra/runs/23_02_02_18_03/results/signoff/ffra.magic.gds
string GDS_START 98782
<< end >>

