magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 224 844
rect 78 386 146 724
rect 78 60 146 237
rect 0 -60 224 60
<< labels >>
rlabel metal1 s 0 724 224 844 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 78 386 146 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 78 60 146 237 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 224 60 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 784
string LEFclass core WELLTAP
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 415834
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 414122
<< end >>
