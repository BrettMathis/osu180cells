magic
tech gf180mcuA
magscale 1 10
timestamp 1669648928
<< checkpaint >>
rect 66400 66400 73000 73000
<< metal3 >>
rect 68400 69678 69678 71000
rect 68400 68779 71000 69678
tri 68400 68400 68779 68779 ne
rect 68779 68400 71000 68779
<< end >>
