magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 3360 844
rect 288 586 356 724
rect 636 601 704 724
rect 56 354 318 426
rect 288 60 356 183
rect 690 354 878 430
rect 656 60 724 215
rect 1541 540 1609 724
rect 2570 656 2638 724
rect 1540 60 1608 162
rect 2969 551 3037 724
rect 2544 60 2612 190
rect 3154 162 3270 597
rect 3000 60 3046 138
rect 0 -60 3360 60
<< obsm1 >>
rect 95 518 141 645
rect 503 542 569 645
rect 766 632 1271 678
rect 766 542 812 632
rect 95 472 433 518
rect 387 275 433 472
rect 75 229 433 275
rect 503 496 812 542
rect 884 529 1058 575
rect 75 147 121 229
rect 503 147 569 496
rect 1011 215 1058 529
rect 880 169 1058 215
rect 1115 410 1183 559
rect 2686 620 2923 666
rect 2686 610 2732 620
rect 1808 478 1876 586
rect 1419 410 1876 478
rect 1115 364 1356 410
rect 1115 158 1161 364
rect 1310 346 1356 364
rect 1218 254 1264 318
rect 1310 300 1740 346
rect 1218 208 1712 254
rect 1666 152 1712 208
rect 1808 198 1876 410
rect 2032 517 2100 586
rect 2358 563 2732 610
rect 2032 471 2726 517
rect 2032 198 2100 471
rect 2658 421 2726 471
rect 2239 152 2285 419
rect 2785 377 2831 570
rect 2877 469 2923 620
rect 2877 423 3092 469
rect 2785 375 3000 377
rect 2435 328 3000 375
rect 2780 300 3000 328
rect 2331 236 2704 282
rect 2331 178 2377 236
rect 1666 106 2285 152
rect 2658 152 2704 236
rect 2780 198 2848 300
rect 3046 230 3092 423
rect 2908 184 3092 230
rect 2908 152 2954 184
rect 2658 106 2954 152
<< labels >>
rlabel metal1 s 690 354 878 430 6 D
port 1 nsew default input
rlabel metal1 s 56 354 318 426 6 CLKN
port 2 nsew clock input
rlabel metal1 s 3154 162 3270 597 6 Q
port 3 nsew default output
rlabel metal1 s 0 724 3360 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 656 3037 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2570 656 2638 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 656 1609 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 656 704 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 656 356 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 601 3037 656 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 601 1609 656 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 601 704 656 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 601 356 656 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 586 3037 601 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 586 1609 601 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 586 356 601 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 551 3037 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 551 1609 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 540 1609 551 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 656 190 724 215 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 183 2612 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 183 724 190 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 162 2612 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 162 724 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 162 356 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 138 2612 162 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1540 138 1608 162 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 138 724 162 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 138 356 162 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3000 60 3046 138 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 60 2612 138 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1540 60 1608 138 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 60 724 138 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 60 356 138 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3360 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 848142
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 840762
<< end >>
