magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1456 844
rect 242 508 310 724
rect 928 506 974 724
rect 141 242 318 322
rect 273 60 319 196
rect 1132 161 1214 676
rect 1357 506 1404 724
rect 909 60 955 138
rect 1357 60 1403 229
rect 0 -60 1456 60
<< obsm1 >>
rect 49 462 95 565
rect 49 415 407 462
rect 49 128 95 415
rect 361 394 407 415
rect 477 358 523 565
rect 621 456 667 542
rect 621 410 1075 456
rect 477 310 811 358
rect 477 128 543 310
rect 1029 250 1075 410
rect 810 204 1075 250
rect 810 153 857 204
rect 629 106 857 153
<< labels >>
rlabel metal1 s 141 242 318 322 6 I
port 1 nsew default input
rlabel metal1 s 1132 161 1214 676 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 1456 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1357 508 1404 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 928 508 974 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 242 508 310 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1357 506 1404 508 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 928 506 974 508 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1357 196 1403 229 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1357 138 1403 196 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 138 319 196 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1357 60 1403 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 909 60 955 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1456 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1064900
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1061040
<< end >>
