magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -2104 -186 2105 299
rect -2105 -300 2105 -186
<< nsubdiff >>
rect -1957 102 1957 157
rect -1957 56 -1900 102
rect -1854 56 -1737 102
rect -1691 56 -1574 102
rect -1528 56 -1411 102
rect -1365 56 -1247 102
rect -1201 56 -1084 102
rect -1038 56 -921 102
rect -875 56 -758 102
rect -712 56 -595 102
rect -549 56 -431 102
rect -385 56 -268 102
rect -222 56 -105 102
rect -59 56 59 102
rect 105 56 222 102
rect 268 56 385 102
rect 431 56 549 102
rect 595 56 712 102
rect 758 56 875 102
rect 921 56 1038 102
rect 1084 56 1201 102
rect 1247 56 1365 102
rect 1411 56 1528 102
rect 1574 56 1691 102
rect 1737 56 1854 102
rect 1900 56 1957 102
rect -1957 -56 1957 56
rect -1957 -102 -1900 -56
rect -1854 -102 -1737 -56
rect -1691 -102 -1574 -56
rect -1528 -102 -1411 -56
rect -1365 -102 -1247 -56
rect -1201 -102 -1084 -56
rect -1038 -102 -921 -56
rect -875 -102 -758 -56
rect -712 -102 -595 -56
rect -549 -102 -431 -56
rect -385 -102 -268 -56
rect -222 -102 -105 -56
rect -59 -102 59 -56
rect 105 -102 222 -56
rect 268 -102 385 -56
rect 431 -102 549 -56
rect 595 -102 712 -56
rect 758 -102 875 -56
rect 921 -102 1038 -56
rect 1084 -102 1201 -56
rect 1247 -102 1365 -56
rect 1411 -102 1528 -56
rect 1574 -102 1691 -56
rect 1737 -102 1854 -56
rect 1900 -102 1957 -56
rect -1957 -157 1957 -102
<< nsubdiffcont >>
rect -1900 56 -1854 102
rect -1737 56 -1691 102
rect -1574 56 -1528 102
rect -1411 56 -1365 102
rect -1247 56 -1201 102
rect -1084 56 -1038 102
rect -921 56 -875 102
rect -758 56 -712 102
rect -595 56 -549 102
rect -431 56 -385 102
rect -268 56 -222 102
rect -105 56 -59 102
rect 59 56 105 102
rect 222 56 268 102
rect 385 56 431 102
rect 549 56 595 102
rect 712 56 758 102
rect 875 56 921 102
rect 1038 56 1084 102
rect 1201 56 1247 102
rect 1365 56 1411 102
rect 1528 56 1574 102
rect 1691 56 1737 102
rect 1854 56 1900 102
rect -1900 -102 -1854 -56
rect -1737 -102 -1691 -56
rect -1574 -102 -1528 -56
rect -1411 -102 -1365 -56
rect -1247 -102 -1201 -56
rect -1084 -102 -1038 -56
rect -921 -102 -875 -56
rect -758 -102 -712 -56
rect -595 -102 -549 -56
rect -431 -102 -385 -56
rect -268 -102 -222 -56
rect -105 -102 -59 -56
rect 59 -102 105 -56
rect 222 -102 268 -56
rect 385 -102 431 -56
rect 549 -102 595 -56
rect 712 -102 758 -56
rect 875 -102 921 -56
rect 1038 -102 1084 -56
rect 1201 -102 1247 -56
rect 1365 -102 1411 -56
rect 1528 -102 1574 -56
rect 1691 -102 1737 -56
rect 1854 -102 1900 -56
<< metal1 >>
rect -1936 102 1937 137
rect -1936 56 -1900 102
rect -1854 56 -1737 102
rect -1691 56 -1574 102
rect -1528 56 -1411 102
rect -1365 56 -1247 102
rect -1201 56 -1084 102
rect -1038 56 -921 102
rect -875 56 -758 102
rect -712 56 -595 102
rect -549 56 -431 102
rect -385 56 -268 102
rect -222 56 -105 102
rect -59 56 59 102
rect 105 56 222 102
rect 268 56 385 102
rect 431 56 549 102
rect 595 56 712 102
rect 758 56 875 102
rect 921 56 1038 102
rect 1084 56 1201 102
rect 1247 56 1365 102
rect 1411 56 1528 102
rect 1574 56 1691 102
rect 1737 56 1854 102
rect 1900 56 1937 102
rect -1936 -56 1937 56
rect -1936 -102 -1900 -56
rect -1854 -102 -1737 -56
rect -1691 -102 -1574 -56
rect -1528 -102 -1411 -56
rect -1365 -102 -1247 -56
rect -1201 -102 -1084 -56
rect -1038 -102 -921 -56
rect -875 -102 -758 -56
rect -712 -102 -595 -56
rect -549 -102 -431 -56
rect -385 -102 -268 -56
rect -222 -102 -105 -56
rect -59 -102 59 -56
rect 105 -102 222 -56
rect 268 -102 385 -56
rect 431 -102 549 -56
rect 595 -102 712 -56
rect 758 -102 875 -56
rect 921 -102 1038 -56
rect 1084 -102 1201 -56
rect 1247 -102 1365 -56
rect 1411 -102 1528 -56
rect 1574 -102 1691 -56
rect 1737 -102 1854 -56
rect 1900 -102 1937 -56
rect -1936 -137 1937 -102
<< properties >>
string GDS_END 845448
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 842084
<< end >>
