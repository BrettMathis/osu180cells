VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adder
  CLASS BLOCK ;
  FOREIGN adder ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN a_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 57.680 0.000 58.240 4.000 ;
    END
  END a_in[0]
  PIN a_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 169.680 0.000 170.240 4.000 ;
    END
  END a_in[1]
  PIN a_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END a_in[2]
  PIN a_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 393.680 0.000 394.240 4.000 ;
    END
  END a_in[3]
  PIN a_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 505.680 0.000 506.240 4.000 ;
    END
  END a_in[4]
  PIN a_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 617.680 0.000 618.240 4.000 ;
    END
  END a_in[5]
  PIN a_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 729.680 0.000 730.240 4.000 ;
    END
  END a_in[6]
  PIN a_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 841.680 0.000 842.240 4.000 ;
    END
  END a_in[7]
  PIN b_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 38.640 900.000 39.200 ;
    END
  END b_in[0]
  PIN b_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 113.120 900.000 113.680 ;
    END
  END b_in[1]
  PIN b_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 187.600 900.000 188.160 ;
    END
  END b_in[2]
  PIN b_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 262.080 900.000 262.640 ;
    END
  END b_in[3]
  PIN b_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 336.560 900.000 337.120 ;
    END
  END b_in[4]
  PIN b_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 411.040 900.000 411.600 ;
    END
  END b_in[5]
  PIN b_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 485.520 900.000 486.080 ;
    END
  END b_in[6]
  PIN b_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 560.000 900.000 560.560 ;
    END
  END b_in[7]
  PIN sum[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 57.680 596.000 58.240 600.000 ;
    END
  END sum[0]
  PIN sum[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 169.680 596.000 170.240 600.000 ;
    END
  END sum[1]
  PIN sum[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 281.680 596.000 282.240 600.000 ;
    END
  END sum[2]
  PIN sum[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 393.680 596.000 394.240 600.000 ;
    END
  END sum[3]
  PIN sum[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 505.680 596.000 506.240 600.000 ;
    END
  END sum[4]
  PIN sum[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 617.680 596.000 618.240 600.000 ;
    END
  END sum[5]
  PIN sum[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 729.680 596.000 730.240 600.000 ;
    END
  END sum[6]
  PIN sum[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 841.680 596.000 842.240 600.000 ;
    END
  END sum[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET4 ;
        RECT 16.720 24.300 18.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 170.320 24.300 171.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 323.920 24.300 325.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 477.520 24.300 479.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 631.120 24.300 632.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 784.720 24.300 786.320 572.250 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET4 ;
        RECT 93.520 24.300 95.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 247.120 24.300 248.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 400.720 24.300 402.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 554.320 24.300 555.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 707.920 24.300 709.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 861.520 24.300 863.120 572.250 ;
    END
  END vss
  OBS
      LAYER MET1 ;
        RECT 1.200 24.300 898.800 572.250 ;
      LAYER MET2 ;
        RECT 16.860 595.700 57.380 596.000 ;
        RECT 58.540 595.700 169.380 596.000 ;
        RECT 170.540 595.700 281.380 596.000 ;
        RECT 282.540 595.700 393.380 596.000 ;
        RECT 394.540 595.700 505.380 596.000 ;
        RECT 506.540 595.700 617.380 596.000 ;
        RECT 618.540 595.700 729.380 596.000 ;
        RECT 730.540 595.700 841.380 596.000 ;
        RECT 842.540 595.700 898.100 596.000 ;
        RECT 16.860 4.300 898.100 595.700 ;
        RECT 16.860 3.500 57.380 4.300 ;
        RECT 58.540 3.500 169.380 4.300 ;
        RECT 170.540 3.500 281.380 4.300 ;
        RECT 282.540 3.500 393.380 4.300 ;
        RECT 394.540 3.500 505.380 4.300 ;
        RECT 506.540 3.500 617.380 4.300 ;
        RECT 618.540 3.500 729.380 4.300 ;
        RECT 730.540 3.500 841.380 4.300 ;
        RECT 842.540 3.500 898.100 4.300 ;
      LAYER MET3 ;
        RECT 16.810 560.860 898.150 572.090 ;
        RECT 16.810 559.700 895.700 560.860 ;
        RECT 16.810 486.380 898.150 559.700 ;
        RECT 16.810 485.220 895.700 486.380 ;
        RECT 16.810 411.900 898.150 485.220 ;
        RECT 16.810 410.740 895.700 411.900 ;
        RECT 16.810 337.420 898.150 410.740 ;
        RECT 16.810 336.260 895.700 337.420 ;
        RECT 16.810 262.940 898.150 336.260 ;
        RECT 16.810 261.780 895.700 262.940 ;
        RECT 16.810 188.460 898.150 261.780 ;
        RECT 16.810 187.300 895.700 188.460 ;
        RECT 16.810 113.980 898.150 187.300 ;
        RECT 16.810 112.820 895.700 113.980 ;
        RECT 16.810 39.500 898.150 112.820 ;
        RECT 16.810 38.340 895.700 39.500 ;
        RECT 16.810 24.460 898.150 38.340 ;
      LAYER MET4 ;
        RECT 391.580 242.010 394.100 256.110 ;
  END
END adder
END LIBRARY

