* NGSPICE file created from gf180mcu_fd_ip_sram__sram256x8m8wm1.ext - technology: gf180mcuB

.subckt dcap_103_novia_256x8m81 w_n203_44# a_n67_185# a_73_103#
X0 a_n67_185# a_73_103# a_n67_185# w_n203_44# pmos_3p3 w=2.275u l=2.365u
.ends

.subckt x018SRAM_cell1_256x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_2x_256x8m81 018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS
X018SRAM_cell1_256x8m81_0 018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_256x8m81
X018SRAM_cell1_256x8m81_1 018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_256x8m81
.ends

.subckt Cell_array32x1_256x8m81 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_246_342# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
X018SRAM_cell1_2x_256x8m81_10 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_11 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_13 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_12 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_14 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_15 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_1 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_0 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_2 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_3 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_4 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_5 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_6 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_7 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_8 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_246_712# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_9 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_246_712#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_246_342# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_246_712# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
.ends

.subckt rarray4_256_256x8m81 WL[23] WL[26] WL[18] WL[11] WL[15] WL[14] WL[19] WL[31]
+ WL[13] WL[16] Cell_array32x1_256x8m81_18/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_30/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_28/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_9/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_27/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_20/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_21/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_17/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[5] Cell_array32x1_256x8m81_25/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[2] Cell_array32x1_256x8m81_26/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_13/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_12/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_26/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_24/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_10/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_8/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_11/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[27] Cell_array32x1_256x8m81_11/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_16/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[0] Cell_array32x1_256x8m81_29/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_22/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_4/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_14/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_15/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_7/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_16/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[8] Cell_array32x1_256x8m81_0/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_20/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_19/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_2/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_25/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_2/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[24] Cell_array32x1_256x8m81_10/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_31/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_23/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[3] Cell_array32x1_256x8m81_15/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_28/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_5/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_30/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_13/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_1/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[6] Cell_array32x1_256x8m81_6/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_7/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_21/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_3/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[1] Cell_array32x1_256x8m81_18/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_6/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[29] Cell_array32x1_256x8m81_4/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[4] WL[12] Cell_array32x1_256x8m81_9/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_24/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_22/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[28] WL[30] Cell_array32x1_256x8m81_29/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_14/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ WL[9] Cell_array32x1_256x8m81_27/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[25] Cell_array32x1_256x8m81_0/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_12/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_19/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_5/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ Cell_array32x1_256x8m81_17/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[20] Cell_array32x1_256x8m81_1/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[21] WL[7] Cell_array32x1_256x8m81_3/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[17] Cell_array32x1_256x8m81_31/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ WL[10] WL[22] Cell_array32x1_256x8m81_8/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81_23/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
XCell_array32x1_256x8m81_30 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_30/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_30/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_0 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_0/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_0/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_20 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_20/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_20/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_31 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_31/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_31/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_1 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_1/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_1/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_21 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_21/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_21/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_10 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_10/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_10/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_2 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_2/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_2/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_22 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_22/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_22/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_11 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_11/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_11/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_3 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_3/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_3/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_23 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_23/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_23/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_12 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_12/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_12/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_4 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_4/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_4/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_24 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_24/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_24/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_13 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_13/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_13/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_5 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_5/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_5/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_25 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_25/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_25/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_14 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_14/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_14/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_6 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_6/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_6/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_26 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_26/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_26/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_15 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_15/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_15/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_7 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_7/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_7/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_27 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_27/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_27/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_16 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_16/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_16/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_8 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_8/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_8/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_17 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_17/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_17/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_28 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_28/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_28/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_9 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_9/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_9/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_18 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_18/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_18/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_29 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_29/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_29/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
XCell_array32x1_256x8m81_19 VSS WL[4] VSS WL[28] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] WL[25] VSS WL[11] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS VSS WL[21] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[0] VSS WL[1] WL[4] VSS VSS WL[5] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[22] WL[6] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[7] WL[2] WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[8] VSS WL[5] VSS WL[29] WL[9] WL[15] WL[10] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[11] VSS VSS WL[12] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[13] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[14] VSS WL[0] WL[15] WL[26] VSS WL[12] WL[16] WL[23] WL[17] WL[9] VSS WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[18] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[19]
+ WL[19] VSS WL[22] WL[20] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[21] WL[23] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[24] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[25] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[6] WL[26]
+ WL[30] VSS WL[16] WL[1] WL[27] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[27] WL[28] WL[13] VSS WL[29] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[30] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS WL[31] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ WL[2] Cell_array32x1_256x8m81_19/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ WL[3] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS WL[24]
+ 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[10] VSS WL[20]
+ VSS WL[7] 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# WL[31]
+ WL[17] VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS
+ VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622# VSS 018SRAM_strap1_2x_256x8m81_9/018SRAM_strap1_256x8m81_1/w_n68_622#
+ VSS Cell_array32x1_256x8m81_19/018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ Cell_array32x1_256x8m81
.ends

.subckt pmos_5p0431059087814_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.61u l=0.6u
.ends

.subckt pmos_1p2$$46887980_256x8m81 pmos_5p0431059087814_256x8m81_0/S a_n31_n74# pmos_5p0431059087814_256x8m81_0/D
+ w_n286_n142#
Xpmos_5p0431059087814_256x8m81_0 w_n286_n142# pmos_5p0431059087814_256x8m81_0/D a_n31_n74#
+ pmos_5p0431059087814_256x8m81_0/S pmos_5p0431059087814_256x8m81
.ends

.subckt pmos_5p0431059087816_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_5p0431059087817_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=13.61u l=0.6u
.ends

.subckt nmos_1p2$$46884908_256x8m81 nmos_5p0431059087817_256x8m81_0/S nmos_5p0431059087817_256x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p0431059087817_256x8m81_0 nmos_5p0431059087817_256x8m81_0/D a_n31_n74# nmos_5p0431059087817_256x8m81_0/S
+ VSUBS nmos_5p0431059087817_256x8m81
.ends

.subckt pmos_5p0431059087810_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.81u l=0.6u
.ends

.subckt pmos_1p2$$46889004_256x8m81 pmos_5p0431059087810_256x8m81_0/D w_n286_n142#
+ a_n31_n74# pmos_5p0431059087810_256x8m81_0/S
Xpmos_5p0431059087810_256x8m81_0 w_n286_n142# pmos_5p0431059087810_256x8m81_0/D a_n31_n74#
+ pmos_5p0431059087810_256x8m81_0/S pmos_5p0431059087810_256x8m81
.ends

.subckt nmos_5p0431059087815_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_1p2$$46883884_256x8m81 nmos_5p0431059087815_256x8m81_0/S a_n31_n73# nmos_5p0431059087815_256x8m81_0/D
+ VSUBS
Xnmos_5p0431059087815_256x8m81_0 nmos_5p0431059087815_256x8m81_0/D a_n31_n73# nmos_5p0431059087815_256x8m81_0/S
+ VSUBS nmos_5p0431059087815_256x8m81
.ends

.subckt nmos_5p04310590878111_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_1p2$$46885932_256x8m81 pmos_5p0431059087816_256x8m81_0/D a_193_n73# a_n31_n74#
+ w_n286_n141# pmos_5p0431059087816_256x8m81_0/S
Xpmos_5p0431059087816_256x8m81_0 w_n286_n141# pmos_5p0431059087816_256x8m81_0/D a_n31_n74#
+ pmos_5p0431059087816_256x8m81_0/S a_193_n73# pmos_5p0431059087816_256x8m81
.ends

.subckt nmos_5p0431059087818_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$46563372_256x8m81 nmos_5p0431059087818_256x8m81_0/D a_n31_n74# nmos_5p0431059087818_256x8m81_0/S
+ VSUBS
Xnmos_5p0431059087818_256x8m81_0 nmos_5p0431059087818_256x8m81_0/D a_n31_n74# nmos_5p0431059087818_256x8m81_0/S
+ VSUBS nmos_5p0431059087818_256x8m81
.ends

.subckt nmos_5p04310590878110_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p0431059087819_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt pmos_5p0431059087813_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_1p2$$46273580_256x8m81 pmos_5p0431059087813_256x8m81_0/S a_193_n74# pmos_5p0431059087813_256x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p0431059087813_256x8m81_0 w_n286_n142# pmos_5p0431059087813_256x8m81_0/D a_n31_n74#
+ pmos_5p0431059087813_256x8m81_0/S a_193_n74# pmos_5p0431059087813_256x8m81
.ends

.subckt din_256x8m81 datain wep men d db m1_164_8068# pmos_5p0431059087810_256x8m81_0/D
+ vdd vss
Xpmos_1p2$$46887980_256x8m81_0 vdd pmos_5p0431059087810_256x8m81_0/S pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ vdd pmos_1p2$$46887980_256x8m81
Xpmos_5p0431059087816_256x8m81_0 vdd vdd datain pmos_5p0431059087816_256x8m81_0/S
+ pmos_5p0431059087816_256x8m81_0/S pmos_5p0431059087816_256x8m81
Xnmos_1p2$$46884908_256x8m81_0 vss pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ pmos_5p0431059087810_256x8m81_0/S vss nmos_1p2$$46884908_256x8m81
Xpmos_1p2$$46889004_256x8m81_1 pmos_5p0431059087819_256x8m81_0/S vdd a_500_6666# db
+ pmos_1p2$$46889004_256x8m81
Xpmos_1p2$$46889004_256x8m81_0 pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ vdd a_500_6666# d pmos_1p2$$46889004_256x8m81
Xpmos_5p0431059087810_256x8m81_0 vdd pmos_5p0431059087810_256x8m81_0/D nmos_5p04310590878111_256x8m81_1/D
+ pmos_5p0431059087810_256x8m81_0/S pmos_5p0431059087810_256x8m81
Xnmos_1p2$$46883884_256x8m81_0 db wep pmos_5p0431059087819_256x8m81_0/S vss nmos_1p2$$46883884_256x8m81
Xnmos_1p2$$46883884_256x8m81_1 pmos_5p0431059087819_256x8m81_0/S pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ vss vss nmos_1p2$$46883884_256x8m81
Xnmos_1p2$$46883884_256x8m81_2 d wep pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ vss nmos_1p2$$46883884_256x8m81
Xnmos_5p04310590878111_256x8m81_0 vss datain pmos_5p0431059087816_256x8m81_0/S pmos_5p0431059087816_256x8m81_0/S
+ vss nmos_5p04310590878111_256x8m81
Xpmos_1p2$$46885932_256x8m81_0 nmos_5p04310590878111_256x8m81_1/D pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ men vdd pmos_5p0431059087816_256x8m81_0/S pmos_1p2$$46885932_256x8m81
Xnmos_5p04310590878111_256x8m81_1 nmos_5p04310590878111_256x8m81_1/D pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ pmos_5p0431059087816_256x8m81_0/S men vss nmos_5p04310590878111_256x8m81
Xnmos_1p2$$46563372_256x8m81_0 pmos_5p0431059087816_256x8m81_0/S pmos_5p0431059087810_256x8m81_0/S
+ vss vss nmos_1p2$$46563372_256x8m81
Xnmos_1p2$$46563372_256x8m81_1 pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ men vss vss nmos_1p2$$46563372_256x8m81
Xnmos_5p04310590878110_256x8m81_0 vss nmos_5p04310590878111_256x8m81_1/D pmos_5p0431059087810_256x8m81_0/S
+ vss nmos_5p04310590878110_256x8m81
Xpmos_5p0431059087819_256x8m81_0 vdd vdd pmos_1p2$$46889004_256x8m81_0/pmos_5p0431059087810_256x8m81_0/D
+ pmos_5p0431059087819_256x8m81_0/S pmos_5p0431059087819_256x8m81
Xpmos_1p2$$46273580_256x8m81_0 vdd men pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ vdd men pmos_1p2$$46273580_256x8m81
Xpmos_1p2$$46273580_256x8m81_1 vdd pmos_5p0431059087810_256x8m81_0/S pmos_5p0431059087816_256x8m81_0/S
+ vdd pmos_5p0431059087810_256x8m81_0/S pmos_1p2$$46273580_256x8m81
X0 vdd wep a_500_6666# vdd pmos_3p3 w=1.485u l=0.6u
X1 a_500_6666# wep vss vss nmos_3p3 w=1.14u l=0.6u
X2 a_500_6666# wep vdd vdd pmos_3p3 w=1.485u l=0.6u
.ends

.subckt nmos_5p04310590878124_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45102124_256x8m81 a_1313_n74# nmos_5p04310590878124_256x8m81_0/S
+ a_193_n74# a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# nmos_5p04310590878124_256x8m81_0/D
+ a_417_n74# VSUBS
Xnmos_5p04310590878124_256x8m81_0 nmos_5p04310590878124_256x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590878124_256x8m81_0/S a_417_n74# a_193_n74# a_1313_n74#
+ a_1089_n74# VSUBS nmos_5p04310590878124_256x8m81
.ends

.subckt pmos_5p04310590878138_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt nmos_5p04310590878126_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_5p04310590878135_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
.ends

.subckt nmos_1p2$$45103148_256x8m81 nmos_5p04310590878135_256x8m81_0/D a_865_n73#
+ a_193_n74# nmos_5p04310590878135_256x8m81_0/S a_1089_n74# a_n31_n74# a_641_n74#
+ a_417_n74# VSUBS
Xnmos_5p04310590878135_256x8m81_0 nmos_5p04310590878135_256x8m81_0/D a_n31_n74# a_865_n73#
+ a_641_n74# nmos_5p04310590878135_256x8m81_0/S a_417_n74# a_193_n74# a_1089_n74#
+ VSUBS nmos_5p04310590878135_256x8m81
.ends

.subckt pmos_5p04310590878136_256x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
.ends

.subckt pmos_1p2$$46283820_256x8m81 a_641_n74# a_1985_n74# a_1761_n74# a_417_n74#
+ a_1537_n74# a_1313_n74# pmos_5p04310590878136_256x8m81_0/D w_n286_n142# a_193_n74#
+ a_1089_n74# a_865_n74# a_n31_n74# pmos_5p04310590878136_256x8m81_0/S
Xpmos_5p04310590878136_256x8m81_0 w_n286_n142# pmos_5p04310590878136_256x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590878136_256x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310590878136_256x8m81
.ends

.subckt nmos_5p04310590878127_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.61u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.61u l=0.6u
.ends

.subckt nmos_1p2$$45100076_256x8m81 nmos_5p04310590878127_256x8m81_0/D a_193_n74#
+ a_n31_n74# nmos_5p04310590878127_256x8m81_0/S VSUBS
Xnmos_5p04310590878127_256x8m81_0 nmos_5p04310590878127_256x8m81_0/D a_n31_n74# nmos_5p04310590878127_256x8m81_0/S
+ a_193_n74# VSUBS nmos_5p04310590878127_256x8m81
.ends

.subckt pmos_5p04310590878125_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt nmos_5p04310590878133_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.44u l=0.6u
.ends

.subckt nmos_5p04310590878123_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.6u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt pmos_5p04310590878129_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.41u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.41u l=0.6u
.ends

.subckt pmos_1p2$$46287916_256x8m81 pmos_5p04310590878129_256x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310590878129_256x8m81_0/S
Xpmos_5p04310590878129_256x8m81_0 w_n286_n142# pmos_5p04310590878129_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878129_256x8m81_0/S a_193_n74# pmos_5p04310590878129_256x8m81
.ends

.subckt pmos_5p04310590878130_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$46284844_256x8m81 a_n31_n74# pmos_5p04310590878130_256x8m81_0/S
+ pmos_5p04310590878130_256x8m81_0/D w_n286_n142# a_193_n74#
Xpmos_5p04310590878130_256x8m81_0 w_n286_n142# pmos_5p04310590878130_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878130_256x8m81_0/S a_193_n74# pmos_5p04310590878130_256x8m81
.ends

.subckt nmos_5p04310590878132_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt pmos_5p04310590878122_256x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$46281772_256x8m81 a_n31_n73# pmos_5p04310590878122_256x8m81_0/S
+ w_n286_n142# pmos_5p04310590878122_256x8m81_0/D a_193_n73# a_417_n73#
Xpmos_5p04310590878122_256x8m81_0 w_n286_n142# pmos_5p04310590878122_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878122_256x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310590878122_256x8m81
.ends

.subckt pmos_5p04310590878128_256x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
.ends

.subckt pmos_1p2$$45095980_256x8m81 pmos_5p04310590878128_256x8m81_0/S a_193_n74#
+ a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# pmos_5p04310590878128_256x8m81_0/D
+ a_1985_n74# a_1761_n74# a_417_n74# w_n286_n142# a_1537_n74# a_1313_n74#
Xpmos_5p04310590878128_256x8m81_0 w_n286_n142# pmos_5p04310590878128_256x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590878128_256x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310590878128_256x8m81
.ends

.subckt nmos_5p04310590878112_256x8m81 D a_0_n44# a_672_n44# S a_448_n44# a_224_n44#
+ VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_5p04310590878131_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_5p04310590878114_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46285868_256x8m81 pmos_5p04310590878114_256x8m81_0/D pmos_5p04310590878114_256x8m81_0/S
+ w_n286_n142# a_n31_n73#
Xpmos_5p04310590878114_256x8m81_0 w_n286_n142# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt pmos_5p04310590878137_256x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46282796_256x8m81 a_193_n74# pmos_5p04310590878137_256x8m81_0/D
+ a_865_n74# a_n31_n74# a_641_n74# a_417_n74# w_n286_n142# pmos_5p04310590878137_256x8m81_0/S
Xpmos_5p04310590878137_256x8m81_0 w_n286_n142# pmos_5p04310590878137_256x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590878137_256x8m81_0/S a_417_n74# a_193_n74#
+ pmos_5p04310590878137_256x8m81
.ends

.subckt nmos_5p04310590878134_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_1p2$$45101100_256x8m81 nmos_5p04310590878134_256x8m81_0/D a_193_n74#
+ a_865_n74# a_n31_n74# a_641_n74# a_417_n74# nmos_5p04310590878134_256x8m81_0/S VSUBS
Xnmos_5p04310590878134_256x8m81_0 nmos_5p04310590878134_256x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590878134_256x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310590878134_256x8m81
.ends

.subckt pmos_5p04310590878113_256x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46286892_256x8m81 a_193_n73# pmos_5p04310590878113_256x8m81_0/D
+ a_n31_n73# a_417_n73# w_n286_n142# pmos_5p04310590878113_256x8m81_0/S
Xpmos_5p04310590878113_256x8m81_0 w_n286_n142# pmos_5p04310590878113_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878113_256x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310590878113_256x8m81
.ends

.subckt sacntl_2_256x8m81 pcb men a_4718_983# pmos_5p04310590878125_256x8m81_1/S nmos_5p04310590878123_256x8m81_1/D
+ pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D a_4560_1922# a_2796_670#
+ pmos_5p04310590878125_256x8m81_2/S se vss vdd
Xnmos_1p2$$45102124_256x8m81_0 pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ vss pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pcb pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ vss nmos_1p2$$45102124_256x8m81
Xpmos_5p04310590878138_256x8m81_0 vdd vdd pmos_5p04310590878125_256x8m81_0/S pmos_5p04310590878138_256x8m81_0/S
+ pmos_5p04310590878138_256x8m81
Xnmos_5p04310590878126_256x8m81_0 nmos_5p04310590878126_256x8m81_1/D nmos_5p04310590878131_256x8m81_0/D
+ nmos_5p04310590878131_256x8m81_0/D nmos_5p04310590878131_256x8m81_0/D vss nmos_5p04310590878131_256x8m81_0/D
+ nmos_5p04310590878131_256x8m81_0/D vss nmos_5p04310590878126_256x8m81
Xnmos_5p04310590878126_256x8m81_1 nmos_5p04310590878126_256x8m81_1/D pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ nmos_5p04310590878126_256x8m81_1/S pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D vss nmos_5p04310590878126_256x8m81
Xnmos_1p2$$45103148_256x8m81_0 pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S
+ nmos_5p04310590878133_256x8m81_0/D nmos_5p04310590878133_256x8m81_0/D vss pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D nmos_5p04310590878126_256x8m81_1/S
+ nmos_5p04310590878126_256x8m81_1/S vss nmos_1p2$$45103148_256x8m81
Xpmos_1p2$$46283820_256x8m81_0 pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pcb vdd pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S vdd pmos_1p2$$46283820_256x8m81
Xnmos_1p2$$45100076_256x8m81_0 pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S
+ vss vss nmos_1p2$$45100076_256x8m81
Xpmos_5p04310590878125_256x8m81_0 vdd vdd a_2796_670# pmos_5p04310590878125_256x8m81_0/S
+ pmos_5p04310590878125_256x8m81_0/S pmos_5p04310590878125_256x8m81
Xpmos_5p04310590878125_256x8m81_1 vdd vdd pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_5p04310590878125_256x8m81_1/S vss pmos_5p04310590878125_256x8m81
Xpmos_5p04310590878125_256x8m81_2 vdd vdd pmos_5p04310590878125_256x8m81_1/S pmos_5p04310590878125_256x8m81_2/S
+ pmos_5p04310590878125_256x8m81_2/S pmos_5p04310590878125_256x8m81
Xnmos_5p04310590878133_256x8m81_0 nmos_5p04310590878133_256x8m81_0/D pmos_5p04310590878125_256x8m81_1/S
+ vss vss nmos_5p04310590878133_256x8m81
Xnmos_5p04310590878123_256x8m81_0 vss a_2796_670# pmos_5p04310590878125_256x8m81_0/S
+ pmos_5p04310590878125_256x8m81_0/S vss nmos_5p04310590878123_256x8m81
Xnmos_5p04310590878123_256x8m81_1 nmos_5p04310590878123_256x8m81_1/D pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_5p04310590878125_256x8m81_1/S vss vss nmos_5p04310590878123_256x8m81
Xpmos_1p2$$46287916_256x8m81_0 nmos_5p04310590878131_256x8m81_0/D nmos_5p04310590878133_256x8m81_0/D
+ vdd nmos_5p04310590878133_256x8m81_0/D vdd pmos_1p2$$46287916_256x8m81
Xnmos_5p04310590878123_256x8m81_2 vss pmos_5p04310590878125_256x8m81_1/S pmos_5p04310590878125_256x8m81_2/S
+ pmos_5p04310590878125_256x8m81_2/S vss nmos_5p04310590878123_256x8m81
Xpmos_1p2$$46284844_256x8m81_0 pmos_5p04310590878125_256x8m81_1/S vdd nmos_5p04310590878133_256x8m81_0/D
+ vdd pmos_5p04310590878125_256x8m81_1/S pmos_1p2$$46284844_256x8m81
Xnmos_5p04310590878132_256x8m81_0 vss pmos_5p04310590878125_256x8m81_0/S pmos_5p04310590878138_256x8m81_0/S
+ vss nmos_5p04310590878132_256x8m81
Xpmos_1p2$$46281772_256x8m81_0 pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_0/pmos_5p04310590878122_256x8m81_0/S vdd vdd pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S
+ pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S pmos_1p2$$46281772_256x8m81
Xpmos_1p2$$46281772_256x8m81_1 pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_1p2$$46281772_256x8m81_1/pmos_5p04310590878122_256x8m81_0/S vdd vdd nmos_5p04310590878133_256x8m81_0/D
+ nmos_5p04310590878126_256x8m81_1/S pmos_1p2$$46281772_256x8m81
Xpmos_1p2$$45095980_256x8m81_0 vdd nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S
+ nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S
+ se nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S
+ vdd nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S pmos_1p2$$45095980_256x8m81
Xnmos_5p04310590878112_256x8m81_0 se nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S
+ vss nmos_5p04310590878126_256x8m81_1/S nmos_5p04310590878126_256x8m81_1/S vss nmos_5p04310590878112_256x8m81
Xnmos_5p04310590878131_256x8m81_0 nmos_5p04310590878131_256x8m81_0/D nmos_5p04310590878133_256x8m81_0/D
+ vss nmos_5p04310590878133_256x8m81_0/D vss nmos_5p04310590878131_256x8m81
Xpmos_1p2$$46285868_256x8m81_0 vdd nmos_5p04310590878126_256x8m81_1/S vdd pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ pmos_1p2$$46285868_256x8m81
Xpmos_1p2$$46282796_256x8m81_0 men pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ men men men men vdd vdd pmos_1p2$$46282796_256x8m81
Xnmos_1p2$$45101100_256x8m81_0 pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ men men men men men vss vss nmos_1p2$$45101100_256x8m81
Xpmos_1p2$$46286892_256x8m81_0 nmos_5p04310590878131_256x8m81_0/D nmos_5p04310590878126_256x8m81_1/S
+ nmos_5p04310590878131_256x8m81_0/D nmos_5p04310590878131_256x8m81_0/D vdd vdd pmos_1p2$$46286892_256x8m81
.ends

.subckt nmos_5p0431059087812_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.81u l=0.6u
.ends

.subckt nmos_1p2$$47119404_256x8m81 nmos_5p0431059087812_256x8m81_0/S nmos_5p0431059087812_256x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p0431059087812_256x8m81_0 nmos_5p0431059087812_256x8m81_0/D a_n31_n74# nmos_5p0431059087812_256x8m81_0/S
+ VSUBS nmos_5p0431059087812_256x8m81
.ends

.subckt nmos_5p0431059087811_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.57u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.57u l=0.6u
.ends

.subckt ypass_gate_a_256x8m81 d pcb b bb db ypass a_222_11191# a_n4_11191# vdd m3_n1_4331#
+ a_447_11191# vss a_n80_n10# a_222_10416# m3_n1_1708# a_n4_10416# m3_n1_1160# m3_n1_2030#
+ pmos_5p0431059087810_256x8m81_1/D m3_n1_3366# a_447_10416# m3_n1_2352# m3_n1_3688#
+ m3_n1_4009# m3_n1_2674#
Xpmos_1p2$$46889004_256x8m81_0 d vdd nmos_5p0431059087811_256x8m81_0/D b pmos_1p2$$46889004_256x8m81
Xpmos_5p0431059087810_256x8m81_0 vdd b pcb bb pmos_5p0431059087810_256x8m81
Xpmos_5p0431059087810_256x8m81_1 vdd pmos_5p0431059087810_256x8m81_1/D nmos_5p0431059087811_256x8m81_0/D
+ bb pmos_5p0431059087810_256x8m81
Xnmos_1p2$$47119404_256x8m81_0 b d ypass vss nmos_1p2$$47119404_256x8m81
Xnmos_1p2$$47119404_256x8m81_1 bb pmos_5p0431059087810_256x8m81_1/D ypass vss nmos_1p2$$47119404_256x8m81
Xnmos_5p0431059087811_256x8m81_0 nmos_5p0431059087811_256x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059087811_256x8m81
X0 nmos_5p0431059087811_256x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd ypass nmos_5p0431059087811_256x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X2 a_447_11191# pcb a_222_11191# vdd pmos_3p3 w=3.41u l=0.6u
X3 a_222_11191# pcb a_n4_11191# vdd pmos_3p3 w=3.41u l=0.6u
X4 a_447_10416# pcb a_222_10416# vdd pmos_3p3 w=3.41u l=0.6u
X5 a_222_10416# pcb a_n4_10416# vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt ypass_gate_256x8m81 d pcb bb db ypass vdd m3_n1_4331# vss b m3_n1_1708# m3_n1_1160#
+ m3_n1_2030# m3_n1_3366# m3_n1_2352# m3_n1_3688# m3_n1_4009# m3_n1_2674#
Xpmos_1p2$$46889004_256x8m81_0 d vdd nmos_5p0431059087811_256x8m81_0/D b pmos_1p2$$46889004_256x8m81
Xpmos_5p0431059087810_256x8m81_0 vdd b pcb bb pmos_5p0431059087810_256x8m81
Xpmos_5p0431059087810_256x8m81_1 vdd db nmos_5p0431059087811_256x8m81_0/D bb pmos_5p0431059087810_256x8m81
Xnmos_1p2$$47119404_256x8m81_0 b d ypass vss nmos_1p2$$47119404_256x8m81
Xnmos_1p2$$47119404_256x8m81_1 bb db ypass vss nmos_1p2$$47119404_256x8m81
Xnmos_5p0431059087811_256x8m81_0 nmos_5p0431059087811_256x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059087811_256x8m81
X0 nmos_5p0431059087811_256x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd ypass nmos_5p0431059087811_256x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt mux821_256x8m81 ypass_gate_a_256x8m81_0/a_447_11191# ypass_gate_256x8m81_4/ypass
+ a_656_7735# ypass_gate_256x8m81_5/ypass ypass_gate_256x8m81_5/d ypass_gate_256x8m81_6/ypass
+ ypass_gate_256x8m81_6/db ypass_gate_a_256x8m81_0/ypass ypass_gate_256x8m81_4/db
+ ypass_gate_256x8m81_6/m3_n1_4331# ypass_gate_a_256x8m81_0/a_222_10416# ypass_gate_256x8m81_0/d
+ ypass_gate_256x8m81_2/d ypass_gate_a_256x8m81_0/a_447_10416# ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_5/db ypass_gate_256x8m81_4/d ypass_gate_256x8m81_6/m3_n1_2030#
+ ypass_gate_256x8m81_6/d ypass_gate_256x8m81_6/m3_n1_3366# ypass_gate_256x8m81_6/m3_n1_2352#
+ ypass_gate_256x8m81_4/b a_4992_424# ypass_gate_a_256x8m81_0/a_222_11191# ypass_gate_256x8m81_6/m3_n1_3688#
+ ypass_gate_a_256x8m81_0/a_n80_n10# ypass_gate_a_256x8m81_0/d ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81_1/db ypass_gate_a_256x8m81_0/b
+ ypass_gate_256x8m81_0/ypass ypass_gate_256x8m81_1/d ypass_gate_256x8m81_1/ypass
+ ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_2/ypass ypass_gate_256x8m81_6/vdd
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_3/ypass ypass_gate_256x8m81_3/d
Xypass_gate_a_256x8m81_0 ypass_gate_a_256x8m81_0/d ypass_gate_256x8m81_6/pcb ypass_gate_a_256x8m81_0/b
+ ypass_gate_a_256x8m81_0/bb ypass_gate_a_256x8m81_0/db ypass_gate_a_256x8m81_0/ypass
+ ypass_gate_a_256x8m81_0/a_222_11191# ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/vdd
+ ypass_gate_256x8m81_6/m3_n1_4331# ypass_gate_a_256x8m81_0/a_447_11191# ypass_gate_256x8m81_6/vss
+ ypass_gate_a_256x8m81_0/a_n80_n10# ypass_gate_a_256x8m81_0/a_222_10416# ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030#
+ ypass_gate_256x8m81_1/db ypass_gate_256x8m81_6/m3_n1_3366# ypass_gate_a_256x8m81_0/a_447_10416#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_a_256x8m81
Xypass_gate_256x8m81_0 ypass_gate_256x8m81_0/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_0/bb
+ ypass_gate_256x8m81_4/db ypass_gate_256x8m81_0/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_0/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_1 ypass_gate_256x8m81_1/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_1/bb
+ ypass_gate_256x8m81_1/db ypass_gate_256x8m81_1/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_1/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_2 ypass_gate_256x8m81_2/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_2/bb
+ ypass_gate_256x8m81_5/db ypass_gate_256x8m81_2/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_2/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_3 ypass_gate_256x8m81_3/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_3/bb
+ ypass_gate_256x8m81_6/db ypass_gate_256x8m81_3/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_3/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_4 ypass_gate_256x8m81_4/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_4/bb
+ ypass_gate_256x8m81_4/db ypass_gate_256x8m81_4/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_4/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_5 ypass_gate_256x8m81_5/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_5/bb
+ ypass_gate_256x8m81_5/db ypass_gate_256x8m81_5/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_5/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
Xypass_gate_256x8m81_6 ypass_gate_256x8m81_6/d ypass_gate_256x8m81_6/pcb ypass_gate_256x8m81_6/bb
+ ypass_gate_256x8m81_6/db ypass_gate_256x8m81_6/ypass ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_4331#
+ ypass_gate_256x8m81_6/vss ypass_gate_256x8m81_6/b ypass_gate_256x8m81_6/m3_n1_1708#
+ ypass_gate_256x8m81_6/vdd ypass_gate_256x8m81_6/m3_n1_2030# ypass_gate_256x8m81_6/m3_n1_3366#
+ ypass_gate_256x8m81_6/m3_n1_2352# ypass_gate_256x8m81_6/m3_n1_3688# ypass_gate_256x8m81_6/m3_n1_4009#
+ ypass_gate_256x8m81_6/m3_n1_2674# ypass_gate_256x8m81
.ends

.subckt nmos_5p04310590878140_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.37u l=0.6u
.ends

.subckt nmos_1p2$$202594348_256x8m81 nmos_5p04310590878140_256x8m81_0/S a_n31_n73#
+ nmos_5p04310590878140_256x8m81_0/D VSUBS
Xnmos_5p04310590878140_256x8m81_0 nmos_5p04310590878140_256x8m81_0/D a_n31_n73# nmos_5p04310590878140_256x8m81_0/S
+ VSUBS nmos_5p04310590878140_256x8m81
.ends

.subckt nmos_1p2$$202598444_256x8m81 nmos_5p04310590878110_256x8m81_0/D a_n31_n74#
+ nmos_5p04310590878110_256x8m81_0/S VSUBS
Xnmos_5p04310590878110_256x8m81_0 nmos_5p04310590878110_256x8m81_0/D a_n31_n74# nmos_5p04310590878110_256x8m81_0/S
+ VSUBS nmos_5p04310590878110_256x8m81
.ends

.subckt nmos_1p2$$202595372_256x8m81 nmos_5p0431059087818_256x8m81_0/D a_n31_n73#
+ nmos_5p0431059087818_256x8m81_0/S VSUBS
Xnmos_5p0431059087818_256x8m81_0 nmos_5p0431059087818_256x8m81_0/D a_n31_n73# nmos_5p0431059087818_256x8m81_0/S
+ VSUBS nmos_5p0431059087818_256x8m81
.ends

.subckt nmos_1p2$$202596396_256x8m81 nmos_5p0431059087818_256x8m81_0/D a_n31_n73#
+ nmos_5p0431059087818_256x8m81_0/S VSUBS
Xnmos_5p0431059087818_256x8m81_0 nmos_5p0431059087818_256x8m81_0/D a_n31_n73# nmos_5p0431059087818_256x8m81_0/S
+ VSUBS nmos_5p0431059087818_256x8m81
.ends

.subckt pmos_1p2$$202584108_256x8m81 pmos_5p04310590878114_256x8m81_0/D a_n31_n74#
+ pmos_5p04310590878114_256x8m81_0/S w_n286_n141#
Xpmos_5p04310590878114_256x8m81_0 w_n286_n141# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt nmos_5p04310590878142_256x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.8u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
.ends

.subckt pmos_5p04310590878143_256x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_1p2$$202585132_256x8m81 pmos_5p04310590878114_256x8m81_0/D w_n256_n141#
+ pmos_5p04310590878114_256x8m81_0/S a_n31_n74#
Xpmos_5p04310590878114_256x8m81_0 w_n256_n141# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt pmos_5p04310590878141_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_1p2$$202586156_256x8m81 pmos_5p04310590878114_256x8m81_0/D pmos_5p04310590878114_256x8m81_0/S
+ w_n286_n141# a_n31_n74#
Xpmos_5p04310590878114_256x8m81_0 w_n286_n141# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt pmos_1p2$$202583084_256x8m81 pmos_5p04310590878130_256x8m81_0/S a_193_n74#
+ pmos_5p04310590878130_256x8m81_0/D w_n286_n142# a_n31_n74#
Xpmos_5p04310590878130_256x8m81_0 w_n286_n142# pmos_5p04310590878130_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878130_256x8m81_0/S a_193_n74# pmos_5p04310590878130_256x8m81
.ends

.subckt pmos_5p04310590878120_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$202587180_256x8m81 pmos_5p04310590878114_256x8m81_0/D pmos_5p04310590878114_256x8m81_0/S
+ w_n286_n141# a_n31_n74#
Xpmos_5p04310590878114_256x8m81_0 w_n286_n141# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt nmos_5p04310590878139_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt wen_wm1_256x8m81 wep wen GWEN men vdd vss
Xnmos_1p2$$202594348_256x8m81_0 pmos_1p2$$202583084_256x8m81_0/pmos_5p04310590878130_256x8m81_0/D
+ nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D vss vss nmos_1p2$$202594348_256x8m81
Xnmos_5p0431059087818_256x8m81_0 vss GWEN nmos_5p0431059087818_256x8m81_2/D vss nmos_5p0431059087818_256x8m81
Xnmos_1p2$$202598444_256x8m81_0 pmos_5p04310590878141_256x8m81_0/S pmos_5p04310590878114_256x8m81_4/D
+ nmos_5p0431059087818_256x8m81_1/D vss nmos_1p2$$202598444_256x8m81
Xnmos_5p0431059087818_256x8m81_1 nmos_5p0431059087818_256x8m81_1/D nmos_5p0431059087818_256x8m81_2/D
+ vss vss nmos_5p0431059087818_256x8m81
Xnmos_1p2$$202595372_256x8m81_0 pmos_5p04310590878141_256x8m81_0/D nmos_5p0431059087818_256x8m81_3/D
+ pmos_5p04310590878141_256x8m81_0/S vss nmos_1p2$$202595372_256x8m81
Xnmos_1p2$$202595372_256x8m81_1 vss pmos_5p04310590878141_256x8m81_0/S nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ vss nmos_1p2$$202595372_256x8m81
Xnmos_5p0431059087818_256x8m81_2 nmos_5p0431059087818_256x8m81_2/D wen vss vss nmos_5p0431059087818_256x8m81
Xnmos_5p0431059087818_256x8m81_3 nmos_5p0431059087818_256x8m81_3/D pmos_5p04310590878114_256x8m81_4/D
+ vss vss nmos_5p0431059087818_256x8m81
Xnmos_1p2$$202596396_256x8m81_0 nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S vss vss nmos_1p2$$202596396_256x8m81
Xnmos_1p2$$202596396_256x8m81_1 vss nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ pmos_5p04310590878141_256x8m81_0/D vss nmos_1p2$$202596396_256x8m81
Xpmos_1p2$$202584108_256x8m81_0 vdd pmos_5p04310590878141_256x8m81_0/S nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ vdd pmos_1p2$$202584108_256x8m81
Xpmos_5p04310590878114_256x8m81_0 vdd pmos_5p04310590878114_256x8m81_2/S wen vdd pmos_5p04310590878114_256x8m81
Xnmos_5p04310590878142_256x8m81_0 wep pmos_5p04310590878130_256x8m81_0/D vss pmos_5p04310590878130_256x8m81_0/D
+ pmos_5p04310590878130_256x8m81_0/D vss nmos_5p04310590878142_256x8m81
Xpmos_5p04310590878143_256x8m81_0 vdd wep pmos_5p04310590878130_256x8m81_0/D vdd pmos_5p04310590878130_256x8m81_0/D
+ pmos_5p04310590878130_256x8m81_0/D pmos_5p04310590878143_256x8m81
Xpmos_5p04310590878114_256x8m81_1 vdd nmos_5p0431059087818_256x8m81_1/D nmos_5p0431059087818_256x8m81_2/D
+ vdd pmos_5p04310590878114_256x8m81
Xpmos_1p2$$202585132_256x8m81_0 nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ vdd vdd nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S pmos_1p2$$202585132_256x8m81
Xpmos_5p04310590878114_256x8m81_2 vdd nmos_5p0431059087818_256x8m81_2/D GWEN pmos_5p04310590878114_256x8m81_2/S
+ pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_3 vdd nmos_5p0431059087818_256x8m81_3/D pmos_5p04310590878114_256x8m81_4/D
+ vdd pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_4 vdd pmos_5p04310590878114_256x8m81_4/D vss pmos_5p04310590878114_256x8m81_5/D
+ pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_5 vdd pmos_5p04310590878114_256x8m81_5/D men vdd pmos_5p04310590878114_256x8m81
Xnmos_5p04310590878140_256x8m81_0 pmos_5p04310590878130_256x8m81_0/D pmos_5p04310590878120_256x8m81_0/S
+ vss vss nmos_5p04310590878140_256x8m81
Xpmos_5p04310590878141_256x8m81_0 vdd pmos_5p04310590878141_256x8m81_0/D pmos_5p04310590878114_256x8m81_4/D
+ pmos_5p04310590878141_256x8m81_0/S pmos_5p04310590878141_256x8m81
Xnmos_5p04310590878140_256x8m81_1 pmos_5p04310590878114_256x8m81_4/D men vss vss nmos_5p04310590878140_256x8m81
Xnmos_5p04310590878140_256x8m81_2 vss vss pmos_5p04310590878114_256x8m81_4/D vss nmos_5p04310590878140_256x8m81
Xpmos_1p2$$202586156_256x8m81_0 vdd pmos_5p04310590878141_256x8m81_0/D vdd nmos_1p2$$202595372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ pmos_1p2$$202586156_256x8m81
Xnmos_5p04310590878110_256x8m81_0 vss nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ pmos_5p04310590878120_256x8m81_0/S vss nmos_5p04310590878110_256x8m81
Xpmos_1p2$$202583084_256x8m81_0 vdd nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ pmos_1p2$$202583084_256x8m81_0/pmos_5p04310590878130_256x8m81_0/D vdd nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ pmos_1p2$$202583084_256x8m81
Xpmos_5p04310590878130_256x8m81_0 vdd pmos_5p04310590878130_256x8m81_0/D pmos_5p04310590878120_256x8m81_0/S
+ vdd pmos_5p04310590878120_256x8m81_0/S pmos_5p04310590878130_256x8m81
Xpmos_5p04310590878120_256x8m81_0 vdd men nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ pmos_5p04310590878120_256x8m81_0/S nmos_1p2$$202596396_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ pmos_5p04310590878120_256x8m81
Xpmos_1p2$$202587180_256x8m81_0 pmos_5p04310590878141_256x8m81_0/S nmos_5p0431059087818_256x8m81_1/D
+ vdd nmos_5p0431059087818_256x8m81_3/D pmos_1p2$$202587180_256x8m81
Xnmos_5p04310590878139_256x8m81_0 men pmos_1p2$$202583084_256x8m81_0/pmos_5p04310590878130_256x8m81_0/D
+ pmos_5p04310590878120_256x8m81_0/S pmos_1p2$$202583084_256x8m81_0/pmos_5p04310590878130_256x8m81_0/D
+ vss nmos_5p04310590878139_256x8m81
.ends

.subckt pmos_5p04310590878148_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.5u l=0.6u
.ends

.subckt nmos_5p04310590878146_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
.ends

.subckt pmos_5p04310590878147_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4u l=0.6u
.ends

.subckt pmos_1p2$$171625516_256x8m81 pmos_5p0431059087813_256x8m81_0/S a_193_n74#
+ w_n286_n142# pmos_5p0431059087813_256x8m81_0/D pmos_5p0431059087813_256x8m81_0/w_n208_n120#
+ a_n31_n74#
Xpmos_5p0431059087813_256x8m81_0 pmos_5p0431059087813_256x8m81_0/w_n208_n120# pmos_5p0431059087813_256x8m81_0/D
+ a_n31_n74# pmos_5p0431059087813_256x8m81_0/S a_193_n74# pmos_5p0431059087813_256x8m81
.ends

.subckt nmos_5p04310590878145_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310590878144_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310590878152_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.6u l=0.6u
.ends

.subckt nmos_5p04310590878150_256x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310590878151_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.67u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_5p04310590878149_256x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
.ends

.subckt outbuf_oe_256x8m81 se q GWE qp qn a_4913_n316# vdd vss
Xpmos_5p04310590878148_256x8m81_0 vdd vdd pmos_5p04310590878147_256x8m81_0/S pmos_5p04310590878148_256x8m81_0/S
+ pmos_5p04310590878148_256x8m81
Xpmos_5p04310590878138_256x8m81_0 vdd pmos_5p04310590878138_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ vdd pmos_5p04310590878138_256x8m81
Xnmos_5p0431059087818_256x8m81_0 nmos_5p0431059087818_256x8m81_0/D se vss vss nmos_5p0431059087818_256x8m81
Xnmos_5p04310590878146_256x8m81_0 vss pmos_5p04310590878151_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ pmos_5p04310590878151_256x8m81_0/D q pmos_5p04310590878151_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ pmos_5p04310590878151_256x8m81_0/D vss nmos_5p04310590878146_256x8m81
Xpmos_5p04310590878147_256x8m81_0 vdd vdd GWE pmos_5p04310590878147_256x8m81_0/S pmos_5p04310590878147_256x8m81
Xnmos_5p0431059087818_256x8m81_1 vss pmos_5p04310590878138_256x8m81_0/D nmos_5p0431059087818_256x8m81_1/S
+ vss nmos_5p0431059087818_256x8m81
Xpmos_1p2$$171625516_256x8m81_0 vdd pmos_5p04310590878138_256x8m81_0/D vdd nmos_5p0431059087818_256x8m81_1/S
+ vdd pmos_5p04310590878138_256x8m81_0/D pmos_1p2$$171625516_256x8m81
Xnmos_5p04310590878145_256x8m81_0 vss pmos_5p04310590878147_256x8m81_0/S nmos_5p04310590878145_256x8m81_1/S
+ pmos_5p04310590878147_256x8m81_0/S vss nmos_5p04310590878145_256x8m81
Xnmos_5p04310590878145_256x8m81_1 pmos_5p04310590878151_256x8m81_0/D qn nmos_5p04310590878145_256x8m81_1/S
+ qn vss nmos_5p04310590878145_256x8m81
Xnmos_5p04310590878144_256x8m81_0 vss pmos_5p04310590878147_256x8m81_0/S pmos_5p04310590878148_256x8m81_0/S
+ vss nmos_5p04310590878144_256x8m81
Xpmos_5p04310590878114_256x8m81_0 vdd nmos_5p0431059087818_256x8m81_0/D se vdd pmos_5p04310590878114_256x8m81
Xnmos_5p04310590878152_256x8m81_0 vss GWE pmos_5p04310590878147_256x8m81_0/S vss nmos_5p04310590878152_256x8m81
Xnmos_5p04310590878132_256x8m81_0 pmos_5p04310590878138_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ vss vss nmos_5p04310590878132_256x8m81
Xpmos_5p04310590878113_256x8m81_0 vdd nmos_5p0431059087818_256x8m81_1/S se pmos_5p04310590878151_256x8m81_0/D
+ se se pmos_5p04310590878113_256x8m81
Xnmos_5p04310590878150_256x8m81_0 nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_0/D
+ pmos_5p04310590878151_256x8m81_0/D nmos_5p0431059087818_256x8m81_0/D nmos_5p0431059087818_256x8m81_0/D
+ vss nmos_5p04310590878150_256x8m81
Xpmos_5p04310590878151_256x8m81_0 vdd pmos_5p04310590878151_256x8m81_0/D qp pmos_5p04310590878151_256x8m81_1/S
+ qp pmos_5p04310590878151_256x8m81
Xpmos_5p04310590878151_256x8m81_1 vdd vdd pmos_5p04310590878148_256x8m81_0/S pmos_5p04310590878151_256x8m81_1/S
+ pmos_5p04310590878148_256x8m81_0/S pmos_5p04310590878151_256x8m81
Xpmos_5p04310590878149_256x8m81_0 vdd vdd pmos_5p04310590878151_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ pmos_5p04310590878151_256x8m81_0/D q pmos_5p04310590878151_256x8m81_0/D pmos_5p04310590878151_256x8m81_0/D
+ pmos_5p04310590878151_256x8m81_0/D pmos_5p04310590878149_256x8m81
.ends

.subckt pmos_5p04310590878119_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46898220_256x8m81 pmos_5p04310590878119_256x8m81_0/D pmos_5p04310590878119_256x8m81_0/S
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310590878119_256x8m81_0 w_n286_n142# pmos_5p04310590878119_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878119_256x8m81_0/S pmos_5p04310590878119_256x8m81
.ends

.subckt pmos_5p04310590878121_256x8m81 w_n208_n120# D a_0_n44# a_672_n44# S a_448_n44#
+ a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46896172_256x8m81 pmos_5p04310590878121_256x8m81_0/D a_668_n74#
+ a_193_n74# pmos_5p04310590878121_256x8m81_0/S w_n286_n142# a_n31_n74# a_417_n74#
Xpmos_5p04310590878121_256x8m81_0 w_n286_n142# pmos_5p04310590878121_256x8m81_0/D
+ a_n31_n74# a_668_n74# pmos_5p04310590878121_256x8m81_0/S a_417_n74# a_193_n74# pmos_5p04310590878121_256x8m81
.ends

.subckt nmos_1p2$$45107244_256x8m81 a_193_n73# a_n31_n73# a_641_n73# nmos_5p04310590878112_256x8m81_0/S
+ a_417_n73# nmos_5p04310590878112_256x8m81_0/D VSUBS
Xnmos_5p04310590878112_256x8m81_0 nmos_5p04310590878112_256x8m81_0/D a_n31_n73# a_641_n73#
+ nmos_5p04310590878112_256x8m81_0/S a_417_n73# a_193_n73# VSUBS nmos_5p04310590878112_256x8m81
.ends

.subckt pmos_5p04310590878118_256x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46549036_256x8m81 pmos_5p04310590878118_256x8m81_0/D a_193_n74#
+ w_n286_n142# a_1089_n74# a_865_n74# a_n31_n74# pmos_5p04310590878118_256x8m81_0/S
+ a_641_n74# a_417_n74#
Xpmos_5p04310590878118_256x8m81_0 w_n286_n142# pmos_5p04310590878118_256x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590878118_256x8m81_0/S a_417_n74# a_193_n74#
+ a_1089_n74# pmos_5p04310590878118_256x8m81
.ends

.subckt pmos_1p2$$46897196_256x8m81 pmos_5p04310590878120_256x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310590878120_256x8m81_0/S
Xpmos_5p04310590878120_256x8m81_0 w_n286_n142# pmos_5p04310590878120_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878120_256x8m81_0/S a_193_n74# pmos_5p04310590878120_256x8m81
.ends

.subckt nmos_5p04310590878116_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46552108_256x8m81 nmos_5p04310590878116_256x8m81_0/D a_1089_n74#
+ a_865_n74# a_641_n74# a_n31_n74# a_1537_n74# a_1313_n74# nmos_5p04310590878116_256x8m81_0/S
+ a_417_n74# a_193_n74# VSUBS
Xnmos_5p04310590878116_256x8m81_0 nmos_5p04310590878116_256x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590878116_256x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310590878116_256x8m81
.ends

.subckt nmos_5p04310590878115_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46553132_256x8m81 nmos_5p04310590878115_256x8m81_0/D a_n31_n74#
+ nmos_5p04310590878115_256x8m81_0/S VSUBS
Xnmos_5p04310590878115_256x8m81_0 nmos_5p04310590878115_256x8m81_0/D a_n31_n74# nmos_5p04310590878115_256x8m81_0/S
+ VSUBS nmos_5p04310590878115_256x8m81
.ends

.subckt nmos_5p04310590878117_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_1p2$$46550060_256x8m81 a_1537_n74# a_1313_n74# nmos_5p04310590878117_256x8m81_0/S
+ a_193_n74# a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# nmos_5p04310590878117_256x8m81_0/D
+ a_417_n74# VSUBS
Xnmos_5p04310590878117_256x8m81_0 nmos_5p04310590878117_256x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590878117_256x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310590878117_256x8m81
.ends

.subckt nmos_1p2$$46551084_256x8m81 nmos_5p04310590878110_256x8m81_0/D a_n31_n73#
+ nmos_5p04310590878110_256x8m81_0/S VSUBS
Xnmos_5p04310590878110_256x8m81_0 nmos_5p04310590878110_256x8m81_0/D a_n31_n73# nmos_5p04310590878110_256x8m81_0/S
+ VSUBS nmos_5p04310590878110_256x8m81
.ends

.subckt sa_256x8m81 wep se pcb qp vss d
Xpmos_1p2$$46898220_256x8m81_0 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ d d d pmos_1p2$$46898220_256x8m81
Xpmos_1p2$$46898220_256x8m81_1 d pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ d d pmos_1p2$$46898220_256x8m81
Xpmos_1p2$$46896172_256x8m81_0 d pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ d pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46896172_256x8m81
Xnmos_1p2$$45107244_256x8m81_0 qp pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ qp qp qp vss vss nmos_1p2$$45107244_256x8m81
Xpmos_1p2$$46549036_256x8m81_0 qp pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ d pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S d qp qp pmos_1p2$$46549036_256x8m81
Xpmos_1p2$$46897196_256x8m81_0 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ se d se d pmos_1p2$$46897196_256x8m81
Xnmos_1p2$$46552108_256x8m81_0 nmos_1p2$$46552108_256x8m81_0/nmos_5p04310590878116_256x8m81_0/D
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S vss nmos_1p2$$46552108_256x8m81
Xpmos_1p2$$46897196_256x8m81_1 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ se d se d pmos_1p2$$46897196_256x8m81
Xpmos_1p2$$46897196_256x8m81_2 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ se d se d pmos_1p2$$46897196_256x8m81
Xpmos_1p2$$46897196_256x8m81_3 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ se d se d pmos_1p2$$46897196_256x8m81
Xnmos_1p2$$46553132_256x8m81_0 vss vss pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ vss nmos_1p2$$46553132_256x8m81
Xnmos_1p2$$46550060_256x8m81_0 se se vss se se se se se nmos_1p2$$46552108_256x8m81_0/nmos_5p04310590878116_256x8m81_0/D
+ se vss nmos_1p2$$46550060_256x8m81
Xnmos_1p2$$46553132_256x8m81_1 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_256x8m81
Xpmos_1p2$$46285868_256x8m81_0 pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S d pcb pmos_1p2$$46285868_256x8m81
Xpmos_1p2$$46286892_256x8m81_0 pcb d pcb pcb d d pmos_1p2$$46286892_256x8m81
Xnmos_1p2$$46551084_256x8m81_0 vss pmos_1p2$$46898220_256x8m81_1/pmos_5p04310590878119_256x8m81_0/S
+ qp vss nmos_1p2$$46551084_256x8m81
.ends

.subckt saout_R_m2_256x8m81 pcb datain WEN ypass[1] ypass[2] ypass[3] ypass[4] ypass[5]
+ ypass[6] ypass[7] ypass[0] GWE GWEN b[7] b[0] bb[5] q wen_wm1_256x8m81_0/wen mux821_256x8m81_0/a_656_7735#
+ mux821_256x8m81_0/ypass_gate_256x8m81_4/b b[2] b[6] bb[1] bb[3] b[5] bb[4] mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b
+ b[4] men a_5189_27169# a_5414_27169# bb[6] a_5189_27944# a_5414_27944# mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass
+ mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass sacntl_2_256x8m81_0/a_4560_1922#
+ outbuf_oe_256x8m81_0/a_4913_n316# bb[7] bb[0] mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass
+ sacntl_2_256x8m81_0/a_4718_983# wen_wm1_256x8m81_0/GWEN mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass wen_wm1_256x8m81_0/vdd sa_256x8m81_0/pcb
+ bb[2] b[3] mux821_256x8m81_0/ypass_gate_256x8m81_6/vdd mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass vdd mux821_256x8m81_0/a_4992_424#
+ sa_256x8m81_0/wep vss sacntl_2_256x8m81_0/vdd b[1] mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass
Xdin_256x8m81_0 datain sa_256x8m81_0/wep men vdd vdd sa_256x8m81_0/pcb vdd vdd vss
+ din_256x8m81
Xsacntl_2_256x8m81_0 sa_256x8m81_0/pcb men sacntl_2_256x8m81_0/a_4718_983# sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_1/S
+ vss sacntl_2_256x8m81_0/pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ sacntl_2_256x8m81_0/a_4560_1922# sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_2/S
+ sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_2/S sa_256x8m81_0/se vss sacntl_2_256x8m81_0/vdd
+ sacntl_2_256x8m81
Xmux821_256x8m81_0 a_5414_27944# mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass mux821_256x8m81_0/a_656_7735#
+ mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass
+ vdd mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass vdd mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass
+ a_5189_27169# vdd vdd a_5414_27169# mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass
+ vdd vdd mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ mux821_256x8m81_0/a_4992_424# a_5189_27944# mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass
+ mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10# vdd mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass vdd mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b
+ mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass
+ sa_256x8m81_0/pcb mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass mux821_256x8m81_0/ypass_gate_256x8m81_6/vdd
+ vss mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass vdd mux821_256x8m81
Xwen_wm1_256x8m81_0 sa_256x8m81_0/wep wen_wm1_256x8m81_0/wen wen_wm1_256x8m81_0/GWEN
+ men wen_wm1_256x8m81_0/vdd vss wen_wm1_256x8m81
Xoutbuf_oe_256x8m81_0 sa_256x8m81_0/se q GWE sa_256x8m81_0/qp sa_256x8m81_0/qp outbuf_oe_256x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_256x8m81
Xsa_256x8m81_0 sa_256x8m81_0/wep sa_256x8m81_0/se sa_256x8m81_0/pcb sa_256x8m81_0/qp
+ vss vdd sa_256x8m81
.ends

.subckt saout_m2_256x8m81 pcb datain WEN ypass[1] ypass[2] ypass[3] ypass[4] ypass[5]
+ ypass[6] ypass[7] ypass[0] GWEN GWE bb[2] b[0] q a_5189_27176# a_5414_27176# a_5189_27951#
+ a_5414_27951# mux821_256x8m81_0/a_656_7735# b[5] b[1] mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass
+ bb[6] bb[4] b[2] mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10# bb[3] b[3]
+ men bb[1] mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass sacntl_2_256x8m81_0/a_4560_1922#
+ outbuf_oe_256x8m81_0/a_4913_n316# bb[0] bb[7] mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass
+ sacntl_2_256x8m81_0/a_4718_983# wen_wm1_256x8m81_0/GWEN mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass wen_wm1_256x8m81_0/vdd b[7] bb[5]
+ sa_256x8m81_0/pcb b[4] mux821_256x8m81_0/ypass_gate_256x8m81_6/vdd sacntl_2_256x8m81_0/vdd
+ mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass
+ sa_256x8m81_0/wep mux821_256x8m81_0/a_4992_424# vss b[6] mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass
Xdin_256x8m81_0 datain sa_256x8m81_0/wep men vdd vdd sa_256x8m81_0/pcb vdd vdd vss
+ din_256x8m81
Xsacntl_2_256x8m81_0 sa_256x8m81_0/pcb men sacntl_2_256x8m81_0/a_4718_983# sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_1/S
+ vss sacntl_2_256x8m81_0/pmos_1p2$$46282796_256x8m81_0/pmos_5p04310590878137_256x8m81_0/D
+ sacntl_2_256x8m81_0/a_4560_1922# sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_2/S
+ sacntl_2_256x8m81_0/pmos_5p04310590878125_256x8m81_2/S sa_256x8m81_0/se vss sacntl_2_256x8m81_0/vdd
+ sacntl_2_256x8m81
Xmux821_256x8m81_0 a_5414_27951# mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass mux821_256x8m81_0/a_656_7735#
+ mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass
+ vdd mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass
+ a_5189_27176# vdd vdd a_5414_27176# mux821_256x8m81_0/ypass_gate_a_256x8m81_0/ypass
+ vdd vdd mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_5/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_4/ypass mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ mux821_256x8m81_0/a_4992_424# a_5189_27951# mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass
+ mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10# vdd mux821_256x8m81_0/ypass_gate_256x8m81_6/ypass
+ mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass vdd mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b
+ mux821_256x8m81_0/ypass_gate_256x8m81_0/ypass vdd mux821_256x8m81_0/ypass_gate_256x8m81_1/ypass
+ sa_256x8m81_0/pcb mux821_256x8m81_0/ypass_gate_256x8m81_2/ypass mux821_256x8m81_0/ypass_gate_256x8m81_6/vdd
+ vss mux821_256x8m81_0/ypass_gate_256x8m81_3/ypass vdd mux821_256x8m81
Xwen_wm1_256x8m81_0 sa_256x8m81_0/wep wen_wm1_256x8m81_0/wen wen_wm1_256x8m81_0/GWEN
+ men wen_wm1_256x8m81_0/vdd vss wen_wm1_256x8m81
Xoutbuf_oe_256x8m81_0 sa_256x8m81_0/se q GWE sa_256x8m81_0/qp sa_256x8m81_0/qp outbuf_oe_256x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_256x8m81
Xsa_256x8m81_0 sa_256x8m81_0/wep sa_256x8m81_0/se sa_256x8m81_0/pcb sa_256x8m81_0/qp
+ vss vdd sa_256x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_256x8m81 a_n36_52# a_444_n42# a_246_342# a_126_298#
+ m3_n36_330# a_36_n42# w_n68_622# VSUBS
X0 a_444_206# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_126_298# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_444_206# a_246_342# a_126_298# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_444_206# a_246_342# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_dummy_256x8m81 a_n36_52# m2_90_n50# a_246_342# m2_390_n50#
+ a_246_712# m3_n36_330# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt nmos_5p04310590878156_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.38u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.38u l=0.6u
.ends

.subckt nmos_5p04310590878154_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=8.5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=8.5u l=0.6u
.ends

.subckt pmos_5p04310590878155_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10.64u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.64u l=0.6u
.ends

.subckt pmos_5p04310590878153_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.51u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.51u l=0.6u
.ends

.subckt ypass_gate_256x8m81_0 pcb vss bb db ypass vdd m3_n1_4331# d pmos_5p0431059087810_256x8m81_2/D
+ m3_n1_1708# m3_n1_1160# m3_n1_2030# m3_n1_3366# m3_n1_2352# m3_n1_3688# m3_n1_4009#
+ m3_n1_2674# b a_66_539#
Xpmos_5p0431059087810_256x8m81_0 vdd d nmos_5p0431059087811_256x8m81_0/D b pmos_5p0431059087810_256x8m81
Xpmos_5p0431059087810_256x8m81_1 vdd b pcb bb pmos_5p0431059087810_256x8m81
Xpmos_5p0431059087810_256x8m81_2 vdd pmos_5p0431059087810_256x8m81_2/D nmos_5p0431059087811_256x8m81_0/D
+ bb pmos_5p0431059087810_256x8m81
Xnmos_5p0431059087812_256x8m81_0 pmos_5p0431059087810_256x8m81_2/D a_66_539# bb vss
+ nmos_5p0431059087812_256x8m81
Xnmos_5p0431059087812_256x8m81_1 d a_66_539# b vss nmos_5p0431059087812_256x8m81
Xnmos_5p0431059087811_256x8m81_0 nmos_5p0431059087811_256x8m81_0/D a_66_539# vss a_66_539#
+ vss nmos_5p0431059087811_256x8m81
X0 nmos_5p0431059087811_256x8m81_0/D a_66_539# vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd a_66_539# nmos_5p0431059087811_256x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt rdummy_256x4_a_256x8m81 pcb tblhl m3_117_16293# m3_117_15650# m3_117_15971#
+ m3_264_359# ypass_gate_256x8m81_0_0/d m3_117_13670# ypass_gate_256x8m81_0_0/bb w_523_3317#
+ ypass_gate_256x8m81_0_0/b m3_117_13992# m3_117_15328# vdd vss m3_117_14314# pmos_5p04310590878155_256x8m81_0/S
+ m3_117_14636#
Xnmos_5p04310590878156_256x8m81_0 pmos_5p04310590878153_256x8m81_0/D ypass_gate_256x8m81_0_0/d
+ vss ypass_gate_256x8m81_0_0/d vss nmos_5p04310590878156_256x8m81
Xnmos_5p04310590878154_256x8m81_0 tblhl pmos_5p04310590878153_256x8m81_0/D vss pmos_5p04310590878153_256x8m81_0/D
+ vss nmos_5p04310590878154_256x8m81
Xpmos_5p04310590878155_256x8m81_0 w_523_3317# tblhl pmos_5p04310590878153_256x8m81_0/D
+ pmos_5p04310590878155_256x8m81_0/S pmos_5p04310590878153_256x8m81_0/D pmos_5p04310590878155_256x8m81
Xpmos_5p04310590878153_256x8m81_0 vdd pmos_5p04310590878153_256x8m81_0/D ypass_gate_256x8m81_0_0/d
+ vdd ypass_gate_256x8m81_0_0/d pmos_5p04310590878153_256x8m81
Xypass_gate_256x8m81_0_0 ypass_gate_256x8m81_0_0/pcb vss ypass_gate_256x8m81_0_0/bb
+ ypass_gate_256x8m81_0_0/db ypass_gate_256x8m81_0_0/ypass vdd m3_117_16293# ypass_gate_256x8m81_0_0/d
+ ypass_gate_256x8m81_0_0/bb m3_117_13670# vdd m3_117_13992# m3_117_15328# m3_117_14314#
+ m3_117_15650# m3_117_15971# m3_117_14636# ypass_gate_256x8m81_0_0/b vdd ypass_gate_256x8m81_0
.ends

.subckt rdummy_256x4_256x8m81 018SRAM_cell1_dummy_R_256x8m81_11/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_41/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_4/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_51/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_12/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_5/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_16/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_13/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_61/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_22/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_5/a_246_342# 018SRAM_cell1_dummy_256x8m81_17/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_7/a_126_298# 018SRAM_cell1_dummy_R_256x8m81_14/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_32/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_7/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_18/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_15/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_42/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_50/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_20/a_246_342# a_28741_1594# 018SRAM_cell1_dummy_R_256x8m81_8/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_19/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_16/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_52/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_51/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_30/a_246_342#
+ 018SRAM_cell1_dummy_R_256x8m81_9/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_17/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_62/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_2/a_126_298#
+ 018SRAM_cell1_dummy_256x8m81_23/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_52/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_28/a_126_298# 018SRAM_cell1_dummy_256x8m81_53/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_18/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_33/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_11/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_19/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_54/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_43/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_21/a_246_342#
+ 018SRAM_cell1_dummy_R_256x8m81_7/w_n68_622# 018SRAM_cell1_dummy_256x8m81_55/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_53/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_31/a_246_342# 018SRAM_cell1_dummy_256x8m81_56/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_63/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_3/a_126_298#
+ 018SRAM_cell1_dummy_256x8m81_24/m2_90_n50# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_7/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_57/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_29/a_126_298#
+ 018SRAM_cell1_dummy_256x8m81_34/m2_90_n50# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_12/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_2/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_58/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_44/m2_90_n50# rdummy_256x4_a_256x8m81_0/tblhl 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_22/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_28/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_59/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_54/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_40/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ rdummy_256x4_a_256x8m81_0/m3_117_13670# 018SRAM_cell1_dummy_R_256x8m81_4/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_32/a_246_342# rdummy_256x4_a_256x8m81_0/m3_264_359#
+ DWL 018SRAM_cell1_dummy_256x8m81_41/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_25/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_8/a_246_342# 018SRAM_cell1_dummy_256x8m81_42/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_35/m2_90_n50# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_13/a_246_342# 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_3/w_n68_622# 018SRAM_cell1_dummy_256x8m81_43/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_45/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_23/a_246_342#
+ 018SRAM_cell1_dummy_R_256x8m81_29/w_n68_622# 018SRAM_cell1_dummy_256x8m81_44/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_55/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_16/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_33/a_246_342# rdummy_256x4_a_256x8m81_0/pmos_5p04310590878155_256x8m81_0/S
+ 018SRAM_cell1_dummy_256x8m81_45/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_26/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_9/a_246_342#
+ rdummy_256x4_a_256x8m81_0/m3_117_13992# 018SRAM_cell1_dummy_R_256x8m81_4/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_46/m2_390_n50# rdummy_256x4_a_256x8m81_0/m3_117_15328#
+ 018SRAM_cell1_dummy_256x8m81_36/m2_90_n50# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_14/a_246_342# 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_47/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_30/a_126_298#
+ 018SRAM_cell1_dummy_256x8m81_46/m2_90_n50# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_24/a_246_342# rdummy_256x4_a_256x8m81_0/m3_117_14314#
+ 018SRAM_cell1_dummy_256x8m81_48/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_56/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_17/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_49/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_30/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_27/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_31/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_21/a_126_298# 018SRAM_cell1_dummy_256x8m81_37/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_15/a_246_342# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/d
+ 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_32/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_31/a_126_298# 018SRAM_cell1_dummy_256x8m81_47/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50#
+ 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_25/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_33/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_18/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_57/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_30/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50#
+ rdummy_256x4_a_256x8m81_0/w_523_3317# 018SRAM_cell1_dummy_R_256x8m81_30/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_34/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_28/m2_90_n50#
+ rdummy_256x4_a_256x8m81_0/m3_117_14636# 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_31/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_35/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_9/a_126_298#
+ 018SRAM_cell1_dummy_256x8m81_38/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_32/m3_n36_330# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_16/a_246_342# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_36/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_32/a_126_298# 018SRAM_cell1_dummy_256x8m81_48/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_33/m3_n36_330#
+ 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_26/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_21/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_37/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_58/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_19/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_31/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_38/m2_390_n50# a_5143_1594# 018SRAM_cell1_dummy_256x8m81_29/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_39/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_20/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_8/a_126_298# 018SRAM_cell1_dummy_256x8m81_39/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_17/a_246_342# 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_21/m2_390_n50# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_5/a_126_298# 018SRAM_cell1_dummy_256x8m81_49/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_27/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_9/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_22/m2_390_n50#
+ rdummy_256x4_a_256x8m81_0/m3_117_16293# 018SRAM_cell1_dummy_256x8m81_59/m2_90_n50#
+ 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_32/w_n68_622# 018SRAM_cell1_dummy_256x8m81_23/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_20/a_126_298# 018SRAM_cell1_dummy_R_256x8m81_20/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_2/a_246_342# 018SRAM_cell1_dummy_256x8m81_24/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_24/a_126_298# VSS 018SRAM_cell1_dummy_R_256x8m81_21/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_18/a_246_342# 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_25/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_22/m3_n36_330#
+ rdummy_256x4_a_256x8m81_0/m3_117_15650# 018SRAM_cell1_dummy_R_256x8m81_28/a_246_342#
+ 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_R_256x8m81_8/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_26/m2_390_n50# a_5143_52# 018SRAM_cell1_dummy_R_256x8m81_23/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_5/w_n68_622# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_27/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_24/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_20/m2_90_n50# a_28741_23194# 018SRAM_cell1_dummy_R_256x8m81_3/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_28/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_30/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_60/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_25/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_19/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_20/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_29/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_26/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_40/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_61/m2_390_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_29/a_246_342# rdummy_256x4_a_256x8m81_0/m3_117_15971#
+ 018SRAM_cell1_dummy_R_256x8m81_24/w_n68_622# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/m3_n36_330#
+ rdummy_256x4_a_256x8m81_0/vdd 018SRAM_cell1_dummy_R_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50#
+ 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_50/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_27/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_62/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50#
+ 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_60/m2_90_n50#
+ 018SRAM_cell1_dummy_R_256x8m81_28/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_21/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_63/m2_390_n50# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_256x8m81_4/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_2/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_R_256x8m81_29/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_31/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_10/m3_n36_330#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_R_256x8m81_3/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
X018SRAM_cell1_2x_256x8m81_10 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_10/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_11 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_11/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_12 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_12/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_13 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_13/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_0 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_0/a_246_342# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_dummy_R_256x8m81_0/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_2x_256x8m81_14 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_14/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_1 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ VSUBS 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_52# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_2x_256x8m81_15 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_15/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_2 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_2/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_2/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_2/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_2/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_0 a_5143_52# 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_60 DWL 018SRAM_cell1_dummy_256x8m81_60/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_60/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_3 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_3/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_3/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_3/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_3/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_1 a_5143_52# 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_61 DWL 018SRAM_cell1_dummy_256x8m81_61/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_61/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_50 DWL 018SRAM_cell1_dummy_256x8m81_50/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_50/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_4 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_4/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_4/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_4/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_4/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_2 a_5143_52# 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_62 DWL 018SRAM_cell1_dummy_256x8m81_62/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_62/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_51 DWL 018SRAM_cell1_dummy_256x8m81_51/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_51/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_40 DWL 018SRAM_cell1_dummy_256x8m81_40/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_40/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_5 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_5/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_5/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_5/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_5/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_30 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_30/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_30/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_30/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_30/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_3 a_5143_52# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_6 DWL rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ VSUBS 018SRAM_cell1_256x8m81_1/w_n68_622# DWL rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_63 DWL 018SRAM_cell1_dummy_256x8m81_63/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_63/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_52 DWL 018SRAM_cell1_dummy_256x8m81_52/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_52/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_41 DWL 018SRAM_cell1_dummy_256x8m81_41/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_41/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_30 a_5143_52# 018SRAM_cell1_dummy_256x8m81_30/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_30/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_31 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_31/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_31/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_31/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_31/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_20 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_20/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_20/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_20/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_20/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_4 a_5143_52# 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_7 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_7/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_7/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_7/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_7/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_53 DWL 018SRAM_cell1_dummy_256x8m81_53/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_53/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_42 DWL 018SRAM_cell1_dummy_256x8m81_42/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_42/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_31 a_5143_52# 018SRAM_cell1_dummy_256x8m81_31/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_31/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_20 a_5143_52# 018SRAM_cell1_dummy_256x8m81_20/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_20/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_5 a_5143_52# 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_32 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_32/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_32/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_32/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_32/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_10 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_10/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_30/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_10/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_30/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_21 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_21/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_21/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_21/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_21/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_54 DWL 018SRAM_cell1_dummy_256x8m81_54/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_54/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_32 DWL 018SRAM_cell1_dummy_256x8m81_32/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_32/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_43 DWL 018SRAM_cell1_dummy_256x8m81_43/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_43/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_8 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_8/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_8/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_8/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_8/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_21 a_5143_52# 018SRAM_cell1_dummy_256x8m81_21/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_21/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_10 a_5143_52# 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_22 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_22/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_9/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_22/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_9/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_11 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_11/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_29/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_11/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_29/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_33 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_33/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_5/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_33/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_5/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_6 a_5143_52# 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_55 DWL 018SRAM_cell1_dummy_256x8m81_55/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_55/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_33 DWL 018SRAM_cell1_dummy_256x8m81_33/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_33/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_44 DWL 018SRAM_cell1_dummy_256x8m81_44/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_44/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_9 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_9/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_9/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_9/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_9/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_22 a_5143_52# 018SRAM_cell1_dummy_256x8m81_22/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_22/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_11 a_5143_52# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_7 a_5143_52# 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_23 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_23/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_8/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_23/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_8/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_12 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_12/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_21/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_12/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_21/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_56 DWL 018SRAM_cell1_dummy_256x8m81_56/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_56/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_34 DWL 018SRAM_cell1_dummy_256x8m81_34/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_34/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_45 DWL 018SRAM_cell1_dummy_256x8m81_45/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_45/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_23 a_5143_52# 018SRAM_cell1_dummy_256x8m81_23/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_23/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_12 a_5143_52# 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_24 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_24/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_24/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_24/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_24/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_13 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_13/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_28/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_13/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_28/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_8 a_5143_52# 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_57 DWL 018SRAM_cell1_dummy_256x8m81_57/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_57/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_35 DWL 018SRAM_cell1_dummy_256x8m81_35/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_35/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_46 DWL 018SRAM_cell1_dummy_256x8m81_46/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_46/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_24 a_5143_52# 018SRAM_cell1_dummy_256x8m81_24/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_24/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_13 a_5143_52# 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_9 a_5143_52# 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_25 DWL rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_25/a_246_342# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_dummy_R_256x8m81_25/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_14 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_14/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_20/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_14/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_20/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_58 DWL 018SRAM_cell1_dummy_256x8m81_58/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_58/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_36 DWL 018SRAM_cell1_dummy_256x8m81_36/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_36/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_47 DWL 018SRAM_cell1_dummy_256x8m81_47/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_47/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_25 a_5143_52# 018SRAM_cell1_dummy_256x8m81_25/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_25/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_14 a_5143_52# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_15 DWL rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_15/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_32/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_15/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_32/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_26 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_26/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_4/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_26/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_4/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_256x8m81_0 a_5143_52# 018SRAM_cell1_256x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS x018SRAM_cell1_256x8m81
X018SRAM_cell1_dummy_256x8m81_59 DWL 018SRAM_cell1_dummy_256x8m81_59/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_59/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_48 DWL 018SRAM_cell1_dummy_256x8m81_48/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_48/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_37 DWL 018SRAM_cell1_dummy_256x8m81_37/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_37/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_26 a_5143_52# 018SRAM_cell1_dummy_256x8m81_26/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_26/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_15 a_5143_52# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_16 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_16/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_24/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_16/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_24/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_256x8m81_1 a_5143_1594# 018SRAM_cell1_256x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS x018SRAM_cell1_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_27 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_27/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_7/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_27/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_7/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_49 DWL 018SRAM_cell1_dummy_256x8m81_49/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_49/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_38 DWL 018SRAM_cell1_dummy_256x8m81_38/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_38/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_16 a_5143_52# 018SRAM_cell1_dummy_256x8m81_16/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_16/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_27 a_5143_52# 018SRAM_cell1_dummy_256x8m81_27/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_27/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_17 a_28741_23194# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_17/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_31/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_17/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_31/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_28 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_28/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_28/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_28/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_28/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_39 DWL 018SRAM_cell1_dummy_256x8m81_39/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_39/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_17 a_5143_52# 018SRAM_cell1_dummy_256x8m81_17/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_17/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_28 a_5143_52# 018SRAM_cell1_dummy_256x8m81_28/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_28/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_2x_256x8m81_0 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_0/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_29 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_29/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_29/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_29/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_29/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_18 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_18/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_2/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_18/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_2/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_18 a_5143_52# 018SRAM_cell1_dummy_256x8m81_18/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_18/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_29 a_5143_52# 018SRAM_cell1_dummy_256x8m81_29/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_29/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_2x_256x8m81_1 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_1/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_dummy_R_256x8m81_19 a_28741_1594# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ 018SRAM_cell1_dummy_R_256x8m81_19/a_246_342# 018SRAM_cell1_dummy_R_256x8m81_3/a_126_298#
+ 018SRAM_cell1_dummy_R_256x8m81_19/m3_n36_330# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ 018SRAM_cell1_dummy_R_256x8m81_3/w_n68_622# VSUBS x018SRAM_cell1_dummy_R_256x8m81
X018SRAM_cell1_dummy_256x8m81_19 a_5143_52# 018SRAM_cell1_dummy_256x8m81_19/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_19/m2_390_n50# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_52# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_2x_256x8m81_2 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_3 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_4 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_5 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_6 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
Xrdummy_256x4_a_256x8m81_0 rdummy_256x4_a_256x8m81_0/pcb rdummy_256x4_a_256x8m81_0/tblhl
+ rdummy_256x4_a_256x8m81_0/m3_117_16293# rdummy_256x4_a_256x8m81_0/m3_117_15650#
+ rdummy_256x4_a_256x8m81_0/m3_117_15971# rdummy_256x4_a_256x8m81_0/m3_264_359# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/d
+ rdummy_256x4_a_256x8m81_0/m3_117_13670# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/bb
+ rdummy_256x4_a_256x8m81_0/w_523_3317# rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/b
+ rdummy_256x4_a_256x8m81_0/m3_117_13992# rdummy_256x4_a_256x8m81_0/m3_117_15328#
+ rdummy_256x4_a_256x8m81_0/vdd VSUBS rdummy_256x4_a_256x8m81_0/m3_117_14314# rdummy_256x4_a_256x8m81_0/pmos_5p04310590878155_256x8m81_0/S
+ rdummy_256x4_a_256x8m81_0/m3_117_14636# rdummy_256x4_a_256x8m81
X018SRAM_cell1_2x_256x8m81_7 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_8 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_9 018SRAM_cell1_256x8m81_1/w_n68_622# a_5143_1594# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ a_5143_1594# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/m3_n36_330# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
.ends

.subckt rcol4_256_256x8m81 pcb[6] pcb[7] pcb[4] vdd PCB[8] WEN[4] WEN[7] pcb[5] WEN[5]
+ WEN[6] men ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] DWL tblhl GWEN
+ ypass[0] WL[23] WL[22] WL[27] WL[30] WL[18] WL[15] WL[12] ypass[7] WL[13] WL[14]
+ WL[16] WL[17] WL[19] WL[28] din[4] din[7] q[5] q[6] q[7] din[5] din[6] q[4] saout_R_m2_256x8m81_1/pcb
+ rdummy_256x4_256x8m81_0/DWL saout_R_m2_256x8m81_1/WEN WL[2] WL[3] WL[6] WL[7] WL[20]
+ WL[21] WL[4] WL[5] WL[8] WL[9] WL[24] GWE WL[29] WL[25] rdummy_256x4_256x8m81_0/VSS
+ WL[26] WL[10] WL[11] WL[31] WL[0] WL[1] VSS VDD
Xdcap_103_novia_256x8m81_0[0] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[1] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[2] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[3] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[4] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[5] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[6] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[7] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[8] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[9] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[10] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[11] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[12] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[13] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[14] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[15] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[16] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[17] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[18] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[19] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[20] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[21] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[22] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[23] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[24] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[25] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[26] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[27] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[28] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[29] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[30] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[31] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[32] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[33] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[34] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[35] VDD VDD VSS dcap_103_novia_256x8m81
Xrarray4_256_256x8m81_0 WL[23] WL[26] WL[18] WL[11] WL[15] WL[14] WL[19] WL[31] WL[13]
+ WL[16] saout_m2_256x8m81_0/bb[7] saout_m2_256x8m81_0/bb[0] saout_m2_256x8m81_0/b[2]
+ saout_R_m2_256x8m81_0/b[5] saout_m2_256x8m81_1/b[0] saout_m2_256x8m81_1/b[7] saout_m2_256x8m81_1/bb[6]
+ saout_m2_256x8m81_0/b[6] WL[5] saout_m2_256x8m81_1/bb[2] WL[2] saout_m2_256x8m81_1/b[1]
+ saout_R_m2_256x8m81_0/b[1] saout_R_m2_256x8m81_0/bb[2] saout_m2_256x8m81_1/bb[1]
+ saout_m2_256x8m81_1/b[3] saout_R_m2_256x8m81_0/b[4] saout_R_m2_256x8m81_0/bb[6]
+ saout_R_m2_256x8m81_0/bb[3] WL[27] saout_R_m2_256x8m81_0/b[3] saout_m2_256x8m81_0/bb[5]
+ WL[0] saout_m2_256x8m81_0/b[1] saout_m2_256x8m81_1/bb[5] saout_R_m2_256x8m81_1/bb[2]
+ saout_R_m2_256x8m81_0/b[0] saout_R_m2_256x8m81_1/bb[7] saout_R_m2_256x8m81_0/b[7]
+ saout_m2_256x8m81_0/b[5] WL[8] saout_R_m2_256x8m81_1/b[6] saout_m2_256x8m81_1/bb[7]
+ saout_m2_256x8m81_0/b[3] saout_R_m2_256x8m81_1/bb[4] saout_m2_256x8m81_1/b[2] saout_R_m2_256x8m81_1/b[4]
+ WL[24] saout_R_m2_256x8m81_0/bb[4] saout_m2_256x8m81_0/b[4] saout_m2_256x8m81_1/bb[4]
+ WL[3] saout_R_m2_256x8m81_1/b[7] saout_m2_256x8m81_0/bb[2] saout_R_m2_256x8m81_1/bb[1]
+ saout_m2_256x8m81_0/b[0] saout_R_m2_256x8m81_0/bb[1] saout_R_m2_256x8m81_1/b[5]
+ WL[6] saout_R_m2_256x8m81_1/b[0] saout_R_m2_256x8m81_0/bb[7] saout_m2_256x8m81_1/b[6]
+ saout_R_m2_256x8m81_1/b[3] WL[1] saout_m2_256x8m81_0/b[7] saout_R_m2_256x8m81_1/bb[0]
+ WL[29] saout_R_m2_256x8m81_1/b[2] WL[4] WL[12] saout_R_m2_256x8m81_0/bb[5] saout_m2_256x8m81_1/bb[3]
+ saout_m2_256x8m81_1/b[5] WL[28] WL[30] saout_m2_256x8m81_0/bb[1] saout_R_m2_256x8m81_0/bb[0]
+ WL[9] saout_m2_256x8m81_1/bb[0] WL[25] saout_R_m2_256x8m81_1/bb[6] saout_R_m2_256x8m81_0/b[2]
+ saout_m2_256x8m81_0/bb[3] saout_R_m2_256x8m81_1/b[1] saout_m2_256x8m81_0/bb[6] WL[20]
+ saout_R_m2_256x8m81_1/bb[5] WL[21] WL[7] saout_R_m2_256x8m81_1/bb[3] WL[17] saout_m2_256x8m81_0/bb[4]
+ WL[10] WL[22] saout_R_m2_256x8m81_0/b[6] saout_m2_256x8m81_1/b[4] VDD VSS rarray4_256_256x8m81
Xsaout_R_m2_256x8m81_0 saout_R_m2_256x8m81_0/pcb saout_R_m2_256x8m81_0/datain saout_R_m2_256x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWE GWEN
+ saout_R_m2_256x8m81_0/b[7] saout_R_m2_256x8m81_0/b[0] saout_R_m2_256x8m81_0/bb[5]
+ saout_R_m2_256x8m81_0/q saout_R_m2_256x8m81_0/wen_wm1_256x8m81_0/wen VDD saout_R_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ saout_R_m2_256x8m81_0/b[2] saout_R_m2_256x8m81_0/b[6] saout_R_m2_256x8m81_0/bb[1]
+ saout_R_m2_256x8m81_0/bb[3] saout_R_m2_256x8m81_0/b[5] saout_R_m2_256x8m81_0/bb[4]
+ saout_R_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b saout_R_m2_256x8m81_0/b[4]
+ men a_6900_27175# a_6434_27175# saout_R_m2_256x8m81_0/bb[6] a_6900_27950# a_6434_27950#
+ ypass[0] ypass[7] VSS VSS saout_R_m2_256x8m81_0/bb[7] saout_R_m2_256x8m81_0/bb[0]
+ ypass[1] saout_R_m2_256x8m81_0/sacntl_2_256x8m81_0/a_4718_983# GWEN ypass[4] ypass[2]
+ VDD saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb saout_R_m2_256x8m81_0/bb[2] saout_R_m2_256x8m81_0/b[3]
+ VDD ypass[5] ypass[6] VDD VSS saout_R_m2_256x8m81_0/sa_256x8m81_0/wep VSS VDD saout_R_m2_256x8m81_0/b[1]
+ ypass[3] saout_R_m2_256x8m81
Xsaout_R_m2_256x8m81_1 saout_R_m2_256x8m81_1/pcb saout_R_m2_256x8m81_1/datain saout_R_m2_256x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWE GWEN
+ saout_R_m2_256x8m81_1/b[7] saout_R_m2_256x8m81_1/b[0] saout_R_m2_256x8m81_1/bb[5]
+ saout_R_m2_256x8m81_1/q saout_R_m2_256x8m81_1/wen_wm1_256x8m81_0/wen VDD saout_R_m2_256x8m81_1/mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ saout_R_m2_256x8m81_1/b[2] saout_R_m2_256x8m81_1/b[6] saout_R_m2_256x8m81_1/bb[1]
+ saout_R_m2_256x8m81_1/bb[3] saout_R_m2_256x8m81_1/b[5] saout_R_m2_256x8m81_1/bb[4]
+ saout_R_m2_256x8m81_1/b[7] saout_R_m2_256x8m81_1/b[4] men a_17700_27175# a_17234_27175#
+ saout_R_m2_256x8m81_1/bb[6] a_17700_27950# a_17234_27950# ypass[0] ypass[7] VSS
+ VSS saout_R_m2_256x8m81_1/bb[7] saout_R_m2_256x8m81_1/bb[0] ypass[1] saout_R_m2_256x8m81_1/sacntl_2_256x8m81_0/a_4718_983#
+ GWEN ypass[4] ypass[2] VDD saout_R_m2_256x8m81_1/pcb saout_R_m2_256x8m81_1/bb[2]
+ saout_R_m2_256x8m81_1/b[3] VDD ypass[5] ypass[6] VDD saout_R_m2_256x8m81_1/mux821_256x8m81_0/a_4992_424#
+ saout_R_m2_256x8m81_1/sa_256x8m81_0/wep VSS VDD saout_R_m2_256x8m81_1/b[1] ypass[3]
+ saout_R_m2_256x8m81
Xsaout_m2_256x8m81_0 saout_m2_256x8m81_0/pcb saout_m2_256x8m81_0/datain saout_m2_256x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWEN GWE
+ saout_m2_256x8m81_0/bb[2] saout_m2_256x8m81_0/b[0] saout_m2_256x8m81_0/q a_17009_27175#
+ a_17234_27175# a_17009_27950# a_17234_27950# VDD saout_m2_256x8m81_0/b[5] saout_m2_256x8m81_0/b[1]
+ ypass[7] saout_m2_256x8m81_0/bb[6] saout_m2_256x8m81_0/bb[4] saout_m2_256x8m81_0/b[2]
+ saout_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10# saout_m2_256x8m81_0/bb[3]
+ saout_m2_256x8m81_0/b[3] men saout_m2_256x8m81_0/bb[1] ypass[0] saout_m2_256x8m81_0/sacntl_2_256x8m81_0/a_4560_1922#
+ VSS saout_m2_256x8m81_0/bb[0] saout_m2_256x8m81_0/bb[7] ypass[1] saout_m2_256x8m81_0/sacntl_2_256x8m81_0/a_4718_983#
+ GWEN ypass[4] ypass[2] VDD saout_m2_256x8m81_0/b[7] saout_m2_256x8m81_0/bb[5] saout_m2_256x8m81_0/sa_256x8m81_0/pcb
+ saout_m2_256x8m81_0/b[4] VDD VDD ypass[5] VDD ypass[6] saout_m2_256x8m81_0/sa_256x8m81_0/wep
+ saout_m2_256x8m81_0/mux821_256x8m81_0/a_4992_424# VSS saout_m2_256x8m81_0/b[6] ypass[3]
+ saout_m2_256x8m81
Xsaout_m2_256x8m81_1 saout_m2_256x8m81_1/pcb saout_m2_256x8m81_1/datain saout_m2_256x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWEN GWE
+ saout_m2_256x8m81_1/bb[2] saout_m2_256x8m81_1/b[0] saout_m2_256x8m81_1/q a_6209_27175#
+ a_6434_27175# a_6209_27950# a_6434_27950# VDD saout_m2_256x8m81_1/b[5] saout_m2_256x8m81_1/b[1]
+ ypass[7] saout_m2_256x8m81_1/bb[6] saout_m2_256x8m81_1/bb[4] saout_m2_256x8m81_1/b[2]
+ saout_m2_256x8m81_1/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10# saout_m2_256x8m81_1/bb[3]
+ saout_m2_256x8m81_1/b[3] men saout_m2_256x8m81_1/bb[1] ypass[0] VSS VSS saout_m2_256x8m81_1/bb[0]
+ saout_m2_256x8m81_1/bb[7] ypass[1] VSS GWEN ypass[4] ypass[2] VDD saout_m2_256x8m81_1/b[7]
+ saout_m2_256x8m81_1/bb[5] saout_m2_256x8m81_1/sa_256x8m81_0/pcb saout_m2_256x8m81_1/b[4]
+ VDD VDD ypass[5] VDD ypass[6] saout_m2_256x8m81_1/sa_256x8m81_0/wep saout_m2_256x8m81_1/mux821_256x8m81_0/a_4992_424#
+ VSS saout_m2_256x8m81_1/b[6] ypass[3] saout_m2_256x8m81
Xrdummy_256x4_256x8m81_0 WL[18] saout_m2_256x8m81_1/b[4] WL[4] saout_m2_256x8m81_0/b[1]
+ saout_m2_256x8m81_0/b[2] WL[16] saout_m2_256x8m81_0/bb[5] WL[2] saout_m2_256x8m81_1/b[5]
+ WL[14] saout_R_m2_256x8m81_1/bb[5] saout_R_m2_256x8m81_0/b[0] VSS saout_m2_256x8m81_1/b[3]
+ VDD WL[12] saout_R_m2_256x8m81_0/bb[7] VSS saout_m2_256x8m81_0/bb[7] WL[10] saout_m2_256x8m81_1/bb[2]
+ WL[30] saout_m2_256x8m81_1/bb[5] saout_m2_256x8m81_0/b[1] VSS VSS WL[24] saout_m2_256x8m81_1/b[1]
+ WL[28] saout_m2_256x8m81_0/bb[3] saout_m2_256x8m81_0/bb[2] saout_m2_256x8m81_0/bb[3]
+ VSS WL[20] WL[26] saout_R_m2_256x8m81_1/b[6] VDD saout_R_m2_256x8m81_0/bb[1] saout_m2_256x8m81_0/b[3]
+ VDD saout_m2_256x8m81_0/b[5] WL[5] saout_R_m2_256x8m81_0/b[6] VSS WL[7] saout_m2_256x8m81_0/bb[4]
+ saout_m2_256x8m81_1/bb[3] WL[15] VSS VDD saout_m2_256x8m81_0/b[7] saout_m2_256x8m81_0/bb[5]
+ saout_m2_256x8m81_0/b[2] VSS saout_R_m2_256x8m81_1/bb[0] saout_R_m2_256x8m81_1/bb[7]
+ VDD saout_R_m2_256x8m81_0/b[2] WL[28] WL[3] VSS saout_R_m2_256x8m81_1/b[1] VDD saout_R_m2_256x8m81_0/b[4]
+ WL[23] VSS VDD saout_m2_256x8m81_0/b[0] saout_R_m2_256x8m81_1/bb[2] saout_m2_256x8m81_1/b[2]
+ tblhl WL[7] VSS VDD saout_R_m2_256x8m81_1/b[3] saout_m2_256x8m81_0/b[4] saout_m2_256x8m81_1/bb[6]
+ saout_m2_256x8m81_0/bb[1] ypass[0] VDD VSS VSS rdummy_256x4_256x8m81_0/DWL saout_m2_256x8m81_1/bb[4]
+ saout_R_m2_256x8m81_0/bb[3] VSS saout_m2_256x8m81_1/b[5] saout_R_m2_256x8m81_0/bb[5]
+ WL[30] VSS saout_R_m2_256x8m81_1/bb[1] VDD saout_m2_256x8m81_1/b[3] saout_m2_256x8m81_1/bb[1]
+ VSS VDD saout_m2_256x8m81_1/bb[2] saout_m2_256x8m81_0/bb[7] saout_m2_256x8m81_1/bb[5]
+ VSS VDD saout_m2_256x8m81_1/b[1] saout_R_m2_256x8m81_0/bb[5] WL[13] VSS ypass[1]
+ VDD saout_m2_256x8m81_1/bb[0] ypass[4] saout_R_m2_256x8m81_0/b[2] WL[4] VSS saout_R_m2_256x8m81_1/b[2]
+ saout_m2_256x8m81_1/b[7] VDD saout_m2_256x8m81_1/b[0] WL[5] VSS ypass[2] saout_m2_256x8m81_0/bb[6]
+ saout_R_m2_256x8m81_1/b[0] saout_m2_256x8m81_1/bb[3] saout_m2_256x8m81_0/bb[0] saout_m2_256x8m81_1/bb[6]
+ saout_R_m2_256x8m81_0/b[4] saout_m2_256x8m81_0/bb[0] saout_m2_256x8m81_1/bb[4] VDD
+ saout_R_m2_256x8m81_0/bb[1] WL[16] saout_R_m2_256x8m81_1/b[1] WL[29] WL[24] VSS
+ rdummy_256x4_256x8m81_0/rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/d saout_R_m2_256x8m81_1/bb[3]
+ saout_R_m2_256x8m81_0/b[7] VDD saout_m2_256x8m81_1/bb[7] WL[8] saout_R_m2_256x8m81_1/bb[2]
+ WL[25] VSS WL[26] saout_R_m2_256x8m81_0/bb[6] saout_m2_256x8m81_1/b[2] saout_R_m2_256x8m81_1/bb[1]
+ WL[21] saout_R_m2_256x8m81_1/b[3] VDD VDD saout_R_m2_256x8m81_0/bb[4] saout_R_m2_256x8m81_0/b[6]
+ ypass[3] saout_R_m2_256x8m81_1/bb[4] WL[25] VSS saout_R_m2_256x8m81_0/b[5] VDD saout_R_m2_256x8m81_0/b[0]
+ saout_R_m2_256x8m81_1/bb[0] WL[29] WL[18] VSS WL[20] saout_R_m2_256x8m81_1/b[4]
+ saout_R_m2_256x8m81_0/bb[2] VDD saout_m2_256x8m81_0/b[6] saout_R_m2_256x8m81_1/b[5]
+ WL[1] WL[19] VSS WL[31] VDD saout_R_m2_256x8m81_0/b[1] saout_R_m2_256x8m81_1/b[2]
+ saout_R_m2_256x8m81_1/bb[6] saout_m2_256x8m81_1/bb[1] WL[10] VDD saout_R_m2_256x8m81_0/bb[0]
+ VSS saout_R_m2_256x8m81_0/bb[7] saout_R_m2_256x8m81_1/b[7] WL[11] saout_R_m2_256x8m81_0/b[3]
+ saout_m2_256x8m81_1/bb[0] VDD saout_R_m2_256x8m81_0/bb[3] saout_m2_256x8m81_0/b[7]
+ rdummy_256x4_256x8m81_0/rdummy_256x4_a_256x8m81_0/ypass_gate_256x8m81_0_0/d VSS
+ saout_R_m2_256x8m81_1/b[0] saout_m2_256x8m81_1/b[7] WL[17] VDD saout_m2_256x8m81_0/b[0]
+ VSS VDD WL[2] saout_R_m2_256x8m81_0/bb[0] ypass[7] saout_R_m2_256x8m81_1/bb[3] WL[12]
+ WL[0] VDD saout_R_m2_256x8m81_0/b[1] VDD WL[11] VSS saout_R_m2_256x8m81_0/bb[2]
+ VDD rdummy_256x4_256x8m81_0/VSS WL[15] VSS saout_R_m2_256x8m81_1/bb[5] saout_R_m2_256x8m81_0/b[3]
+ WL[19] ypass[5] VSS WL[14] VDD saout_R_m2_256x8m81_0/b[5] VSS WL[23] saout_m2_256x8m81_0/b[6]
+ WL[9] VDD WL[27] saout_R_m2_256x8m81_0/bb[4] WL[27] saout_m2_256x8m81_1/b[0] VSS
+ VSS saout_R_m2_256x8m81_0/bb[6] saout_m2_256x8m81_1/b[6] saout_R_m2_256x8m81_1/bb[4]
+ WL[31] VSS VDD saout_R_m2_256x8m81_1/b[6] saout_m2_256x8m81_0/bb[6] saout_R_m2_256x8m81_0/b[7]
+ WL[3] saout_m2_256x8m81_1/b[6] saout_R_m2_256x8m81_1/b[5] VSS ypass[6] VDD WL[21]
+ VDD WL[0] saout_m2_256x8m81_0/bb[4] WL[1] saout_m2_256x8m81_0/bb[1] WL[9] saout_m2_256x8m81_0/b[4]
+ saout_R_m2_256x8m81_1/bb[6] saout_m2_256x8m81_0/b[5] WL[6] saout_R_m2_256x8m81_1/b[4]
+ WL[13] saout_m2_256x8m81_1/bb[7] saout_R_m2_256x8m81_1/b[7] WL[22] VSS WL[6] saout_m2_256x8m81_0/b[3]
+ WL[17] saout_m2_256x8m81_1/b[4] WL[22] VSS saout_R_m2_256x8m81_1/bb[7] WL[8] VDD
+ saout_m2_256x8m81_0/bb[2] rdummy_256x4_256x8m81
.ends

.subckt pmos_5p043105908781101_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.59u l=0.6u
.ends

.subckt pmoscap_W2_5_477_R270_256x8m81 m3_489_n1# m3_1409_n1# w_n60_n407# a_81_507#
X0 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
X1 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_5p043105908781102_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.63u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.63u l=0.6u
.ends

.subckt pmos_1p2$$204216364_256x8m81 pmos_5p043105908781102_256x8m81_0/D w_n296_n137#
+ a_193_n71# pmos_5p043105908781102_256x8m81_0/S a_n31_n71#
Xpmos_5p043105908781102_256x8m81_0 w_n296_n137# pmos_5p043105908781102_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781102_256x8m81_0/S a_193_n71# pmos_5p043105908781102_256x8m81
.ends

.subckt pmos_5p043105908781104_256x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
.ends

.subckt pmos_5p043105908781103_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.5u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.5u l=0.6u
.ends

.subckt pmos_1p2$$49272876_R270_256x8m81 w_n296_n137# pmos_5p043105908781103_256x8m81_0/S
+ a_n31_n71# pmos_5p043105908781103_256x8m81_0/D a_193_n71#
Xpmos_5p043105908781103_256x8m81_0 w_n296_n137# pmos_5p043105908781103_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781103_256x8m81_0/S a_193_n71# pmos_5p043105908781103_256x8m81
.ends

.subckt nmos_5p043105908781109_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=3.3u l=0.6u
.ends

.subckt nmos_1p2$$49277996_R270_256x8m81 nmos_5p04310590878144_256x8m81_0/S a_n31_n71#
+ nmos_5p04310590878144_256x8m81_0/D VSUBS
Xnmos_5p04310590878144_256x8m81_0 nmos_5p04310590878144_256x8m81_0/D a_n31_n71# nmos_5p04310590878144_256x8m81_0/S
+ VSUBS nmos_5p04310590878144_256x8m81
.ends

.subckt nmos_5p043105908781108_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=5u l=0.6u
.ends

.subckt nmos_5p043105908781107_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.66u l=0.6u
.ends

.subckt pmos_5p043105908781110_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.59u l=0.6u
.ends

.subckt pmos_5p043105908781105_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_1p2$$49271852_R270_256x8m81 pmos_5p043105908781105_256x8m81_0/S w_n296_n137#
+ pmos_5p043105908781105_256x8m81_0/D a_193_n71# a_n31_n71#
Xpmos_5p043105908781105_256x8m81_0 w_n296_n137# pmos_5p043105908781105_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781105_256x8m81_0/S a_193_n71# pmos_5p043105908781105_256x8m81
.ends

.subckt pmos_1p2$$49270828_R270_256x8m81 w_n296_n137# pmos_5p043105908781104_256x8m81_0/S
+ a_193_n71# pmos_5p043105908781104_256x8m81_0/D a_n31_n71# a_417_n71#
Xpmos_5p043105908781104_256x8m81_0 w_n296_n137# pmos_5p043105908781104_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781104_256x8m81_0/S a_417_n71# a_193_n71# pmos_5p043105908781104_256x8m81
.ends

.subckt pmos_5p043105908781106_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.62u l=0.6u
.ends

.subckt xdec_256x8m81 xc xb xa RWL m2_16621_n223# m2_17754_n223# m2_11825_n223# m2_12202_n223#
+ m2_12958_n223# m2_15487_n223# m2_12580_n223# m2_15110_n223# m2_11069_n223# m2_15865_n223#
+ m2_16243_n223# LWL m2_10314_n223# m2_16998_n223# m2_17376_n223# men m2_11447_n223#
+ vdd vss m2_10691_n223#
Xpmos_5p043105908781104_256x8m81_0 vdd vdd pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D
+ RWL pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D
+ pmos_5p043105908781104_256x8m81
Xpmos_1p2$$49272876_R270_256x8m81_0 vdd vdd nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D
+ nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81
Xnmos_5p043105908781109_256x8m81_0 men pmos_5p043105908781110_256x8m81_0/S nmos_5p043105908781109_256x8m81_0/S
+ pmos_5p043105908781110_256x8m81_0/S vss nmos_5p043105908781109_256x8m81
Xnmos_1p2$$49277996_R270_256x8m81_0 nmos_5p043105908781109_256x8m81_0/S pmos_5p043105908781106_256x8m81_2/S
+ vss vss nmos_1p2$$49277996_R270_256x8m81
Xpmos_1p2$$49272876_R270_256x8m81_1 vdd vdd nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D
+ nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81
Xnmos_5p043105908781108_256x8m81_0 LWL pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D
+ vss pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D vss nmos_5p043105908781108_256x8m81
Xnmos_5p043105908781108_256x8m81_1 RWL pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D
+ vss pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D vss nmos_5p043105908781108_256x8m81
Xnmos_5p043105908781107_256x8m81_0 vss pmos_5p043105908781106_256x8m81_2/S pmos_5p043105908781110_256x8m81_0/S
+ vss nmos_5p043105908781107_256x8m81
Xpmos_5p043105908781110_256x8m81_0 vdd vdd pmos_5p043105908781106_256x8m81_2/S pmos_5p043105908781110_256x8m81_0/S
+ pmos_5p043105908781110_256x8m81
Xpmos_1p2$$49271852_R270_256x8m81_0 nmos_5p043105908781109_256x8m81_0/S vdd men pmos_5p043105908781106_256x8m81_2/S
+ pmos_5p043105908781106_256x8m81_2/S pmos_1p2$$49271852_R270_256x8m81
Xpmos_1p2$$49270828_R270_256x8m81_0 vdd LWL pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D
+ vdd pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D
+ pmos_1p2$$49270828_R270_256x8m81
Xpmos_5p043105908781106_256x8m81_0 vdd pmos_5p043105908781106_256x8m81_2/S xb vdd
+ pmos_5p043105908781106_256x8m81
Xpmos_5p043105908781106_256x8m81_1 vdd vdd xc pmos_5p043105908781106_256x8m81_2/S
+ pmos_5p043105908781106_256x8m81
Xpmos_5p043105908781106_256x8m81_2 vdd vdd xa pmos_5p043105908781106_256x8m81_2/S
+ pmos_5p043105908781106_256x8m81
X0 a_13291_624# xb a_13291_400# vss nmos_3p3 w=3.15u l=0.6u
X1 vss xc a_13291_624# vss nmos_3p3 w=3.15u l=0.6u
X2 a_13291_400# xa pmos_5p043105908781106_256x8m81_2/S vss nmos_3p3 w=3.15u l=0.6u
X3 vss nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81_0/pmos_5p043105908781103_256x8m81_0/D vss nmos_3p3 w=5u l=0.6u
X4 vss nmos_5p043105908781109_256x8m81_0/S pmos_1p2$$49272876_R270_256x8m81_1/pmos_5p043105908781103_256x8m81_0/D vss nmos_3p3 w=5u l=0.6u
.ends

.subckt xdec8_256x8m81 xa[5] xa[2] RWL[0] LWL[5] LWL[4] RWL[2] RWL[1] RWL[7] RWL[6]
+ LWL[1] LWL[7] LWL[6] LWL[0] LWL[3] RWL[3] xa[1] xa[7] xa[4] xa[3] xb xa[0] xa[6]
+ RWL[5] xdec_256x8m81_7/m2_16243_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_10314_n223#
+ xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_16621_n223#
+ xdec_256x8m81_7/m2_11069_n223# RWL[4] xdec_256x8m81_7/m2_12958_n223# xdec_256x8m81_7/m2_17376_n223#
+ xdec_256x8m81_7/m2_15110_n223# xdec_256x8m81_7/m2_11447_n223# LWL[2] men xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_15865_n223#
+ vss xdec_256x8m81_7/m2_12202_n223# vdd xc
Xxdec_256x8m81_7 xc xb xa[1] RWL[1] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[1] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_0 xc xb xa[6] RWL[6] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[6] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_1 xc xb xa[4] RWL[4] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[4] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_3 xc xb xa[0] xdec_256x8m81_3/RWL xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[0] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_2 xc xb xa[2] RWL[2] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[2] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_4 xc xb xa[7] RWL[7] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[7] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_5 xc xb xa[5] RWL[5] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[5] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
Xxdec_256x8m81_6 xc xb xa[3] RWL[3] xdec_256x8m81_7/m2_16621_n223# xdec_256x8m81_7/m2_17754_n223#
+ xdec_256x8m81_7/m2_11825_n223# xdec_256x8m81_7/m2_12202_n223# xdec_256x8m81_7/m2_12958_n223#
+ xdec_256x8m81_7/m2_15487_n223# xdec_256x8m81_7/m2_12580_n223# xdec_256x8m81_7/m2_15110_n223#
+ xdec_256x8m81_7/m2_11069_n223# xdec_256x8m81_7/m2_15865_n223# xdec_256x8m81_7/m2_16243_n223#
+ LWL[3] xdec_256x8m81_7/m2_10314_n223# xdec_256x8m81_7/m2_16998_n223# xdec_256x8m81_7/m2_17376_n223#
+ men xdec_256x8m81_7/m2_11447_n223# vdd vss xdec_256x8m81_7/m2_10691_n223# xdec_256x8m81
.ends

.subckt xdec32_256x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[16] RWL[15] RWL[14] RWL[13]
+ RWL[12] LWL[9] LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10]
+ RWL[9] RWL[8] RWL[7] RWL[5] RWL[3] RWL[1] RWL[0] RWL[2] LWL[18] LWL[17] LWL[16]
+ LWL[15] LWL[14] LWL[13] LWL[11] LWL[10] RWL[4] RWL[6] LWL[28] LWL[25] LWL[24] LWL[23]
+ LWL[22] LWL[21] LWL[20] LWL[19] RWL[20] RWL[21] RWL[22] RWL[23] RWL[24] RWL[25]
+ RWL[28] RWL[29] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[0] xa[3]
+ xa[4] xa[5] xa[6] xa[7] xb[3] xb[2] xb[1] xb[0] xc xdec8_256x8m81_3/xdec_256x8m81_7/m2_10314_n223#
+ xdec8_256x8m81_3/xdec_256x8m81_7/m2_10691_n223# LWL[27] xdec8_256x8m81_3/xdec_256x8m81_7/m2_11069_n223#
+ LWL[26] RWL[27] men xa[1] RWL[26] LWL[12] vss vdd
Xxdec8_256x8m81_0 xa[5] xa[2] RWL[24] LWL[29] LWL[28] RWL[26] RWL[25] RWL[31] RWL[30]
+ LWL[25] LWL[31] LWL[30] LWL[24] LWL[27] RWL[27] xa[1] xa[7] xa[4] xa[3] xb[3] xa[0]
+ xa[6] RWL[29] xa[4] xb[1] xdec8_256x8m81_3/xdec_256x8m81_7/m2_10314_n223# xdec8_256x8m81_3/xdec_256x8m81_7/m2_10691_n223#
+ xa[2] xa[3] xdec8_256x8m81_3/xdec_256x8m81_7/m2_11069_n223# RWL[28] xb[0] xa[1]
+ xa[7] xc LWL[26] men xa[0] xa[6] xb[3] xa[5] vss xb[2] vdd xc xdec8_256x8m81
Xxdec8_256x8m81_1 xa[5] xa[2] xdec8_256x8m81_1/RWL[0] LWL[5] LWL[4] RWL[2] RWL[1]
+ RWL[7] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0] LWL[3] RWL[3] xa[1] xa[7] xa[4] xa[3]
+ xb[0] xa[0] xa[6] RWL[5] xa[4] xb[1] xdec8_256x8m81_3/xdec_256x8m81_7/m2_10314_n223#
+ xdec8_256x8m81_3/xdec_256x8m81_7/m2_10691_n223# xa[2] xa[3] xdec8_256x8m81_3/xdec_256x8m81_7/m2_11069_n223#
+ RWL[4] xb[0] xa[1] xa[7] xc LWL[2] men xa[0] xa[6] xb[3] xa[5] vss xb[2] vdd xc
+ xdec8_256x8m81
Xxdec8_256x8m81_2 xa[5] xa[2] RWL[8] LWL[13] LWL[12] RWL[10] RWL[9] RWL[15] RWL[14]
+ LWL[9] LWL[15] LWL[14] LWL[8] LWL[11] RWL[11] xa[1] xa[7] xa[4] xa[3] xb[1] xa[0]
+ xa[6] RWL[13] xa[4] xb[1] xdec8_256x8m81_3/xdec_256x8m81_7/m2_10314_n223# xdec8_256x8m81_3/xdec_256x8m81_7/m2_10691_n223#
+ xa[2] xa[3] xdec8_256x8m81_3/xdec_256x8m81_7/m2_11069_n223# RWL[12] xb[0] xa[1]
+ xa[7] xc LWL[10] men xa[0] xa[6] xb[3] xa[5] vss xb[2] vdd xc xdec8_256x8m81
Xxdec8_256x8m81_3 xa[5] xa[2] RWL[16] LWL[21] LWL[20] RWL[18] RWL[17] RWL[23] RWL[22]
+ LWL[17] LWL[23] LWL[22] LWL[16] LWL[19] RWL[19] xa[1] xa[7] xa[4] xa[3] xb[2] xa[0]
+ xa[6] RWL[21] xa[4] xb[1] xdec8_256x8m81_3/xdec_256x8m81_7/m2_10314_n223# xdec8_256x8m81_3/xdec_256x8m81_7/m2_10691_n223#
+ xa[2] xa[3] xdec8_256x8m81_3/xdec_256x8m81_7/m2_11069_n223# RWL[20] xb[0] xa[1]
+ xa[7] xc LWL[18] men xa[0] xa[6] xb[3] xa[5] vss xb[2] vdd xc xdec8_256x8m81
.ends

.subckt pmoscap_W2_5_R270_256x8m81 w_n60_n407# a_81_507# m3_509_n1#
X0 a_81_507# M1_POLY2$$204395564_256x8m81_0/VSUBS a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_1p2$$204217388_256x8m81 w_n295_n137# pmos_5p043105908781101_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781101_256x8m81_0/S
Xpmos_5p043105908781101_256x8m81_0 w_n295_n137# pmos_5p043105908781101_256x8m81_0/D
+ a_n31_n71# pmos_5p043105908781101_256x8m81_0/S pmos_5p043105908781101_256x8m81
.ends

.subckt nmos_5p04310590878199_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=10.11u l=0.6u
.ends

.subckt nmos_5p043105908781111_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.64u l=0.6u
.ends

.subckt nmos_5p043105908781100_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.59u l=0.6u
.ends

.subckt nmos_1p2$$204215340_256x8m81 nmos_5p043105908781100_256x8m81_0/S nmos_5p043105908781100_256x8m81_0/D
+ a_n31_n71# VSUBS
Xnmos_5p043105908781100_256x8m81_0 nmos_5p043105908781100_256x8m81_0/D a_n31_n71#
+ nmos_5p043105908781100_256x8m81_0/S VSUBS nmos_5p043105908781100_256x8m81
.ends

.subckt nmos_1p2$$204213292_R90_256x8m81 nmos_5p04310590878199_256x8m81_0/S nmos_5p04310590878199_256x8m81_0/D
+ a_n31_n71# VSUBS
Xnmos_5p04310590878199_256x8m81_0 nmos_5p04310590878199_256x8m81_0/D a_n31_n71# nmos_5p04310590878199_256x8m81_0/S
+ VSUBS nmos_5p04310590878199_256x8m81
.ends

.subckt xdec32_256_256x8m81 DRWL RWL[31] RWL[29] RWL[6] RWL[2] RWL[0] RWL[5] RWL[7]
+ RWL[8] RWL[9] RWL[10] RWL[11] RWL[12] RWL[13] RWL[14] RWL[15] RWL[16] RWL[17] RWL[18]
+ LWL[30] LWL[31] LWL[20] LWL[21] LWL[22] LWL[13] LWL[15] LWL[16] LWL[18] LWL[5] LWL[4]
+ LWL[3] LWL[1] LWL[8] LWL[9] LWL[6] DLWL xb[0] xb[2] xb[3] xa[7] xa[6] xa[5] xa[4]
+ xa[0] xa[3] xa[2] xc[1] LWL[28] LWL[26] LWL[29] LWL[24] RWL[22] RWL[20] RWL[27]
+ LWL[27] LWL[14] xa[1] LWL[12] RWL[25] LWL[25] RWL[4] LWL[10] LWL[23] LWL[2] LWL[0]
+ LWL[11] xc[0] RWL[30] RWL[23] RWL[3] RWL[28] RWL[26] RWL[24] LWL[19] RWL[21] RWL[1]
+ xb[1] LWL[7] LWL[17] RWL[19] men vss vdd
Xpmos_5p043105908781101_256x8m81_0 vdd pmos_5p043105908781101_256x8m81_0/D vss men
+ pmos_5p043105908781101_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_30 RWL[3] RWL[2] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmos_5p043105908781101_256x8m81_1 vdd vdd pmos_5p043105908781101_256x8m81_0/D pmos_5p043105908781101_256x8m81_1/S
+ pmos_5p043105908781101_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_20 RWL[23] RWL[22] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_31 RWL[1] RWL[0] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_21 RWL[21] RWL[20] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_10 LWL[11] LWL[10] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmos_1p2$$204216364_256x8m81_0 DRWL vdd pmos_5p043105908781101_256x8m81_1/S vdd pmos_5p043105908781101_256x8m81_1/S
+ pmos_1p2$$204216364_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_22 RWL[19] RWL[18] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_23 RWL[17] RWL[16] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_12 LWL[7] LWL[6] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_11 LWL[9] LWL[8] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmos_1p2$$204216364_256x8m81_1 DLWL vdd nmos_5p043105908781111_256x8m81_1/S vdd nmos_5p043105908781111_256x8m81_1/S
+ pmos_1p2$$204216364_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_24 RWL[15] RWL[14] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_13 LWL[5] LWL[4] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_25 RWL[13] RWL[12] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_14 LWL[3] LWL[2] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xxdec32_256x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[16] RWL[15] RWL[14] RWL[13] RWL[12]
+ LWL[9] LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8]
+ RWL[7] RWL[5] RWL[3] RWL[1] RWL[0] RWL[2] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14]
+ LWL[13] LWL[11] LWL[10] RWL[4] RWL[6] LWL[28] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21]
+ LWL[20] LWL[19] RWL[20] RWL[21] RWL[22] RWL[23] RWL[24] RWL[25] RWL[28] RWL[29]
+ RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[0] xa[3] xa[4] xa[5] xa[6]
+ xa[7] xb[3] xb[2] xb[1] xb[0] xc[0] vdd vdd LWL[27] xc[1] LWL[26] RWL[27] men xa[1]
+ RWL[26] LWL[12] vss vdd xdec32_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_26 RWL[11] RWL[10] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_15 LWL[1] LWL[0] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_16 RWL[31] RWL[30] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_27 RWL[9] RWL[8] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_17 RWL[29] RWL[28] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_28 RWL[7] RWL[6] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_R270_256x8m81_1 vdd vdd DRWL pmoscap_W2_5_R270_256x8m81
Xpmoscap_W2_5_R270_256x8m81_0 vdd vdd DLWL pmoscap_W2_5_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_0 LWL[31] LWL[30] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_18 RWL[27] RWL[26] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_29 RWL[5] RWL[4] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmos_1p2$$204217388_256x8m81_0 vdd vdd pmos_5p043105908781101_256x8m81_0/D nmos_5p043105908781111_256x8m81_1/S
+ pmos_1p2$$204217388_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_1 LWL[29] LWL[28] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_19 RWL[25] RWL[24] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_2 LWL[27] LWL[26] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_3 LWL[25] LWL[24] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_4 LWL[23] LWL[22] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xnmos_5p04310590878199_256x8m81_0 vss pmos_5p043105908781101_256x8m81_1/S DRWL vss
+ nmos_5p04310590878199_256x8m81
Xnmos_5p043105908781111_256x8m81_0 vss pmos_5p043105908781101_256x8m81_0/D pmos_5p043105908781101_256x8m81_1/S
+ vss nmos_5p043105908781111_256x8m81
Xnmos_1p2$$204215340_256x8m81_0 pmos_5p043105908781101_256x8m81_0/D men vdd vss nmos_1p2$$204215340_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_5 LWL[21] LWL[20] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xnmos_5p043105908781111_256x8m81_1 vss pmos_5p043105908781101_256x8m81_0/D nmos_5p043105908781111_256x8m81_1/S
+ vss nmos_5p043105908781111_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_6 LWL[19] LWL[18] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_7 LWL[17] LWL[16] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xnmos_1p2$$204213292_R90_256x8m81_0 DLWL vss nmos_5p043105908781111_256x8m81_1/S vss
+ nmos_1p2$$204213292_R90_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_9 LWL[13] LWL[12] vdd vdd pmoscap_W2_5_477_R270_256x8m81
Xpmoscap_W2_5_477_R270_256x8m81_8 LWL[15] LWL[14] vdd vdd pmoscap_W2_5_477_R270_256x8m81
.ends

.subckt nmos_5p04310590878157_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.36u l=0.6u
.ends

.subckt nmos_1p2$$47342636_256x8m81 nmos_5p04310590878157_256x8m81_0/D a_n31_n73#
+ nmos_5p04310590878157_256x8m81_0/S VSUBS
Xnmos_5p04310590878157_256x8m81_0 nmos_5p04310590878157_256x8m81_0/D a_n31_n73# nmos_5p04310590878157_256x8m81_0/S
+ VSUBS nmos_5p04310590878157_256x8m81
.ends

.subckt pmos_5p04310590878165_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.77u l=0.6u
.ends

.subckt pmos_1p2$$47820844_256x8m81 pmos_5p04310590878165_256x8m81_0/S w_n286_n141#
+ pmos_5p04310590878165_256x8m81_0/D a_n30_n74#
Xpmos_5p04310590878165_256x8m81_0 w_n286_n141# pmos_5p04310590878165_256x8m81_0/D
+ a_n30_n74# pmos_5p04310590878165_256x8m81_0/S pmos_5p04310590878165_256x8m81
.ends

.subckt pmos_5p04310590878164_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$47821868_256x8m81 pmos_5p04310590878164_256x8m81_0/S w_n286_n142#
+ a_n31_n74# pmos_5p04310590878164_256x8m81_0/D
Xpmos_5p04310590878164_256x8m81_0 w_n286_n142# pmos_5p04310590878164_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878164_256x8m81_0/S pmos_5p04310590878164_256x8m81
.ends

.subckt ypredec1_xa_256x8m81 m1_n58_n4290# m1_n58_n4895# m1_n58_n5097# m3_n1_n7124#
+ a_644_n6680# m1_n58_n4492# m1_n58_n4088# a_421_n4311# a_n1_81# pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_197_n5120# m1_n58_n4694# pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ M3_M2$$47819820_256x8m81_0/VSUBS
Xpmos_1p2$$47820844_256x8m81_0 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D pmos_1p2$$47820844_256x8m81
Xpmos_1p2$$47820844_256x8m81_1 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D pmos_1p2$$47820844_256x8m81
Xpmos_1p2$$47820844_256x8m81_2 pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D pmos_1p2$$47820844_256x8m81
Xpmos_1p2$$47821868_256x8m81_0 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S a_197_n5120# pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D
+ pmos_1p2$$47821868_256x8m81
Xpmos_1p2$$47821868_256x8m81_1 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S a_421_n4311# pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81
Xpmos_1p2$$47821868_256x8m81_2 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S a_644_n6680# pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D
+ pmos_1p2$$47821868_256x8m81
Xnmos_1p2$$46551084_256x8m81_0 pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D M3_M2$$47819820_256x8m81_0/VSUBS
+ M3_M2$$47819820_256x8m81_0/VSUBS nmos_1p2$$46551084_256x8m81
Xnmos_1p2$$46551084_256x8m81_1 M3_M2$$47819820_256x8m81_0/VSUBS pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D
+ pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S M3_M2$$47819820_256x8m81_0/VSUBS
+ nmos_1p2$$46551084_256x8m81
Xnmos_1p2$$46551084_256x8m81_2 pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D M3_M2$$47819820_256x8m81_0/VSUBS
+ M3_M2$$47819820_256x8m81_0/VSUBS nmos_1p2$$46551084_256x8m81
X0 pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/D a_644_n6680# a_542_n6607# M3_M2$$47819820_256x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X1 a_318_n6607# a_197_n5120# M3_M2$$47819820_256x8m81_0/VSUBS M3_M2$$47819820_256x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X2 a_542_n6607# a_421_n4311# a_318_n6607# M3_M2$$47819820_256x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
.ends

.subckt ypredec1_xax8_256x8m81 ypredec1_xa_256x8m81_6/a_n1_81# ypredec1_xa_256x8m81_3/a_n1_81#
+ ypredec1_xa_256x8m81_7/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_0/a_n1_81# ypredec1_xa_256x8m81_6/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_5/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_7/a_n1_81# a_527_2758# ypredec1_xa_256x8m81_4/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_2/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_6100_2150# a_975_1949# ypredec1_xa_256x8m81_1/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_0/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xa_256x8m81_3/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_6324_2352# a_751_2554# a_303_2957# VSUBS ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
Xypredec1_xa_256x8m81_0 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_256x8m81_0/a_n1_81# ypredec1_xa_256x8m81_0/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_751_2554# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_1 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS ypredec1_xa_256x8m81_1/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_751_2554# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_2 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS ypredec1_xa_256x8m81_2/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_751_2554# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_3 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_256x8m81_3/a_n1_81# ypredec1_xa_256x8m81_3/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_751_2554# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_5 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS ypredec1_xa_256x8m81_5/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_975_1949# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_4 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_256x8m81_4/a_n1_81# ypredec1_xa_256x8m81_4/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_975_1949# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_6 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_256x8m81_6/a_n1_81# ypredec1_xa_256x8m81_6/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_975_1949# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
Xypredec1_xa_256x8m81_7 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_256x8m81_7/a_n1_81# ypredec1_xa_256x8m81_7/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ a_975_1949# a_6324_2352# ypredec1_xa_256x8m81_7/pmos_1p2$$47821868_256x8m81_2/pmos_5p04310590878164_256x8m81_0/S
+ VSUBS ypredec1_xa_256x8m81
.ends

.subckt nmos_5p04310590878158_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=9.08u l=0.6u
.ends

.subckt pmos_5p04310590878159_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=20u l=0.6u
.ends

.subckt ypredec1_ys_256x8m81 a_254_2184# pmos_5p04310590878159_256x8m81_3/S pmos_5p04310590878159_256x8m81_1/S
+ pmos_5p04310590878159_256x8m81_3/D nmos_5p04310590878158_256x8m81_1/D nmos_5p04310590878158_256x8m81_3/D
+ nmos_5p04310590878158_256x8m81_2/S VSUBS
Xnmos_5p04310590878158_256x8m81_3 nmos_5p04310590878158_256x8m81_3/D pmos_5p04310590878159_256x8m81_0/D
+ pmos_5p04310590878159_256x8m81_3/S VSUBS nmos_5p04310590878158_256x8m81
Xnmos_5p04310590878158_256x8m81_2 pmos_5p04310590878159_256x8m81_0/D a_254_2184# nmos_5p04310590878158_256x8m81_2/S
+ VSUBS nmos_5p04310590878158_256x8m81
Xpmos_5p04310590878159_256x8m81_2 pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81_3/S
+ pmos_5p04310590878159_256x8m81_0/D pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81
Xpmos_5p04310590878159_256x8m81_3 pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81_3/D
+ pmos_5p04310590878159_256x8m81_0/D pmos_5p04310590878159_256x8m81_3/S pmos_5p04310590878159_256x8m81
Xnmos_5p04310590878158_256x8m81_0 pmos_5p04310590878159_256x8m81_3/S pmos_5p04310590878159_256x8m81_0/D
+ nmos_5p04310590878158_256x8m81_1/D VSUBS nmos_5p04310590878158_256x8m81
Xpmos_5p04310590878159_256x8m81_0 pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81_0/D
+ a_254_2184# pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81
Xnmos_5p04310590878158_256x8m81_1 nmos_5p04310590878158_256x8m81_1/D pmos_5p04310590878159_256x8m81_0/D
+ pmos_5p04310590878159_256x8m81_1/S VSUBS nmos_5p04310590878158_256x8m81
Xpmos_5p04310590878159_256x8m81_1 pmos_5p04310590878159_256x8m81_3/D pmos_5p04310590878159_256x8m81_3/D
+ pmos_5p04310590878159_256x8m81_0/D pmos_5p04310590878159_256x8m81_1/S pmos_5p04310590878159_256x8m81
.ends

.subckt nmos_5p04310590878161_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=4.54u l=0.6u
.ends

.subckt nmos_1p2$$47514668_256x8m81 nmos_5p04310590878161_256x8m81_0/S a_n30_n73#
+ VSUBS nmos_5p04310590878161_256x8m81_0/D
Xnmos_5p04310590878161_256x8m81_0 nmos_5p04310590878161_256x8m81_0/D a_n30_n73# nmos_5p04310590878161_256x8m81_0/S
+ VSUBS nmos_5p04310590878161_256x8m81
.ends

.subckt pmos_1p2$$46285868_160_256x8m81 pmos_5p04310590878114_256x8m81_0/D a_n31_n74#
+ pmos_5p04310590878114_256x8m81_0/S w_n286_n142#
Xpmos_5p04310590878114_256x8m81_0 w_n286_n142# pmos_5p04310590878114_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878114_256x8m81_0/S pmos_5p04310590878114_256x8m81
.ends

.subckt pmos_1p2$$47330348_161_256x8m81 pmos_5p04310590878141_256x8m81_0/S a_n31_191#
+ w_n286_n141# pmos_5p04310590878141_256x8m81_0/D
Xpmos_5p04310590878141_256x8m81_0 w_n286_n141# pmos_5p04310590878141_256x8m81_0/D
+ a_n31_191# pmos_5p04310590878141_256x8m81_0/S pmos_5p04310590878141_256x8m81
.ends

.subckt nmos_5p04310590878162_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.82u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.82u l=0.6u
.ends

.subckt nmos_1p2$$47329324_256x8m81 a_194_n74# nmos_5p04310590878162_256x8m81_0/S
+ nmos_5p04310590878162_256x8m81_0/D a_n30_n74# VSUBS
Xnmos_5p04310590878162_256x8m81_0 nmos_5p04310590878162_256x8m81_0/D a_n30_n74# nmos_5p04310590878162_256x8m81_0/S
+ a_194_n74# VSUBS nmos_5p04310590878162_256x8m81
.ends

.subckt nmos_1p2$$46551084_157_256x8m81 nmos_5p04310590878110_256x8m81_0/D a_n31_n74#
+ nmos_5p04310590878110_256x8m81_0/S VSUBS
Xnmos_5p04310590878110_256x8m81_0 nmos_5p04310590878110_256x8m81_0/D a_n31_n74# nmos_5p04310590878110_256x8m81_0/S
+ VSUBS nmos_5p04310590878110_256x8m81
.ends

.subckt pmos_5p04310590878163_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$47331372_256x8m81 pmos_5p04310590878163_256x8m81_0/D a_n30_n74#
+ w_n286_n142# pmos_5p04310590878163_256x8m81_0/S a_194_n74#
Xpmos_5p04310590878163_256x8m81_0 w_n286_n142# pmos_5p04310590878163_256x8m81_0/D
+ a_n30_n74# pmos_5p04310590878163_256x8m81_0/S a_194_n74# pmos_5p04310590878163_256x8m81
.ends

.subckt alatch_256x8m81 enb en ab a vss vdd
Xpmos_1p2$$46285868_160_256x8m81_0 a enb nmos_5p0431059087818_256x8m81_1/S vdd pmos_1p2$$46285868_160_256x8m81
Xpmos_1p2$$47330348_161_256x8m81_0 nmos_5p0431059087818_256x8m81_1/S en vdd nmos_5p0431059087818_256x8m81_1/D
+ pmos_1p2$$47330348_161_256x8m81
Xpmos_1p2$$47330348_161_256x8m81_1 nmos_5p0431059087818_256x8m81_1/D ab vdd vdd pmos_1p2$$47330348_161_256x8m81
Xnmos_5p0431059087818_256x8m81_0 vss ab nmos_5p0431059087818_256x8m81_1/D vss nmos_5p0431059087818_256x8m81
Xnmos_5p0431059087818_256x8m81_1 nmos_5p0431059087818_256x8m81_1/D enb nmos_5p0431059087818_256x8m81_1/S
+ vss nmos_5p0431059087818_256x8m81
Xnmos_1p2$$47329324_256x8m81_0 nmos_5p0431059087818_256x8m81_1/S vss ab nmos_5p0431059087818_256x8m81_1/S
+ vss nmos_1p2$$47329324_256x8m81
Xnmos_1p2$$46551084_157_256x8m81_0 a en nmos_5p0431059087818_256x8m81_1/S vss nmos_1p2$$46551084_157_256x8m81
Xpmos_1p2$$47331372_256x8m81_0 ab nmos_5p0431059087818_256x8m81_1/S vdd vdd nmos_5p0431059087818_256x8m81_1/S
+ pmos_1p2$$47331372_256x8m81
.ends

.subckt ypredec1_bot_256x8m81 m1_n14_3279# m1_n14_2674# alatch_256x8m81_0/a pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ m1_n14_2876# m1_n14_3078# m1_n14_3481# pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ m1_n14_2472# pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D alatch_256x8m81_0/vdd
+ alatch_256x8m81_0/vss alatch_256x8m81_0/en alatch_256x8m81_0/enb
Xpmos_1p2$$46887980_256x8m81_0 pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S pmos_1p2$$46887980_256x8m81
Xpmos_1p2$$46887980_256x8m81_1 pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ alatch_256x8m81_0/ab pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S pmos_1p2$$46887980_256x8m81
Xnmos_1p2$$47514668_256x8m81_0 alatch_256x8m81_0/vss pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ alatch_256x8m81_0/vss pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ nmos_1p2$$47514668_256x8m81
Xnmos_1p2$$47514668_256x8m81_1 alatch_256x8m81_0/vss alatch_256x8m81_0/ab alatch_256x8m81_0/vss
+ pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D nmos_1p2$$47514668_256x8m81
Xalatch_256x8m81_0 alatch_256x8m81_0/enb alatch_256x8m81_0/en alatch_256x8m81_0/ab
+ alatch_256x8m81_0/a alatch_256x8m81_0/vss alatch_256x8m81_0/vdd alatch_256x8m81
.ends

.subckt pmos_5p04310590878166_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$47109164_256x8m81 pmos_5p04310590878166_256x8m81_0/S a_n31_341#
+ pmos_5p04310590878166_256x8m81_0/D pmos_5p04310590878166_256x8m81_0/w_n208_n120#
+ a_193_341#
Xpmos_5p04310590878166_256x8m81_0 pmos_5p04310590878166_256x8m81_0/w_n208_n120# pmos_5p04310590878166_256x8m81_0/D
+ a_n31_341# pmos_5p04310590878166_256x8m81_0/S a_193_341# pmos_5p04310590878166_256x8m81
.ends

.subckt nmos_5p04310590878160_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.91u l=0.6u
.ends

.subckt ypredec1_256x8m81 ly[5] ly[4] ly[7] ly[3] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd
+ pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120# ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ ypredec1_ys_256x8m81_9/VSUBS pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S
Xnmos_1p2$$47342636_256x8m81_0 ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81_1/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/enb ypredec1_ys_256x8m81_9/VSUBS nmos_1p2$$47342636_256x8m81
Xypredec1_xax8_256x8m81_0 ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_7/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_6/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_5/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_4/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_2/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_1/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_0/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_3/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ ypredec1_xax8_256x8m81
Xypredec1_ys_256x8m81_0 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_5/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[0] ly[0] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_1 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_1/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[1] ly[1] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_2 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_4/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[2] ly[2] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_bot_256x8m81_0 ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ A[0] ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81_1/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/enb ypredec1_bot_256x8m81
Xpmos_1p2$$47109164_256x8m81_0 pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S
+ nmos_5p04310590878160_256x8m81_1/D ypredec1_bot_256x8m81_2/alatch_256x8m81_0/enb
+ pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120# nmos_5p04310590878160_256x8m81_1/D
+ pmos_1p2$$47109164_256x8m81
Xypredec1_bot_256x8m81_1 ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ A[2] ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81_1/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/enb ypredec1_bot_256x8m81
Xypredec1_ys_256x8m81_3 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_0/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[3] ly[3] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_4 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_6/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[4] ly[4] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_bot_256x8m81_2 ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ A[1] ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/S
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_1/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_1/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_0/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/pmos_1p2$$46887980_256x8m81_0/pmos_5p0431059087814_256x8m81_0/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81_1/D
+ ypredec1_bot_256x8m81_2/alatch_256x8m81_0/enb ypredec1_bot_256x8m81
Xypredec1_ys_256x8m81_5 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_2/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[5] ly[5] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_6 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_7/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[6] ly[6] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_10 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_6/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[4] ry[4] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xnmos_5p04310590878160_256x8m81_0 ypredec1_ys_256x8m81_9/VSUBS clk nmos_5p04310590878160_256x8m81_1/D
+ ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81
Xnmos_5p04310590878160_256x8m81_1 nmos_5p04310590878160_256x8m81_1/D men ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS nmos_5p04310590878160_256x8m81
Xypredec1_ys_256x8m81_7 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_1/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[1] ry[1] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_11 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_2/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[5] ry[5] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_12 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_7/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[6] ry[6] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_8 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_4/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[2] ry[2] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_13 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_3/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[7] ry[7] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_9 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_0/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[3] ry[3] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_14 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_5/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ry[0] ry[0] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
Xypredec1_ys_256x8m81_15 ypredec1_xax8_256x8m81_0/ypredec1_xa_256x8m81_3/pmos_1p2$$47820844_256x8m81_2/pmos_5p04310590878165_256x8m81_0/S
+ ly[7] ly[7] ypredec1_ys_256x8m81_9/pmos_5p04310590878159_256x8m81_3/D ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS ypredec1_ys_256x8m81_9/VSUBS
+ ypredec1_ys_256x8m81
X0 a_7843_267# clk nmos_5p04310590878160_256x8m81_1/D pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X1 nmos_5p04310590878160_256x8m81_1/D clk a_7395_267# pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X2 a_7395_267# men pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X3 pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S men a_7843_267# pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/S pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310590878176_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.43u l=0.6u
.ends

.subckt pmos_1p2$$47512620_256x8m81 pmos_5p04310590878176_256x8m81_0/S a_n30_n74#
+ w_n286_n142# pmos_5p04310590878176_256x8m81_0/D
Xpmos_5p04310590878176_256x8m81_0 w_n286_n142# pmos_5p04310590878176_256x8m81_0/D
+ a_n30_n74# pmos_5p04310590878176_256x8m81_0/S pmos_5p04310590878176_256x8m81
.ends

.subckt pmos_5p04310590878168_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt pmos_1p2$$47513644_256x8m81 pmos_5p04310590878168_256x8m81_0/D a_n30_n74#
+ w_n286_n141# pmos_5p04310590878168_256x8m81_0/S
Xpmos_5p04310590878168_256x8m81_0 w_n286_n141# pmos_5p04310590878168_256x8m81_0/D
+ a_n30_n74# pmos_5p04310590878168_256x8m81_0/S pmos_5p04310590878168_256x8m81
.ends

.subckt xpredec1_xa_256x8m81 a_197_n10255# m1_n58_n7539# a_421_n10255# m1_n58_n6933#
+ a_645_n10255# m1_n58_n7135# m1_n58_n6530# m1_n58_n7337# a_n1_81# pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ m1_n58_n6732# M3_M2$$47333420_256x8m81_1/VSUBS pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
Xpmos_1p2$$47512620_256x8m81_0 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ a_645_n10255# pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D
+ pmos_1p2$$47512620_256x8m81
Xpmos_1p2$$47512620_256x8m81_2 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ a_197_n10255# pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D
+ pmos_1p2$$47512620_256x8m81
Xpmos_1p2$$47512620_256x8m81_1 pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D
+ a_421_n10255# pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47512620_256x8m81
Xnmos_1p2$$47514668_256x8m81_0 M3_M2$$47333420_256x8m81_1/VSUBS pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D
+ M3_M2$$47333420_256x8m81_1/VSUBS pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ nmos_1p2$$47514668_256x8m81
Xnmos_1p2$$47514668_256x8m81_1 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D M3_M2$$47333420_256x8m81_1/VSUBS
+ M3_M2$$47333420_256x8m81_1/VSUBS nmos_1p2$$47514668_256x8m81
Xnmos_1p2$$47514668_256x8m81_2 M3_M2$$47333420_256x8m81_1/VSUBS pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D
+ M3_M2$$47333420_256x8m81_1/VSUBS pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ nmos_1p2$$47514668_256x8m81
Xpmos_1p2$$47513644_256x8m81_0 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47513644_256x8m81_1 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47513644_256x8m81_2 pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/D
+ pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47513644_256x8m81_2/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47513644_256x8m81
X0 pmos_1p2$$47512620_256x8m81_2/pmos_5p04310590878176_256x8m81_0/D a_645_n10255# a_541_n10182# M3_M2$$47333420_256x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X1 a_317_n10182# a_197_n10255# M3_M2$$47333420_256x8m81_1/VSUBS M3_M2$$47333420_256x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X2 a_541_n10182# a_421_n10255# a_317_n10182# M3_M2$$47333420_256x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
.ends

.subckt nmos_5p04310590878175_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.58u l=0.6u
.ends

.subckt nmos_1p2$$47336492_256x8m81 nmos_5p04310590878175_256x8m81_0/S nmos_5p04310590878175_256x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p04310590878175_256x8m81_0 nmos_5p04310590878175_256x8m81_0/D a_n31_n74# nmos_5p04310590878175_256x8m81_0/S
+ VSUBS nmos_5p04310590878175_256x8m81
.ends

.subckt pmos_5p04310590878174_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=16.33u l=0.6u
.ends

.subckt pmos_1p2$$47337516_256x8m81 pmos_5p04310590878174_256x8m81_0/D a_n31_n73#
+ w_n286_n141# pmos_5p04310590878174_256x8m81_0/S
Xpmos_5p04310590878174_256x8m81_0 w_n286_n141# pmos_5p04310590878174_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878174_256x8m81_0/S pmos_5p04310590878174_256x8m81
.ends

.subckt xpredec1_bot_256x8m81 m1_n106_2472# m1_n106_3279# alatch_256x8m81_0/a m1_n106_2674#
+ pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D alatch_256x8m81_0/vdd
+ m1_n106_2876# alatch_256x8m81_0/enb pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ alatch_256x8m81_0/en m1_n106_3078# m1_n106_3481# VSUBS pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/S
Xnmos_1p2$$47336492_256x8m81_0 VSUBS pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D VSUBS nmos_1p2$$47336492_256x8m81
Xpmos_1p2$$47337516_256x8m81_0 pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/S
+ pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/S pmos_1p2$$47337516_256x8m81
Xnmos_1p2$$47336492_256x8m81_1 VSUBS pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ alatch_256x8m81_0/ab VSUBS nmos_1p2$$47336492_256x8m81
Xpmos_1p2$$47337516_256x8m81_1 pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ alatch_256x8m81_0/ab pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/S
+ pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/S pmos_1p2$$47337516_256x8m81
Xalatch_256x8m81_0 alatch_256x8m81_0/enb alatch_256x8m81_0/en alatch_256x8m81_0/ab
+ alatch_256x8m81_0/a VSUBS alatch_256x8m81_0/vdd alatch_256x8m81
.ends

.subckt xpredec1_256x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1] A[0]
+ clk w_7178_9364# pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120#
+ vdd vss
Xnmos_1p2$$47342636_256x8m81_0 vss nmos_5p04310590878160_256x8m81_1/D xpredec1_bot_256x8m81_2/alatch_256x8m81_0/enb
+ vss nmos_1p2$$47342636_256x8m81
Xpmos_1p2$$47109164_256x8m81_0 vdd nmos_5p04310590878160_256x8m81_1/D xpredec1_bot_256x8m81_2/alatch_256x8m81_0/enb
+ pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120# nmos_5p04310590878160_256x8m81_1/D
+ pmos_1p2$$47109164_256x8m81
Xnmos_5p04310590878160_256x8m81_0 vss clk nmos_5p04310590878160_256x8m81_1/D vss nmos_5p04310590878160_256x8m81
Xxpredec1_xa_256x8m81_0 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ vss x[3] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xnmos_5p04310590878160_256x8m81_1 nmos_5p04310590878160_256x8m81_1/D men vss vss nmos_5p04310590878160_256x8m81
Xxpredec1_xa_256x8m81_1 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_xa_256x8m81_1/a_n1_81# x[1] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_xa_256x8m81_2 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ vss x[5] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_bot_256x8m81_0 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ A[0] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vdd xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/alatch_256x8m81_0/enb xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ nmos_5p04310590878160_256x8m81_1/D xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_bot_256x8m81
Xxpredec1_xa_256x8m81_3 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_xa_256x8m81_3/a_n1_81# x[7] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_bot_256x8m81_1 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ A[2] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vdd xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/alatch_256x8m81_0/enb xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ nmos_5p04310590878160_256x8m81_1/D xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_bot_256x8m81
Xxpredec1_xa_256x8m81_5 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ vss x[0] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_xa_256x8m81_4 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ vss x[2] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_bot_256x8m81_2 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ A[1] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vdd xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/alatch_256x8m81_0/enb xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ nmos_5p04310590878160_256x8m81_1/D xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_bot_256x8m81
Xxpredec1_xa_256x8m81_6 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ vss x[4] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
Xxpredec1_xa_256x8m81_7 xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_0/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_1/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_0/pmos_5p04310590878174_256x8m81_0/D
+ xpredec1_xa_256x8m81_7/a_n1_81# x[6] xpredec1_bot_256x8m81_2/pmos_1p2$$47337516_256x8m81_1/pmos_5p04310590878174_256x8m81_0/D
+ vss vdd xpredec1_xa_256x8m81
X0 nmos_5p04310590878160_256x8m81_1/D clk a_7553_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X1 a_7553_9505# men vdd w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X2 a_8001_9505# clk nmos_5p04310590878160_256x8m81_1/D w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X3 vdd men a_8001_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
.ends

.subckt nmos_5p04310590878170_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=5.22u l=0.6u
.ends

.subckt nmos_1p2$$47502380_256x8m81 nmos_5p04310590878170_256x8m81_0/S nmos_5p04310590878170_256x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p04310590878170_256x8m81_0 nmos_5p04310590878170_256x8m81_0/D a_n31_n74# nmos_5p04310590878170_256x8m81_0/S
+ VSUBS nmos_5p04310590878170_256x8m81
.ends

.subckt pmos_5p04310590878169_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=17.69u l=0.6u
.ends

.subckt pmos_1p2$$47503404_256x8m81 a_n31_n73# pmos_5p04310590878169_256x8m81_0/S
+ w_n286_n141# pmos_5p04310590878169_256x8m81_0/D
Xpmos_5p04310590878169_256x8m81_0 w_n286_n141# pmos_5p04310590878169_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878169_256x8m81_0/S pmos_5p04310590878169_256x8m81
.ends

.subckt nmos_5p04310590878172_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=7.04u l=0.6u
.ends

.subckt pmos_5p04310590878171_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.16u l=0.6u
.ends

.subckt pmos_1p2$$47504428_256x8m81 pmos_5p04310590878171_256x8m81_0/S w_n286_n142#
+ pmos_5p04310590878171_256x8m81_0/w_n208_n120# pmos_5p04310590878171_256x8m81_0/D
+ a_n31_n73#
Xpmos_5p04310590878171_256x8m81_0 pmos_5p04310590878171_256x8m81_0/w_n208_n120# pmos_5p04310590878171_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878171_256x8m81_0/S pmos_5p04310590878171_256x8m81
.ends

.subckt xpredec0_bot_256x8m81 m1_n106_2472# pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ alatch_256x8m81_0/a nmos_5p04310590878172_256x8m81_0/D pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S
+ m1_n106_2674# alatch_256x8m81_0/vdd m1_n106_2876# alatch_256x8m81_0/enb alatch_256x8m81_0/en
+ m1_n106_3078# VSUBS
Xnmos_1p2$$47502380_256x8m81_0 VSUBS pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ nmos_5p04310590878172_256x8m81_0/D VSUBS nmos_1p2$$47502380_256x8m81
Xpmos_1p2$$47503404_256x8m81_0 alatch_256x8m81_0/ab pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S
+ pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S nmos_5p04310590878172_256x8m81_0/D
+ pmos_1p2$$47503404_256x8m81
Xnmos_5p04310590878172_256x8m81_0 nmos_5p04310590878172_256x8m81_0/D alatch_256x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310590878172_256x8m81
Xpmos_1p2$$47504428_256x8m81_0 pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S
+ pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/S
+ pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D nmos_5p04310590878172_256x8m81_0/D
+ pmos_1p2$$47504428_256x8m81
Xalatch_256x8m81_0 alatch_256x8m81_0/enb alatch_256x8m81_0/en alatch_256x8m81_0/ab
+ alatch_256x8m81_0/a VSUBS alatch_256x8m81_0/vdd alatch_256x8m81
.ends

.subckt nmos_1p2$$47641644_256x8m81 a_n31_n73# nmos_5p04310590878161_256x8m81_0/S
+ VSUBS nmos_5p04310590878161_256x8m81_0/D
Xnmos_5p04310590878161_256x8m81_0 nmos_5p04310590878161_256x8m81_0/D a_n31_n73# nmos_5p04310590878161_256x8m81_0/S
+ VSUBS nmos_5p04310590878161_256x8m81
.ends

.subckt pmos_5p04310590878167_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=15.2u l=0.6u
.ends

.subckt pmos_1p2$$47642668_256x8m81 w_n546_n142# pmos_5p04310590878167_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878167_256x8m81_0/S
Xpmos_5p04310590878167_256x8m81_0 w_n546_n142# pmos_5p04310590878167_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878167_256x8m81_0/S pmos_5p04310590878167_256x8m81
.ends

.subckt pmos_1p2$$47643692_256x8m81 pmos_5p04310590878167_256x8m81_0/D w_n286_n142#
+ a_n31_n74# pmos_5p04310590878167_256x8m81_0/S
Xpmos_5p04310590878167_256x8m81_0 w_n286_n142# pmos_5p04310590878167_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878167_256x8m81_0/S pmos_5p04310590878167_256x8m81
.ends

.subckt xpredec0_xa_256x8m81 m1_342_3273# a_875_414# m3_855_1044# a_651_414# nmos_1p2$$47641644_256x8m81_3/nmos_5p04310590878161_256x8m81_0/D
+ nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S m1_342_3474# pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D
+ m3_153_8117# m1_342_3071# m1_342_3676# M3_M2$$47644716_256x8m81_2/VSUBS pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/S
Xnmos_1p2$$47641644_256x8m81_0 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S
+ nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S M3_M2$$47644716_256x8m81_2/VSUBS
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D nmos_1p2$$47641644_256x8m81
Xnmos_1p2$$47641644_256x8m81_1 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S
+ nmos_1p2$$47641644_256x8m81_3/nmos_5p04310590878161_256x8m81_0/D M3_M2$$47644716_256x8m81_2/VSUBS
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D nmos_1p2$$47641644_256x8m81
Xnmos_1p2$$47641644_256x8m81_2 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D M3_M2$$47644716_256x8m81_2/VSUBS
+ nmos_1p2$$47641644_256x8m81_3/nmos_5p04310590878161_256x8m81_0/D nmos_1p2$$47641644_256x8m81
Xnmos_1p2$$47641644_256x8m81_3 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D M3_M2$$47644716_256x8m81_2/VSUBS
+ nmos_1p2$$47641644_256x8m81_3/nmos_5p04310590878161_256x8m81_0/D nmos_1p2$$47641644_256x8m81
Xpmos_1p2$$47513644_256x8m81_0 pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47513644_256x8m81_1 pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47513644_256x8m81_3 pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/S pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47513644_256x8m81_2 pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/S
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47513644_256x8m81_3/pmos_5p04310590878168_256x8m81_0/D pmos_1p2$$47513644_256x8m81
Xpmos_1p2$$47642668_256x8m81_0 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S a_875_414# pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47642668_256x8m81
Xpmos_1p2$$47643692_256x8m81_0 pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D
+ pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/D a_651_414# pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S
+ pmos_1p2$$47643692_256x8m81
X0 a_771_486# a_651_414# pmos_1p2$$47643692_256x8m81_0/pmos_5p04310590878167_256x8m81_0/S M3_M2$$47644716_256x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
X1 M3_M2$$47644716_256x8m81_2/VSUBS a_875_414# a_771_486# M3_M2$$47644716_256x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
.ends

.subckt pmos_5p04310590878173_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt xpredec0_256x8m81 A[0] men x[1] x[3] A[1] clk xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ x[2] x[0] xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ vss vdd
Xxpredec0_bot_256x8m81_1 xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ A[1] xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vdd xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ vdd xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ pmos_5p04310590878173_256x8m81_0/D nmos_5p04310590878140_256x8m81_1/S xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D
+ vss xpredec0_bot_256x8m81
Xxpredec0_xa_256x8m81_0 xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ vdd xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ vss xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ x[0] vss xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vss vdd vdd xpredec0_xa_256x8m81
Xxpredec0_xa_256x8m81_1 xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ vdd xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vss xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ x[2] vss xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vss vdd vdd xpredec0_xa_256x8m81
Xxpredec0_xa_256x8m81_2 xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D vdd xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ vss xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ x[1] vss xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vss vdd vdd xpredec0_xa_256x8m81
Xxpredec0_xa_256x8m81_3 xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D vdd xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D
+ vss xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ x[3] vss xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D vss vdd vdd xpredec0_xa_256x8m81
Xpmos_5p04310590878173_256x8m81_0 vdd pmos_5p04310590878173_256x8m81_0/D nmos_5p04310590878140_256x8m81_1/S
+ vdd nmos_5p04310590878140_256x8m81_1/S pmos_5p04310590878173_256x8m81
Xnmos_5p04310590878140_256x8m81_0 nmos_5p04310590878140_256x8m81_1/S men vss vss nmos_5p04310590878140_256x8m81
Xnmos_1p2$$46563372_256x8m81_0 vss nmos_5p04310590878140_256x8m81_1/S pmos_5p04310590878173_256x8m81_0/D
+ vss nmos_1p2$$46563372_256x8m81
Xnmos_5p04310590878140_256x8m81_1 vss clk nmos_5p04310590878140_256x8m81_1/S vss nmos_5p04310590878140_256x8m81
Xxpredec0_bot_256x8m81_0 xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ xpredec0_bot_256x8m81_0/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ A[0] xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D vdd xpredec0_bot_256x8m81_0/nmos_5p04310590878172_256x8m81_0/D
+ vdd xpredec0_bot_256x8m81_1/pmos_1p2$$47504428_256x8m81_0/pmos_5p04310590878171_256x8m81_0/D
+ pmos_5p04310590878173_256x8m81_0/D nmos_5p04310590878140_256x8m81_1/S xpredec0_bot_256x8m81_1/nmos_5p04310590878172_256x8m81_0/D
+ vss xpredec0_bot_256x8m81
X0 vdd men a_4894_9505# vdd pmos_3p3 w=1.705u l=0.6u
X1 a_4446_9505# men vdd vdd pmos_3p3 w=1.705u l=0.6u
X2 a_4894_9505# clk nmos_5p04310590878140_256x8m81_1/S vdd pmos_3p3 w=1.705u l=0.6u
X3 nmos_5p04310590878140_256x8m81_1/S clk a_4446_9505# vdd pmos_3p3 w=1.705u l=0.6u
.ends

.subckt prexdec_top_256x8m81 clk A[2] A[6] A[4] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1]
+ xb[2] xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1] xpredec1_256x8m81_0/pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120#
+ xpredec0_256x8m81_0/xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_256x8m81_0/xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_256x8m81_1/xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xpredec0_256x8m81_1/xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xc[0] xpredec1_256x8m81_0/w_7178_9364# men xpredec1_256x8m81_0/vdd VSUBS
Xxpredec1_256x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] clk xpredec1_256x8m81_0/w_7178_9364# xpredec1_256x8m81_0/pmos_1p2$$47109164_256x8m81_0/pmos_5p04310590878166_256x8m81_0/w_n208_n120#
+ xpredec1_256x8m81_0/vdd VSUBS xpredec1_256x8m81
Xxpredec0_256x8m81_0 A[3] men xb[1] xb[3] A[4] clk xpredec0_256x8m81_0/xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xb[2] xb[0] xpredec0_256x8m81_0/xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ VSUBS xpredec1_256x8m81_0/vdd xpredec0_256x8m81
Xxpredec0_256x8m81_1 A[5] men xc[1] xc[3] A[6] clk xpredec0_256x8m81_1/xpredec0_xa_256x8m81_3/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ xc[2] xc[0] xpredec0_256x8m81_1/xpredec0_xa_256x8m81_2/nmos_1p2$$47641644_256x8m81_0/nmos_5p04310590878161_256x8m81_0/S
+ VSUBS xpredec1_256x8m81_0/vdd xpredec0_256x8m81
.ends

.subckt pmos_5p04310590878178_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1.2u
.ends

.subckt pmos_5p04310590878196_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1u
.ends

.subckt pmos_5p04310590878195_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=19.5u l=0.6u
.ends

.subckt pmos_1p2$$48624684_256x8m81 pmos_5p04310590878195_256x8m81_0/S w_n286_n141#
+ a_n31_n74# pmos_5p04310590878195_256x8m81_0/D
Xpmos_5p04310590878195_256x8m81_0 w_n286_n141# pmos_5p04310590878195_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878195_256x8m81_0/S pmos_5p04310590878195_256x8m81
.ends

.subckt nmos_5p04310590878188_256x8m81 a_2464_n44# D a_2240_n44# a_3584_n44# a_2016_n44#
+ a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44# a_3808_n44#
+ a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44#
+ a_1120_n44# a_2688_n44# VSUBS
X0 S a_4256_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X1 S a_224_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X2 D a_448_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X3 D a_0_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X4 S a_2912_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X5 D a_3136_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X6 S a_672_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X7 D a_896_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X8 S a_3360_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X9 S a_2016_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X10 D a_3584_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X11 D a_2240_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X12 S a_2464_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X13 D a_2688_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X14 S a_1120_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X15 D a_1344_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X16 S a_1568_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X17 D a_1792_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X18 S a_3808_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X19 D a_4032_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
.ends

.subckt nmos_1p2$$48308268_256x8m81 nmos_5p04310590878188_256x8m81_0/a_3136_n44# nmos_5p04310590878188_256x8m81_0/a_2912_n44#
+ nmos_5p04310590878188_256x8m81_0/a_4256_n44# nmos_5p04310590878188_256x8m81_0/D
+ nmos_5p04310590878188_256x8m81_0/a_4032_n44# nmos_5p04310590878188_256x8m81_0/a_3808_n44#
+ nmos_5p04310590878188_256x8m81_0/a_0_n44# nmos_5p04310590878188_256x8m81_0/a_1792_n44#
+ nmos_5p04310590878188_256x8m81_0/a_1568_n44# nmos_5p04310590878188_256x8m81_0/a_896_n44#
+ nmos_5p04310590878188_256x8m81_0/a_672_n44# nmos_5p04310590878188_256x8m81_0/a_1344_n44#
+ nmos_5p04310590878188_256x8m81_0/a_1120_n44# nmos_5p04310590878188_256x8m81_0/a_448_n44#
+ nmos_5p04310590878188_256x8m81_0/a_2688_n44# nmos_5p04310590878188_256x8m81_0/a_224_n44#
+ nmos_5p04310590878188_256x8m81_0/a_2464_n44# nmos_5p04310590878188_256x8m81_0/a_2240_n44#
+ nmos_5p04310590878188_256x8m81_0/S nmos_5p04310590878188_256x8m81_0/a_2016_n44#
+ nmos_5p04310590878188_256x8m81_0/a_3584_n44# VSUBS nmos_5p04310590878188_256x8m81_0/a_3360_n44#
Xnmos_5p04310590878188_256x8m81_0 nmos_5p04310590878188_256x8m81_0/a_2464_n44# nmos_5p04310590878188_256x8m81_0/D
+ nmos_5p04310590878188_256x8m81_0/a_2240_n44# nmos_5p04310590878188_256x8m81_0/a_3584_n44#
+ nmos_5p04310590878188_256x8m81_0/a_2016_n44# nmos_5p04310590878188_256x8m81_0/a_3360_n44#
+ nmos_5p04310590878188_256x8m81_0/a_3136_n44# nmos_5p04310590878188_256x8m81_0/a_2912_n44#
+ nmos_5p04310590878188_256x8m81_0/a_0_n44# nmos_5p04310590878188_256x8m81_0/a_4256_n44#
+ nmos_5p04310590878188_256x8m81_0/a_4032_n44# nmos_5p04310590878188_256x8m81_0/a_3808_n44#
+ nmos_5p04310590878188_256x8m81_0/a_896_n44# nmos_5p04310590878188_256x8m81_0/a_672_n44#
+ nmos_5p04310590878188_256x8m81_0/S nmos_5p04310590878188_256x8m81_0/a_1792_n44#
+ nmos_5p04310590878188_256x8m81_0/a_448_n44# nmos_5p04310590878188_256x8m81_0/a_224_n44#
+ nmos_5p04310590878188_256x8m81_0/a_1568_n44# nmos_5p04310590878188_256x8m81_0/a_1344_n44#
+ nmos_5p04310590878188_256x8m81_0/a_1120_n44# nmos_5p04310590878188_256x8m81_0/a_2688_n44#
+ VSUBS nmos_5p04310590878188_256x8m81
.ends

.subckt nmos_5p04310590878194_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1u
.ends

.subckt pmos_5p04310590878191_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=22.68u l=0.6u
.ends

.subckt pmos_1p2$$47815724_256x8m81 pmos_5p04310590878191_256x8m81_0/S pmos_5p04310590878191_256x8m81_0/D
+ w_n286_n141# a_n31_n74#
Xpmos_5p04310590878191_256x8m81_0 w_n286_n141# pmos_5p04310590878191_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878191_256x8m81_0/S pmos_5p04310590878191_256x8m81
.ends

.subckt pmos_5p04310590878193_256x8m81 a_2464_n44# w_n208_n120# D a_2240_n44# a_3584_n44#
+ a_2016_n44# a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44#
+ a_3808_n44# a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44#
+ a_1344_n44# a_1120_n44# a_2688_n44#
X0 D a_4032_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X1 S a_4256_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X2 S a_224_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X3 D a_448_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X4 D a_0_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X5 S a_2912_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X6 D a_3136_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X7 S a_672_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X8 D a_896_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X9 S a_3360_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X10 S a_2016_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X11 D a_3584_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X12 D a_2240_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X13 S a_2464_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X14 D a_2688_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X15 S a_1120_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X16 D a_1344_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X17 S a_1568_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X18 D a_1792_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X19 S a_3808_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
.ends

.subckt nmos_5p04310590878185_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
.ends

.subckt pmos_5p04310590878186_256x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
.ends

.subckt pmos_5p04310590878184_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310590878182_256x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_5p04310590878183_256x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X6 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310590878180_256x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310590878181_256x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
.ends

.subckt nmos_5p04310590878179_256x8m81 D a_2016_n44# a_0_n44# a_896_n44# a_672_n44#
+ S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X5 S a_2016_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X6 S a_1120_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X7 D a_1344_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X8 S a_1568_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X9 D a_1792_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
.ends

.subckt wen_v2_256x8m81 wen GWE IGWEN clk vss vdd
Xnmos_5p0431059087818_256x8m81_0 vss pmos_5p04310590878183_256x8m81_0/D nmos_5p0431059087818_256x8m81_1/D
+ vss nmos_5p0431059087818_256x8m81
Xnmos_5p04310590878185_256x8m81_0 pmos_5p04310590878183_256x8m81_0/D nmos_5p0431059087818_256x8m81_1/S
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S vss nmos_5p0431059087818_256x8m81_1/S
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S
+ vss nmos_5p04310590878185_256x8m81
Xpmos_5p04310590878186_256x8m81_0 vdd pmos_5p04310590878186_256x8m81_0/D wen wen wen
+ vdd wen wen wen pmos_5p04310590878186_256x8m81
Xnmos_1p2$$202595372_256x8m81_0 vss pmos_5p04310590878141_256x8m81_1/S pmos_5p04310590878114_256x8m81_2/S
+ vss nmos_1p2$$202595372_256x8m81
Xnmos_5p0431059087818_256x8m81_1 nmos_5p0431059087818_256x8m81_1/D nmos_5p0431059087818_256x8m81_3/D
+ nmos_5p0431059087818_256x8m81_1/S vss nmos_5p0431059087818_256x8m81
Xnmos_1p2$$202595372_256x8m81_1 pmos_5p04310590878141_256x8m81_1/D nmos_5p0431059087818_256x8m81_4/D
+ pmos_5p04310590878141_256x8m81_1/S vss nmos_1p2$$202595372_256x8m81
Xnmos_5p0431059087818_256x8m81_2 vss wen nmos_5p0431059087818_256x8m81_2/S vss nmos_5p0431059087818_256x8m81
Xnmos_5p0431059087818_256x8m81_3 nmos_5p0431059087818_256x8m81_3/D clk vss vss nmos_5p0431059087818_256x8m81
Xnmos_5p0431059087818_256x8m81_4 nmos_5p0431059087818_256x8m81_4/D nmos_5p0431059087818_256x8m81_3/D
+ vss vss nmos_5p0431059087818_256x8m81
Xpmos_5p04310590878184_256x8m81_0 vdd pmos_5p04310590878184_256x8m81_0/D pmos_5p04310590878114_256x8m81_2/S
+ vdd pmos_5p04310590878114_256x8m81_2/S pmos_5p04310590878184_256x8m81
Xnmos_1p2$$202596396_256x8m81_0 vss pmos_5p04310590878114_256x8m81_2/S pmos_5p04310590878141_256x8m81_1/D
+ vss nmos_1p2$$202596396_256x8m81
Xnmos_5p04310590878182_256x8m81_0 pmos_5p04310590878186_256x8m81_0/D wen vss wen wen
+ vss nmos_5p04310590878182_256x8m81
Xpmos_5p04310590878183_256x8m81_0 vdd pmos_5p04310590878183_256x8m81_0/D nmos_5p0431059087818_256x8m81_1/S
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S vdd nmos_5p0431059087818_256x8m81_1/S
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_1/S
+ pmos_5p04310590878183_256x8m81
Xpmos_5p04310590878114_256x8m81_0 vdd vdd pmos_5p04310590878183_256x8m81_0/D nmos_5p0431059087818_256x8m81_1/D
+ pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_1 vdd nmos_5p0431059087818_256x8m81_3/D clk vdd pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_2 vdd vdd pmos_5p04310590878141_256x8m81_1/S pmos_5p04310590878114_256x8m81_2/S
+ pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_3 vdd vdd wen nmos_5p0431059087818_256x8m81_2/S pmos_5p04310590878114_256x8m81
Xpmos_5p04310590878114_256x8m81_4 vdd nmos_5p0431059087818_256x8m81_4/D nmos_5p0431059087818_256x8m81_3/D
+ vdd pmos_5p04310590878114_256x8m81
Xnmos_5p04310590878180_256x8m81_0 pmos_5p04310590878184_256x8m81_0/D pmos_5p04310590878114_256x8m81_2/S
+ vss pmos_5p04310590878114_256x8m81_2/S vss nmos_5p04310590878180_256x8m81
Xpmos_5p04310590878181_256x8m81_0 vdd GWE pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D vdd pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878181_256x8m81
Xpmos_5p04310590878181_256x8m81_1 vdd IGWEN pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D vdd pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878181_256x8m81
Xpmos_5p04310590878141_256x8m81_0 vdd nmos_5p0431059087818_256x8m81_1/D nmos_5p0431059087818_256x8m81_4/D
+ nmos_5p0431059087818_256x8m81_1/S pmos_5p04310590878141_256x8m81
Xpmos_5p04310590878141_256x8m81_1 vdd pmos_5p04310590878141_256x8m81_1/D nmos_5p0431059087818_256x8m81_3/D
+ pmos_5p04310590878141_256x8m81_1/S pmos_5p04310590878141_256x8m81
Xnmos_5p04310590878110_256x8m81_0 pmos_5p04310590878141_256x8m81_1/S nmos_5p0431059087818_256x8m81_3/D
+ nmos_5p0431059087818_256x8m81_2/S vss nmos_5p04310590878110_256x8m81
Xpmos_1p2$$202586156_256x8m81_0 vdd pmos_5p04310590878141_256x8m81_1/D vdd pmos_5p04310590878114_256x8m81_2/S
+ pmos_1p2$$202586156_256x8m81
Xnmos_5p04310590878179_256x8m81_0 GWE pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D vss pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D
+ pmos_5p04310590878183_256x8m81_0/D pmos_5p04310590878183_256x8m81_0/D vss nmos_5p04310590878179_256x8m81
Xnmos_5p04310590878179_256x8m81_1 IGWEN pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D vss pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D
+ pmos_5p04310590878186_256x8m81_0/D pmos_5p04310590878186_256x8m81_0/D vss nmos_5p04310590878179_256x8m81
Xpmos_5p04310590878120_256x8m81_0 vdd pmos_5p04310590878184_256x8m81_0/D nmos_5p0431059087818_256x8m81_3/D
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_3/D pmos_5p04310590878120_256x8m81
Xpmos_1p2$$202587180_256x8m81_0 pmos_5p04310590878141_256x8m81_1/S nmos_5p0431059087818_256x8m81_2/S
+ vdd nmos_5p0431059087818_256x8m81_4/D pmos_1p2$$202587180_256x8m81
Xnmos_5p04310590878139_256x8m81_0 pmos_5p04310590878184_256x8m81_0/D nmos_5p0431059087818_256x8m81_4/D
+ nmos_5p0431059087818_256x8m81_1/S nmos_5p0431059087818_256x8m81_4/D vss nmos_5p04310590878139_256x8m81
.ends

.subckt pmos_5p04310590878192_256x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
.ends

.subckt pmos_1p2$$47330348_256x8m81 pmos_5p04310590878141_256x8m81_0/S a_n31_n73#
+ w_n286_n141# pmos_5p04310590878141_256x8m81_0/D
Xpmos_5p04310590878141_256x8m81_0 w_n286_n141# pmos_5p04310590878141_256x8m81_0/D
+ a_n31_n73# pmos_5p04310590878141_256x8m81_0/S pmos_5p04310590878141_256x8m81
.ends

.subckt nmos_1p2$$48629804_256x8m81 a_193_n73# nmos_5p04310590878139_256x8m81_0/D
+ a_n31_n73# nmos_5p04310590878139_256x8m81_0/S VSUBS
Xnmos_5p04310590878139_256x8m81_0 nmos_5p04310590878139_256x8m81_0/D a_n31_n73# nmos_5p04310590878139_256x8m81_0/S
+ a_193_n73# VSUBS nmos_5p04310590878139_256x8m81
.ends

.subckt nmos_5p04310590878190_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.02u l=0.6u
.ends

.subckt nmos_1p2$$48302124_256x8m81 a_n31_n74# nmos_5p04310590878190_256x8m81_0/D
+ nmos_5p04310590878190_256x8m81_0/S VSUBS
Xnmos_5p04310590878190_256x8m81_0 nmos_5p04310590878190_256x8m81_0/D a_n31_n74# nmos_5p04310590878190_256x8m81_0/S
+ VSUBS nmos_5p04310590878190_256x8m81
.ends

.subckt nmos_5p04310590878189_256x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
.ends

.subckt nmos_1p2$$48306220_256x8m81 nmos_5p04310590878189_256x8m81_0/D a_n31_n74#
+ nmos_5p04310590878189_256x8m81_0/S a_865_n74# a_641_n74# a_417_n74# VSUBS a_193_n74#
Xnmos_5p04310590878189_256x8m81_0 nmos_5p04310590878189_256x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590878189_256x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310590878189_256x8m81
.ends

.subckt nmos_5p04310590878197_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1.2u
.ends

.subckt pmos_5p04310590878198_256x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.89u l=0.6u
.ends

.subckt pmos_5p04310590878177_256x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.77u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.77u l=0.6u
.ends

.subckt pmos_1p2$$48623660_256x8m81 pmos_5p04310590878177_256x8m81_0/S a_193_n74#
+ w_n286_n142# pmos_5p04310590878177_256x8m81_0/D a_n31_n74#
Xpmos_5p04310590878177_256x8m81_0 w_n286_n142# pmos_5p04310590878177_256x8m81_0/D
+ a_n31_n74# pmos_5p04310590878177_256x8m81_0/S a_193_n74# pmos_5p04310590878177_256x8m81
.ends

.subckt nmos_5p04310590878187_256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.75u l=0.6u
.ends

.subckt gen_512x8_256x8m81 WEN GWE tblhl IGWEN cen clk pmos_5p04310590878192_256x8m81_0/D
+ men VSS VDD
Xnmos_1p2$$47342636_256x8m81_0 VSS men nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D
+ VSS nmos_1p2$$47342636_256x8m81
Xpmos_5p04310590878178_256x8m81_1 VDD pmos_5p04310590878178_256x8m81_1/D pmos_5p04310590878178_256x8m81_0/D
+ VDD pmos_5p04310590878178_256x8m81
Xnmos_1p2$$47342636_256x8m81_1 nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D
+ clk VSS VSS nmos_1p2$$47342636_256x8m81
Xpmos_5p04310590878196_256x8m81_0 VDD pmos_5p04310590878196_256x8m81_0/D pmos_5p04310590878178_256x8m81_1/D
+ VDD pmos_5p04310590878196_256x8m81
Xpmos_1p2$$48624684_256x8m81_0 VDD VDD pmos_5p04310590878151_256x8m81_0/D pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S
+ pmos_1p2$$48624684_256x8m81
Xnmos_1p2$$48308268_256x8m81_0 pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D men pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ VSS pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D VSS pmos_5p04310590878192_256x8m81_0/D
+ nmos_1p2$$48308268_256x8m81
Xpmos_1p2$$48624684_256x8m81_1 VDD VDD pmos_1p2$$48623660_256x8m81_0/pmos_5p04310590878177_256x8m81_0/D
+ pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S pmos_1p2$$48624684_256x8m81
Xnmos_5p04310590878194_256x8m81_0 pmos_5p04310590878196_256x8m81_0/D pmos_5p04310590878178_256x8m81_1/D
+ VSS VSS nmos_5p04310590878194_256x8m81
Xpmos_1p2$$48624684_256x8m81_2 pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S
+ VDD clk VDD pmos_1p2$$48624684_256x8m81
Xpmos_1p2$$47815724_256x8m81_0 pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S
+ VDD VDD tblhl pmos_1p2$$47815724_256x8m81
Xpmos_5p04310590878193_256x8m81_0 pmos_5p04310590878192_256x8m81_0/D VDD men pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D VDD pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D pmos_5p04310590878192_256x8m81_0/D
+ pmos_5p04310590878193_256x8m81
Xwen_v2_256x8m81_0 wen_v2_256x8m81_0/wen wen_v2_256x8m81_0/GWE wen_v2_256x8m81_0/IGWEN
+ clk VSS VDD wen_v2_256x8m81
Xpmos_1p2$$47815724_256x8m81_1 VDD pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S
+ VDD pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xpmos_1p2$$47815724_256x8m81_2 VDD pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S
+ VDD tblhl pmos_1p2$$47815724_256x8m81
Xpmos_1p2$$47815724_256x8m81_3 pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S
+ VDD VDD pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xpmos_5p04310590878192_256x8m81_0 VDD pmos_5p04310590878192_256x8m81_0/D pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S VDD pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_5p04310590878192_256x8m81
Xpmos_1p2$$47815724_256x8m81_4 VDD pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ VDD pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xpmos_1p2$$47815724_256x8m81_5 VDD pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ VDD pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xpmos_1p2$$47330348_256x8m81_0 nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D VDD pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ pmos_1p2$$47330348_256x8m81
Xpmos_1p2$$47815724_256x8m81_6 pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ VDD VDD pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xnmos_1p2$$48629804_256x8m81_0 nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ pmos_5p04310590878151_256x8m81_0/D nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ VSS VSS nmos_1p2$$48629804_256x8m81
Xpmos_1p2$$47815724_256x8m81_7 pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ VDD VDD pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S pmos_1p2$$47815724_256x8m81
Xnmos_1p2$$48302124_256x8m81_0 pmos_5p04310590878198_256x8m81_0/D pmos_1p2$$48623660_256x8m81_0/pmos_5p04310590878177_256x8m81_0/D
+ VSS VSS nmos_1p2$$48302124_256x8m81
Xpmos_5p04310590878151_256x8m81_0 VDD pmos_5p04310590878151_256x8m81_0/D nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ VDD nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S pmos_5p04310590878151_256x8m81
Xpmos_1p2$$46285868_256x8m81_0 nmos_1p2$$46563372_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ VDD VDD nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D pmos_1p2$$46285868_256x8m81
Xnmos_1p2$$48306220_256x8m81_0 pmos_5p04310590878192_256x8m81_0/D pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ VSS pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S VSS pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S
+ nmos_1p2$$48306220_256x8m81
Xnmos_1p2$$46563372_256x8m81_0 nmos_1p2$$46563372_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D
+ nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D VSS VSS nmos_1p2$$46563372_256x8m81
Xpmos_1p2$$46285868_256x8m81_1 cen nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ VDD nmos_1p2$$46563372_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D pmos_1p2$$46285868_256x8m81
Xnmos_1p2$$46563372_256x8m81_1 pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ nmos_1p2$$46563372_256x8m81_0/nmos_5p0431059087818_256x8m81_0/D nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S
+ VSS nmos_1p2$$46563372_256x8m81
Xnmos_1p2$$46563372_256x8m81_2 VSS pmos_5p04310590878151_256x8m81_0/D pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ VSS nmos_1p2$$46563372_256x8m81
Xpmos_1p2$$46273580_256x8m81_0 VDD pmos_5p04310590878151_256x8m81_0/D pmos_1p2$$46273580_256x8m81_0/pmos_5p0431059087813_256x8m81_0/D
+ VDD pmos_5p04310590878151_256x8m81_0/D pmos_1p2$$46273580_256x8m81
Xnmos_1p2$$46551084_256x8m81_0 cen nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D
+ nmos_1p2$$46563372_256x8m81_1/nmos_5p0431059087818_256x8m81_0/S VSS nmos_1p2$$46551084_256x8m81
Xnmos_5p04310590878197_256x8m81_0 pmos_5p04310590878178_256x8m81_0/D clk VSS VSS nmos_5p04310590878197_256x8m81
Xpmos_5p04310590878198_256x8m81_0 VDD pmos_5p04310590878198_256x8m81_0/D pmos_5p04310590878196_256x8m81_0/D
+ VDD pmos_5p04310590878198_256x8m81
Xpmos_1p2$$48623660_256x8m81_0 VDD pmos_5p04310590878198_256x8m81_0/D VDD pmos_1p2$$48623660_256x8m81_0/pmos_5p04310590878177_256x8m81_0/D
+ pmos_5p04310590878198_256x8m81_0/D pmos_1p2$$48623660_256x8m81
Xnmos_5p04310590878187_256x8m81_0 pmos_5p04310590878198_256x8m81_0/D pmos_5p04310590878196_256x8m81_0/D
+ VSS VSS nmos_5p04310590878187_256x8m81
Xnmos_5p04310590878197_256x8m81_1 pmos_5p04310590878178_256x8m81_1/D pmos_5p04310590878178_256x8m81_0/D
+ VSS VSS nmos_5p04310590878197_256x8m81
Xpmos_5p04310590878178_256x8m81_0 VDD pmos_5p04310590878178_256x8m81_0/D clk VDD pmos_5p04310590878178_256x8m81
X0 VSS pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S a_11293_484# VSS nmos_6p0 w=18.145u l=0.6u
X1 a_9646_262# pmos_1p2$$48623660_256x8m81_0/pmos_5p04310590878177_256x8m81_0/D VSS VSS nmos_6p0 w=22.68u l=0.6u
X2 pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S a_10845_484# VSS nmos_6p0 w=18.145u l=0.6u
X3 a_12578_3205# tblhl pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S VSS nmos_6p0 w=4.54u l=0.6u
X4 pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S pmos_5p04310590878151_256x8m81_0/D a_9870_262# VSS nmos_6p0 w=22.68u l=0.6u
X5 a_11293_484# pmos_1p2$$48624684_256x8m81_2/pmos_5p04310590878195_256x8m81_0/S pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S VSS nmos_6p0 w=18.145u l=0.6u
X6 a_12130_3205# pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S VSS VSS nmos_6p0 w=4.54u l=0.6u
X7 a_10845_484# pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S VSS VSS nmos_6p0 w=18.145u l=0.6u
X8 pmos_1p2$$47815724_256x8m81_3/pmos_5p04310590878191_256x8m81_0/S tblhl a_12130_3205# VSS nmos_6p0 w=4.54u l=0.6u
X9 nmos_1p2$$47342636_256x8m81_1/nmos_5p04310590878157_256x8m81_0/D clk a_5174_6131# VDD pmos_6p0 w=2.28u l=0.595u
X10 VSS pmos_1p2$$47815724_256x8m81_7/pmos_5p04310590878191_256x8m81_0/S a_12578_3205# VSS nmos_6p0 w=4.54u l=0.6u
X11 a_9870_262# clk a_9646_262# VSS nmos_6p0 w=22.68u l=0.6u
X12 a_5174_6131# men VDD VDD pmos_6p0 w=2.28u l=0.595u
.ends

.subckt control_512x8_256x8m81 GWE GWEN VSS VDD RYS[7] RYS[6] RYS[5] RYS[4] RYS[3]
+ RYS[2] RYS[1] RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl
+ IGWEN xb[3] xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xb[1] xc[3] xc[1] xc[2]
+ xc[0] xa[0] xa[1] A[9] A[7] CLK A[2] A[6] A[3] A[4] A[5] A[8] ypredec1_256x8m81_0/ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd
+ ypredec1_256x8m81_0/ly[2] gen_512x8_256x8m81_0/tblhl A[0] CEN men A[1] prexdec_top_256x8m81_0/xpredec1_256x8m81_0/vdd
+ VSUBS gen_512x8_256x8m81_0/VDD
Xypredec1_256x8m81_0 ypredec1_256x8m81_0/ly[5] ypredec1_256x8m81_0/ly[4] ypredec1_256x8m81_0/ly[7]
+ ypredec1_256x8m81_0/ly[3] ypredec1_256x8m81_0/ly[2] ypredec1_256x8m81_0/ly[1] ypredec1_256x8m81_0/ly[0]
+ RYS[0] RYS[1] RYS[2] RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_256x8m81_0/ly[6]
+ men A[0] A[1] A[2] CLK ypredec1_256x8m81_0/ypredec1_bot_256x8m81_2/alatch_256x8m81_0/vdd
+ gen_512x8_256x8m81_0/VDD gen_512x8_256x8m81_0/VDD gen_512x8_256x8m81_0/VDD VSUBS
+ gen_512x8_256x8m81_0/VDD ypredec1_256x8m81
Xprexdec_top_256x8m81_0 CLK A[5] A[9] A[7] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1] xb[2]
+ xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] prexdec_top_256x8m81_0/xpredec1_256x8m81_0/vdd
+ VSUBS VSUBS VSUBS VSUBS xc[0] prexdec_top_256x8m81_0/xpredec1_256x8m81_0/vdd men
+ prexdec_top_256x8m81_0/xpredec1_256x8m81_0/vdd VSUBS prexdec_top_256x8m81
Xgen_512x8_256x8m81_0 GWEN GWE gen_512x8_256x8m81_0/tblhl IGWEN CEN CLK gen_512x8_256x8m81_0/pmos_5p04310590878192_256x8m81_0/D
+ men VSUBS gen_512x8_256x8m81_0/VDD gen_512x8_256x8m81
.ends

.subckt x018SRAM_cell1_cutPC_256x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt new_dummyrow_unit_256x8m81 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50# 018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
X018SRAM_cell1_dummy_256x8m81_0 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_1 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_2 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_3 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_4 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_5 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_10 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_6 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_7 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_11 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_8 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_12 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_9 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_13 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_14 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_15 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
.ends

.subckt new_dummyrow_unit_01_256x8m81 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50#
+ VSUBS 018SRAM_strap1_256x8m81_1/w_n68_622# 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
X018SRAM_cell1_dummy_256x8m81_0 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_1 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_2 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_3 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_4 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_5 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_10 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_6 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_7 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_11 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_8 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_12 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_9 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_13 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_14 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_15 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_strap1_256x8m81_1/w_n68_622#
+ 018SRAM_strap1_256x8m81_1/a_n36_52# 018SRAM_strap1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
.ends

.subckt ldummy_256x4_256x8m81 018SRAM_cell1_cutPC_256x8m81_30/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_16/a_246_342#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_31/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_5/w_n68_622#
+ 018SRAM_cell1_cutPC_256x8m81_29/a_246_712# 018SRAM_cell1_dummy_256x8m81_22/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_16/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_26/a_246_342# 018SRAM_cell1_cutPC_256x8m81_26/w_n68_622#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_17/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_18/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_19/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_6/a_246_342#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_9/a_246_712# 018SRAM_cell1_cutPC_256x8m81_4/w_n68_622#
+ 018SRAM_cell1_cutPC_256x8m81_17/a_246_342# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_23/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_27/a_246_342# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_7/a_246_342# 018SRAM_cell1_cutPC_256x8m81_18/a_246_342#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_20/m3_n36_330#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_7/a_246_712# 018SRAM_cell1_cutPC_256x8m81_27/a_246_712#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_28/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_21/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_24/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_23/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_28/a_246_712#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_22/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_23/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_8/a_246_342# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_19/a_246_342# 018SRAM_cell1_cutPC_256x8m81_24/m3_n36_330#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_8/w_n68_622# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_25/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_29/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_25/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_24/w_n68_622# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_26/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_27/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_2/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_9/a_246_342#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_28/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_16/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_3/m3_n36_330#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_4/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_10/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_26/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_29/m3_n36_330# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_11/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_5/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_12/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_6/m3_n36_330# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_10/a_246_342# 018SRAM_cell1_cutPC_256x8m81_13/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_17/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_7/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_29/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_30/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_20/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_27/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_14/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_8/m3_n36_330#
+ 018SRAM_cell1_cutPC_256x8m81_25/a_246_712# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_31/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_30/a_246_342# 018SRAM_cell1_cutPC_256x8m81_15/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_31/a_246_712#
+ 018SRAM_cell1_cutPC_256x8m81_9/m3_n36_330# 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_16/m3_n36_330#
+ 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_18/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_17/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_9/w_n68_622#
+ 018SRAM_cell1_cutPC_256x8m81_1/a_246_712# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_11/a_246_342# 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_5/a_246_712#
+ 018SRAM_cell1_dummy_256x8m81_28/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_18/m3_n36_330#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_21/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_26/a_246_712#
+ 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_19/m3_n36_330# 018SRAM_cell1_cutPC_256x8m81_31/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_7/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_1/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_19/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_27/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_12/a_246_342#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_4/a_246_712#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_22/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_29/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_28/w_n68_622# 018SRAM_cell1_dummy_256x8m81_20/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_21/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_2/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_22/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_13/a_246_342# 018SRAM_cell1_cutPC_256x8m81_13/a_246_712#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_23/m2_390_n50#
+ 018SRAM_cell1_cutPC_256x8m81_23/a_246_342# 018SRAM_cell1_cutPC_256x8m81_23/a_246_712#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_24/m2_390_n50#
+ VSS new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_25/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_3/a_246_342#
+ 018SRAM_cell1_dummy_256x8m81_26/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_14/a_246_342#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_8/a_246_712#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_27/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_20/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_24/a_246_342# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_24/a_246_712#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_28/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_256x8m81_30/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_29/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_4/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_15/a_246_342# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_13/w_n68_622# 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ 018SRAM_cell1_cutPC_256x8m81_25/a_246_342# 018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_dummy_256x8m81_21/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_cell1_cutPC_256x8m81_25/w_n68_622#
+ 018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_256x8m81_31/m2_90_n50# 018SRAM_cell1_cutPC_256x8m81_31/w_n68_622#
+ 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50# VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
X018SRAM_cell1_cutPC_256x8m81_23 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_23/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_23/a_246_712# 018SRAM_cell1_cutPC_256x8m81_23/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_23/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_12 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_12/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_4/a_246_712# 018SRAM_cell1_cutPC_256x8m81_12/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_24 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_24/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_24/a_246_712# 018SRAM_cell1_cutPC_256x8m81_24/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_24/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_13 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_13/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_13/a_246_712# 018SRAM_cell1_cutPC_256x8m81_13/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_13/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_25 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_25/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_25/a_246_712# 018SRAM_cell1_cutPC_256x8m81_25/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_25/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_14 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_14/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_8/a_246_712# 018SRAM_cell1_cutPC_256x8m81_14/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_8/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_26 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_26/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_26/a_246_712# 018SRAM_cell1_cutPC_256x8m81_26/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_26/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_15 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_15/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_23/a_246_712# 018SRAM_cell1_cutPC_256x8m81_15/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_23/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_27 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_27/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_27/a_246_712# 018SRAM_cell1_cutPC_256x8m81_27/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_27/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_16 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_16/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_29/a_246_712# 018SRAM_cell1_cutPC_256x8m81_16/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_29/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_28 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_28/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_28/a_246_712# 018SRAM_cell1_cutPC_256x8m81_28/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_28/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_17 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_17/a_246_342#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_17/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_29 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_29/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_29/a_246_712# 018SRAM_cell1_cutPC_256x8m81_29/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_29/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_18 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_18/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_27/a_246_712# 018SRAM_cell1_cutPC_256x8m81_18/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_27/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_19 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_19/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_28/a_246_712# 018SRAM_cell1_cutPC_256x8m81_19/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_28/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_dummy_256x8m81_0 VSUBS 018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_0/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_1 VSUBS 018SRAM_cell1_dummy_256x8m81_1/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_2 VSUBS 018SRAM_cell1_dummy_256x8m81_2/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
Xnew_dummyrow_unit_256x8m81_0 new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# VSUBS new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_90_n50#
+ 018SRAM_cell1_256x8m81_1/w_n68_622# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# VSUBS new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
+ new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# new_dummyrow_unit_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ new_dummyrow_unit_256x8m81
X018SRAM_cell1_dummy_256x8m81_3 VSUBS 018SRAM_cell1_dummy_256x8m81_3/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_30 VSUBS 018SRAM_cell1_dummy_256x8m81_30/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_30/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_4 VSUBS 018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_31 VSUBS 018SRAM_cell1_dummy_256x8m81_31/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_31/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_20 VSUBS 018SRAM_cell1_dummy_256x8m81_20/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_20/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_5 VSUBS 018SRAM_cell1_dummy_256x8m81_5/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_5/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_10 VSUBS 018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_10/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_21 VSUBS 018SRAM_cell1_dummy_256x8m81_21/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_21/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_6 VSUBS 018SRAM_cell1_dummy_256x8m81_6/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_6/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_11 VSUBS 018SRAM_cell1_dummy_256x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_11/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_22 VSUBS 018SRAM_cell1_dummy_256x8m81_22/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_22/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_7 VSUBS 018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_12 VSUBS 018SRAM_cell1_dummy_256x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_23 VSUBS 018SRAM_cell1_dummy_256x8m81_23/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_23/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_8 VSUBS 018SRAM_cell1_dummy_256x8m81_8/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_8/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_13 VSUBS 018SRAM_cell1_dummy_256x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_24 VSUBS 018SRAM_cell1_dummy_256x8m81_24/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_24/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_9 VSUBS 018SRAM_cell1_dummy_256x8m81_9/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_0 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_0/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_1/a_246_712# 018SRAM_cell1_cutPC_256x8m81_0/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_dummy_256x8m81_14 VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_14/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_25 VSUBS 018SRAM_cell1_dummy_256x8m81_25/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_25/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_1 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_1/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_1/a_246_712# 018SRAM_cell1_cutPC_256x8m81_1/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_256x8m81_0 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS
+ x018SRAM_cell1_256x8m81
X018SRAM_cell1_dummy_256x8m81_15 VSUBS 018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_15/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_26 VSUBS 018SRAM_cell1_dummy_256x8m81_26/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_26/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_2 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_2/a_246_342#
+ 018SRAM_cell1_256x8m81_0/w_n68_622# 018SRAM_cell1_cutPC_256x8m81_2/m3_n36_330# 018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_256x8m81_1 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_256x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_256x8m81
X018SRAM_cell1_dummy_256x8m81_16 VSUBS 018SRAM_cell1_dummy_256x8m81_16/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_16/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_27 VSUBS 018SRAM_cell1_dummy_256x8m81_27/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_27/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_3 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_3/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_7/a_246_712# 018SRAM_cell1_cutPC_256x8m81_3/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_7/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_dummy_256x8m81_17 VSUBS 018SRAM_cell1_dummy_256x8m81_17/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_17/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_28 VSUBS 018SRAM_cell1_dummy_256x8m81_28/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_28/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_4 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_4/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_4/a_246_712# 018SRAM_cell1_cutPC_256x8m81_4/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_dummy_256x8m81_18 VSUBS 018SRAM_cell1_dummy_256x8m81_18/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_18/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_dummy_256x8m81_29 VSUBS 018SRAM_cell1_dummy_256x8m81_29/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_29/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_5 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_5/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_5/a_246_712# 018SRAM_cell1_cutPC_256x8m81_5/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_dummy_256x8m81_19 VSUBS 018SRAM_cell1_dummy_256x8m81_19/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_256x8m81_19/m2_390_n50# 018SRAM_cell1_256x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_256x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_256x8m81
X018SRAM_cell1_cutPC_256x8m81_6 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_6/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_9/a_246_712# 018SRAM_cell1_cutPC_256x8m81_6/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_9/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_7 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_7/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_7/a_246_712# 018SRAM_cell1_cutPC_256x8m81_7/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_7/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_8 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_8/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_8/a_246_712# 018SRAM_cell1_cutPC_256x8m81_8/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_8/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
Xnew_dummyrow_unit_01_256x8m81_0 new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_15/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_1/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_0/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_2/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_3/m2_390_n50# VSUBS
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_4/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_9/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_5/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_6/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_7/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_10/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_90_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_11/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_12/m2_390_n50# VSUBS
+ 018SRAM_cell1_256x8m81_1/w_n68_622# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_8/m2_90_n50#
+ new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_13/m2_390_n50# new_dummyrow_unit_01_256x8m81_0/018SRAM_cell1_dummy_256x8m81_14/m2_390_n50#
+ new_dummyrow_unit_01_256x8m81
X018SRAM_cell1_cutPC_256x8m81_9 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_9/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_9/a_246_712# 018SRAM_cell1_cutPC_256x8m81_9/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_9/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_30 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_30/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_31/a_246_712# 018SRAM_cell1_cutPC_256x8m81_30/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_31/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_31 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_31/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_31/a_246_712# 018SRAM_cell1_cutPC_256x8m81_31/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_31/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_20 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_20/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_25/a_246_712# 018SRAM_cell1_cutPC_256x8m81_20/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_25/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_21 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_21/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_26/a_246_712# 018SRAM_cell1_cutPC_256x8m81_21/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_26/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_10 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_10/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_13/a_246_712# 018SRAM_cell1_cutPC_256x8m81_10/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_13/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_22 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_22/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_24/a_246_712# 018SRAM_cell1_cutPC_256x8m81_22/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_24/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
X018SRAM_cell1_cutPC_256x8m81_11 VSUBS 018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_256x8m81_11/a_246_342#
+ 018SRAM_cell1_cutPC_256x8m81_5/a_246_712# 018SRAM_cell1_cutPC_256x8m81_11/m3_n36_330#
+ 018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_256x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_256x8m81
.ends

.subckt Cell_array8x8x4_256x8m81 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622# 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42#
+ VSUBS
X018SRAM_cell1_2x_256x8m81_378 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_301 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_389 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_323 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_334 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_312 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_356 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_367 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_345 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_120 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_131 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_153 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_142 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_197 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_175 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_164 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_186 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_40 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_84 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_95 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_51 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_73 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_62 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_505 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_379 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_368 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_302 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_324 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_335 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_313 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_357 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_346 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_121 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_132 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_154 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_143 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_198 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_110 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_165 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_176 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_187 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_41 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_30 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_85 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_96 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_74 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_63 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_52 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_506 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_369 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_303 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_325 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_314 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_358 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_336 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_347 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_122 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_133 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_144 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_155 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_199 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_100 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_111 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_166 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_177 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_188 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_31 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_42 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_20 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_86 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_97 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_75 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_53 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_64 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_507 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_326 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_315 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_304 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_337 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_359 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_348 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_156 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_123 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_134 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_112 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_145 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_101 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_178 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_189 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_167 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_10 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_32 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_21 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_43 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_87 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_98 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_76 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_54 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_65 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_508 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_327 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_316 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_305 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_338 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_349 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_157 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_135 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_124 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_113 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_146 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_102 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_179 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_168 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_11 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_44 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_33 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_22 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_99 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_88 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_55 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_66 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_77 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_509 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_328 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_317 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_306 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_339 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_114 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_158 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_136 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_125 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_147 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_103 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_169 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_23 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_12 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_45 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_34 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_89 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_56 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_67 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_78 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_329 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_318 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_307 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_115 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_137 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_159 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_126 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_148 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_104 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_490 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_13 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_24 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_46 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_35 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_57 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_68 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_79 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_319 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_308 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_116 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_149 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_138 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_127 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_105 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_480 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_491 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_36 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_14 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_25 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_47 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_58 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_69 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_309 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_117 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_128 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_139 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_106 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_481 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_470 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_492 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_26 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_37 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_15 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_48 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_59 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_118 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_129 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_107 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_482 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_471 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_493 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_460 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_290 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_27 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_38 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_16 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_49 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_119 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_108 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_483 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_450 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_494 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_461 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_472 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_280 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_291 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_28 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_39 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_17 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_109 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_440 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_484 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_451 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_495 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_462 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_473 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_281 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_270 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_292 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_29 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_18 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_441 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_430 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_485 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_452 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_496 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_463 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_474 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_282 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_271 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_293 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_260 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_19 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_36/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_442 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_431 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_420 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_486 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_453 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_497 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_464 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_475 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_283 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_272 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_261 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_294 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_250 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_410 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_443 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_432 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_421 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_487 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_454 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_498 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_465 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_476 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_262 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_251 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_240 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_284 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_273 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_295 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_400 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_411 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_444 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_433 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_422 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_455 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_499 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_466 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_488 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_477 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_285 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_274 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_263 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_296 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_230 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_252 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_241 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_401 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_412 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_445 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_434 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_423 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_467 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_489 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_456 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_478 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_297 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_286 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_264 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_275 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_220 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_253 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_242 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_231 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_402 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_413 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_446 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_424 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_435 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_468 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_457 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_479 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_298 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_287 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_265 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_276 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_221 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_210 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_254 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_243 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_232 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_403 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_414 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_447 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_425 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_436 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_469 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_458 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_299 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_288 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_266 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_277 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_211 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_200 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_222 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_255 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_244 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_233 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_404 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_415 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_426 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_437 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_448 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_459 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_267 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_278 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_256 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_212 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_201 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_223 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_245 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_234 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_289 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_405 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_427 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_438 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_416 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_449 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_268 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_279 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_257 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_213 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_202 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_224 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_235 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_246 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_406 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_439 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_428 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_417 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_269 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_258 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_214 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_203 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_225 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_236 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_247 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_407 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_429 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_418 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_259 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_0 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_215 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_204 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_248 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_226 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_463/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_237 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_408 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_419 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_227 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_1 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_216 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_205 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_249 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_238 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_409 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_228 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_2 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_217 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_206 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_239 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_229 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_3 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_218 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_207 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_390 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_4 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_219 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_208 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_380 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_391 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_5 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_209 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_462/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_392 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_381 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_370 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_6 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_6/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_371 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_360 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_393 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_382 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_190 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_7 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_394 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_383 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_372 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_361 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_350 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_191 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_180 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_8 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_510 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_395 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_373 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_384 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_340 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_362 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_351 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_192 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_170 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_181 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_9 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_90 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_500 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_511 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_396 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_374 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_385 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_330 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_341 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_2/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_363 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_352 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_193 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_160 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_171 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_182 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_80 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_91 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_501 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_397 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_375 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_386 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_320 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_331 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_342 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_3/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_364 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_353 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_150 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_489/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_194 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_161 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_490/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_172 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_183 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_81 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_92 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_92/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_70 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_7/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_502 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_376 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_387 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_321 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_332 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_310 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_343 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_365 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_354 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_398 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_4/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_151 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_140 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_488/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_195 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_456/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_162 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_173 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_184 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_460/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_82 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_93 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_93/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_60 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_71 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_8/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_503 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_503/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_399 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_377 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_407/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_89/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_300 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_399/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_459/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_388 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_415/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_322 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_458/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_333 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_447/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_493/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_311 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_438/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_344 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_363/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_366 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_355 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_367/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_130 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_152 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_5/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_494/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_141 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_491/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_196 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_457/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_163 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_492/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_174 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_495/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_185 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_79/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_461/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_83 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_99/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_91/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_94 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_94/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_50 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_90/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_61 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_95/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_72 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_76/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
X018SRAM_cell1_2x_256x8m81_504 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52# 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_256x8m81_511/018SRAM_cell1_256x8m81_0/a_n36_52# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_444_n42# 018SRAM_cell1_2x_256x8m81_9/018SRAM_cell1_256x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_2x_256x8m81_88/018SRAM_cell1_256x8m81_1/a_36_n42# VSUBS x018SRAM_cell1_2x_256x8m81
.ends

.subckt col_256a_256x8m81 pcb[0] pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1] WEN[0]
+ WL[3] ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] GWE WL[2] WL[1] WL[31] WL[30]
+ WL[29] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[12] WL[11] WL[10] WL[9] WL[8]
+ WL[7] WL[6] WL[5] WL[4] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[28] WL[27]
+ WL[26] WL[0] ypass[2] WL[25] b[13] b[16] b[25] din[1] din[3] din[2] din[0] q[0]
+ q[1] q[2] q[3] b[17] b[14] bb[10] bb[11] bb[12] bb[13] bb[14] bb[15] bb[16] bb[20]
+ bb[29] bb[30] bb[31] b[30] b[15] b[12] b[0] b[18] a_15501_29383# m3_n1102_31970#
+ b[3] a_15261_28608# bb[19] b[21] a_4701_29383# ypass[6] ypass[7] b[27] a_4461_28608#
+ a_15501_28608# bb[22] bb[5] b[6] bb[3] b[5] bb[23] bb[0] saout_m2_256x8m81_1/GWEN
+ bb[4] saout_R_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_256x8m81_4/b b[26] b[28]
+ b[8] a_15261_29383# b[10] b[2] bb[26] b[7] saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735#
+ b[1] bb[6] saout_R_m2_256x8m81_0/wen_wm1_256x8m81_0/wen b[20] bb[25] bb[27] bb[28]
+ b[11] a_4701_28608# bb[18] bb[9] b[31] saout_m2_256x8m81_1/sa_256x8m81_0/pcb bb[21]
+ bb[7] saout_m2_256x8m81_0/pcb bb[2] b[4] bb[1] saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb
+ bb[17] b[24] saout_m2_256x8m81_0/WEN b[23] bb[8] b[22] saout_R_m2_256x8m81_1/sa_256x8m81_0/pcb
+ a_4461_29383# VDD b[29] bb[24] b[19] b[9] VSS men
Xsaout_R_m2_256x8m81_0 saout_R_m2_256x8m81_0/pcb saout_R_m2_256x8m81_0/datain saout_R_m2_256x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWE saout_m2_256x8m81_1/GWEN
+ b[7] b[0] bb[5] saout_R_m2_256x8m81_0/q saout_R_m2_256x8m81_0/wen_wm1_256x8m81_0/wen
+ saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735# saout_R_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ b[2] b[6] bb[1] bb[3] b[5] bb[4] saout_R_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b
+ b[4] men a_15727_28608# a_15501_28608# bb[6] a_15727_29383# a_15501_29383# ypass[0]
+ ypass[7] VSS VSS bb[7] bb[0] ypass[1] saout_R_m2_256x8m81_0/sacntl_2_256x8m81_0/a_4718_983#
+ saout_m2_256x8m81_1/GWEN ypass[4] ypass[2] VDD saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb
+ bb[2] b[3] VDD ypass[5] ypass[6] VDD saout_R_m2_256x8m81_0/mux821_256x8m81_0/a_4992_424#
+ saout_R_m2_256x8m81_0/sa_256x8m81_0/wep VSS VDD b[1] ypass[3] saout_R_m2_256x8m81
Xsaout_R_m2_256x8m81_1 saout_R_m2_256x8m81_1/pcb saout_R_m2_256x8m81_1/datain saout_R_m2_256x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] GWE saout_m2_256x8m81_1/GWEN
+ b[23] b[16] bb[21] saout_R_m2_256x8m81_1/q saout_R_m2_256x8m81_1/wen_wm1_256x8m81_0/wen
+ saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735# saout_R_m2_256x8m81_1/mux821_256x8m81_0/ypass_gate_256x8m81_4/b
+ b[18] b[22] bb[17] bb[19] b[21] bb[20] saout_R_m2_256x8m81_1/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/b
+ b[20] men a_4927_28608# a_4701_28608# bb[22] a_4927_29383# a_4701_29383# ypass[0]
+ ypass[7] VSS saout_R_m2_256x8m81_1/outbuf_oe_256x8m81_0/a_4913_n316# bb[23] bb[16]
+ ypass[1] VSS saout_m2_256x8m81_1/GWEN ypass[4] ypass[2] VDD saout_R_m2_256x8m81_1/sa_256x8m81_0/pcb
+ bb[18] b[19] VDD ypass[5] ypass[6] VDD saout_R_m2_256x8m81_1/mux821_256x8m81_0/a_4992_424#
+ saout_R_m2_256x8m81_1/sa_256x8m81_0/wep VSS VDD b[17] ypass[3] saout_R_m2_256x8m81
Xsaout_m2_256x8m81_0 saout_m2_256x8m81_0/pcb saout_m2_256x8m81_0/datain saout_m2_256x8m81_0/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] saout_m2_256x8m81_1/GWEN
+ GWE bb[26] b[24] saout_m2_256x8m81_0/q a_4236_28608# a_4461_28608# a_4236_29383#
+ a_4461_29383# saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735# b[29] b[25] ypass[7]
+ bb[30] bb[28] b[26] saout_m2_256x8m81_0/mux821_256x8m81_0/ypass_gate_a_256x8m81_0/a_n80_n10#
+ bb[27] b[27] men bb[25] ypass[0] VSS VSS bb[24] bb[31] ypass[1] VSS saout_m2_256x8m81_1/GWEN
+ ypass[4] ypass[2] VDD b[31] bb[29] saout_m2_256x8m81_0/pcb b[28] VDD VDD ypass[5]
+ VDD ypass[6] saout_m2_256x8m81_0/sa_256x8m81_0/wep saout_m2_256x8m81_0/mux821_256x8m81_0/a_4992_424#
+ VSS b[30] ypass[3] saout_m2_256x8m81
Xsaout_m2_256x8m81_1 saout_m2_256x8m81_1/pcb saout_m2_256x8m81_1/datain saout_m2_256x8m81_1/WEN
+ ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] ypass[0] saout_m2_256x8m81_1/GWEN
+ GWE bb[10] b[8] saout_m2_256x8m81_1/q a_15036_28608# a_15261_28608# a_15036_29383#
+ a_15261_29383# saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735# b[13] b[9] ypass[7]
+ bb[14] bb[12] b[10] VSS bb[11] b[11] men bb[9] ypass[0] VSS VSS bb[8] bb[15] ypass[1]
+ VSS saout_m2_256x8m81_1/GWEN ypass[4] ypass[2] VDD b[15] bb[13] saout_m2_256x8m81_1/sa_256x8m81_0/pcb
+ b[12] VDD VDD ypass[5] VDD ypass[6] saout_m2_256x8m81_1/sa_256x8m81_0/wep VSS VSS
+ b[14] ypass[3] saout_m2_256x8m81
XCell_array8x8x4_256x8m81_0 b[18] bb[23] bb[15] bb[11] bb[20] b[2] bb[7] bb[4] b[20]
+ b[14] bb[28] b[11] b[10] b[21] bb[14] b[31] b[30] b[4] b[5] bb[13] bb[17] WL[2]
+ bb[29] b[22] bb[9] bb[24] b[9] bb[22] WL[22] bb[16] bb[12] WL[21] WL[13] bb[6] bb[0]
+ WL[4] b[28] b[6] b[8] bb[19] b[23] b[17] bb[30] WL[15] WL[3] WL[30] b[29] bb[31]
+ WL[23] b[15] b[7] b[1] bb[25] WL[6] WL[17] bb[27] bb[3] bb[18] b[16] bb[21] WL[5]
+ WL[18] b[27] bb[10] WL[29] WL[9] b[26] bb[8] WL[14] b[25] WL[24] bb[26] WL[20] WL[26]
+ bb[2] WL[25] b[3] WL[11] WL[31] b[12] b[13] WL[8] b[24] bb[1] WL[1] WL[7] WL[12]
+ WL[19] WL[10] WL[0] bb[5] WL[27] WL[28] VDD b[0] WL[16] b[19] VSS Cell_array8x8x4_256x8m81
.ends

.subckt lcol4_256_256x8m81 pcb[2] pcb[3] pcb[0] pcb[1] vdd WEN[3] WEN[2] WEN[1] WEN[0]
+ WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+ WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+ WL[0] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] men ypass[0] ypass[1] ypass[2] ypass[3]
+ ypass[4] ypass[5] ypass[6] ypass[7] GWEN GWE din[0] din[1] din[3] din[2] q[0] q[1]
+ q[2] q[3] col_256a_256x8m81_0/WL[7] col_256a_256x8m81_0/saout_m2_256x8m81_1/GWEN
+ ldummy_256x4_256x8m81_0/VSS col_256a_256x8m81_0/WL[8] col_256a_256x8m81_0/WL[9]
+ col_256a_256x8m81_0/a_15501_28608# col_256a_256x8m81_0/a_4461_29383# col_256a_256x8m81_0/WL[20]
+ col_256a_256x8m81_0/WL[21] col_256a_256x8m81_0/WL[22] col_256a_256x8m81_0/WL[23]
+ col_256a_256x8m81_0/a_15261_29383# col_256a_256x8m81_0/WL[24] col_256a_256x8m81_0/saout_R_m2_256x8m81_0/wen_wm1_256x8m81_0/wen
+ col_256a_256x8m81_0/WL[25] col_256a_256x8m81_0/WL[26] col_256a_256x8m81_0/WL[27]
+ col_256a_256x8m81_0/WL[28] col_256a_256x8m81_0/WL[29] col_256a_256x8m81_0/a_4701_29383#
+ col_256a_256x8m81_0/saout_m2_256x8m81_0/WEN col_256a_256x8m81_0/a_4461_28608# col_256a_256x8m81_0/WL[10]
+ col_256a_256x8m81_0/a_15501_29383# col_256a_256x8m81_0/men col_256a_256x8m81_0/WL[11]
+ col_256a_256x8m81_0/GWE col_256a_256x8m81_0/WL[12] col_256a_256x8m81_0/WL[13] col_256a_256x8m81_0/WL[30]
+ col_256a_256x8m81_0/saout_m2_256x8m81_0/pcb col_256a_256x8m81_0/ypass[0] col_256a_256x8m81_0/a_15261_28608#
+ col_256a_256x8m81_0/WL[14] col_256a_256x8m81_0/WL[31] col_256a_256x8m81_0/ypass[1]
+ col_256a_256x8m81_0/WL[0] col_256a_256x8m81_0/WL[15] col_256a_256x8m81_0/ypass[2]
+ col_256a_256x8m81_0/WL[1] col_256a_256x8m81_0/WL[16] col_256a_256x8m81_0/ypass[3]
+ col_256a_256x8m81_0/WL[2] col_256a_256x8m81_0/WL[17] col_256a_256x8m81_0/ypass[4]
+ col_256a_256x8m81_0/WL[3] col_256a_256x8m81_0/saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735#
+ col_256a_256x8m81_0/WL[18] col_256a_256x8m81_0/ypass[5] col_256a_256x8m81_0/WL[4]
+ col_256a_256x8m81_0/saout_R_m2_256x8m81_1/sa_256x8m81_0/pcb col_256a_256x8m81_0/WL[19]
+ col_256a_256x8m81_0/ypass[6] col_256a_256x8m81_0/WL[5] col_256a_256x8m81_0/saout_m2_256x8m81_1/sa_256x8m81_0/pcb
+ col_256a_256x8m81_0/saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb VDD col_256a_256x8m81_0/ypass[7]
+ col_256a_256x8m81_0/a_4701_28608# col_256a_256x8m81_0/WL[6] VSS
Xldummy_256x4_256x8m81_0 col_256a_256x8m81_0/WL[15] VSS col_256a_256x8m81_0/bb[26]
+ col_256a_256x8m81_0/bb[19] VDD VSS col_256a_256x8m81_0/bb[5] col_256a_256x8m81_0/WL[16]
+ col_256a_256x8m81_0/bb[13] VDD VDD col_256a_256x8m81_0/b[22] col_256a_256x8m81_0/b[27]
+ col_256a_256x8m81_0/b[28] VSS VDD col_256a_256x8m81_0/bb[11] col_256a_256x8m81_0/b[29]
+ col_256a_256x8m81_0/bb[28] col_256a_256x8m81_0/bb[9] col_256a_256x8m81_0/bb[30]
+ VSS col_256a_256x8m81_0/b[18] col_256a_256x8m81_0/b[12] VDD VDD VSS col_256a_256x8m81_0/bb[3]
+ col_256a_256x8m81_0/b[30] col_256a_256x8m81_0/b[20] VSS col_256a_256x8m81_0/bb[13]
+ VSS VSS col_256a_256x8m81_0/bb[17] col_256a_256x8m81_0/WL[25] col_256a_256x8m81_0/b[2]
+ col_256a_256x8m81_0/b[14] VDD VDD col_256a_256x8m81_0/bb[31] VSS col_256a_256x8m81_0/WL[23]
+ col_256a_256x8m81_0/bb[21] VDD VDD col_256a_256x8m81_0/b[12] col_256a_256x8m81_0/WL[21]
+ col_256a_256x8m81_0/bb[7] col_256a_256x8m81_0/WL[19] VSS col_256a_256x8m81_0/b[16]
+ VSS col_256a_256x8m81_0/WL[22] col_256a_256x8m81_0/bb[1] col_256a_256x8m81_0/b[26]
+ VDD col_256a_256x8m81_0/bb[23] col_256a_256x8m81_0/bb[19] VSS col_256a_256x8m81_0/WL[26]
+ col_256a_256x8m81_0/WL[3] VDD col_256a_256x8m81_0/b[14] col_256a_256x8m81_0/WL[24]
+ col_256a_256x8m81_0/WL[4] col_256a_256x8m81_0/b[6] col_256a_256x8m81_0/WL[28] col_256a_256x8m81_0/WL[0]
+ VSS col_256a_256x8m81_0/b[24] col_256a_256x8m81_0/WL[30] col_256a_256x8m81_0/bb[27]
+ col_256a_256x8m81_0/WL[14] col_256a_256x8m81_0/b[0] col_256a_256x8m81_0/WL[12] col_256a_256x8m81_0/WL[8]
+ col_256a_256x8m81_0/b[18] col_256a_256x8m81_0/WL[18] col_256a_256x8m81_0/bb[15]
+ col_256a_256x8m81_0/WL[9] col_256a_256x8m81_0/WL[10] col_256a_256x8m81_0/b[4] col_256a_256x8m81_0/WL[11]
+ col_256a_256x8m81_0/WL[5] col_256a_256x8m81_0/bb[25] VSS col_256a_256x8m81_0/WL[7]
+ col_256a_256x8m81_0/bb[29] col_256a_256x8m81_0/b[8] col_256a_256x8m81_0/WL[13] VDD
+ col_256a_256x8m81_0/b[25] VSS col_256a_256x8m81_0/b[7] col_256a_256x8m81_0/bb[17]
+ col_256a_256x8m81_0/WL[1] col_256a_256x8m81_0/WL[2] VDD col_256a_256x8m81_0/bb[7]
+ col_256a_256x8m81_0/b[15] col_256a_256x8m81_0/bb[22] VSS col_256a_256x8m81_0/WL[20]
+ col_256a_256x8m81_0/bb[6] VDD col_256a_256x8m81_0/WL[6] col_256a_256x8m81_0/bb[5]
+ col_256a_256x8m81_0/bb[20] col_256a_256x8m81_0/WL[17] col_256a_256x8m81_0/bb[4]
+ VSS col_256a_256x8m81_0/b[28] col_256a_256x8m81_0/b[21] col_256a_256x8m81_0/WL[31]
+ VDD VDD col_256a_256x8m81_0/b[26] VSS col_256a_256x8m81_0/b[5] col_256a_256x8m81_0/bb[9]
+ VDD col_256a_256x8m81_0/b[16] col_256a_256x8m81_0/WL[27] col_256a_256x8m81_0/b[19]
+ VSS col_256a_256x8m81_0/b[3] VDD col_256a_256x8m81_0/bb[2] col_256a_256x8m81_0/bb[18]
+ col_256a_256x8m81_0/WL[29] VSS col_256a_256x8m81_0/bb[3] col_256a_256x8m81_0/b[1]
+ col_256a_256x8m81_0/b[17] col_256a_256x8m81_0/bb[16] VDD VSS col_256a_256x8m81_0/bb[0]
+ col_256a_256x8m81_0/b[30] VDD VSS col_256a_256x8m81_0/b[10] VDD col_256a_256x8m81_0/bb[24]
+ VSS col_256a_256x8m81_0/b[24] col_256a_256x8m81_0/bb[8] VDD col_256a_256x8m81_0/b[31]
+ col_256a_256x8m81_0/b[25] col_256a_256x8m81_0/b[9] col_256a_256x8m81_0/b[2] col_256a_256x8m81_0/bb[26]
+ col_256a_256x8m81_0/bb[6] col_256a_256x8m81_0/b[23] col_256a_256x8m81_0/bb[4] VSS
+ col_256a_256x8m81_0/bb[22] col_256a_256x8m81_0/b[22] VSS VDD col_256a_256x8m81_0/b[5]
+ col_256a_256x8m81_0/bb[20] VSS VDD col_256a_256x8m81_0/b[3] col_256a_256x8m81_0/b[21]
+ ldummy_256x4_256x8m81_0/VSS col_256a_256x8m81_0/b[27] col_256a_256x8m81_0/bb[1]
+ col_256a_256x8m81_0/bb[2] col_256a_256x8m81_0/b[19] col_256a_256x8m81_0/b[29] col_256a_256x8m81_0/b[1]
+ VSS col_256a_256x8m81_0/bb[18] col_256a_256x8m81_0/b[20] col_256a_256x8m81_0/b[10]
+ VSS col_256a_256x8m81_0/b[11] col_256a_256x8m81_0/bb[28] col_256a_256x8m81_0/b[6]
+ VDD col_256a_256x8m81_0/bb[0] col_256a_256x8m81_0/b[17] col_256a_256x8m81_0/bb[27]
+ col_256a_256x8m81_0/bb[31] VSS col_256a_256x8m81_0/b[13] col_256a_256x8m81_0/bb[30]
+ VDD col_256a_256x8m81_0/bb[8] col_256a_256x8m81_0/bb[16] col_256a_256x8m81_0/bb[12]
+ col_256a_256x8m81_0/bb[25] col_256a_256x8m81_0/b[31] col_256a_256x8m81_0/b[9] col_256a_256x8m81_0/b[0]
+ col_256a_256x8m81_0/bb[10] col_256a_256x8m81_0/bb[24] col_256a_256x8m81_0/bb[14]
+ col_256a_256x8m81_0/b[23] col_256a_256x8m81_0/bb[10] col_256a_256x8m81_0/b[11] VSS
+ VSS col_256a_256x8m81_0/b[4] col_256a_256x8m81_0/b[15] col_256a_256x8m81_0/bb[21]
+ VDD col_256a_256x8m81_0/bb[11] col_256a_256x8m81_0/b[13] col_256a_256x8m81_0/bb[29]
+ VSS VDD col_256a_256x8m81_0/bb[23] col_256a_256x8m81_0/b[7] VDD VDD col_256a_256x8m81_0/bb[12]
+ col_256a_256x8m81_0/bb[15] VDD col_256a_256x8m81_0/b[8] VSS col_256a_256x8m81_0/bb[14]
+ ldummy_256x4_256x8m81
Xdcap_103_novia_256x8m81_0[0] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[1] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[2] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[3] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[4] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[5] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[6] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[7] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[8] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[9] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[10] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[11] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[12] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[13] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[14] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[15] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[16] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[17] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[18] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[19] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[20] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[21] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[22] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[23] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[24] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[25] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[26] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[27] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[28] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[29] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[30] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[31] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[32] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[33] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[34] VDD VDD VSS dcap_103_novia_256x8m81
Xdcap_103_novia_256x8m81_0[35] VDD VDD VSS dcap_103_novia_256x8m81
Xcol_256a_256x8m81_0 col_256a_256x8m81_0/pcb[0] col_256a_256x8m81_0/pcb[1] col_256a_256x8m81_0/pcb[3]
+ col_256a_256x8m81_0/pcb[2] col_256a_256x8m81_0/WEN[3] col_256a_256x8m81_0/WEN[2]
+ col_256a_256x8m81_0/WEN[1] col_256a_256x8m81_0/WEN[0] col_256a_256x8m81_0/WL[3]
+ col_256a_256x8m81_0/ypass[0] col_256a_256x8m81_0/ypass[1] col_256a_256x8m81_0/ypass[3]
+ col_256a_256x8m81_0/ypass[4] col_256a_256x8m81_0/ypass[5] col_256a_256x8m81_0/GWE
+ col_256a_256x8m81_0/WL[2] col_256a_256x8m81_0/WL[1] col_256a_256x8m81_0/WL[31] col_256a_256x8m81_0/WL[30]
+ col_256a_256x8m81_0/WL[29] col_256a_256x8m81_0/WL[24] col_256a_256x8m81_0/WL[23]
+ col_256a_256x8m81_0/WL[22] col_256a_256x8m81_0/WL[21] col_256a_256x8m81_0/WL[20]
+ col_256a_256x8m81_0/WL[19] col_256a_256x8m81_0/WL[12] col_256a_256x8m81_0/WL[11]
+ col_256a_256x8m81_0/WL[10] col_256a_256x8m81_0/WL[9] col_256a_256x8m81_0/WL[8] col_256a_256x8m81_0/WL[7]
+ col_256a_256x8m81_0/WL[6] col_256a_256x8m81_0/WL[5] col_256a_256x8m81_0/WL[4] col_256a_256x8m81_0/WL[18]
+ col_256a_256x8m81_0/WL[17] col_256a_256x8m81_0/WL[16] col_256a_256x8m81_0/WL[15]
+ col_256a_256x8m81_0/WL[14] col_256a_256x8m81_0/WL[13] col_256a_256x8m81_0/WL[28]
+ col_256a_256x8m81_0/WL[27] col_256a_256x8m81_0/WL[26] col_256a_256x8m81_0/WL[0]
+ col_256a_256x8m81_0/ypass[2] col_256a_256x8m81_0/WL[25] col_256a_256x8m81_0/b[13]
+ col_256a_256x8m81_0/b[16] col_256a_256x8m81_0/b[25] col_256a_256x8m81_0/din[1] col_256a_256x8m81_0/din[3]
+ col_256a_256x8m81_0/din[2] col_256a_256x8m81_0/din[0] col_256a_256x8m81_0/q[0] col_256a_256x8m81_0/q[1]
+ col_256a_256x8m81_0/q[2] col_256a_256x8m81_0/q[3] col_256a_256x8m81_0/b[17] col_256a_256x8m81_0/b[14]
+ col_256a_256x8m81_0/bb[10] col_256a_256x8m81_0/bb[11] col_256a_256x8m81_0/bb[12]
+ col_256a_256x8m81_0/bb[13] col_256a_256x8m81_0/bb[14] col_256a_256x8m81_0/bb[15]
+ col_256a_256x8m81_0/bb[16] col_256a_256x8m81_0/bb[20] col_256a_256x8m81_0/bb[29]
+ col_256a_256x8m81_0/bb[30] col_256a_256x8m81_0/bb[31] col_256a_256x8m81_0/b[30]
+ col_256a_256x8m81_0/b[15] col_256a_256x8m81_0/b[12] col_256a_256x8m81_0/b[0] col_256a_256x8m81_0/b[18]
+ col_256a_256x8m81_0/a_15501_29383# VSS col_256a_256x8m81_0/b[3] col_256a_256x8m81_0/a_15261_28608#
+ col_256a_256x8m81_0/bb[19] col_256a_256x8m81_0/b[21] col_256a_256x8m81_0/a_4701_29383#
+ col_256a_256x8m81_0/ypass[6] col_256a_256x8m81_0/ypass[7] col_256a_256x8m81_0/b[27]
+ col_256a_256x8m81_0/a_4461_28608# col_256a_256x8m81_0/a_15501_28608# col_256a_256x8m81_0/bb[22]
+ col_256a_256x8m81_0/bb[5] col_256a_256x8m81_0/b[6] col_256a_256x8m81_0/bb[3] col_256a_256x8m81_0/b[5]
+ col_256a_256x8m81_0/bb[23] col_256a_256x8m81_0/bb[0] col_256a_256x8m81_0/saout_m2_256x8m81_1/GWEN
+ col_256a_256x8m81_0/bb[4] col_256a_256x8m81_0/b[5] col_256a_256x8m81_0/b[26] col_256a_256x8m81_0/b[28]
+ col_256a_256x8m81_0/b[8] col_256a_256x8m81_0/a_15261_29383# col_256a_256x8m81_0/b[10]
+ col_256a_256x8m81_0/b[2] col_256a_256x8m81_0/bb[26] col_256a_256x8m81_0/b[7] col_256a_256x8m81_0/saout_m2_256x8m81_1/mux821_256x8m81_0/a_656_7735#
+ col_256a_256x8m81_0/b[1] col_256a_256x8m81_0/bb[6] col_256a_256x8m81_0/saout_R_m2_256x8m81_0/wen_wm1_256x8m81_0/wen
+ col_256a_256x8m81_0/b[20] col_256a_256x8m81_0/bb[25] col_256a_256x8m81_0/bb[27]
+ col_256a_256x8m81_0/bb[28] col_256a_256x8m81_0/b[11] col_256a_256x8m81_0/a_4701_28608#
+ col_256a_256x8m81_0/bb[18] col_256a_256x8m81_0/bb[9] col_256a_256x8m81_0/b[31] col_256a_256x8m81_0/saout_m2_256x8m81_1/sa_256x8m81_0/pcb
+ col_256a_256x8m81_0/bb[21] col_256a_256x8m81_0/bb[7] col_256a_256x8m81_0/saout_m2_256x8m81_0/pcb
+ col_256a_256x8m81_0/bb[2] col_256a_256x8m81_0/b[4] col_256a_256x8m81_0/bb[1] col_256a_256x8m81_0/saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb
+ col_256a_256x8m81_0/bb[17] col_256a_256x8m81_0/b[24] col_256a_256x8m81_0/saout_m2_256x8m81_0/WEN
+ col_256a_256x8m81_0/b[23] col_256a_256x8m81_0/bb[8] col_256a_256x8m81_0/b[22] col_256a_256x8m81_0/saout_R_m2_256x8m81_1/sa_256x8m81_0/pcb
+ col_256a_256x8m81_0/a_4461_29383# VDD col_256a_256x8m81_0/b[29] col_256a_256x8m81_0/bb[24]
+ col_256a_256x8m81_0/b[19] col_256a_256x8m81_0/b[9] VSS col_256a_256x8m81_0/men col_256a_256x8m81
.ends

.subckt gf180mcu_fd_ip_sram__sram256x8m8wm1 VSS CLK D[0] A[7] A[2] A[1] A[0] Q[2]
+ Q[3] CEN A[5] A[6] A[4] WEN[3] D[3] D[1] D[2] A[3] Q[1] Q[6] D[5] Q[4] WEN[5] WEN[2]
+ WEN[1] WEN[4] WEN[7] WEN[6] D[6] Q[5] Q[0] GWEN WEN[0] D[4] D[7] Q[7]
Xrcol4_256_256x8m81_0 rcol4_256_256x8m81_0/pcb[6] rcol4_256_256x8m81_0/pcb[7] rcol4_256_256x8m81_0/pcb[4]
+ VSS rcol4_256_256x8m81_0/PCB[8] WEN[7] WEN[4] rcol4_256_256x8m81_0/pcb[5] WEN[6]
+ WEN[5] rcol4_256_256x8m81_0/men rcol4_256_256x8m81_0/ypass[1] rcol4_256_256x8m81_0/ypass[2]
+ rcol4_256_256x8m81_0/ypass[3] rcol4_256_256x8m81_0/ypass[4] rcol4_256_256x8m81_0/ypass[5]
+ rcol4_256_256x8m81_0/ypass[6] rcol4_256_256x8m81_0/DWL rcol4_256_256x8m81_0/tblhl
+ rcol4_256_256x8m81_0/GWEN rcol4_256_256x8m81_0/ypass[0] rcol4_256_256x8m81_0/WL[23]
+ rcol4_256_256x8m81_0/WL[22] rcol4_256_256x8m81_0/WL[27] rcol4_256_256x8m81_0/WL[30]
+ rcol4_256_256x8m81_0/WL[18] rcol4_256_256x8m81_0/WL[15] rcol4_256_256x8m81_0/WL[12]
+ rcol4_256_256x8m81_0/ypass[7] rcol4_256_256x8m81_0/WL[13] rcol4_256_256x8m81_0/WL[14]
+ rcol4_256_256x8m81_0/WL[16] rcol4_256_256x8m81_0/WL[17] rcol4_256_256x8m81_0/WL[19]
+ rcol4_256_256x8m81_0/WL[28] D[4] D[7] Q[5] Q[6] Q[7] D[5] D[6] Q[4] rcol4_256_256x8m81_0/PCB[8]
+ rcol4_256_256x8m81_0/DWL WEN[7] rcol4_256_256x8m81_0/WL[2] rcol4_256_256x8m81_0/WL[3]
+ rcol4_256_256x8m81_0/WL[6] rcol4_256_256x8m81_0/WL[7] rcol4_256_256x8m81_0/WL[20]
+ rcol4_256_256x8m81_0/WL[21] rcol4_256_256x8m81_0/WL[4] rcol4_256_256x8m81_0/WL[5]
+ rcol4_256_256x8m81_0/WL[8] rcol4_256_256x8m81_0/WL[9] rcol4_256_256x8m81_0/WL[24]
+ rcol4_256_256x8m81_0/GWE rcol4_256_256x8m81_0/WL[29] rcol4_256_256x8m81_0/WL[25]
+ VSS rcol4_256_256x8m81_0/WL[26] rcol4_256_256x8m81_0/WL[10] rcol4_256_256x8m81_0/WL[11]
+ rcol4_256_256x8m81_0/WL[31] rcol4_256_256x8m81_0/WL[0] rcol4_256_256x8m81_0/WL[1]
+ VSS VSS rcol4_256_256x8m81
Xxdec32_256_256x8m81_0 rcol4_256_256x8m81_0/DWL rcol4_256_256x8m81_0/WL[31] rcol4_256_256x8m81_0/WL[29]
+ rcol4_256_256x8m81_0/WL[6] rcol4_256_256x8m81_0/WL[2] rcol4_256_256x8m81_0/WL[0]
+ rcol4_256_256x8m81_0/WL[5] rcol4_256_256x8m81_0/WL[7] rcol4_256_256x8m81_0/WL[8]
+ rcol4_256_256x8m81_0/WL[9] rcol4_256_256x8m81_0/WL[10] rcol4_256_256x8m81_0/WL[11]
+ rcol4_256_256x8m81_0/WL[12] rcol4_256_256x8m81_0/WL[13] rcol4_256_256x8m81_0/WL[14]
+ rcol4_256_256x8m81_0/WL[15] rcol4_256_256x8m81_0/WL[16] rcol4_256_256x8m81_0/WL[17]
+ rcol4_256_256x8m81_0/WL[18] xdec32_256_256x8m81_0/LWL[30] xdec32_256_256x8m81_0/LWL[31]
+ xdec32_256_256x8m81_0/LWL[20] xdec32_256_256x8m81_0/LWL[21] xdec32_256_256x8m81_0/LWL[22]
+ xdec32_256_256x8m81_0/LWL[13] xdec32_256_256x8m81_0/LWL[15] xdec32_256_256x8m81_0/LWL[16]
+ xdec32_256_256x8m81_0/LWL[18] xdec32_256_256x8m81_0/LWL[5] xdec32_256_256x8m81_0/LWL[4]
+ xdec32_256_256x8m81_0/LWL[3] xdec32_256_256x8m81_0/LWL[1] xdec32_256_256x8m81_0/LWL[8]
+ xdec32_256_256x8m81_0/LWL[9] xdec32_256_256x8m81_0/LWL[6] xdec32_256_256x8m81_0/DLWL
+ xdec32_256_256x8m81_0/xb[0] xdec32_256_256x8m81_0/xb[2] xdec32_256_256x8m81_0/xb[3]
+ xdec32_256_256x8m81_0/xa[7] xdec32_256_256x8m81_0/xa[6] xdec32_256_256x8m81_0/xa[5]
+ xdec32_256_256x8m81_0/xa[4] xdec32_256_256x8m81_0/xa[0] xdec32_256_256x8m81_0/xa[3]
+ xdec32_256_256x8m81_0/xa[2] xdec32_256_256x8m81_0/xc[1] xdec32_256_256x8m81_0/LWL[28]
+ xdec32_256_256x8m81_0/LWL[26] xdec32_256_256x8m81_0/LWL[29] xdec32_256_256x8m81_0/LWL[24]
+ rcol4_256_256x8m81_0/WL[22] rcol4_256_256x8m81_0/WL[20] rcol4_256_256x8m81_0/WL[27]
+ xdec32_256_256x8m81_0/LWL[27] xdec32_256_256x8m81_0/LWL[14] xdec32_256_256x8m81_0/xa[1]
+ xdec32_256_256x8m81_0/LWL[12] rcol4_256_256x8m81_0/WL[25] xdec32_256_256x8m81_0/LWL[25]
+ rcol4_256_256x8m81_0/WL[4] xdec32_256_256x8m81_0/LWL[10] xdec32_256_256x8m81_0/LWL[23]
+ xdec32_256_256x8m81_0/LWL[2] xdec32_256_256x8m81_0/LWL[0] xdec32_256_256x8m81_0/LWL[11]
+ VSS rcol4_256_256x8m81_0/WL[30] rcol4_256_256x8m81_0/WL[23] rcol4_256_256x8m81_0/WL[3]
+ rcol4_256_256x8m81_0/WL[28] rcol4_256_256x8m81_0/WL[26] rcol4_256_256x8m81_0/WL[24]
+ xdec32_256_256x8m81_0/LWL[19] rcol4_256_256x8m81_0/WL[21] rcol4_256_256x8m81_0/WL[1]
+ xdec32_256_256x8m81_0/xb[1] xdec32_256_256x8m81_0/LWL[7] xdec32_256_256x8m81_0/LWL[17]
+ rcol4_256_256x8m81_0/WL[19] rcol4_256_256x8m81_0/men VSS VSS xdec32_256_256x8m81
Xcontrol_512x8_256x8m81_0 rcol4_256_256x8m81_0/GWE GWEN VSS VSS rcol4_256_256x8m81_0/ypass[7]
+ rcol4_256_256x8m81_0/ypass[6] rcol4_256_256x8m81_0/ypass[5] rcol4_256_256x8m81_0/ypass[4]
+ rcol4_256_256x8m81_0/ypass[3] rcol4_256_256x8m81_0/ypass[2] rcol4_256_256x8m81_0/ypass[1]
+ rcol4_256_256x8m81_0/ypass[0] control_512x8_256x8m81_0/LYS[0] control_512x8_256x8m81_0/LYS[1]
+ control_512x8_256x8m81_0/LYS[2] control_512x8_256x8m81_0/LYS[3] control_512x8_256x8m81_0/LYS[6]
+ control_512x8_256x8m81_0/LYS[5] control_512x8_256x8m81_0/LYS[4] control_512x8_256x8m81_0/LYS[7]
+ rcol4_256_256x8m81_0/tblhl rcol4_256_256x8m81_0/GWEN xdec32_256_256x8m81_0/xb[3]
+ xdec32_256_256x8m81_0/xb[2] xdec32_256_256x8m81_0/xb[0] xdec32_256_256x8m81_0/xa[7]
+ xdec32_256_256x8m81_0/xa[6] xdec32_256_256x8m81_0/xa[5] xdec32_256_256x8m81_0/xa[4]
+ xdec32_256_256x8m81_0/xa[3] xdec32_256_256x8m81_0/xa[2] xdec32_256_256x8m81_0/xb[1]
+ control_512x8_256x8m81_0/xc[3] xdec32_256_256x8m81_0/xc[1] control_512x8_256x8m81_0/xc[2]
+ control_512x8_256x8m81_0/xc[0] xdec32_256_256x8m81_0/xa[0] xdec32_256_256x8m81_0/xa[1]
+ VSS A[7] CLK A[2] A[6] A[3] A[4] A[5] VSS VSS control_512x8_256x8m81_0/LYS[2] rcol4_256_256x8m81_0/tblhl
+ A[0] CEN rcol4_256_256x8m81_0/men A[1] VSS VSS VSS control_512x8_256x8m81
Xlcol4_256_256x8m81_0 lcol4_256_256x8m81_0/pcb[2] lcol4_256_256x8m81_0/pcb[3] lcol4_256_256x8m81_0/pcb[0]
+ lcol4_256_256x8m81_0/pcb[1] VSS WEN[0] WEN[1] WEN[2] WEN[3] lcol4_256_256x8m81_0/WL[25]
+ lcol4_256_256x8m81_0/WL[24] lcol4_256_256x8m81_0/WL[23] lcol4_256_256x8m81_0/WL[22]
+ lcol4_256_256x8m81_0/WL[21] lcol4_256_256x8m81_0/WL[20] lcol4_256_256x8m81_0/WL[19]
+ lcol4_256_256x8m81_0/WL[18] lcol4_256_256x8m81_0/WL[17] lcol4_256_256x8m81_0/WL[16]
+ lcol4_256_256x8m81_0/WL[15] lcol4_256_256x8m81_0/WL[14] lcol4_256_256x8m81_0/WL[13]
+ lcol4_256_256x8m81_0/WL[12] lcol4_256_256x8m81_0/WL[11] lcol4_256_256x8m81_0/WL[10]
+ lcol4_256_256x8m81_0/WL[9] lcol4_256_256x8m81_0/WL[8] lcol4_256_256x8m81_0/WL[7]
+ lcol4_256_256x8m81_0/WL[6] lcol4_256_256x8m81_0/WL[5] lcol4_256_256x8m81_0/WL[4]
+ lcol4_256_256x8m81_0/WL[3] lcol4_256_256x8m81_0/WL[2] lcol4_256_256x8m81_0/WL[1]
+ lcol4_256_256x8m81_0/WL[0] lcol4_256_256x8m81_0/WL[31] lcol4_256_256x8m81_0/WL[30]
+ lcol4_256_256x8m81_0/WL[29] lcol4_256_256x8m81_0/WL[28] lcol4_256_256x8m81_0/WL[27]
+ lcol4_256_256x8m81_0/WL[26] lcol4_256_256x8m81_0/men lcol4_256_256x8m81_0/ypass[0]
+ lcol4_256_256x8m81_0/ypass[1] lcol4_256_256x8m81_0/ypass[2] lcol4_256_256x8m81_0/ypass[3]
+ lcol4_256_256x8m81_0/ypass[4] lcol4_256_256x8m81_0/ypass[5] lcol4_256_256x8m81_0/ypass[6]
+ lcol4_256_256x8m81_0/ypass[7] lcol4_256_256x8m81_0/GWEN lcol4_256_256x8m81_0/GWE
+ D[0] D[1] D[3] D[2] Q[0] Q[1] Q[2] Q[3] xdec32_256_256x8m81_0/LWL[7] rcol4_256_256x8m81_0/GWEN
+ VSS xdec32_256_256x8m81_0/LWL[8] xdec32_256_256x8m81_0/LWL[9] VSS VSS xdec32_256_256x8m81_0/LWL[20]
+ xdec32_256_256x8m81_0/LWL[21] xdec32_256_256x8m81_0/LWL[22] xdec32_256_256x8m81_0/LWL[23]
+ VSS xdec32_256_256x8m81_0/LWL[24] WEN[3] xdec32_256_256x8m81_0/LWL[25] xdec32_256_256x8m81_0/LWL[26]
+ xdec32_256_256x8m81_0/LWL[27] xdec32_256_256x8m81_0/LWL[28] xdec32_256_256x8m81_0/LWL[29]
+ VSS WEN[0] VSS xdec32_256_256x8m81_0/LWL[10] VSS rcol4_256_256x8m81_0/men xdec32_256_256x8m81_0/LWL[11]
+ rcol4_256_256x8m81_0/GWE xdec32_256_256x8m81_0/LWL[12] xdec32_256_256x8m81_0/LWL[13]
+ xdec32_256_256x8m81_0/LWL[30] lcol4_256_256x8m81_0/col_256a_256x8m81_0/saout_m2_256x8m81_0/pcb
+ control_512x8_256x8m81_0/LYS[0] VSS xdec32_256_256x8m81_0/LWL[14] xdec32_256_256x8m81_0/LWL[31]
+ control_512x8_256x8m81_0/LYS[1] xdec32_256_256x8m81_0/LWL[0] xdec32_256_256x8m81_0/LWL[15]
+ control_512x8_256x8m81_0/LYS[2] xdec32_256_256x8m81_0/LWL[1] xdec32_256_256x8m81_0/LWL[16]
+ control_512x8_256x8m81_0/LYS[3] xdec32_256_256x8m81_0/LWL[2] xdec32_256_256x8m81_0/LWL[17]
+ control_512x8_256x8m81_0/LYS[4] xdec32_256_256x8m81_0/LWL[3] VSS xdec32_256_256x8m81_0/LWL[18]
+ control_512x8_256x8m81_0/LYS[5] xdec32_256_256x8m81_0/LWL[4] lcol4_256_256x8m81_0/col_256a_256x8m81_0/saout_R_m2_256x8m81_1/sa_256x8m81_0/pcb
+ xdec32_256_256x8m81_0/LWL[19] control_512x8_256x8m81_0/LYS[6] xdec32_256_256x8m81_0/LWL[5]
+ lcol4_256_256x8m81_0/col_256a_256x8m81_0/saout_m2_256x8m81_1/sa_256x8m81_0/pcb lcol4_256_256x8m81_0/col_256a_256x8m81_0/saout_R_m2_256x8m81_0/sa_256x8m81_0/pcb
+ VSS control_512x8_256x8m81_0/LYS[7] VSS xdec32_256_256x8m81_0/LWL[6] VSS lcol4_256_256x8m81
.ends

