magic
tech gf180mcuC
magscale 1 10
timestamp 1669650257
<< checkpaint >>
rect 66400 66400 73000 73000
<< metal4 >>
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68400 68769 68769 ne
rect 68769 68400 71000 68769
<< end >>
