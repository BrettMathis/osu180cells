magic
tech gf180mcuB
magscale 1 10
timestamp 1669648930
<< checkpaint >>
rect 11108 11108 48414 47051
<< metal1 >>
rect 13108 44848 13280 45051
tri 13280 44848 13352 44920 sw
tri 13108 44828 13128 44848 ne
rect 13128 44828 13352 44848
tri 13352 44828 13372 44848 sw
tri 13128 44584 13372 44828 ne
tri 13372 44584 13616 44828 sw
tri 13372 44340 13616 44584 ne
tri 13616 44340 13860 44584 sw
tri 13616 44096 13860 44340 ne
tri 13860 44096 14104 44340 sw
tri 13860 43852 14104 44096 ne
tri 14104 43852 14348 44096 sw
tri 14104 43608 14348 43852 ne
tri 14348 43608 14592 43852 sw
tri 14348 43364 14592 43608 ne
tri 14592 43364 14836 43608 sw
tri 14592 43120 14836 43364 ne
tri 14836 43120 15080 43364 sw
tri 14836 42876 15080 43120 ne
tri 15080 42876 15324 43120 sw
tri 15080 42632 15324 42876 ne
tri 15324 42632 15568 42876 sw
tri 15324 42388 15568 42632 ne
tri 15568 42388 15812 42632 sw
tri 15568 42144 15812 42388 ne
tri 15812 42144 16056 42388 sw
tri 15812 41900 16056 42144 ne
tri 16056 41900 16300 42144 sw
tri 16056 41656 16300 41900 ne
tri 16300 41656 16544 41900 sw
tri 16300 41412 16544 41656 ne
tri 16544 41412 16788 41656 sw
tri 16544 41168 16788 41412 ne
tri 16788 41168 17032 41412 sw
tri 16788 40924 17032 41168 ne
tri 17032 40924 17276 41168 sw
tri 17032 40680 17276 40924 ne
tri 17276 40680 17520 40924 sw
tri 17276 40436 17520 40680 ne
tri 17520 40436 17764 40680 sw
tri 17520 40192 17764 40436 ne
tri 17764 40192 18008 40436 sw
tri 17764 39948 18008 40192 ne
tri 18008 39948 18252 40192 sw
tri 18008 39704 18252 39948 ne
tri 18252 39704 18496 39948 sw
tri 18252 39460 18496 39704 ne
tri 18496 39460 18740 39704 sw
tri 18496 39216 18740 39460 ne
tri 18740 39216 18984 39460 sw
tri 18740 38972 18984 39216 ne
tri 18984 38972 19228 39216 sw
tri 18984 38728 19228 38972 ne
tri 19228 38728 19472 38972 sw
tri 19228 38484 19472 38728 ne
tri 19472 38484 19716 38728 sw
tri 19472 38240 19716 38484 ne
tri 19716 38240 19960 38484 sw
tri 19716 37996 19960 38240 ne
tri 19960 37996 20204 38240 sw
tri 19960 37752 20204 37996 ne
tri 20204 37752 20448 37996 sw
tri 20204 37508 20448 37752 ne
tri 20448 37508 20692 37752 sw
tri 20448 37264 20692 37508 ne
tri 20692 37264 20936 37508 sw
tri 20692 37020 20936 37264 ne
tri 20936 37020 21180 37264 sw
tri 20936 36776 21180 37020 ne
tri 21180 36776 21424 37020 sw
tri 21180 36532 21424 36776 ne
tri 21424 36532 21668 36776 sw
tri 21424 36288 21668 36532 ne
tri 21668 36288 21912 36532 sw
tri 21668 36044 21912 36288 ne
tri 21912 36044 22156 36288 sw
tri 21912 35800 22156 36044 ne
tri 22156 35800 22400 36044 sw
tri 22156 35556 22400 35800 ne
tri 22400 35556 22644 35800 sw
tri 22400 35312 22644 35556 ne
tri 22644 35312 22888 35556 sw
tri 22644 35068 22888 35312 ne
tri 22888 35068 23132 35312 sw
tri 22888 34824 23132 35068 ne
tri 23132 34824 23376 35068 sw
tri 23132 34580 23376 34824 ne
tri 23376 34580 23620 34824 sw
tri 23376 34336 23620 34580 ne
tri 23620 34336 23864 34580 sw
tri 23620 34092 23864 34336 ne
tri 23864 34092 24108 34336 sw
tri 23864 33848 24108 34092 ne
tri 24108 33848 24352 34092 sw
tri 24108 33604 24352 33848 ne
tri 24352 33604 24596 33848 sw
tri 24352 33360 24596 33604 ne
tri 24596 33360 24840 33604 sw
tri 24596 33116 24840 33360 ne
tri 24840 33116 25084 33360 sw
tri 24840 32872 25084 33116 ne
tri 25084 32872 25328 33116 sw
tri 25084 32628 25328 32872 ne
tri 25328 32628 25572 32872 sw
tri 25328 32384 25572 32628 ne
tri 25572 32384 25816 32628 sw
tri 25572 32140 25816 32384 ne
tri 25816 32140 26060 32384 sw
tri 25816 31896 26060 32140 ne
tri 26060 31896 26304 32140 sw
tri 26060 31652 26304 31896 ne
tri 26304 31652 26548 31896 sw
tri 26304 31408 26548 31652 ne
tri 26548 31408 26792 31652 sw
tri 26548 31164 26792 31408 ne
tri 26792 31164 27036 31408 sw
tri 26792 30920 27036 31164 ne
tri 27036 30920 27280 31164 sw
tri 27036 30676 27280 30920 ne
tri 27280 30676 27524 30920 sw
tri 27280 30432 27524 30676 ne
tri 27524 30432 27768 30676 sw
tri 27524 30188 27768 30432 ne
tri 27768 30188 28012 30432 sw
tri 27768 29944 28012 30188 ne
tri 28012 29944 28256 30188 sw
tri 28012 29700 28256 29944 ne
tri 28256 29700 28500 29944 sw
tri 28256 29456 28500 29700 ne
tri 28500 29456 28744 29700 sw
tri 28500 29212 28744 29456 ne
tri 28744 29212 28988 29456 sw
tri 28744 28968 28988 29212 ne
tri 28988 28968 29232 29212 sw
tri 28988 28724 29232 28968 ne
tri 29232 28724 29476 28968 sw
tri 29232 28480 29476 28724 ne
tri 29476 28480 29720 28724 sw
tri 29476 28236 29720 28480 ne
tri 29720 28236 29964 28480 sw
tri 29720 27992 29964 28236 ne
tri 29964 27992 30208 28236 sw
tri 29964 27748 30208 27992 ne
tri 30208 27748 30452 27992 sw
tri 30208 27504 30452 27748 ne
tri 30452 27504 30696 27748 sw
tri 30452 27260 30696 27504 ne
tri 30696 27260 30940 27504 sw
tri 30696 27016 30940 27260 ne
tri 30940 27016 31184 27260 sw
tri 30940 26772 31184 27016 ne
tri 31184 26772 31428 27016 sw
tri 31184 26528 31428 26772 ne
tri 31428 26528 31672 26772 sw
tri 31428 26284 31672 26528 ne
tri 31672 26284 31916 26528 sw
tri 31672 26040 31916 26284 ne
tri 31916 26040 32160 26284 sw
tri 31916 25796 32160 26040 ne
tri 32160 25796 32404 26040 sw
tri 32160 25552 32404 25796 ne
tri 32404 25552 32648 25796 sw
tri 32404 25308 32648 25552 ne
tri 32648 25308 32892 25552 sw
tri 32648 25064 32892 25308 ne
tri 32892 25064 33136 25308 sw
tri 32892 24820 33136 25064 ne
tri 33136 24820 33380 25064 sw
tri 33136 24576 33380 24820 ne
tri 33380 24576 33624 24820 sw
tri 33380 24332 33624 24576 ne
tri 33624 24332 33868 24576 sw
tri 33624 24088 33868 24332 ne
tri 33868 24088 34112 24332 sw
tri 33868 23844 34112 24088 ne
tri 34112 23844 34356 24088 sw
tri 34112 23600 34356 23844 ne
tri 34356 23600 34600 23844 sw
tri 34356 23356 34600 23600 ne
tri 34600 23356 34844 23600 sw
tri 34600 23112 34844 23356 ne
tri 34844 23112 35088 23356 sw
tri 34844 22868 35088 23112 ne
tri 35088 22868 35332 23112 sw
tri 35088 22624 35332 22868 ne
tri 35332 22624 35576 22868 sw
tri 35332 22380 35576 22624 ne
tri 35576 22380 35820 22624 sw
tri 35576 22136 35820 22380 ne
tri 35820 22136 36064 22380 sw
tri 35820 21892 36064 22136 ne
tri 36064 21892 36308 22136 sw
tri 36064 21648 36308 21892 ne
tri 36308 21648 36552 21892 sw
tri 36308 21404 36552 21648 ne
tri 36552 21404 36796 21648 sw
tri 36552 21160 36796 21404 ne
tri 36796 21160 37040 21404 sw
tri 36796 20916 37040 21160 ne
tri 37040 20916 37284 21160 sw
tri 37040 20672 37284 20916 ne
tri 37284 20672 37528 20916 sw
tri 37284 20428 37528 20672 ne
tri 37528 20428 37772 20672 sw
tri 37528 20184 37772 20428 ne
tri 37772 20184 38016 20428 sw
tri 37772 19940 38016 20184 ne
tri 38016 19940 38260 20184 sw
tri 38016 19696 38260 19940 ne
tri 38260 19696 38504 19940 sw
tri 38260 19452 38504 19696 ne
tri 38504 19452 38748 19696 sw
tri 38504 19208 38748 19452 ne
tri 38748 19208 38992 19452 sw
tri 38748 18964 38992 19208 ne
tri 38992 18964 39236 19208 sw
tri 38992 18720 39236 18964 ne
tri 39236 18720 39480 18964 sw
tri 39236 18476 39480 18720 ne
tri 39480 18476 39724 18720 sw
tri 39480 18232 39724 18476 ne
tri 39724 18232 39968 18476 sw
tri 39724 17988 39968 18232 ne
tri 39968 17988 40212 18232 sw
tri 39968 17744 40212 17988 ne
tri 40212 17744 40456 17988 sw
tri 40212 17500 40456 17744 ne
tri 40456 17500 40700 17744 sw
tri 40456 17256 40700 17500 ne
tri 40700 17256 40944 17500 sw
tri 40700 17012 40944 17256 ne
tri 40944 17012 41188 17256 sw
tri 40944 16768 41188 17012 ne
tri 41188 16768 41432 17012 sw
tri 41188 16524 41432 16768 ne
tri 41432 16524 41676 16768 sw
tri 41432 16280 41676 16524 ne
tri 41676 16280 41920 16524 sw
tri 41676 16036 41920 16280 ne
tri 41920 16036 42164 16280 sw
tri 41920 15792 42164 16036 ne
tri 42164 15792 42408 16036 sw
tri 42164 15548 42408 15792 ne
tri 42408 15548 42652 15792 sw
tri 42408 15304 42652 15548 ne
tri 42652 15304 42896 15548 sw
tri 42652 15060 42896 15304 ne
tri 42896 15060 43140 15304 sw
tri 42896 14816 43140 15060 ne
tri 43140 14816 43384 15060 sw
tri 43140 14572 43384 14816 ne
tri 43384 14572 43628 14816 sw
tri 43384 14328 43628 14572 ne
tri 43628 14328 43872 14572 sw
tri 43628 14084 43872 14328 ne
tri 43872 14084 44116 14328 sw
tri 43872 13840 44116 14084 ne
tri 44116 13840 44360 14084 sw
tri 44116 13596 44360 13840 ne
tri 44360 13596 44604 13840 sw
tri 44360 13352 44604 13596 ne
tri 44604 13352 44848 13596 sw
tri 44604 13108 44848 13352 ne
tri 44848 13280 44920 13352 sw
rect 44848 13108 46414 13280
<< end >>
