magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4342 1094
<< pwell >>
rect -86 -86 4342 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 215 836 333
rect 1016 215 1136 333
rect 1240 215 1360 333
rect 1408 215 1528 333
rect 1640 215 1760 333
rect 1968 215 2088 333
rect 2136 215 2256 333
rect 2360 215 2480 333
rect 2584 215 2704 333
rect 3072 175 3192 333
rect 3240 175 3360 333
rect 3464 175 3584 333
rect 3632 175 3752 333
rect 4012 69 4132 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 736 573 836 773
rect 940 573 1040 773
rect 1144 573 1244 773
rect 1348 573 1448 773
rect 1640 667 1740 867
rect 1988 667 2088 867
rect 2280 573 2380 773
rect 2484 573 2584 773
rect 2688 573 2788 773
rect 3056 573 3156 849
rect 3260 573 3360 849
rect 3464 573 3564 849
rect 3668 573 3768 849
rect 4016 573 4116 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 274 716 333
rect 628 228 641 274
rect 687 228 716 274
rect 628 215 716 228
rect 836 320 1016 333
rect 836 274 865 320
rect 911 274 1016 320
rect 836 215 1016 274
rect 1136 320 1240 333
rect 1136 274 1165 320
rect 1211 274 1240 320
rect 1136 215 1240 274
rect 1360 215 1408 333
rect 1528 215 1640 333
rect 1760 274 1968 333
rect 1760 228 1789 274
rect 1835 228 1968 274
rect 1760 215 1968 228
rect 2088 215 2136 333
rect 2256 320 2360 333
rect 2256 274 2285 320
rect 2331 274 2360 320
rect 2256 215 2360 274
rect 2480 320 2584 333
rect 2480 274 2509 320
rect 2555 274 2584 320
rect 2480 215 2584 274
rect 2704 320 2792 333
rect 2704 274 2733 320
rect 2779 274 2792 320
rect 2704 215 2792 274
rect 2984 320 3072 333
rect 2984 274 2997 320
rect 3043 274 3072 320
rect 2984 175 3072 274
rect 3192 175 3240 333
rect 3360 234 3464 333
rect 3360 188 3389 234
rect 3435 188 3464 234
rect 3360 175 3464 188
rect 3584 175 3632 333
rect 3752 320 3840 333
rect 3752 274 3781 320
rect 3827 274 3840 320
rect 3752 175 3840 274
rect 3924 320 4012 333
rect 3924 180 3937 320
rect 3983 180 4012 320
rect 3924 69 4012 180
rect 4132 222 4220 333
rect 4132 82 4161 222
rect 4207 82 4220 222
rect 4132 69 4220 82
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 1508 932 1580 945
rect 1508 886 1521 932
rect 1567 886 1580 932
rect 2148 932 2220 945
rect 1508 867 1580 886
rect 2148 886 2161 932
rect 2207 886 2220 932
rect 2148 867 2220 886
rect 1508 773 1640 867
rect 448 586 477 726
rect 523 586 536 726
rect 448 573 536 586
rect 648 760 736 773
rect 648 714 661 760
rect 707 714 736 760
rect 648 573 736 714
rect 836 726 940 773
rect 836 586 865 726
rect 911 586 940 726
rect 836 573 940 586
rect 1040 726 1144 773
rect 1040 586 1069 726
rect 1115 586 1144 726
rect 1040 573 1144 586
rect 1244 726 1348 773
rect 1244 680 1273 726
rect 1319 680 1348 726
rect 1244 573 1348 680
rect 1448 667 1640 773
rect 1740 726 1828 867
rect 1740 680 1769 726
rect 1815 680 1828 726
rect 1740 667 1828 680
rect 1900 726 1988 867
rect 1900 680 1913 726
rect 1959 680 1988 726
rect 1900 667 1988 680
rect 2088 773 2220 867
rect 2968 836 3056 849
rect 2968 790 2981 836
rect 3027 790 3056 836
rect 2088 667 2280 773
rect 1448 573 1528 667
rect 2200 573 2280 667
rect 2380 726 2484 773
rect 2380 586 2409 726
rect 2455 586 2484 726
rect 2380 573 2484 586
rect 2584 726 2688 773
rect 2584 586 2613 726
rect 2659 586 2688 726
rect 2584 573 2688 586
rect 2788 632 2876 773
rect 2788 586 2817 632
rect 2863 586 2876 632
rect 2788 573 2876 586
rect 2968 573 3056 790
rect 3156 632 3260 849
rect 3156 586 3185 632
rect 3231 586 3260 632
rect 3156 573 3260 586
rect 3360 836 3464 849
rect 3360 790 3389 836
rect 3435 790 3464 836
rect 3360 573 3464 790
rect 3564 634 3668 849
rect 3564 588 3593 634
rect 3639 588 3668 634
rect 3564 573 3668 588
rect 3768 836 3856 849
rect 3768 696 3797 836
rect 3843 696 3856 836
rect 3768 573 3856 696
rect 3928 726 4016 939
rect 3928 586 3941 726
rect 3987 586 4016 726
rect 3928 573 4016 586
rect 4116 926 4204 939
rect 4116 786 4145 926
rect 4191 786 4204 926
rect 4116 573 4204 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 228 687 274
rect 865 274 911 320
rect 1165 274 1211 320
rect 1789 228 1835 274
rect 2285 274 2331 320
rect 2509 274 2555 320
rect 2733 274 2779 320
rect 2997 274 3043 320
rect 3389 188 3435 234
rect 3781 274 3827 320
rect 3937 180 3983 320
rect 4161 82 4207 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 1521 886 1567 932
rect 2161 886 2207 932
rect 477 586 523 726
rect 661 714 707 760
rect 865 586 911 726
rect 1069 586 1115 726
rect 1273 680 1319 726
rect 1769 680 1815 726
rect 1913 680 1959 726
rect 2981 790 3027 836
rect 2409 586 2455 726
rect 2613 586 2659 726
rect 2817 586 2863 632
rect 3185 586 3231 632
rect 3389 790 3435 836
rect 3593 588 3639 634
rect 3797 696 3843 836
rect 3941 586 3987 726
rect 4145 786 4191 926
<< polysilicon >>
rect 348 909 1040 949
rect 144 849 244 893
rect 348 849 448 909
rect 736 773 836 817
rect 940 773 1040 909
rect 1640 867 1740 911
rect 1988 867 2088 911
rect 1144 852 1244 865
rect 1144 806 1157 852
rect 1203 806 1244 852
rect 1144 773 1244 806
rect 1348 773 1448 817
rect 2280 913 3156 953
rect 4016 939 4116 983
rect 2280 773 2380 913
rect 2484 852 2584 865
rect 2484 806 2497 852
rect 2543 806 2584 852
rect 3056 849 3156 913
rect 3260 849 3360 893
rect 3464 849 3564 893
rect 3668 849 3768 893
rect 2484 773 2584 806
rect 2688 773 2788 817
rect 144 504 244 573
rect 144 458 157 504
rect 203 458 244 504
rect 144 377 244 458
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 736 523 836 573
rect 940 529 1040 573
rect 736 477 749 523
rect 795 477 836 523
rect 1144 513 1244 573
rect 1348 513 1448 573
rect 736 377 836 477
rect 1096 473 1244 513
rect 1408 480 1528 513
rect 1096 377 1136 473
rect 1408 434 1421 480
rect 1467 434 1528 480
rect 407 366 468 377
rect 348 333 468 366
rect 716 333 836 377
rect 1016 333 1136 377
rect 1240 412 1360 425
rect 1240 366 1257 412
rect 1303 366 1360 412
rect 1240 333 1360 366
rect 1408 333 1528 434
rect 1640 377 1740 667
rect 1988 572 2088 667
rect 1988 526 2001 572
rect 2047 526 2088 572
rect 1988 377 2088 526
rect 2280 513 2380 573
rect 1640 333 1760 377
rect 1968 333 2088 377
rect 2136 473 2380 513
rect 2484 513 2584 573
rect 2688 529 2788 573
rect 2484 473 2624 513
rect 2136 333 2256 473
rect 2584 377 2624 473
rect 2748 437 2788 529
rect 3056 540 3156 573
rect 3056 494 3069 540
rect 3115 494 3156 540
rect 2748 397 2924 437
rect 2360 333 2480 377
rect 2584 333 2704 377
rect 2852 317 2924 397
rect 3056 393 3156 494
rect 3072 377 3156 393
rect 3260 412 3360 573
rect 3260 377 3301 412
rect 3072 333 3192 377
rect 3240 366 3301 377
rect 3347 366 3360 412
rect 3240 333 3360 366
rect 3464 497 3564 573
rect 3464 451 3502 497
rect 3548 451 3564 497
rect 3464 377 3564 451
rect 3668 540 3768 573
rect 3668 494 3692 540
rect 3738 494 3768 540
rect 3668 481 3768 494
rect 3668 377 3708 481
rect 4016 465 4116 573
rect 3836 452 4116 465
rect 3836 406 3849 452
rect 3895 406 4116 452
rect 3836 393 4116 406
rect 4012 377 4116 393
rect 3464 333 3584 377
rect 3632 333 3752 377
rect 4012 333 4132 377
rect 2852 271 2865 317
rect 2911 271 2924 317
rect 2852 258 2924 271
rect 124 131 244 175
rect 348 115 468 175
rect 716 171 836 215
rect 1016 171 1136 215
rect 1240 115 1360 215
rect 1408 171 1528 215
rect 348 75 1360 115
rect 1640 75 1760 215
rect 1968 171 2088 215
rect 2136 171 2256 215
rect 2360 182 2480 215
rect 2360 136 2373 182
rect 2419 136 2480 182
rect 2584 171 2704 215
rect 2360 123 2480 136
rect 3072 131 3192 175
rect 3240 131 3360 175
rect 3464 75 3584 175
rect 3632 131 3752 175
rect 1640 35 3584 75
rect 4012 25 4132 69
<< polycontact >>
rect 1157 806 1203 852
rect 2497 806 2543 852
rect 157 458 203 504
rect 361 366 407 412
rect 749 477 795 523
rect 1421 434 1467 480
rect 1257 366 1303 412
rect 2001 526 2047 572
rect 3069 494 3115 540
rect 3301 366 3347 412
rect 3502 451 3548 497
rect 3692 494 3738 540
rect 3849 406 3895 452
rect 2865 271 2911 317
rect 2373 136 2419 182
<< metal1 >>
rect 0 932 4256 1098
rect 0 918 1521 932
rect 273 836 319 918
rect 69 739 115 750
rect 661 760 707 918
rect 1567 918 2161 932
rect 1521 875 1567 886
rect 2207 926 4256 932
rect 2207 918 4145 926
rect 2161 875 2207 886
rect 2497 852 2543 863
rect 273 685 319 696
rect 477 726 523 737
rect 115 599 407 634
rect 69 588 407 599
rect 142 504 315 542
rect 142 458 157 504
rect 203 458 315 504
rect 142 447 315 458
rect 361 412 407 588
rect 361 348 407 366
rect 49 320 407 348
rect 95 302 407 320
rect 661 703 707 714
rect 753 806 1157 852
rect 1203 829 1214 852
rect 1203 806 2497 829
rect 753 783 2543 806
rect 2970 836 3038 918
rect 2970 790 2981 836
rect 3027 790 3038 836
rect 3378 836 3446 918
rect 3378 790 3389 836
rect 3435 790 3446 836
rect 3797 836 3843 918
rect 753 657 799 783
rect 523 611 799 657
rect 865 726 911 737
rect 523 586 543 611
rect 477 320 543 586
rect 589 523 795 542
rect 589 477 749 523
rect 589 466 795 477
rect 95 274 131 302
rect 49 263 131 274
rect 477 274 497 320
rect 865 320 911 586
rect 1069 726 1115 737
rect 1273 726 1815 737
rect 1319 680 1769 726
rect 1273 669 1815 680
rect 1913 726 2455 737
rect 1959 689 2409 726
rect 1959 680 2331 689
rect 1913 669 2331 680
rect 1069 583 1115 586
rect 1069 572 2047 583
rect 1069 537 2001 572
rect 477 263 543 274
rect 641 274 687 285
rect 273 234 319 245
rect 273 90 319 188
rect 865 263 911 274
rect 1165 320 1211 537
rect 2001 515 2047 526
rect 1421 480 1467 491
rect 2278 469 2331 669
rect 2409 575 2455 586
rect 2613 726 3738 737
rect 2659 691 3738 726
rect 1467 434 2331 469
rect 1421 423 2331 434
rect 1257 412 1303 423
rect 1303 366 2239 377
rect 1257 331 2239 366
rect 1165 263 1211 274
rect 1789 274 1835 285
rect 641 90 687 228
rect 1789 90 1835 228
rect 2193 182 2239 331
rect 2285 320 2331 423
rect 2613 331 2659 586
rect 2817 632 2863 643
rect 2817 423 2863 586
rect 3185 632 3231 643
rect 2909 540 3115 561
rect 2909 494 3069 540
rect 2909 466 3115 494
rect 2285 263 2331 274
rect 2509 320 2659 331
rect 2555 274 2659 320
rect 2509 263 2659 274
rect 2733 420 2863 423
rect 3185 420 3231 586
rect 3593 634 3646 645
rect 3639 588 3646 634
rect 3593 577 3646 588
rect 3393 497 3554 552
rect 3393 451 3502 497
rect 3548 451 3554 497
rect 3393 440 3554 451
rect 2733 374 3231 420
rect 3301 412 3347 423
rect 2733 320 2779 374
rect 2733 263 2779 274
rect 2865 317 2911 328
rect 2865 182 2911 271
rect 2997 320 3043 374
rect 3600 405 3646 577
rect 3692 540 3738 691
rect 4191 918 4256 926
rect 4145 775 4191 786
rect 3797 685 3843 696
rect 3941 726 4002 737
rect 3692 483 3738 494
rect 3987 586 4002 726
rect 3782 452 3895 463
rect 3782 406 3849 452
rect 3782 405 3895 406
rect 3600 395 3895 405
rect 3600 394 3827 395
rect 3347 366 3827 394
rect 3301 348 3827 366
rect 2997 263 3043 274
rect 3781 320 3827 348
rect 3941 331 4002 586
rect 3781 263 3827 274
rect 3937 320 4002 331
rect 2193 136 2373 182
rect 2419 136 2911 182
rect 3389 234 3435 245
rect 3389 90 3435 188
rect 3983 180 4002 320
rect 3937 169 4002 180
rect 4161 222 4207 233
rect 0 82 4161 90
rect 4207 82 4256 90
rect 0 -90 4256 82
<< labels >>
flabel metal1 s 142 447 315 542 0 FreeSans 200 0 0 0 CLKN
port 4 nsew clock input
flabel metal1 s 589 466 795 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3941 331 4002 737 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3393 440 3554 552 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 2909 466 3115 561 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 4256 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1789 245 1835 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 169 4002 331 1 Q
port 5 nsew default output
rlabel metal1 s 4145 875 4191 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3797 875 3843 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3378 875 3446 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2970 875 3038 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2161 875 2207 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1521 875 1567 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 661 875 707 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 875 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4145 790 4191 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3797 790 3843 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3378 790 3446 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2970 790 3038 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 661 790 707 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 790 319 875 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4145 775 4191 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3797 775 3843 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 661 775 707 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3797 703 3843 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 661 703 707 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 703 319 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3797 685 3843 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 245 687 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3389 233 3435 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1789 233 1835 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4161 90 4207 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3389 90 3435 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1789 90 1835 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4256 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 1008
string GDS_END 520620
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 511064
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
