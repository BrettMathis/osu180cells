magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3446 1094
<< pwell >>
rect -86 -86 3446 453
<< mvnmos >>
rect 124 97 244 333
rect 392 215 512 333
rect 560 215 680 333
rect 728 215 848 333
rect 952 215 1072 333
rect 1176 215 1296 333
rect 1400 215 1520 333
rect 1624 215 1744 333
rect 1992 215 2112 333
rect 2216 215 2336 333
rect 2440 215 2560 333
rect 2664 215 2784 333
rect 2832 215 2952 333
rect 3100 69 3220 333
<< mvpmos >>
rect 144 573 244 939
rect 412 594 512 792
rect 580 594 680 792
rect 748 594 848 792
rect 972 594 1072 792
rect 1196 594 1296 792
rect 1400 594 1500 792
rect 1604 594 1704 792
rect 2012 573 2112 771
rect 2216 573 2316 771
rect 2440 573 2540 771
rect 2664 573 2764 771
rect 2832 573 2932 771
rect 3100 573 3200 939
<< mvndiff >>
rect 36 320 124 333
rect 36 180 49 320
rect 95 180 124 320
rect 36 97 124 180
rect 244 250 392 333
rect 244 110 273 250
rect 319 215 392 250
rect 512 215 560 333
rect 680 215 728 333
rect 848 320 952 333
rect 848 274 877 320
rect 923 274 952 320
rect 848 215 952 274
rect 1072 320 1176 333
rect 1072 274 1101 320
rect 1147 274 1176 320
rect 1072 215 1176 274
rect 1296 274 1400 333
rect 1296 228 1325 274
rect 1371 228 1400 274
rect 1296 215 1400 228
rect 1520 320 1624 333
rect 1520 274 1549 320
rect 1595 274 1624 320
rect 1520 215 1624 274
rect 1744 274 1832 333
rect 1744 228 1773 274
rect 1819 228 1832 274
rect 1744 215 1832 228
rect 1904 320 1992 333
rect 1904 274 1917 320
rect 1963 274 1992 320
rect 1904 215 1992 274
rect 2112 274 2216 333
rect 2112 228 2141 274
rect 2187 228 2216 274
rect 2112 215 2216 228
rect 2336 308 2440 333
rect 2336 262 2365 308
rect 2411 262 2440 308
rect 2336 215 2440 262
rect 2560 320 2664 333
rect 2560 274 2589 320
rect 2635 274 2664 320
rect 2560 215 2664 274
rect 2784 215 2832 333
rect 2952 222 3100 333
rect 2952 215 3025 222
rect 319 110 332 215
rect 244 97 332 110
rect 3012 82 3025 215
rect 3071 82 3100 222
rect 3012 69 3100 82
rect 3220 320 3308 333
rect 3220 180 3249 320
rect 3295 180 3308 320
rect 3220 69 3308 180
<< mvpdiff >>
rect 56 726 144 939
rect 56 586 69 726
rect 115 586 144 726
rect 56 573 144 586
rect 244 926 332 939
rect 244 786 273 926
rect 319 792 332 926
rect 3012 926 3100 939
rect 319 786 412 792
rect 244 594 412 786
rect 512 594 580 792
rect 680 594 748 792
rect 848 747 972 792
rect 848 607 877 747
rect 923 607 972 747
rect 848 594 972 607
rect 1072 758 1196 792
rect 1072 618 1121 758
rect 1167 618 1196 758
rect 1072 594 1196 618
rect 1296 779 1400 792
rect 1296 733 1325 779
rect 1371 733 1400 779
rect 1296 594 1400 733
rect 1500 653 1604 792
rect 1500 607 1529 653
rect 1575 607 1604 653
rect 1500 594 1604 607
rect 1704 779 1792 792
rect 1704 639 1733 779
rect 1779 639 1792 779
rect 3012 786 3025 926
rect 3071 786 3100 926
rect 3012 771 3100 786
rect 1704 594 1792 639
rect 1924 758 2012 771
rect 1924 618 1937 758
rect 1983 618 2012 758
rect 244 573 324 594
rect 1924 573 2012 618
rect 2112 758 2216 771
rect 2112 712 2141 758
rect 2187 712 2216 758
rect 2112 573 2216 712
rect 2316 758 2440 771
rect 2316 618 2345 758
rect 2391 618 2440 758
rect 2316 573 2440 618
rect 2540 726 2664 771
rect 2540 586 2569 726
rect 2615 586 2664 726
rect 2540 573 2664 586
rect 2764 573 2832 771
rect 2932 573 3100 771
rect 3200 726 3288 939
rect 3200 586 3229 726
rect 3275 586 3288 726
rect 3200 573 3288 586
<< mvndiffc >>
rect 49 180 95 320
rect 273 110 319 250
rect 877 274 923 320
rect 1101 274 1147 320
rect 1325 228 1371 274
rect 1549 274 1595 320
rect 1773 228 1819 274
rect 1917 274 1963 320
rect 2141 228 2187 274
rect 2365 262 2411 308
rect 2589 274 2635 320
rect 3025 82 3071 222
rect 3249 180 3295 320
<< mvpdiffc >>
rect 69 586 115 726
rect 273 786 319 926
rect 877 607 923 747
rect 1121 618 1167 758
rect 1325 733 1371 779
rect 1529 607 1575 653
rect 1733 639 1779 779
rect 3025 786 3071 926
rect 1937 618 1983 758
rect 2141 712 2187 758
rect 2345 618 2391 758
rect 2569 586 2615 726
rect 3229 586 3275 726
<< polysilicon >>
rect 144 939 244 983
rect 3100 939 3200 983
rect 580 884 2764 924
rect 412 792 512 836
rect 580 792 680 884
rect 748 792 848 836
rect 972 792 1072 836
rect 1196 792 1296 836
rect 1400 792 1500 884
rect 1604 792 1704 836
rect 2012 771 2112 884
rect 2216 771 2316 815
rect 2440 771 2540 815
rect 2664 771 2764 884
rect 2832 771 2932 815
rect 144 412 244 573
rect 144 377 185 412
rect 124 366 185 377
rect 231 366 244 412
rect 412 523 512 594
rect 412 477 453 523
rect 499 477 512 523
rect 412 377 512 477
rect 580 377 680 594
rect 748 469 848 594
rect 748 423 789 469
rect 835 423 848 469
rect 748 377 848 423
rect 972 561 1072 594
rect 972 515 1013 561
rect 1059 515 1072 561
rect 972 377 1072 515
rect 1196 377 1296 594
rect 124 333 244 366
rect 392 333 512 377
rect 560 333 680 377
rect 728 333 848 377
rect 952 333 1072 377
rect 1176 333 1296 377
rect 1400 377 1500 594
rect 1604 469 1704 594
rect 1604 423 1617 469
rect 1663 423 1704 469
rect 1604 393 1704 423
rect 1400 333 1520 377
rect 1624 333 1744 393
rect 2012 377 2112 573
rect 1992 333 2112 377
rect 2216 377 2316 573
rect 2440 469 2540 573
rect 2440 423 2453 469
rect 2499 423 2540 469
rect 2440 377 2540 423
rect 2664 510 2764 573
rect 2664 464 2705 510
rect 2751 464 2764 510
rect 2664 377 2764 464
rect 2832 377 2932 573
rect 3100 412 3200 573
rect 2216 333 2336 377
rect 2440 333 2560 377
rect 2664 333 2784 377
rect 2832 333 2952 377
rect 3100 366 3113 412
rect 3159 377 3200 412
rect 3159 366 3220 377
rect 3100 333 3220 366
rect 392 123 512 215
rect 560 171 680 215
rect 728 171 848 215
rect 952 171 1072 215
rect 1176 123 1296 215
rect 1400 171 1520 215
rect 1624 171 1744 215
rect 1992 171 2112 215
rect 2216 123 2336 215
rect 2440 171 2560 215
rect 2664 171 2784 215
rect 2832 123 2952 215
rect 124 53 244 97
rect 392 83 2952 123
rect 3100 25 3220 69
<< polycontact >>
rect 185 366 231 412
rect 453 477 499 523
rect 789 423 835 469
rect 1013 515 1059 561
rect 1617 423 1663 469
rect 2453 423 2499 469
rect 2705 464 2751 510
rect 3113 366 3159 412
<< metal1 >>
rect 0 926 3360 1098
rect 0 918 273 926
rect 319 918 3025 926
rect 273 775 319 786
rect 1325 779 1371 918
rect 30 726 115 766
rect 1121 758 1167 769
rect 30 586 69 726
rect 877 747 923 758
rect 30 320 115 586
rect 361 607 877 634
rect 1325 722 1371 733
rect 1733 779 1779 918
rect 1167 618 1529 653
rect 1121 607 1529 618
rect 1575 607 1586 653
rect 1733 628 1779 639
rect 1937 758 1983 769
rect 2141 758 2187 918
rect 3071 918 3360 926
rect 3025 775 3071 786
rect 2141 701 2187 712
rect 2345 758 2391 769
rect 1983 618 2345 653
rect 1937 607 2391 618
rect 2569 726 2615 737
rect 361 588 923 607
rect 361 412 407 588
rect 3166 726 3295 737
rect 2615 588 2862 634
rect 2569 561 2615 586
rect 453 523 691 542
rect 499 477 691 523
rect 1002 515 1013 561
rect 1059 515 2615 561
rect 453 466 691 477
rect 2705 510 2770 542
rect 778 423 789 469
rect 835 423 1617 469
rect 1663 423 2453 469
rect 2499 423 2510 469
rect 2751 464 2770 510
rect 2705 453 2770 464
rect 2816 423 2862 588
rect 3166 586 3229 726
rect 3275 586 3295 726
rect 3166 578 3295 586
rect 174 366 185 412
rect 231 377 407 412
rect 231 366 923 377
rect 174 331 923 366
rect 30 180 49 320
rect 95 180 115 320
rect 877 320 923 331
rect 877 263 923 274
rect 1101 331 1595 377
rect 1101 320 1147 331
rect 1549 320 1595 331
rect 1101 263 1147 274
rect 1325 274 1371 285
rect 30 169 115 180
rect 273 250 319 261
rect 273 90 319 110
rect 1917 331 2336 377
rect 2382 354 2434 423
rect 2816 412 3159 423
rect 2816 401 3113 412
rect 2589 366 3113 401
rect 2589 355 3159 366
rect 1917 320 1963 331
rect 1549 263 1595 274
rect 1773 274 1819 285
rect 1325 90 1371 228
rect 2290 308 2336 331
rect 2589 320 2635 355
rect 1917 263 1963 274
rect 2141 274 2187 285
rect 1773 90 1819 228
rect 2290 262 2365 308
rect 2411 262 2422 308
rect 2589 263 2635 274
rect 3229 320 3295 578
rect 2141 90 2187 228
rect 3025 222 3071 233
rect 0 82 3025 90
rect 3229 180 3249 320
rect 3229 169 3295 180
rect 3071 82 3360 90
rect 0 -90 3360 82
<< labels >>
flabel metal1 s 453 466 691 542 0 FreeSans 200 0 0 0 A
port 1 nsew default input
flabel metal1 s 2705 453 2770 542 0 FreeSans 200 0 0 0 B
port 2 nsew default input
flabel metal1 s 778 423 2510 469 0 FreeSans 200 0 0 0 CI
port 3 nsew default input
flabel metal1 s 3166 578 3295 737 0 FreeSans 200 0 0 0 CO
port 4 nsew default output
flabel metal1 s 30 169 115 766 0 FreeSans 200 0 0 0 S
port 5 nsew default output
flabel metal1 s 0 918 3360 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2141 261 2187 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2382 354 2434 423 1 CI
port 3 nsew default input
rlabel metal1 s 3229 169 3295 578 1 CO
port 4 nsew default output
rlabel metal1 s 3025 775 3071 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2141 775 2187 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1733 775 1779 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1325 775 1371 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2141 722 2187 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1733 722 1779 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1325 722 1371 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2141 701 2187 722 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1733 701 1779 722 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1733 628 1779 701 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1773 261 1819 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1325 261 1371 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2141 233 2187 261 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1773 233 1819 261 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1325 233 1371 261 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 261 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3025 90 3071 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2141 90 2187 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1773 90 1819 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1325 90 1371 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3360 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 1008
string GDS_END 1065294
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1058206
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
