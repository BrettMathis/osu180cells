magic
tech gf180mcuB
magscale 1 5
timestamp 1669648930
<< checkpaint >>
rect 7600 7600 36500 36500
<< metal3 >>
rect 8600 23702 10100 35500
tri 10100 23702 10722 24324 sw
tri 8600 23454 8848 23702 ne
rect 8848 23454 10722 23702
tri 10722 23454 10970 23702 sw
tri 8848 21332 10970 23454 ne
tri 10970 21332 13092 23454 sw
tri 10970 19210 13092 21332 ne
tri 13092 19210 15214 21332 sw
tri 13092 17088 15214 19210 ne
tri 15214 17088 17336 19210 sw
tri 15214 14966 17336 17088 ne
tri 17336 14966 19458 17088 sw
tri 17336 12844 19458 14966 ne
tri 19458 12844 21580 14966 sw
tri 19458 10722 21580 12844 ne
tri 21580 10722 23702 12844 sw
tri 21580 8600 23702 10722 ne
tri 23702 10100 24324 10722 sw
rect 23702 8600 35500 10100
<< end >>
