magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 384
rect 224 0 344 384
rect 448 0 568 384
rect 672 0 792 384
rect 896 0 1016 384
rect 1120 0 1240 384
rect 1344 0 1464 384
rect 1568 0 1688 384
rect 1792 0 1912 384
rect 2016 0 2136 384
<< mvndiff >>
rect -88 371 0 384
rect -88 325 -75 371
rect -29 325 0 371
rect -88 267 0 325
rect -88 221 -75 267
rect -29 221 0 267
rect -88 163 0 221
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 371 224 384
rect 120 325 149 371
rect 195 325 224 371
rect 120 267 224 325
rect 120 221 149 267
rect 195 221 224 267
rect 120 163 224 221
rect 120 117 149 163
rect 195 117 224 163
rect 120 59 224 117
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 371 448 384
rect 344 325 373 371
rect 419 325 448 371
rect 344 267 448 325
rect 344 221 373 267
rect 419 221 448 267
rect 344 163 448 221
rect 344 117 373 163
rect 419 117 448 163
rect 344 59 448 117
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 371 672 384
rect 568 325 597 371
rect 643 325 672 371
rect 568 267 672 325
rect 568 221 597 267
rect 643 221 672 267
rect 568 163 672 221
rect 568 117 597 163
rect 643 117 672 163
rect 568 59 672 117
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 371 896 384
rect 792 325 821 371
rect 867 325 896 371
rect 792 267 896 325
rect 792 221 821 267
rect 867 221 896 267
rect 792 163 896 221
rect 792 117 821 163
rect 867 117 896 163
rect 792 59 896 117
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 371 1120 384
rect 1016 325 1045 371
rect 1091 325 1120 371
rect 1016 267 1120 325
rect 1016 221 1045 267
rect 1091 221 1120 267
rect 1016 163 1120 221
rect 1016 117 1045 163
rect 1091 117 1120 163
rect 1016 59 1120 117
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 371 1344 384
rect 1240 325 1269 371
rect 1315 325 1344 371
rect 1240 267 1344 325
rect 1240 221 1269 267
rect 1315 221 1344 267
rect 1240 163 1344 221
rect 1240 117 1269 163
rect 1315 117 1344 163
rect 1240 59 1344 117
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 371 1568 384
rect 1464 325 1493 371
rect 1539 325 1568 371
rect 1464 267 1568 325
rect 1464 221 1493 267
rect 1539 221 1568 267
rect 1464 163 1568 221
rect 1464 117 1493 163
rect 1539 117 1568 163
rect 1464 59 1568 117
rect 1464 13 1493 59
rect 1539 13 1568 59
rect 1464 0 1568 13
rect 1688 371 1792 384
rect 1688 325 1717 371
rect 1763 325 1792 371
rect 1688 267 1792 325
rect 1688 221 1717 267
rect 1763 221 1792 267
rect 1688 163 1792 221
rect 1688 117 1717 163
rect 1763 117 1792 163
rect 1688 59 1792 117
rect 1688 13 1717 59
rect 1763 13 1792 59
rect 1688 0 1792 13
rect 1912 371 2016 384
rect 1912 325 1941 371
rect 1987 325 2016 371
rect 1912 267 2016 325
rect 1912 221 1941 267
rect 1987 221 2016 267
rect 1912 163 2016 221
rect 1912 117 1941 163
rect 1987 117 2016 163
rect 1912 59 2016 117
rect 1912 13 1941 59
rect 1987 13 2016 59
rect 1912 0 2016 13
rect 2136 371 2224 384
rect 2136 325 2165 371
rect 2211 325 2224 371
rect 2136 267 2224 325
rect 2136 221 2165 267
rect 2211 221 2224 267
rect 2136 163 2224 221
rect 2136 117 2165 163
rect 2211 117 2224 163
rect 2136 59 2224 117
rect 2136 13 2165 59
rect 2211 13 2224 59
rect 2136 0 2224 13
<< mvndiffc >>
rect -75 325 -29 371
rect -75 221 -29 267
rect -75 117 -29 163
rect -75 13 -29 59
rect 149 325 195 371
rect 149 221 195 267
rect 149 117 195 163
rect 149 13 195 59
rect 373 325 419 371
rect 373 221 419 267
rect 373 117 419 163
rect 373 13 419 59
rect 597 325 643 371
rect 597 221 643 267
rect 597 117 643 163
rect 597 13 643 59
rect 821 325 867 371
rect 821 221 867 267
rect 821 117 867 163
rect 821 13 867 59
rect 1045 325 1091 371
rect 1045 221 1091 267
rect 1045 117 1091 163
rect 1045 13 1091 59
rect 1269 325 1315 371
rect 1269 221 1315 267
rect 1269 117 1315 163
rect 1269 13 1315 59
rect 1493 325 1539 371
rect 1493 221 1539 267
rect 1493 117 1539 163
rect 1493 13 1539 59
rect 1717 325 1763 371
rect 1717 221 1763 267
rect 1717 117 1763 163
rect 1717 13 1763 59
rect 1941 325 1987 371
rect 1941 221 1987 267
rect 1941 117 1987 163
rect 1941 13 1987 59
rect 2165 325 2211 371
rect 2165 221 2211 267
rect 2165 117 2211 163
rect 2165 13 2211 59
<< polysilicon >>
rect 0 384 120 428
rect 224 384 344 428
rect 448 384 568 428
rect 672 384 792 428
rect 896 384 1016 428
rect 1120 384 1240 428
rect 1344 384 1464 428
rect 1568 384 1688 428
rect 1792 384 1912 428
rect 2016 384 2136 428
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
<< metal1 >>
rect -75 371 -29 384
rect -75 267 -29 325
rect -75 163 -29 221
rect -75 59 -29 117
rect -75 0 -29 13
rect 149 371 195 384
rect 149 267 195 325
rect 149 163 195 221
rect 149 59 195 117
rect 149 0 195 13
rect 373 371 419 384
rect 373 267 419 325
rect 373 163 419 221
rect 373 59 419 117
rect 373 0 419 13
rect 597 371 643 384
rect 597 267 643 325
rect 597 163 643 221
rect 597 59 643 117
rect 597 0 643 13
rect 821 371 867 384
rect 821 267 867 325
rect 821 163 867 221
rect 821 59 867 117
rect 821 0 867 13
rect 1045 371 1091 384
rect 1045 267 1091 325
rect 1045 163 1091 221
rect 1045 59 1091 117
rect 1045 0 1091 13
rect 1269 371 1315 384
rect 1269 267 1315 325
rect 1269 163 1315 221
rect 1269 59 1315 117
rect 1269 0 1315 13
rect 1493 371 1539 384
rect 1493 267 1539 325
rect 1493 163 1539 221
rect 1493 59 1539 117
rect 1493 0 1539 13
rect 1717 371 1763 384
rect 1717 267 1763 325
rect 1717 163 1763 221
rect 1717 59 1763 117
rect 1717 0 1763 13
rect 1941 371 1987 384
rect 1941 267 1987 325
rect 1941 163 1987 221
rect 1941 59 1987 117
rect 1941 0 1987 13
rect 2165 371 2211 384
rect 2165 267 2211 325
rect 2165 163 2211 221
rect 2165 59 2211 117
rect 2165 0 2211 13
<< labels >>
flabel metal1 s -52 192 -52 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 2188 192 2188 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 192 172 192 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 192 396 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 192 620 192 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 192 844 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 192 1068 192 0 FreeSans 200 0 0 0 D
flabel metal1 s 1292 192 1292 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 1516 192 1516 192 0 FreeSans 200 0 0 0 D
flabel metal1 s 1740 192 1740 192 0 FreeSans 200 0 0 0 S
flabel metal1 s 1964 192 1964 192 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 386676
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 379526
<< end >>
