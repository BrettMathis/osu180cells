magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 1280 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 490 190 550 360
rect 720 190 780 360
rect 850 190 910 360
rect 1020 190 1080 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 490 700 550 1040
rect 720 700 780 1040
rect 850 700 910 1040
rect 1020 700 1080 1040
<< ndiff >>
rect 580 360 680 370
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 490 360
rect 550 350 720 360
rect 550 210 612 350
rect 658 210 720 350
rect 550 190 720 210
rect 780 190 850 360
rect 910 298 1020 360
rect 910 252 942 298
rect 988 252 1020 298
rect 910 190 1020 252
rect 1080 298 1180 360
rect 1080 252 1112 298
rect 1158 252 1180 298
rect 1080 190 1180 252
<< pdiff >>
rect 90 1003 190 1040
rect 90 957 112 1003
rect 158 957 190 1003
rect 90 700 190 957
rect 250 1003 360 1040
rect 250 957 282 1003
rect 328 957 360 1003
rect 250 700 360 957
rect 420 700 490 1040
rect 550 1003 720 1040
rect 550 957 612 1003
rect 658 957 720 1003
rect 550 700 720 957
rect 780 700 850 1040
rect 910 1003 1020 1040
rect 910 957 942 1003
rect 988 957 1020 1003
rect 910 700 1020 957
rect 1080 1003 1180 1040
rect 1080 957 1112 1003
rect 1158 957 1180 1003
rect 1080 700 1180 957
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 612 210 658 350
rect 942 252 988 298
rect 1112 252 1158 298
<< pdiffc >>
rect 112 957 158 1003
rect 282 957 328 1003
rect 612 957 658 1003
rect 942 957 988 1003
rect 1112 957 1158 1003
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 490 1040 550 1090
rect 720 1040 780 1090
rect 850 1040 910 1090
rect 1020 1040 1080 1090
rect 190 520 250 700
rect 360 680 420 700
rect 310 653 420 680
rect 310 607 337 653
rect 383 607 420 653
rect 310 580 420 607
rect 490 680 550 700
rect 720 680 780 700
rect 850 680 910 700
rect 1020 680 1080 700
rect 490 653 630 680
rect 490 607 557 653
rect 603 607 630 653
rect 490 580 630 607
rect 700 653 800 680
rect 700 607 727 653
rect 773 607 800 653
rect 850 630 1080 680
rect 700 580 800 607
rect 190 493 350 520
rect 190 447 277 493
rect 323 490 350 493
rect 323 447 420 490
rect 190 420 420 447
rect 190 360 250 420
rect 360 360 420 420
rect 490 360 550 580
rect 1020 520 1080 630
rect 600 500 700 520
rect 600 493 780 500
rect 600 447 627 493
rect 673 447 780 493
rect 910 493 1080 520
rect 910 470 937 493
rect 600 420 780 447
rect 720 360 780 420
rect 850 447 937 470
rect 983 447 1080 493
rect 850 420 1080 447
rect 850 360 910 420
rect 1020 360 1080 420
rect 190 140 250 190
rect 360 140 420 190
rect 490 140 550 190
rect 720 140 780 190
rect 850 140 910 190
rect 1020 140 1080 190
<< polycontact >>
rect 337 607 383 653
rect 557 607 603 653
rect 727 607 773 653
rect 277 447 323 493
rect 627 447 673 493
rect 937 447 983 493
<< metal1 >>
rect 0 1178 1280 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1280 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1280 1176
rect 0 1110 1280 1124
rect 110 1003 160 1040
rect 110 957 112 1003
rect 158 957 160 1003
rect 110 660 160 957
rect 280 1003 330 1110
rect 280 957 282 1003
rect 328 957 330 1003
rect 280 920 330 957
rect 610 1003 660 1040
rect 610 957 612 1003
rect 658 957 660 1003
rect 610 950 660 957
rect 600 886 660 950
rect 940 1003 990 1110
rect 940 957 942 1003
rect 988 957 990 1003
rect 940 920 990 957
rect 1110 1003 1160 1040
rect 1110 957 1112 1003
rect 1158 957 1160 1003
rect 600 834 604 886
rect 656 834 660 886
rect 600 810 660 834
rect 1110 760 1160 957
rect 550 710 1160 760
rect 110 653 480 660
rect 110 607 337 653
rect 383 607 480 653
rect 110 600 480 607
rect 110 298 160 600
rect 420 500 480 600
rect 550 653 610 710
rect 550 607 557 653
rect 603 607 610 653
rect 550 580 610 607
rect 700 656 800 660
rect 700 604 724 656
rect 776 604 800 656
rect 700 600 800 604
rect 250 496 350 500
rect 250 444 274 496
rect 326 444 350 496
rect 250 440 350 444
rect 420 493 700 500
rect 420 447 627 493
rect 673 447 700 493
rect 420 440 700 447
rect 910 496 1010 500
rect 910 444 934 496
rect 986 444 1010 496
rect 910 440 1010 444
rect 600 366 660 390
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 280 252 282 298
rect 328 252 330 298
rect 600 314 604 366
rect 656 350 660 366
rect 600 280 612 314
rect 280 120 330 252
rect 610 210 612 280
rect 658 210 660 350
rect 610 190 660 210
rect 940 298 990 360
rect 940 252 942 298
rect 988 252 990 298
rect 940 120 990 252
rect 1110 298 1160 710
rect 1110 252 1112 298
rect 1158 252 1160 298
rect 1110 190 1160 252
rect 0 106 1280 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1280 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1280 54
rect 0 0 1280 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 604 834 656 886
rect 724 653 776 656
rect 724 607 727 653
rect 727 607 773 653
rect 773 607 776 653
rect 724 604 776 607
rect 274 493 326 496
rect 274 447 277 493
rect 277 447 323 493
rect 323 447 326 493
rect 274 444 326 447
rect 934 493 986 496
rect 934 447 937 493
rect 937 447 983 493
rect 983 447 986 493
rect 934 444 986 447
rect 604 350 656 366
rect 604 314 612 350
rect 612 314 656 350
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 600 900 660 950
rect 590 886 670 900
rect 590 834 604 886
rect 656 834 670 886
rect 590 820 670 834
rect 590 810 660 820
rect 270 510 330 520
rect 260 496 340 510
rect 260 444 274 496
rect 326 444 340 496
rect 260 430 340 444
rect 270 240 330 430
rect 590 380 650 810
rect 720 670 790 680
rect 710 656 800 670
rect 710 604 724 656
rect 776 604 800 656
rect 710 590 800 604
rect 720 580 800 590
rect 580 366 680 380
rect 580 314 604 366
rect 656 314 680 366
rect 580 300 680 314
rect 740 240 800 580
rect 930 510 990 520
rect 920 500 1000 510
rect 910 496 1010 500
rect 910 444 934 496
rect 986 444 1010 496
rect 910 440 1010 444
rect 920 430 1000 440
rect 930 420 990 430
rect 270 180 800 240
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 270 180 330 520 4 A
port 1 nsew signal input
rlabel metal2 s 590 300 650 900 4 Y
port 2 nsew signal output
rlabel metal2 s 930 420 990 520 4 B
port 3 nsew signal input
rlabel metal2 s 260 430 340 510 1 A
port 1 nsew signal input
rlabel metal2 s 270 180 800 240 1 A
port 1 nsew signal input
rlabel metal2 s 720 580 790 680 1 A
port 1 nsew signal input
rlabel metal2 s 740 180 800 670 1 A
port 1 nsew signal input
rlabel metal2 s 710 590 800 670 1 A
port 1 nsew signal input
rlabel metal1 s 250 440 350 500 1 A
port 1 nsew signal input
rlabel metal1 s 700 600 800 660 1 A
port 1 nsew signal input
rlabel metal2 s 920 430 1000 510 1 B
port 3 nsew signal input
rlabel metal2 s 910 440 1010 500 1 B
port 3 nsew signal input
rlabel metal1 s 910 440 1010 500 1 B
port 3 nsew signal input
rlabel metal2 s 90 1120 190 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 280 920 330 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 940 920 990 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1110 1280 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 280 0 330 360 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 940 0 990 360 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 0 1280 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 600 810 660 950 1 Y
port 2 nsew signal output
rlabel metal2 s 590 820 670 900 1 Y
port 2 nsew signal output
rlabel metal2 s 580 300 680 380 1 Y
port 2 nsew signal output
rlabel metal1 s 600 810 660 950 1 Y
port 2 nsew signal output
rlabel metal1 s 610 810 660 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 610 190 660 390 1 Y
port 2 nsew signal output
rlabel metal1 s 600 280 660 390 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1280 1230
string GDS_END 456236
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 445158
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
