magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 147 44 159
rect 11 106 16 147
rect 11 93 21 99
rect 28 73 33 140
rect 26 67 36 73
rect 11 9 16 33
rect 28 16 33 67
rect 0 -3 44 9
<< metal2 >>
rect 10 154 18 155
rect 9 148 19 154
rect 10 147 18 148
rect 11 92 21 100
rect 26 66 36 74
rect 10 8 18 9
rect 9 2 19 8
rect 10 1 18 2
<< labels >>
rlabel metal2 s 11 92 21 100 6 A
port 1 nsew signal input
rlabel metal1 s 11 93 21 99 6 A
port 1 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 147 44 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 -3 44 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 26 66 36 74 6 Y
port 2 nsew signal output
rlabel metal1 s 28 16 33 140 6 Y
port 2 nsew signal output
rlabel metal1 s 26 67 36 73 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 44 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 346036
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 342804
<< end >>
