magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 3446 870
rect -86 352 1453 377
rect 2924 352 3446 377
<< pwell >>
rect 1453 352 2924 377
rect -86 -86 3446 352
<< mvnmos >>
rect 150 124 270 217
rect 374 124 494 217
rect 742 156 862 228
rect 966 156 1086 228
rect 1190 156 1310 228
rect 1358 156 1478 228
rect 1670 185 1790 257
rect 1894 185 2014 257
rect 2118 185 2238 257
rect 2406 131 2526 257
rect 2642 131 2762 257
rect 3075 68 3195 232
<< mvpmos >>
rect 170 472 270 645
rect 374 472 474 645
rect 766 500 866 599
rect 970 500 1070 599
rect 1201 500 1301 599
rect 1378 500 1478 599
rect 1670 500 1770 599
rect 1893 500 1993 599
rect 2204 500 2304 599
rect 2452 500 2552 715
rect 2656 500 2756 715
rect 3075 490 3175 716
<< mvndiff >>
rect 1538 228 1670 257
rect 62 204 150 217
rect 62 158 75 204
rect 121 158 150 204
rect 62 124 150 158
rect 270 183 374 217
rect 270 137 299 183
rect 345 137 374 183
rect 270 124 374 137
rect 494 204 582 217
rect 494 158 523 204
rect 569 158 582 204
rect 494 124 582 158
rect 654 215 742 228
rect 654 169 667 215
rect 713 169 742 215
rect 654 156 742 169
rect 862 215 966 228
rect 862 169 891 215
rect 937 169 966 215
rect 862 156 966 169
rect 1086 215 1190 228
rect 1086 169 1115 215
rect 1161 169 1190 215
rect 1086 156 1190 169
rect 1310 156 1358 228
rect 1478 185 1670 228
rect 1790 244 1894 257
rect 1790 198 1819 244
rect 1865 198 1894 244
rect 1790 185 1894 198
rect 2014 244 2118 257
rect 2014 198 2043 244
rect 2089 198 2118 244
rect 2014 185 2118 198
rect 2238 244 2406 257
rect 2238 198 2331 244
rect 2377 198 2406 244
rect 2238 185 2406 198
rect 1478 162 1610 185
rect 1478 156 1551 162
rect 1538 116 1551 156
rect 1597 116 1610 162
rect 1538 103 1610 116
rect 2318 131 2406 185
rect 2526 190 2642 257
rect 2526 144 2555 190
rect 2601 144 2642 190
rect 2526 131 2642 144
rect 2762 244 2850 257
rect 2762 198 2791 244
rect 2837 198 2850 244
rect 2762 131 2850 198
rect 2987 127 3075 232
rect 2987 81 3000 127
rect 3046 81 3075 127
rect 2987 68 3075 81
rect 3195 219 3283 232
rect 3195 173 3224 219
rect 3270 173 3283 219
rect 3195 68 3283 173
<< mvpdiff >>
rect 634 647 706 660
rect 82 632 170 645
rect 82 492 95 632
rect 141 492 170 632
rect 82 472 170 492
rect 270 632 374 645
rect 270 586 299 632
rect 345 586 374 632
rect 270 472 374 586
rect 474 632 562 645
rect 474 492 503 632
rect 549 492 562 632
rect 634 601 647 647
rect 693 601 706 647
rect 634 599 706 601
rect 2364 609 2452 715
rect 2364 599 2377 609
rect 634 500 766 599
rect 866 575 970 599
rect 866 529 895 575
rect 941 529 970 575
rect 866 500 970 529
rect 1070 559 1201 599
rect 1070 513 1126 559
rect 1172 513 1201 559
rect 1070 500 1201 513
rect 1301 500 1378 599
rect 1478 586 1670 599
rect 1478 540 1552 586
rect 1598 540 1670 586
rect 1478 500 1670 540
rect 1770 575 1893 599
rect 1770 529 1818 575
rect 1864 529 1893 575
rect 1770 500 1893 529
rect 1993 575 2204 599
rect 1993 529 2043 575
rect 2089 529 2204 575
rect 1993 500 2204 529
rect 2304 563 2377 599
rect 2423 563 2452 609
rect 2304 500 2452 563
rect 2552 702 2656 715
rect 2552 656 2581 702
rect 2627 656 2656 702
rect 2552 500 2656 656
rect 2756 559 2844 715
rect 2756 513 2785 559
rect 2831 513 2844 559
rect 2756 500 2844 513
rect 2967 703 3075 716
rect 2967 657 2980 703
rect 3026 657 3075 703
rect 2967 597 3075 657
rect 2967 551 2980 597
rect 3026 551 3075 597
rect 474 472 562 492
rect 2967 490 3075 551
rect 3175 585 3263 716
rect 3175 539 3204 585
rect 3250 539 3263 585
rect 3175 490 3263 539
<< mvndiffc >>
rect 75 158 121 204
rect 299 137 345 183
rect 523 158 569 204
rect 667 169 713 215
rect 891 169 937 215
rect 1115 169 1161 215
rect 1819 198 1865 244
rect 2043 198 2089 244
rect 2331 198 2377 244
rect 1551 116 1597 162
rect 2555 144 2601 190
rect 2791 198 2837 244
rect 3000 81 3046 127
rect 3224 173 3270 219
<< mvpdiffc >>
rect 95 492 141 632
rect 299 586 345 632
rect 503 492 549 632
rect 647 601 693 647
rect 895 529 941 575
rect 1126 513 1172 559
rect 1552 540 1598 586
rect 1818 529 1864 575
rect 2043 529 2089 575
rect 2377 563 2423 609
rect 2581 656 2627 702
rect 2785 513 2831 559
rect 2980 657 3026 703
rect 2980 551 3026 597
rect 3204 539 3250 585
<< polysilicon >>
rect 374 720 1070 760
rect 170 645 270 690
rect 374 645 474 720
rect 766 599 866 643
rect 970 599 1070 720
rect 1201 720 1993 760
rect 1201 678 1301 720
rect 1201 632 1214 678
rect 1260 632 1301 678
rect 1201 599 1301 632
rect 1378 599 1478 643
rect 1670 599 1770 643
rect 1893 599 1993 720
rect 2452 715 2552 760
rect 2656 715 2756 760
rect 3075 716 3175 760
rect 2204 599 2304 643
rect 170 412 270 472
rect 170 366 183 412
rect 229 366 270 412
rect 170 261 270 366
rect 150 217 270 261
rect 374 326 474 472
rect 374 280 387 326
rect 433 280 474 326
rect 374 261 474 280
rect 766 415 866 500
rect 970 456 1070 500
rect 766 369 807 415
rect 853 369 866 415
rect 1201 408 1301 500
rect 766 288 866 369
rect 966 368 1301 408
rect 1378 467 1478 500
rect 1378 421 1419 467
rect 1465 421 1478 467
rect 766 272 862 288
rect 374 217 494 261
rect 742 228 862 272
rect 966 228 1086 368
rect 1190 307 1310 320
rect 1190 261 1218 307
rect 1264 261 1310 307
rect 1378 272 1478 421
rect 1190 228 1310 261
rect 1358 228 1478 272
rect 1670 346 1770 500
rect 1893 399 1993 500
rect 2204 456 2304 500
rect 2226 408 2304 456
rect 2452 440 2552 500
rect 1893 359 2158 399
rect 1670 300 1683 346
rect 1729 301 1770 346
rect 2118 301 2158 359
rect 2226 362 2239 408
rect 2285 362 2304 408
rect 2226 349 2304 362
rect 2406 400 2552 440
rect 2656 467 2756 500
rect 2656 421 2669 467
rect 2715 421 2756 467
rect 2406 375 2526 400
rect 2656 399 2756 421
rect 2406 329 2446 375
rect 2492 329 2526 375
rect 1729 300 1790 301
rect 1670 257 1790 300
rect 1894 257 2014 301
rect 2118 257 2238 301
rect 2406 257 2526 329
rect 2642 319 2756 399
rect 3075 370 3175 490
rect 2941 357 3175 370
rect 2642 257 2762 319
rect 2941 311 2954 357
rect 3000 344 3175 357
rect 3000 311 3195 344
rect 2941 298 3195 311
rect 150 80 270 124
rect 374 64 494 124
rect 742 112 862 156
rect 966 112 1086 156
rect 1190 64 1310 156
rect 1358 112 1478 156
rect 1670 141 1790 185
rect 1894 152 2014 185
rect 1894 106 1907 152
rect 1953 106 2014 152
rect 2118 141 2238 185
rect 3075 232 3195 298
rect 1894 93 2014 106
rect 374 24 1310 64
rect 2406 24 2526 131
rect 2642 24 2762 131
rect 3075 24 3195 68
<< polycontact >>
rect 1214 632 1260 678
rect 183 366 229 412
rect 387 280 433 326
rect 807 369 853 415
rect 1419 421 1465 467
rect 1218 261 1264 307
rect 1683 300 1729 346
rect 2239 362 2285 408
rect 2669 421 2715 467
rect 2446 329 2492 375
rect 2954 311 3000 357
rect 1907 106 1953 152
<< metal1 >>
rect 0 724 3360 844
rect 95 632 141 645
rect 288 632 356 724
rect 636 647 704 724
rect 288 586 299 632
rect 345 586 356 632
rect 503 632 569 645
rect 141 492 433 518
rect 95 472 433 492
rect 56 412 318 426
rect 56 366 183 412
rect 229 366 318 412
rect 56 354 318 366
rect 387 326 433 472
rect 387 275 433 280
rect 75 229 433 275
rect 549 542 569 632
rect 636 601 647 647
rect 693 601 704 647
rect 766 632 1214 678
rect 1260 632 1271 678
rect 766 542 812 632
rect 1541 586 1609 724
rect 2570 702 2638 724
rect 2570 656 2581 702
rect 2627 656 2638 702
rect 2969 703 3037 724
rect 2686 620 2923 666
rect 2686 610 2732 620
rect 2358 609 2732 610
rect 549 496 812 542
rect 884 529 895 575
rect 941 529 1058 575
rect 549 492 569 496
rect 75 204 121 229
rect 503 204 569 492
rect 690 415 878 430
rect 690 369 807 415
rect 853 369 878 415
rect 690 354 878 369
rect 1011 215 1058 529
rect 75 147 121 158
rect 288 137 299 183
rect 345 137 356 183
rect 503 158 523 204
rect 503 147 569 158
rect 656 169 667 215
rect 713 169 724 215
rect 880 169 891 215
rect 937 169 1058 215
rect 1115 513 1126 559
rect 1172 513 1183 559
rect 1541 540 1552 586
rect 1598 540 1609 586
rect 1808 575 1876 586
rect 1115 410 1183 513
rect 1808 529 1818 575
rect 1864 529 1876 575
rect 1808 478 1876 529
rect 1419 467 1876 478
rect 1465 421 1876 467
rect 1419 410 1876 421
rect 1115 364 1356 410
rect 1115 215 1161 364
rect 1310 346 1356 364
rect 1218 307 1264 318
rect 1310 300 1683 346
rect 1729 300 1740 346
rect 1218 254 1264 261
rect 1218 208 1712 254
rect 288 60 356 137
rect 656 60 724 169
rect 1115 158 1161 169
rect 1540 116 1551 162
rect 1597 116 1608 162
rect 1540 60 1608 116
rect 1666 152 1712 208
rect 1808 244 1876 410
rect 1808 198 1819 244
rect 1865 198 1876 244
rect 2032 575 2100 586
rect 2032 529 2043 575
rect 2089 529 2100 575
rect 2358 563 2377 609
rect 2423 563 2732 609
rect 2032 517 2100 529
rect 2785 559 2831 570
rect 2032 471 2726 517
rect 2032 244 2100 471
rect 2658 467 2726 471
rect 2658 421 2669 467
rect 2715 421 2726 467
rect 2032 198 2043 244
rect 2089 198 2100 244
rect 2239 408 2285 419
rect 2785 377 2831 513
rect 2877 469 2923 620
rect 2969 657 2980 703
rect 3026 657 3037 703
rect 2969 597 3037 657
rect 2969 551 2980 597
rect 3026 551 3037 597
rect 3154 585 3270 597
rect 3154 539 3204 585
rect 3250 539 3270 585
rect 2877 423 3092 469
rect 2785 375 3000 377
rect 2239 152 2285 362
rect 2435 329 2446 375
rect 2492 357 3000 375
rect 2492 329 2954 357
rect 2435 328 2954 329
rect 2780 311 2954 328
rect 2780 300 3000 311
rect 2331 244 2704 282
rect 2377 236 2704 244
rect 2331 178 2377 198
rect 1666 106 1907 152
rect 1953 106 2285 152
rect 2544 144 2555 190
rect 2601 144 2612 190
rect 2544 60 2612 144
rect 2658 152 2704 236
rect 2780 244 2848 300
rect 2780 198 2791 244
rect 2837 198 2848 244
rect 3046 230 3092 423
rect 2908 184 3092 230
rect 3154 219 3270 539
rect 2908 152 2954 184
rect 3154 173 3224 219
rect 3154 162 3270 173
rect 2658 106 2954 152
rect 3000 127 3046 138
rect 3000 60 3046 81
rect 0 -60 3360 60
<< labels >>
flabel metal1 s 56 354 318 426 0 FreeSans 600 0 0 0 CLKN
port 2 nsew clock input
flabel metal1 s 0 724 3360 844 0 FreeSans 600 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 656 190 724 215 0 FreeSans 600 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 690 354 878 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 3154 162 3270 597 0 FreeSans 600 0 0 0 Q
port 3 nsew default output
rlabel metal1 s 2969 656 3037 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2570 656 2638 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 656 1609 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 656 704 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 656 356 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 601 3037 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 601 1609 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 636 601 704 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 601 356 656 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 586 3037 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 586 1609 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 288 586 356 601 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2969 551 3037 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 551 1609 586 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 540 1609 551 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2544 183 2612 190 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 183 724 190 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 162 2612 183 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 162 724 183 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 162 356 183 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 138 2612 162 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1540 138 1608 162 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 138 724 162 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 138 356 162 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3000 60 3046 138 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2544 60 2612 138 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1540 60 1608 138 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 656 60 724 138 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 288 60 356 138 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3360 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 784
string GDS_END 848142
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 840762
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
