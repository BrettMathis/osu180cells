magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 2550 870
rect -86 352 931 377
rect 1151 352 2550 377
<< pwell >>
rect 931 352 1151 377
rect -86 -86 2550 352
<< mvnmos >>
rect 157 93 277 165
rect 341 93 461 165
rect 601 68 721 232
rect 825 68 945 232
rect 1137 68 1257 232
rect 1505 68 1625 232
rect 1729 68 1849 232
rect 1953 68 2073 232
rect 2177 68 2297 232
<< mvpmos >>
rect 157 543 257 620
rect 361 543 461 620
rect 621 497 721 716
rect 845 497 945 716
rect 1137 497 1237 716
rect 1525 472 1625 716
rect 1739 472 1839 716
rect 1963 472 2063 716
rect 2177 472 2277 716
<< mvndiff >>
rect 1005 244 1077 257
rect 1005 232 1018 244
rect 521 165 601 232
rect 69 152 157 165
rect 69 106 82 152
rect 128 106 157 152
rect 69 93 157 106
rect 277 93 341 165
rect 461 152 601 165
rect 461 106 526 152
rect 572 106 601 152
rect 461 93 601 106
rect 521 68 601 93
rect 721 152 825 232
rect 721 106 750 152
rect 796 106 825 152
rect 721 68 825 106
rect 945 198 1018 232
rect 1064 232 1077 244
rect 1064 198 1137 232
rect 945 68 1137 198
rect 1257 152 1345 232
rect 1257 106 1286 152
rect 1332 106 1345 152
rect 1257 68 1345 106
rect 1417 142 1505 232
rect 1417 96 1430 142
rect 1476 96 1505 142
rect 1417 68 1505 96
rect 1625 218 1729 232
rect 1625 172 1654 218
rect 1700 172 1729 218
rect 1625 68 1729 172
rect 1849 171 1953 232
rect 1849 125 1878 171
rect 1924 125 1953 171
rect 1849 68 1953 125
rect 2073 218 2177 232
rect 2073 172 2102 218
rect 2148 172 2177 218
rect 2073 68 2177 172
rect 2297 176 2385 232
rect 2297 130 2326 176
rect 2372 130 2385 176
rect 2297 68 2385 130
<< mvpdiff >>
rect 541 620 621 716
rect 69 605 157 620
rect 69 559 82 605
rect 128 559 157 605
rect 69 543 157 559
rect 257 603 361 620
rect 257 557 286 603
rect 332 557 361 603
rect 257 543 361 557
rect 461 603 621 620
rect 461 557 490 603
rect 536 557 621 603
rect 461 543 621 557
rect 541 497 621 543
rect 721 639 845 716
rect 721 593 760 639
rect 806 593 845 639
rect 721 497 845 593
rect 945 497 1137 716
rect 1237 703 1325 716
rect 1237 563 1266 703
rect 1312 563 1325 703
rect 1237 497 1325 563
rect 1437 665 1525 716
rect 1437 525 1450 665
rect 1496 525 1525 665
rect 1437 472 1525 525
rect 1625 665 1739 716
rect 1625 525 1654 665
rect 1700 525 1739 665
rect 1625 472 1739 525
rect 1839 665 1963 716
rect 1839 619 1868 665
rect 1914 619 1963 665
rect 1839 472 1963 619
rect 2063 665 2177 716
rect 2063 525 2092 665
rect 2138 525 2177 665
rect 2063 472 2177 525
rect 2277 665 2365 716
rect 2277 619 2306 665
rect 2352 619 2365 665
rect 2277 472 2365 619
<< mvndiffc >>
rect 82 106 128 152
rect 526 106 572 152
rect 750 106 796 152
rect 1018 198 1064 244
rect 1286 106 1332 152
rect 1430 96 1476 142
rect 1654 172 1700 218
rect 1878 125 1924 171
rect 2102 172 2148 218
rect 2326 130 2372 176
<< mvpdiffc >>
rect 82 559 128 605
rect 286 557 332 603
rect 490 557 536 603
rect 760 593 806 639
rect 1266 563 1312 703
rect 1450 525 1496 665
rect 1654 525 1700 665
rect 1868 619 1914 665
rect 2092 525 2138 665
rect 2306 619 2352 665
<< polysilicon >>
rect 621 716 721 760
rect 845 716 945 760
rect 1137 716 1237 760
rect 1525 716 1625 760
rect 1739 716 1839 760
rect 1963 716 2063 760
rect 2177 716 2277 760
rect 157 620 257 684
rect 361 620 461 684
rect 157 416 257 543
rect 157 370 190 416
rect 236 370 257 416
rect 157 209 257 370
rect 361 416 461 543
rect 361 370 399 416
rect 445 370 461 416
rect 621 381 721 497
rect 845 381 945 497
rect 361 209 461 370
rect 601 311 721 381
rect 601 265 645 311
rect 691 265 721 311
rect 601 232 721 265
rect 825 344 945 381
rect 825 298 848 344
rect 894 298 945 344
rect 825 232 945 298
rect 1137 415 1237 497
rect 1137 369 1165 415
rect 1211 369 1237 415
rect 1137 276 1237 369
rect 1525 415 1625 472
rect 1525 369 1551 415
rect 1597 369 1625 415
rect 1525 357 1625 369
rect 1739 415 1839 472
rect 1739 369 1767 415
rect 1813 369 1839 415
rect 1739 357 1839 369
rect 1963 415 2063 472
rect 1963 369 1990 415
rect 2036 369 2063 415
rect 1963 357 2063 369
rect 2177 415 2277 472
rect 2177 369 2196 415
rect 2242 369 2277 415
rect 2177 357 2277 369
rect 1525 311 2277 357
rect 1525 288 1625 311
rect 157 165 277 209
rect 341 165 461 209
rect 157 49 277 93
rect 341 49 461 93
rect 1137 232 1257 276
rect 1505 232 1625 288
rect 1729 232 1849 311
rect 1953 232 2073 311
rect 2177 288 2277 311
rect 2177 232 2297 288
rect 601 24 721 68
rect 825 24 945 68
rect 1137 24 1257 68
rect 1505 24 1625 68
rect 1729 24 1849 68
rect 1953 24 2073 68
rect 2177 24 2297 68
<< polycontact >>
rect 190 370 236 416
rect 399 370 445 416
rect 645 265 691 311
rect 848 298 894 344
rect 1165 369 1211 415
rect 1551 369 1597 415
rect 1767 369 1813 415
rect 1990 369 2036 415
rect 2196 369 2242 415
<< metal1 >>
rect 0 724 2464 844
rect 71 605 139 724
rect 71 559 82 605
rect 128 559 139 605
rect 479 603 547 724
rect 1255 703 1323 724
rect 186 557 286 603
rect 332 557 361 603
rect 479 557 490 603
rect 536 557 547 603
rect 732 593 760 639
rect 806 593 1136 639
rect 186 513 238 557
rect 71 466 238 513
rect 600 511 1005 536
rect 71 244 117 466
rect 285 465 1005 511
rect 1090 517 1136 593
rect 1255 563 1266 703
rect 1312 563 1323 703
rect 1450 665 1496 724
rect 1090 470 1345 517
rect 1450 506 1496 525
rect 1654 665 1700 676
rect 1868 665 1914 724
rect 1868 600 1914 619
rect 2092 665 2138 676
rect 1700 525 2092 536
rect 2306 665 2352 724
rect 2306 600 2352 619
rect 2138 525 2356 536
rect 1654 472 2356 525
rect 285 420 340 465
rect 172 416 340 420
rect 959 424 1005 465
rect 172 370 190 416
rect 236 370 340 416
rect 172 362 340 370
rect 387 416 905 419
rect 387 370 399 416
rect 445 370 905 416
rect 387 365 905 370
rect 845 344 905 365
rect 959 415 1236 424
rect 959 369 1165 415
rect 1211 369 1236 415
rect 959 360 1236 369
rect 1299 421 1345 470
rect 1299 415 2255 421
rect 1299 369 1551 415
rect 1597 369 1767 415
rect 1813 369 1990 415
rect 2036 369 2196 415
rect 2242 369 2255 415
rect 1299 363 2255 369
rect 634 265 645 311
rect 691 265 702 311
rect 634 244 702 265
rect 845 298 848 344
rect 894 298 905 344
rect 845 246 905 298
rect 1299 244 1345 363
rect 2302 312 2356 472
rect 71 198 702 244
rect 984 198 1018 244
rect 1064 198 1345 244
rect 1654 248 2356 312
rect 1654 218 1700 248
rect 71 152 139 198
rect 71 106 82 152
rect 128 106 139 152
rect 515 106 526 152
rect 572 106 583 152
rect 721 106 750 152
rect 796 106 1286 152
rect 1332 106 1345 152
rect 1430 142 1476 181
rect 515 60 583 106
rect 2102 218 2148 248
rect 1654 131 1700 172
rect 1878 171 1924 197
rect 1430 60 1476 96
rect 2102 131 2148 172
rect 2326 176 2372 197
rect 1878 60 1924 125
rect 2326 60 2372 130
rect 0 -60 2464 60
<< labels >>
flabel metal1 s 0 724 2464 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2326 181 2372 197 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2092 536 2138 676 0 FreeSans 400 0 0 0 Z
port 3 nsew default output
flabel metal1 s 387 365 905 419 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 600 511 1005 536 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
rlabel metal1 s 845 246 905 365 1 A1
port 1 nsew default input
rlabel metal1 s 285 465 1005 511 1 A2
port 2 nsew default input
rlabel metal1 s 959 424 1005 465 1 A2
port 2 nsew default input
rlabel metal1 s 285 424 340 465 1 A2
port 2 nsew default input
rlabel metal1 s 959 420 1236 424 1 A2
port 2 nsew default input
rlabel metal1 s 285 420 340 424 1 A2
port 2 nsew default input
rlabel metal1 s 959 362 1236 420 1 A2
port 2 nsew default input
rlabel metal1 s 172 362 340 420 1 A2
port 2 nsew default input
rlabel metal1 s 959 360 1236 362 1 A2
port 2 nsew default input
rlabel metal1 s 1654 536 1700 676 1 Z
port 3 nsew default output
rlabel metal1 s 1654 472 2356 536 1 Z
port 3 nsew default output
rlabel metal1 s 2302 312 2356 472 1 Z
port 3 nsew default output
rlabel metal1 s 1654 248 2356 312 1 Z
port 3 nsew default output
rlabel metal1 s 2102 131 2148 248 1 Z
port 3 nsew default output
rlabel metal1 s 1654 131 1700 248 1 Z
port 3 nsew default output
rlabel metal1 s 2306 600 2352 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1868 600 1914 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1450 600 1496 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1255 600 1323 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 479 600 547 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 71 600 139 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1450 563 1496 600 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1255 563 1323 600 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 479 563 547 600 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 71 563 139 600 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1450 559 1496 563 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 479 559 547 563 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 71 559 139 563 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1450 557 1496 559 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 479 557 547 559 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1450 506 1496 557 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1878 181 1924 197 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2326 152 2372 181 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1878 152 1924 181 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1430 152 1476 181 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2326 60 2372 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1878 60 1924 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1430 60 1476 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 515 60 583 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string GDS_END 363730
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 358112
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
