magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 4584 3794
<< mvpmos >>
rect 0 0 120 3674
rect 224 0 344 3674
rect 448 0 568 3674
rect 672 0 792 3674
rect 896 0 1016 3674
rect 1120 0 1240 3674
rect 1344 0 1464 3674
rect 1568 0 1688 3674
rect 1792 0 1912 3674
rect 2016 0 2136 3674
rect 2240 0 2360 3674
rect 2464 0 2584 3674
rect 2688 0 2808 3674
rect 2912 0 3032 3674
rect 3136 0 3256 3674
rect 3360 0 3480 3674
rect 3584 0 3704 3674
rect 3808 0 3928 3674
rect 4032 0 4152 3674
rect 4256 0 4376 3674
<< mvpdiff >>
rect -88 3661 0 3674
rect -88 13 -75 3661
rect -29 13 0 3661
rect -88 0 0 13
rect 120 3661 224 3674
rect 120 13 149 3661
rect 195 13 224 3661
rect 120 0 224 13
rect 344 3661 448 3674
rect 344 13 373 3661
rect 419 13 448 3661
rect 344 0 448 13
rect 568 3661 672 3674
rect 568 13 597 3661
rect 643 13 672 3661
rect 568 0 672 13
rect 792 3661 896 3674
rect 792 13 821 3661
rect 867 13 896 3661
rect 792 0 896 13
rect 1016 3661 1120 3674
rect 1016 13 1045 3661
rect 1091 13 1120 3661
rect 1016 0 1120 13
rect 1240 3661 1344 3674
rect 1240 13 1269 3661
rect 1315 13 1344 3661
rect 1240 0 1344 13
rect 1464 3661 1568 3674
rect 1464 13 1493 3661
rect 1539 13 1568 3661
rect 1464 0 1568 13
rect 1688 3661 1792 3674
rect 1688 13 1717 3661
rect 1763 13 1792 3661
rect 1688 0 1792 13
rect 1912 3661 2016 3674
rect 1912 13 1941 3661
rect 1987 13 2016 3661
rect 1912 0 2016 13
rect 2136 3661 2240 3674
rect 2136 13 2165 3661
rect 2211 13 2240 3661
rect 2136 0 2240 13
rect 2360 3661 2464 3674
rect 2360 13 2389 3661
rect 2435 13 2464 3661
rect 2360 0 2464 13
rect 2584 3661 2688 3674
rect 2584 13 2613 3661
rect 2659 13 2688 3661
rect 2584 0 2688 13
rect 2808 3661 2912 3674
rect 2808 13 2837 3661
rect 2883 13 2912 3661
rect 2808 0 2912 13
rect 3032 3661 3136 3674
rect 3032 13 3061 3661
rect 3107 13 3136 3661
rect 3032 0 3136 13
rect 3256 3661 3360 3674
rect 3256 13 3285 3661
rect 3331 13 3360 3661
rect 3256 0 3360 13
rect 3480 3661 3584 3674
rect 3480 13 3509 3661
rect 3555 13 3584 3661
rect 3480 0 3584 13
rect 3704 3661 3808 3674
rect 3704 13 3733 3661
rect 3779 13 3808 3661
rect 3704 0 3808 13
rect 3928 3661 4032 3674
rect 3928 13 3957 3661
rect 4003 13 4032 3661
rect 3928 0 4032 13
rect 4152 3661 4256 3674
rect 4152 13 4181 3661
rect 4227 13 4256 3661
rect 4152 0 4256 13
rect 4376 3661 4464 3674
rect 4376 13 4405 3661
rect 4451 13 4464 3661
rect 4376 0 4464 13
<< mvpdiffc >>
rect -75 13 -29 3661
rect 149 13 195 3661
rect 373 13 419 3661
rect 597 13 643 3661
rect 821 13 867 3661
rect 1045 13 1091 3661
rect 1269 13 1315 3661
rect 1493 13 1539 3661
rect 1717 13 1763 3661
rect 1941 13 1987 3661
rect 2165 13 2211 3661
rect 2389 13 2435 3661
rect 2613 13 2659 3661
rect 2837 13 2883 3661
rect 3061 13 3107 3661
rect 3285 13 3331 3661
rect 3509 13 3555 3661
rect 3733 13 3779 3661
rect 3957 13 4003 3661
rect 4181 13 4227 3661
rect 4405 13 4451 3661
<< polysilicon >>
rect 0 3674 120 3718
rect 224 3674 344 3718
rect 448 3674 568 3718
rect 672 3674 792 3718
rect 896 3674 1016 3718
rect 1120 3674 1240 3718
rect 1344 3674 1464 3718
rect 1568 3674 1688 3718
rect 1792 3674 1912 3718
rect 2016 3674 2136 3718
rect 2240 3674 2360 3718
rect 2464 3674 2584 3718
rect 2688 3674 2808 3718
rect 2912 3674 3032 3718
rect 3136 3674 3256 3718
rect 3360 3674 3480 3718
rect 3584 3674 3704 3718
rect 3808 3674 3928 3718
rect 4032 3674 4152 3718
rect 4256 3674 4376 3718
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
rect 2240 -44 2360 0
rect 2464 -44 2584 0
rect 2688 -44 2808 0
rect 2912 -44 3032 0
rect 3136 -44 3256 0
rect 3360 -44 3480 0
rect 3584 -44 3704 0
rect 3808 -44 3928 0
rect 4032 -44 4152 0
rect 4256 -44 4376 0
<< metal1 >>
rect -75 3661 -29 3674
rect -75 0 -29 13
rect 149 3661 195 3674
rect 149 0 195 13
rect 373 3661 419 3674
rect 373 0 419 13
rect 597 3661 643 3674
rect 597 0 643 13
rect 821 3661 867 3674
rect 821 0 867 13
rect 1045 3661 1091 3674
rect 1045 0 1091 13
rect 1269 3661 1315 3674
rect 1269 0 1315 13
rect 1493 3661 1539 3674
rect 1493 0 1539 13
rect 1717 3661 1763 3674
rect 1717 0 1763 13
rect 1941 3661 1987 3674
rect 1941 0 1987 13
rect 2165 3661 2211 3674
rect 2165 0 2211 13
rect 2389 3661 2435 3674
rect 2389 0 2435 13
rect 2613 3661 2659 3674
rect 2613 0 2659 13
rect 2837 3661 2883 3674
rect 2837 0 2883 13
rect 3061 3661 3107 3674
rect 3061 0 3107 13
rect 3285 3661 3331 3674
rect 3285 0 3331 13
rect 3509 3661 3555 3674
rect 3509 0 3555 13
rect 3733 3661 3779 3674
rect 3733 0 3779 13
rect 3957 3661 4003 3674
rect 3957 0 4003 13
rect 4181 3661 4227 3674
rect 4181 0 4227 13
rect 4405 3661 4451 3674
rect 4405 0 4451 13
<< labels >>
flabel metal1 s -52 1837 -52 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 4428 1837 4428 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1837 172 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 1837 396 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 1837 620 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 1837 844 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 1837 1068 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 1837 1292 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 1837 1516 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 1740 1837 1740 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 1964 1837 1964 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 2188 1837 2188 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 2412 1837 2412 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 2636 1837 2636 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 2860 1837 2860 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 3084 1837 3084 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 3308 1837 3308 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 3532 1837 3532 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 3756 1837 3756 1837 0 FreeSans 400 0 0 0 D
flabel metal1 s 3980 1837 3980 1837 0 FreeSans 400 0 0 0 S
flabel metal1 s 4204 1837 4204 1837 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 920800
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 864134
<< end >>
