magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect 495 6371 719 7462
rect 495 6315 516 6371
rect 572 6315 640 6371
rect 696 6315 719 6371
rect 495 6247 719 6315
rect 495 6191 516 6247
rect 572 6191 640 6247
rect 696 6191 719 6247
rect 495 6123 719 6191
rect 495 6067 516 6123
rect 572 6067 640 6123
rect 696 6067 719 6123
rect -8 5681 216 5708
rect -8 5625 16 5681
rect 72 5625 140 5681
rect 196 5625 216 5681
rect -8 5557 216 5625
rect -8 5501 16 5557
rect 72 5501 140 5557
rect 196 5501 216 5557
rect -8 5433 216 5501
rect -8 5377 16 5433
rect 72 5377 140 5433
rect 196 5377 216 5433
rect -8 4667 216 5377
rect -8 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 216 4667
rect -8 4543 216 4611
rect -8 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 216 4543
rect -8 4419 216 4487
rect -8 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 216 4419
rect -8 3065 216 4363
rect 495 3313 719 6067
rect 1011 5681 1235 5708
rect 1011 5625 1033 5681
rect 1089 5625 1157 5681
rect 1213 5625 1235 5681
rect 1011 5557 1235 5625
rect 1011 5501 1033 5557
rect 1089 5501 1157 5557
rect 1213 5501 1235 5557
rect 1011 5433 1235 5501
rect 1011 5377 1033 5433
rect 1089 5377 1157 5433
rect 1213 5377 1235 5433
rect 1011 4667 1235 5377
rect 1011 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1235 4667
rect 1011 4543 1235 4611
rect 1011 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1235 4543
rect 1011 4419 1235 4487
rect 1011 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1235 4419
rect 1011 3065 1235 4363
<< via2 >>
rect 516 6315 572 6371
rect 640 6315 696 6371
rect 516 6191 572 6247
rect 640 6191 696 6247
rect 516 6067 572 6123
rect 640 6067 696 6123
rect 16 5625 72 5681
rect 140 5625 196 5681
rect 16 5501 72 5557
rect 140 5501 196 5557
rect 16 5377 72 5433
rect 140 5377 196 5433
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 1033 5625 1089 5681
rect 1157 5625 1213 5681
rect 1033 5501 1089 5557
rect 1157 5501 1213 5557
rect 1033 5377 1089 5433
rect 1157 5377 1213 5433
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 506 6371 706 6381
rect 506 6315 516 6371
rect 572 6315 640 6371
rect 696 6315 706 6371
rect 506 6247 706 6315
rect 506 6191 516 6247
rect 572 6191 640 6247
rect 696 6191 706 6247
rect 506 6123 706 6191
rect 506 6067 516 6123
rect 572 6067 640 6123
rect 696 6067 706 6123
rect 506 6057 706 6067
rect 6 5681 206 5691
rect 6 5625 16 5681
rect 72 5625 140 5681
rect 196 5625 206 5681
rect 6 5557 206 5625
rect 6 5501 16 5557
rect 72 5501 140 5557
rect 196 5501 206 5557
rect 6 5433 206 5501
rect 6 5377 16 5433
rect 72 5377 140 5433
rect 196 5377 206 5433
rect 6 5367 206 5377
rect 1023 5681 1223 5691
rect 1023 5625 1033 5681
rect 1089 5625 1157 5681
rect 1213 5625 1223 5681
rect 1023 5557 1223 5625
rect 1023 5501 1033 5557
rect 1089 5501 1157 5557
rect 1213 5501 1223 5557
rect 1023 5433 1223 5501
rect 1023 5377 1033 5433
rect 1089 5377 1157 5433
rect 1213 5377 1223 5433
rect 1023 5367 1223 5377
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
use M2_M14310589983294_64x8m81  M2_M14310589983294_64x8m81_0
timestamp 1669390400
transform 1 0 1120 0 1 3728
box -100 -472 100 472
use M2_M14310589983294_64x8m81  M2_M14310589983294_64x8m81_1
timestamp 1669390400
transform 1 0 103 0 1 3728
box -100 -472 100 472
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 6219
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_1
timestamp 1669390400
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_2
timestamp 1669390400
transform 1 0 1123 0 1 5529
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_3
timestamp 1669390400
transform 1 0 106 0 1 5529
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_4
timestamp 1669390400
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M24310589983299_64x8m81  M3_M24310589983299_64x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 3696
box -100 -348 100 348
<< properties >>
string GDS_END 1098056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1097460
<< end >>
