magic
tech gf180mcuC
magscale 1 5
timestamp 1675911052
<< obsm1 >>
rect 120 2430 89880 57225
<< metal2 >>
rect 5768 59600 5824 60000
rect 16968 59600 17024 60000
rect 28168 59600 28224 60000
rect 39368 59600 39424 60000
rect 50568 59600 50624 60000
rect 61768 59600 61824 60000
rect 72968 59600 73024 60000
rect 84168 59600 84224 60000
rect 4648 0 4704 400
rect 13608 0 13664 400
rect 22568 0 22624 400
rect 31528 0 31584 400
rect 40488 0 40544 400
rect 49448 0 49504 400
rect 58408 0 58464 400
rect 67368 0 67424 400
rect 76328 0 76384 400
rect 85288 0 85344 400
<< obsm2 >>
rect 336 59570 5738 59682
rect 5854 59570 16938 59682
rect 17054 59570 28138 59682
rect 28254 59570 39338 59682
rect 39454 59570 50538 59682
rect 50654 59570 61738 59682
rect 61854 59570 72938 59682
rect 73054 59570 84138 59682
rect 84254 59570 89759 59682
rect 336 430 89759 59570
rect 336 400 4618 430
rect 4734 400 13578 430
rect 13694 400 22538 430
rect 22654 400 31498 430
rect 31614 400 40458 430
rect 40574 400 49418 430
rect 49534 400 58378 430
rect 58494 400 67338 430
rect 67454 400 76298 430
rect 76414 400 85258 430
rect 85374 400 89759 430
<< metal3 >>
rect 0 52360 400 52416
rect 89600 52360 90000 52416
rect 0 37408 400 37464
rect 89600 37408 90000 37464
rect 0 22456 400 22512
rect 89600 22456 90000 22512
rect 0 7504 400 7560
rect 89600 7504 90000 7560
<< obsm3 >>
rect 345 52446 89759 57209
rect 430 52330 89570 52446
rect 345 37494 89759 52330
rect 430 37378 89570 37494
rect 345 22542 89759 37378
rect 430 22426 89570 22542
rect 345 7590 89759 22426
rect 430 7474 89570 7590
rect 345 2446 89759 7474
<< metal4 >>
rect 1672 2430 1832 57225
rect 9352 2430 9512 57225
rect 17032 2430 17192 57225
rect 24712 2430 24872 57225
rect 32392 2430 32552 57225
rect 40072 2430 40232 57225
rect 47752 2430 47912 57225
rect 55432 2430 55592 57225
rect 63112 2430 63272 57225
rect 70792 2430 70952 57225
rect 78472 2430 78632 57225
rect 86152 2430 86312 57225
<< obsm4 >>
rect 33278 14681 40042 28607
rect 40262 14681 47722 28607
rect 47942 14681 55402 28607
rect 55622 14681 58898 28607
<< labels >>
rlabel metal3 s 89600 7504 90000 7560 6 a[0]
port 1 nsew signal input
rlabel metal3 s 89600 22456 90000 22512 6 a[1]
port 2 nsew signal input
rlabel metal3 s 89600 37408 90000 37464 6 a[2]
port 3 nsew signal input
rlabel metal3 s 89600 52360 90000 52416 6 a[3]
port 4 nsew signal input
rlabel metal3 s 0 7504 400 7560 6 b[0]
port 5 nsew signal input
rlabel metal3 s 0 22456 400 22512 6 b[1]
port 6 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 b[2]
port 7 nsew signal input
rlabel metal3 s 0 52360 400 52416 6 b[3]
port 8 nsew signal input
rlabel metal2 s 22568 0 22624 400 6 ci[0]
port 9 nsew signal input
rlabel metal2 s 31528 0 31584 400 6 ci[1]
port 10 nsew signal input
rlabel metal2 s 40488 0 40544 400 6 ci[2]
port 11 nsew signal input
rlabel metal2 s 49448 0 49504 400 6 ci[3]
port 12 nsew signal input
rlabel metal2 s 58408 0 58464 400 6 ci[4]
port 13 nsew signal input
rlabel metal2 s 67368 0 67424 400 6 ci[5]
port 14 nsew signal input
rlabel metal2 s 76328 0 76384 400 6 ci[6]
port 15 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 ci[7]
port 16 nsew signal input
rlabel metal2 s 4648 0 4704 400 6 clk
port 17 nsew signal input
rlabel metal2 s 5768 59600 5824 60000 6 o[0]
port 18 nsew signal output
rlabel metal2 s 16968 59600 17024 60000 6 o[1]
port 19 nsew signal output
rlabel metal2 s 28168 59600 28224 60000 6 o[2]
port 20 nsew signal output
rlabel metal2 s 39368 59600 39424 60000 6 o[3]
port 21 nsew signal output
rlabel metal2 s 50568 59600 50624 60000 6 o[4]
port 22 nsew signal output
rlabel metal2 s 61768 59600 61824 60000 6 o[5]
port 23 nsew signal output
rlabel metal2 s 72968 59600 73024 60000 6 o[6]
port 24 nsew signal output
rlabel metal2 s 84168 59600 84224 60000 6 o[7]
port 25 nsew signal output
rlabel metal2 s 13608 0 13664 400 6 rst
port 26 nsew signal input
rlabel metal4 s 1672 2430 1832 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 17032 2430 17192 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 32392 2430 32552 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 47752 2430 47912 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 63112 2430 63272 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 78472 2430 78632 57225 6 vdd
port 27 nsew power bidirectional
rlabel metal4 s 9352 2430 9512 57225 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 24712 2430 24872 57225 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 40072 2430 40232 57225 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 55432 2430 55592 57225 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 70792 2430 70952 57225 6 vss
port 28 nsew ground bidirectional
rlabel metal4 s 86152 2430 86312 57225 6 vss
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4890294
string GDS_FILE /Users/lrburle/Library/CloudStorage/OneDrive-Personal/PhD/projects/osu180cells/openlane/ffra/runs/23_02_08_20_47/results/signoff/ffra.magic.gds
string GDS_START 90054
<< end >>

