magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -64 897 65 937
rect -64 845 -26 897
rect 26 845 65 897
rect -64 679 65 845
rect -64 627 -26 679
rect 26 627 65 679
rect -64 461 65 627
rect -64 409 -26 461
rect 26 409 65 461
rect -64 244 65 409
rect -64 192 -26 244
rect 26 192 65 244
rect -64 26 65 192
rect -64 -26 -26 26
rect 26 -26 65 26
rect -64 -192 65 -26
rect -64 -244 -26 -192
rect 26 -244 65 -192
rect -64 -409 65 -244
rect -64 -461 -26 -409
rect 26 -461 65 -409
rect -64 -627 65 -461
rect -64 -679 -26 -627
rect 26 -679 65 -627
rect -64 -845 65 -679
rect -64 -897 -26 -845
rect 26 -897 65 -845
rect -64 -937 65 -897
<< via1 >>
rect -26 845 26 897
rect -26 627 26 679
rect -26 409 26 461
rect -26 192 26 244
rect -26 -26 26 26
rect -26 -244 26 -192
rect -26 -461 26 -409
rect -26 -679 26 -627
rect -26 -897 26 -845
<< metal2 >>
rect -64 897 65 937
rect -64 845 -26 897
rect 26 845 65 897
rect -64 679 65 845
rect -64 627 -26 679
rect 26 627 65 679
rect -64 461 65 627
rect -64 409 -26 461
rect 26 409 65 461
rect -64 244 65 409
rect -64 192 -26 244
rect 26 192 65 244
rect -64 26 65 192
rect -64 -26 -26 26
rect 26 -26 65 26
rect -64 -192 65 -26
rect -64 -244 -26 -192
rect 26 -244 65 -192
rect -64 -409 65 -244
rect -64 -461 -26 -409
rect 26 -461 65 -409
rect -64 -627 65 -461
rect -64 -679 -26 -627
rect 26 -679 65 -627
rect -64 -845 65 -679
rect -64 -897 -26 -845
rect 26 -897 65 -845
rect -64 -937 65 -897
<< properties >>
string GDS_END 1095004
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1094296
<< end >>
