magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 560 844
rect 50 506 96 724
rect 254 460 300 676
rect 458 506 504 724
rect 127 212 200 438
rect 254 414 536 460
rect 248 288 411 364
rect 50 60 96 161
rect 248 111 321 288
rect 458 106 536 414
rect 0 -60 560 60
<< labels >>
rlabel metal1 s 248 288 411 364 6 A1
port 1 nsew default input
rlabel metal1 s 248 111 321 288 6 A1
port 1 nsew default input
rlabel metal1 s 127 212 200 438 6 A2
port 2 nsew default input
rlabel metal1 s 254 460 300 676 6 ZN
port 3 nsew default output
rlabel metal1 s 254 414 536 460 6 ZN
port 3 nsew default output
rlabel metal1 s 458 106 536 414 6 ZN
port 3 nsew default output
rlabel metal1 s 0 724 560 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 458 506 504 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 50 506 96 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 50 60 96 161 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 560 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 560 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 688252
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 685706
<< end >>
