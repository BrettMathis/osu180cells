magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3894 1094
<< pwell >>
rect -86 -86 3894 453
<< mvnmos >>
rect 124 187 244 333
rect 348 187 468 333
rect 572 187 692 333
rect 796 187 916 333
rect 1020 187 1140 333
rect 1244 187 1364 333
rect 1468 187 1588 333
rect 1692 187 1812 333
rect 1916 187 2036 333
rect 2140 187 2260 333
rect 2364 187 2484 333
rect 2588 187 2708 333
rect 2812 187 2932 333
rect 3036 187 3156 333
rect 3260 187 3380 333
rect 3484 187 3604 333
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
rect 572 573 672 939
rect 796 573 896 939
rect 1020 573 1120 939
rect 1244 573 1344 939
rect 1468 573 1568 939
rect 1692 573 1792 939
rect 1916 573 2016 939
rect 2140 573 2240 939
rect 2364 573 2464 939
rect 2588 573 2688 939
rect 2812 573 2912 939
rect 3036 573 3136 939
rect 3260 573 3360 939
rect 3484 573 3584 939
<< mvndiff >>
rect 36 246 124 333
rect 36 200 49 246
rect 95 200 124 246
rect 36 187 124 200
rect 244 246 348 333
rect 244 200 273 246
rect 319 200 348 246
rect 244 187 348 200
rect 468 246 572 333
rect 468 200 497 246
rect 543 200 572 246
rect 468 187 572 200
rect 692 246 796 333
rect 692 200 721 246
rect 767 200 796 246
rect 692 187 796 200
rect 916 246 1020 333
rect 916 200 945 246
rect 991 200 1020 246
rect 916 187 1020 200
rect 1140 246 1244 333
rect 1140 200 1169 246
rect 1215 200 1244 246
rect 1140 187 1244 200
rect 1364 246 1468 333
rect 1364 200 1393 246
rect 1439 200 1468 246
rect 1364 187 1468 200
rect 1588 246 1692 333
rect 1588 200 1617 246
rect 1663 200 1692 246
rect 1588 187 1692 200
rect 1812 246 1916 333
rect 1812 200 1841 246
rect 1887 200 1916 246
rect 1812 187 1916 200
rect 2036 246 2140 333
rect 2036 200 2065 246
rect 2111 200 2140 246
rect 2036 187 2140 200
rect 2260 246 2364 333
rect 2260 200 2289 246
rect 2335 200 2364 246
rect 2260 187 2364 200
rect 2484 246 2588 333
rect 2484 200 2513 246
rect 2559 200 2588 246
rect 2484 187 2588 200
rect 2708 246 2812 333
rect 2708 200 2737 246
rect 2783 200 2812 246
rect 2708 187 2812 200
rect 2932 246 3036 333
rect 2932 200 2961 246
rect 3007 200 3036 246
rect 2932 187 3036 200
rect 3156 246 3260 333
rect 3156 200 3185 246
rect 3231 200 3260 246
rect 3156 187 3260 200
rect 3380 246 3484 333
rect 3380 200 3409 246
rect 3455 200 3484 246
rect 3380 187 3484 200
rect 3604 246 3692 333
rect 3604 200 3633 246
rect 3679 200 3692 246
rect 3604 187 3692 200
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 572 939
rect 448 721 477 861
rect 523 721 572 861
rect 448 573 572 721
rect 672 861 796 939
rect 672 721 701 861
rect 747 721 796 861
rect 672 573 796 721
rect 896 861 1020 939
rect 896 721 925 861
rect 971 721 1020 861
rect 896 573 1020 721
rect 1120 861 1244 939
rect 1120 721 1149 861
rect 1195 721 1244 861
rect 1120 573 1244 721
rect 1344 861 1468 939
rect 1344 721 1373 861
rect 1419 721 1468 861
rect 1344 573 1468 721
rect 1568 861 1692 939
rect 1568 721 1597 861
rect 1643 721 1692 861
rect 1568 573 1692 721
rect 1792 861 1916 939
rect 1792 721 1821 861
rect 1867 721 1916 861
rect 1792 573 1916 721
rect 2016 861 2140 939
rect 2016 721 2045 861
rect 2091 721 2140 861
rect 2016 573 2140 721
rect 2240 861 2364 939
rect 2240 721 2269 861
rect 2315 721 2364 861
rect 2240 573 2364 721
rect 2464 861 2588 939
rect 2464 721 2493 861
rect 2539 721 2588 861
rect 2464 573 2588 721
rect 2688 861 2812 939
rect 2688 721 2717 861
rect 2763 721 2812 861
rect 2688 573 2812 721
rect 2912 861 3036 939
rect 2912 721 2941 861
rect 2987 721 3036 861
rect 2912 573 3036 721
rect 3136 861 3260 939
rect 3136 721 3165 861
rect 3211 721 3260 861
rect 3136 573 3260 721
rect 3360 861 3484 939
rect 3360 721 3389 861
rect 3435 721 3484 861
rect 3360 573 3484 721
rect 3584 861 3672 939
rect 3584 721 3613 861
rect 3659 721 3672 861
rect 3584 573 3672 721
<< mvndiffc >>
rect 49 200 95 246
rect 273 200 319 246
rect 497 200 543 246
rect 721 200 767 246
rect 945 200 991 246
rect 1169 200 1215 246
rect 1393 200 1439 246
rect 1617 200 1663 246
rect 1841 200 1887 246
rect 2065 200 2111 246
rect 2289 200 2335 246
rect 2513 200 2559 246
rect 2737 200 2783 246
rect 2961 200 3007 246
rect 3185 200 3231 246
rect 3409 200 3455 246
rect 3633 200 3679 246
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
rect 701 721 747 861
rect 925 721 971 861
rect 1149 721 1195 861
rect 1373 721 1419 861
rect 1597 721 1643 861
rect 1821 721 1867 861
rect 2045 721 2091 861
rect 2269 721 2315 861
rect 2493 721 2539 861
rect 2717 721 2763 861
rect 2941 721 2987 861
rect 3165 721 3211 861
rect 3389 721 3435 861
rect 3613 721 3659 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 572 939 672 983
rect 796 939 896 983
rect 1020 939 1120 983
rect 1244 939 1344 983
rect 1468 939 1568 983
rect 1692 939 1792 983
rect 1916 939 2016 983
rect 2140 939 2240 983
rect 2364 939 2464 983
rect 2588 939 2688 983
rect 2812 939 2912 983
rect 3036 939 3136 983
rect 3260 939 3360 983
rect 3484 939 3584 983
rect 124 513 224 573
rect 348 513 448 573
rect 572 513 672 573
rect 796 513 896 573
rect 1020 513 1120 573
rect 1244 513 1344 573
rect 1468 513 1568 573
rect 1692 513 1792 573
rect 1916 513 2016 573
rect 2140 513 2240 573
rect 2364 513 2464 573
rect 2588 513 2688 573
rect 2812 513 2912 573
rect 3036 513 3136 573
rect 3260 513 3360 573
rect 124 512 3360 513
rect 3484 512 3584 573
rect 124 500 3584 512
rect 124 454 137 500
rect 1593 454 1870 500
rect 3326 454 3584 500
rect 124 441 3584 454
rect 124 333 244 441
rect 348 333 468 441
rect 572 333 692 441
rect 796 333 916 441
rect 1020 333 1140 441
rect 1244 333 1364 441
rect 1468 333 1588 441
rect 1692 333 1812 441
rect 1916 333 2036 441
rect 2140 333 2260 441
rect 2364 333 2484 441
rect 2588 333 2708 441
rect 2812 333 2932 441
rect 3036 333 3156 441
rect 3260 333 3380 441
rect 3484 377 3584 441
rect 3484 333 3604 377
rect 124 143 244 187
rect 348 143 468 187
rect 572 143 692 187
rect 796 143 916 187
rect 1020 143 1140 187
rect 1244 143 1364 187
rect 1468 143 1588 187
rect 1692 143 1812 187
rect 1916 143 2036 187
rect 2140 143 2260 187
rect 2364 143 2484 187
rect 2588 143 2708 187
rect 2812 143 2932 187
rect 3036 143 3156 187
rect 3260 143 3380 187
rect 3484 143 3604 187
<< polycontact >>
rect 137 454 1593 500
rect 1870 454 3326 500
<< metal1 >>
rect 0 918 3808 1098
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 273 664 319 721
rect 477 861 523 918
rect 477 710 523 721
rect 701 861 747 872
rect 701 664 747 721
rect 925 861 971 918
rect 925 710 971 721
rect 1149 861 1195 872
rect 1149 664 1195 721
rect 1373 861 1419 918
rect 1373 710 1419 721
rect 1597 861 1643 872
rect 1597 664 1643 721
rect 1821 861 1867 918
rect 1821 710 1867 721
rect 2045 861 2091 872
rect 2045 664 2091 721
rect 2269 861 2315 918
rect 2269 710 2315 721
rect 2493 861 2539 872
rect 2493 664 2539 721
rect 2717 861 2763 918
rect 2717 710 2763 721
rect 2941 861 2987 872
rect 2941 664 2987 721
rect 3165 861 3211 918
rect 3165 710 3211 721
rect 3389 861 3435 872
rect 3389 664 3435 721
rect 3613 861 3659 918
rect 3613 710 3659 721
rect 273 618 3435 664
rect 126 500 1604 530
rect 126 454 137 500
rect 1593 454 1604 500
rect 1653 349 1813 618
rect 1859 500 3337 530
rect 1859 454 1870 500
rect 3326 454 3337 500
rect 273 303 3455 349
rect 49 246 95 257
rect 49 90 95 200
rect 273 246 325 303
rect 319 200 325 246
rect 273 189 325 200
rect 497 246 543 257
rect 497 90 543 200
rect 721 246 767 303
rect 721 189 767 200
rect 945 246 991 257
rect 945 90 991 200
rect 1169 246 1215 303
rect 1169 189 1215 200
rect 1393 246 1439 257
rect 1393 90 1439 200
rect 1617 246 1663 303
rect 1617 189 1663 200
rect 1841 246 1887 257
rect 1841 90 1887 200
rect 2065 246 2111 303
rect 2065 189 2111 200
rect 2289 246 2335 257
rect 2289 90 2335 200
rect 2513 246 2559 303
rect 2513 189 2559 200
rect 2737 246 2783 257
rect 2737 90 2783 200
rect 2961 246 3007 303
rect 2961 189 3007 200
rect 3185 246 3231 257
rect 3185 90 3231 200
rect 3409 246 3455 303
rect 3409 189 3455 200
rect 3633 246 3679 257
rect 3633 90 3679 200
rect 0 -90 3808 90
<< labels >>
flabel metal1 s 126 454 1604 530 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 3808 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 3633 90 3679 257 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3389 664 3435 872 0 FreeSans 200 0 0 0 ZN
port 2 nsew default output
rlabel metal1 s 1859 454 3337 530 1 I
port 1 nsew default input
rlabel metal1 s 2941 664 2987 872 1 ZN
port 2 nsew default output
rlabel metal1 s 2493 664 2539 872 1 ZN
port 2 nsew default output
rlabel metal1 s 2045 664 2091 872 1 ZN
port 2 nsew default output
rlabel metal1 s 1597 664 1643 872 1 ZN
port 2 nsew default output
rlabel metal1 s 1149 664 1195 872 1 ZN
port 2 nsew default output
rlabel metal1 s 701 664 747 872 1 ZN
port 2 nsew default output
rlabel metal1 s 273 664 319 872 1 ZN
port 2 nsew default output
rlabel metal1 s 273 618 3435 664 1 ZN
port 2 nsew default output
rlabel metal1 s 1653 349 1813 618 1 ZN
port 2 nsew default output
rlabel metal1 s 273 303 3455 349 1 ZN
port 2 nsew default output
rlabel metal1 s 3409 189 3455 303 1 ZN
port 2 nsew default output
rlabel metal1 s 2961 189 3007 303 1 ZN
port 2 nsew default output
rlabel metal1 s 2513 189 2559 303 1 ZN
port 2 nsew default output
rlabel metal1 s 2065 189 2111 303 1 ZN
port 2 nsew default output
rlabel metal1 s 1617 189 1663 303 1 ZN
port 2 nsew default output
rlabel metal1 s 1169 189 1215 303 1 ZN
port 2 nsew default output
rlabel metal1 s 721 189 767 303 1 ZN
port 2 nsew default output
rlabel metal1 s 273 189 325 303 1 ZN
port 2 nsew default output
rlabel metal1 s 3613 710 3659 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 710 3211 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 710 2763 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 710 2315 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 710 1867 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 710 1419 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3185 90 3231 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2737 90 2783 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 257 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3808 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 1008
string GDS_END 1446494
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1437576
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
