magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 918 1120 1098
rect 49 710 95 918
rect 273 670 319 872
rect 477 716 523 918
rect 701 670 767 872
rect 925 710 971 918
rect 273 624 767 670
rect 116 454 466 530
rect 667 378 767 624
rect 273 332 767 378
rect 49 90 95 286
rect 273 136 319 332
rect 497 90 543 286
rect 721 136 767 332
rect 945 90 991 286
rect 0 -90 1120 90
<< labels >>
rlabel metal1 s 116 454 466 530 6 I
port 1 nsew default input
rlabel metal1 s 701 670 767 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 670 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 624 767 670 6 ZN
port 2 nsew default output
rlabel metal1 s 667 378 767 624 6 ZN
port 2 nsew default output
rlabel metal1 s 273 332 767 378 6 ZN
port 2 nsew default output
rlabel metal1 s 721 136 767 332 6 ZN
port 2 nsew default output
rlabel metal1 s 273 136 319 332 6 ZN
port 2 nsew default output
rlabel metal1 s 0 918 1120 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 716 971 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 716 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 716 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 716 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 716 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 945 90 991 286 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 286 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 286 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1120 90 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 864052
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 860510
<< end >>
