magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4790 1094
<< pwell >>
rect -86 -86 4790 453
<< mvnmos >>
rect 140 69 260 333
rect 364 69 484 333
rect 588 69 708 333
rect 812 69 932 333
rect 1080 173 1200 333
rect 1248 173 1368 333
rect 1416 173 1536 333
rect 1640 173 1760 333
rect 1864 173 1984 333
rect 2088 173 2208 333
rect 2312 173 2432 333
rect 2680 173 2800 333
rect 2904 173 3024 333
rect 3128 173 3248 333
rect 3352 173 3472 333
rect 3520 173 3640 333
rect 3788 69 3908 333
rect 4012 69 4132 333
rect 4236 69 4356 333
rect 4460 69 4580 333
<< mvpmos >>
rect 140 573 240 939
rect 364 573 464 939
rect 589 573 689 939
rect 832 573 932 939
rect 1100 573 1200 851
rect 1268 573 1368 851
rect 1436 573 1536 851
rect 1660 573 1760 851
rect 1884 573 1984 851
rect 2088 573 2188 851
rect 2312 573 2412 851
rect 2700 573 2800 851
rect 2904 573 3004 851
rect 3128 573 3228 851
rect 3352 573 3452 851
rect 3520 573 3620 851
rect 3788 573 3888 939
rect 4012 573 4112 939
rect 4236 573 4336 939
rect 4460 573 4560 939
<< mvndiff >>
rect 52 222 140 333
rect 52 82 65 222
rect 111 82 140 222
rect 52 69 140 82
rect 260 320 364 333
rect 260 180 289 320
rect 335 180 364 320
rect 260 69 364 180
rect 484 222 588 333
rect 484 82 513 222
rect 559 82 588 222
rect 484 69 588 82
rect 708 320 812 333
rect 708 180 737 320
rect 783 180 812 320
rect 708 69 812 180
rect 932 222 1080 333
rect 932 82 961 222
rect 1007 173 1080 222
rect 1200 173 1248 333
rect 1368 173 1416 333
rect 1536 309 1640 333
rect 1536 263 1565 309
rect 1611 263 1640 309
rect 1536 173 1640 263
rect 1760 320 1864 333
rect 1760 274 1789 320
rect 1835 274 1864 320
rect 1760 173 1864 274
rect 1984 232 2088 333
rect 1984 186 2013 232
rect 2059 186 2088 232
rect 1984 173 2088 186
rect 2208 320 2312 333
rect 2208 274 2237 320
rect 2283 274 2312 320
rect 2208 173 2312 274
rect 2432 232 2520 333
rect 2432 186 2461 232
rect 2507 186 2520 232
rect 2432 173 2520 186
rect 2592 320 2680 333
rect 2592 274 2605 320
rect 2651 274 2680 320
rect 2592 173 2680 274
rect 2800 232 2904 333
rect 2800 186 2829 232
rect 2875 186 2904 232
rect 2800 173 2904 186
rect 3024 320 3128 333
rect 3024 274 3053 320
rect 3099 274 3128 320
rect 3024 173 3128 274
rect 3248 320 3352 333
rect 3248 274 3277 320
rect 3323 274 3352 320
rect 3248 173 3352 274
rect 3472 173 3520 333
rect 3640 222 3788 333
rect 3640 173 3713 222
rect 1007 82 1020 173
rect 932 69 1020 82
rect 3700 82 3713 173
rect 3759 82 3788 222
rect 3700 69 3788 82
rect 3908 320 4012 333
rect 3908 180 3937 320
rect 3983 180 4012 320
rect 3908 69 4012 180
rect 4132 222 4236 333
rect 4132 82 4161 222
rect 4207 82 4236 222
rect 4132 69 4236 82
rect 4356 320 4460 333
rect 4356 180 4385 320
rect 4431 180 4460 320
rect 4356 69 4460 180
rect 4580 222 4668 333
rect 4580 82 4609 222
rect 4655 82 4668 222
rect 4580 69 4668 82
<< mvpdiff >>
rect 52 926 140 939
rect 52 786 65 926
rect 111 786 140 926
rect 52 573 140 786
rect 240 726 364 939
rect 240 586 289 726
rect 335 586 364 726
rect 240 573 364 586
rect 464 926 589 939
rect 464 786 511 926
rect 557 786 589 926
rect 464 573 589 786
rect 689 726 832 939
rect 689 586 757 726
rect 803 586 832 726
rect 689 573 832 586
rect 932 926 1040 939
rect 932 786 981 926
rect 1027 851 1040 926
rect 3680 926 3788 939
rect 3680 851 3693 926
rect 1027 786 1100 851
rect 932 573 1100 786
rect 1200 573 1268 851
rect 1368 573 1436 851
rect 1536 726 1660 851
rect 1536 586 1565 726
rect 1611 586 1660 726
rect 1536 573 1660 586
rect 1760 737 1884 851
rect 1760 597 1809 737
rect 1855 597 1884 737
rect 1760 573 1884 597
rect 1984 838 2088 851
rect 1984 792 2013 838
rect 2059 792 2088 838
rect 1984 573 2088 792
rect 2188 632 2312 851
rect 2188 586 2217 632
rect 2263 586 2312 632
rect 2188 573 2312 586
rect 2412 838 2500 851
rect 2412 698 2441 838
rect 2487 698 2500 838
rect 2412 573 2500 698
rect 2612 737 2700 851
rect 2612 597 2625 737
rect 2671 597 2700 737
rect 2612 573 2700 597
rect 2800 838 2904 851
rect 2800 698 2829 838
rect 2875 698 2904 838
rect 2800 573 2904 698
rect 3004 737 3128 851
rect 3004 597 3033 737
rect 3079 597 3128 737
rect 3004 573 3128 597
rect 3228 739 3352 851
rect 3228 599 3257 739
rect 3303 599 3352 739
rect 3228 573 3352 599
rect 3452 573 3520 851
rect 3620 786 3693 851
rect 3739 786 3788 926
rect 3620 573 3788 786
rect 3888 726 4012 939
rect 3888 586 3927 726
rect 3973 586 4012 726
rect 3888 573 4012 586
rect 4112 926 4236 939
rect 4112 786 4150 926
rect 4196 786 4236 926
rect 4112 573 4236 786
rect 4336 726 4460 939
rect 4336 586 4375 726
rect 4421 586 4460 726
rect 4336 573 4460 586
rect 4560 926 4668 939
rect 4560 786 4589 926
rect 4635 786 4668 926
rect 4560 573 4668 786
<< mvndiffc >>
rect 65 82 111 222
rect 289 180 335 320
rect 513 82 559 222
rect 737 180 783 320
rect 961 82 1007 222
rect 1565 263 1611 309
rect 1789 274 1835 320
rect 2013 186 2059 232
rect 2237 274 2283 320
rect 2461 186 2507 232
rect 2605 274 2651 320
rect 2829 186 2875 232
rect 3053 274 3099 320
rect 3277 274 3323 320
rect 3713 82 3759 222
rect 3937 180 3983 320
rect 4161 82 4207 222
rect 4385 180 4431 320
rect 4609 82 4655 222
<< mvpdiffc >>
rect 65 786 111 926
rect 289 586 335 726
rect 511 786 557 926
rect 757 586 803 726
rect 981 786 1027 926
rect 1565 586 1611 726
rect 1809 597 1855 737
rect 2013 792 2059 838
rect 2217 586 2263 632
rect 2441 698 2487 838
rect 2625 597 2671 737
rect 2829 698 2875 838
rect 3033 597 3079 737
rect 3257 599 3303 739
rect 3693 786 3739 926
rect 3927 586 3973 726
rect 4150 786 4196 926
rect 4375 586 4421 726
rect 4589 786 4635 926
<< polysilicon >>
rect 140 939 240 983
rect 364 939 464 983
rect 589 939 689 983
rect 832 939 932 983
rect 1268 943 3452 983
rect 1100 851 1200 895
rect 1268 851 1368 943
rect 1436 851 1536 895
rect 1660 851 1760 895
rect 1884 851 1984 895
rect 2088 851 2188 943
rect 2312 851 2412 895
rect 2700 851 2800 943
rect 2904 851 3004 895
rect 3128 851 3228 895
rect 3352 851 3452 943
rect 3788 939 3888 983
rect 4012 939 4112 983
rect 4236 939 4336 983
rect 4460 939 4560 983
rect 3520 851 3620 895
rect 140 513 240 573
rect 364 513 464 573
rect 589 513 689 573
rect 832 513 932 573
rect 140 506 932 513
rect 140 441 873 506
rect 140 333 260 441
rect 364 333 484 441
rect 588 333 708 441
rect 812 366 873 441
rect 919 366 932 506
rect 1100 523 1200 573
rect 1100 383 1141 523
rect 1187 383 1200 523
rect 1100 377 1200 383
rect 1268 377 1368 573
rect 1436 430 1536 573
rect 1436 384 1477 430
rect 1523 384 1536 430
rect 1436 377 1536 384
rect 1660 540 1760 573
rect 1660 494 1701 540
rect 1747 494 1760 540
rect 1660 377 1760 494
rect 1884 377 1984 573
rect 812 333 932 366
rect 1080 333 1200 377
rect 1248 333 1368 377
rect 1416 333 1536 377
rect 1640 333 1760 377
rect 1864 333 1984 377
rect 2088 377 2188 573
rect 2312 430 2412 573
rect 2312 384 2325 430
rect 2371 384 2412 430
rect 2312 377 2412 384
rect 2700 377 2800 573
rect 2088 333 2208 377
rect 2312 333 2432 377
rect 2680 333 2800 377
rect 2904 377 3004 573
rect 3128 430 3228 573
rect 3128 384 3141 430
rect 3187 384 3228 430
rect 3128 377 3228 384
rect 3352 523 3452 573
rect 3352 477 3393 523
rect 3439 477 3452 523
rect 3352 377 3452 477
rect 3520 377 3620 573
rect 3788 513 3888 573
rect 4012 513 4112 573
rect 4236 513 4336 573
rect 4460 513 4560 573
rect 3788 508 4560 513
rect 3788 506 4580 508
rect 2904 333 3024 377
rect 3128 333 3248 377
rect 3352 333 3472 377
rect 3520 333 3640 377
rect 3788 366 3801 506
rect 3847 454 4580 506
rect 3847 453 4132 454
rect 3847 366 3908 453
rect 3788 333 3908 366
rect 4012 333 4132 453
rect 4236 333 4356 454
rect 4460 333 4580 454
rect 1080 81 1200 173
rect 1248 129 1368 173
rect 1416 129 1536 173
rect 1640 129 1760 173
rect 1864 81 1984 173
rect 2088 129 2208 173
rect 2312 129 2432 173
rect 2680 129 2800 173
rect 2904 81 3024 173
rect 3128 129 3248 173
rect 3352 129 3472 173
rect 3520 81 3640 173
rect 140 25 260 69
rect 364 25 484 69
rect 588 25 708 69
rect 812 25 932 69
rect 1080 41 3640 81
rect 3788 25 3908 69
rect 4012 25 4132 69
rect 4236 25 4356 69
rect 4460 25 4580 69
<< polycontact >>
rect 873 366 919 506
rect 1141 383 1187 523
rect 1477 384 1523 430
rect 1701 494 1747 540
rect 2325 384 2371 430
rect 3141 384 3187 430
rect 3393 477 3439 523
rect 3801 366 3847 506
<< metal1 >>
rect 0 926 4704 1098
rect 0 918 65 926
rect 111 918 511 926
rect 65 775 111 786
rect 557 918 981 926
rect 511 775 557 786
rect 1027 918 3693 926
rect 981 775 1027 786
rect 2013 838 2059 918
rect 2013 781 2059 792
rect 2441 838 2487 918
rect 1809 737 1855 748
rect 289 726 335 737
rect 757 726 803 737
rect 335 586 757 621
rect 1565 726 1611 737
rect 289 575 803 586
rect 1049 588 1565 634
rect 476 331 568 575
rect 862 506 919 517
rect 862 366 873 506
rect 1049 412 1095 588
rect 2829 838 2875 918
rect 2441 687 2487 698
rect 2625 737 2671 748
rect 1855 597 2217 632
rect 1809 586 2217 597
rect 2263 586 2274 632
rect 3739 918 4150 926
rect 3693 775 3739 786
rect 4196 918 4589 926
rect 4150 775 4196 786
rect 4635 918 4704 926
rect 4589 775 4635 786
rect 2829 687 2875 698
rect 3033 737 3079 748
rect 2671 597 3033 632
rect 3257 739 3303 750
rect 2625 586 3079 597
rect 3125 599 3257 634
rect 3927 726 3973 737
rect 3303 599 3847 634
rect 3125 588 3847 599
rect 1565 575 1611 586
rect 919 366 1095 412
rect 1141 523 1357 542
rect 3125 540 3171 588
rect 1187 383 1357 523
rect 1690 494 1701 540
rect 1747 494 3171 540
rect 3393 523 3706 542
rect 3439 477 3706 523
rect 3393 466 3706 477
rect 3801 506 3847 588
rect 4375 726 4421 737
rect 3973 586 4375 621
rect 3927 575 4421 586
rect 1466 384 1477 430
rect 1523 384 2325 430
rect 2371 384 3141 430
rect 3187 384 3198 430
rect 1141 372 1357 383
rect 289 320 783 331
rect 65 222 111 233
rect 0 82 65 90
rect 335 285 737 320
rect 289 169 335 180
rect 513 222 559 233
rect 111 82 513 90
rect 1049 309 1095 366
rect 2382 354 2434 384
rect 3277 366 3801 401
rect 3277 355 3847 366
rect 1789 320 2283 335
rect 1049 263 1565 309
rect 1611 263 1622 309
rect 1835 289 2237 320
rect 1789 263 1835 274
rect 2237 263 2283 274
rect 2605 320 3099 335
rect 2651 289 3053 320
rect 2605 263 2651 274
rect 3053 263 3099 274
rect 3277 320 3323 355
rect 4145 331 4237 575
rect 3277 263 3323 274
rect 3937 320 4431 331
rect 737 169 783 180
rect 961 222 1007 233
rect 559 82 961 90
rect 2013 232 2059 243
rect 2013 90 2059 186
rect 2461 232 2507 243
rect 2461 90 2507 186
rect 2829 232 2875 243
rect 2829 90 2875 186
rect 3713 222 3759 233
rect 1007 82 3713 90
rect 3983 285 4385 320
rect 3937 169 3983 180
rect 4161 222 4207 233
rect 3759 82 4161 90
rect 4385 169 4431 180
rect 4609 222 4655 233
rect 4207 82 4609 90
rect 4655 82 4704 90
rect 0 -90 4704 82
<< labels >>
flabel metal1 s 1141 372 1357 542 0 FreeSans 200 0 0 0 A
port 1 nsew default input
flabel metal1 s 3393 466 3706 542 0 FreeSans 200 0 0 0 B
port 2 nsew default input
flabel metal1 s 1466 384 3198 430 0 FreeSans 200 0 0 0 CI
port 3 nsew default input
flabel metal1 s 4375 621 4421 737 0 FreeSans 200 0 0 0 CO
port 4 nsew default output
flabel metal1 s 757 621 803 737 0 FreeSans 200 0 0 0 S
port 5 nsew default output
flabel metal1 s 0 918 4704 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2829 233 2875 243 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2382 354 2434 384 1 CI
port 3 nsew default input
rlabel metal1 s 3927 621 3973 737 1 CO
port 4 nsew default output
rlabel metal1 s 3927 575 4421 621 1 CO
port 4 nsew default output
rlabel metal1 s 4145 331 4237 575 1 CO
port 4 nsew default output
rlabel metal1 s 3937 285 4431 331 1 CO
port 4 nsew default output
rlabel metal1 s 4385 169 4431 285 1 CO
port 4 nsew default output
rlabel metal1 s 3937 169 3983 285 1 CO
port 4 nsew default output
rlabel metal1 s 289 621 335 737 1 S
port 5 nsew default output
rlabel metal1 s 289 575 803 621 1 S
port 5 nsew default output
rlabel metal1 s 476 331 568 575 1 S
port 5 nsew default output
rlabel metal1 s 289 285 783 331 1 S
port 5 nsew default output
rlabel metal1 s 737 169 783 285 1 S
port 5 nsew default output
rlabel metal1 s 289 169 335 285 1 S
port 5 nsew default output
rlabel metal1 s 4589 781 4635 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4150 781 4196 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 781 3739 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2829 781 2875 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2441 781 2487 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2013 781 2059 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 981 781 1027 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 511 781 557 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 65 781 111 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4589 775 4635 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4150 775 4196 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 775 3739 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2829 775 2875 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2441 775 2487 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 981 775 1027 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 511 775 557 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 65 775 111 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2829 687 2875 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2441 687 2487 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2461 233 2507 243 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2013 233 2059 243 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4609 90 4655 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4161 90 4207 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3713 90 3759 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2829 90 2875 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2461 90 2507 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2013 90 2059 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 961 90 1007 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 513 90 559 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 65 90 111 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4704 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 1008
string GDS_END 1082910
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1073182
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
