magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 5936 844
rect 252 569 320 724
rect 1050 661 1118 724
rect 1620 670 1688 724
rect 2702 672 2770 724
rect 141 119 206 430
rect 273 60 319 232
rect 365 119 430 430
rect 682 354 886 430
rect 1242 354 1558 430
rect 3197 586 3243 724
rect 3986 532 4054 724
rect 4457 506 4503 724
rect 1090 60 1158 95
rect 1614 60 1682 95
rect 2770 60 2838 183
rect 4865 506 4911 724
rect 5062 458 5128 676
rect 5276 506 5322 724
rect 5488 458 5582 676
rect 5714 506 5760 724
rect 5062 411 5582 458
rect 4015 242 4246 318
rect 4390 60 4436 204
rect 5488 269 5582 411
rect 4838 60 4884 229
rect 5062 223 5582 269
rect 5062 161 5108 223
rect 5275 60 5343 150
rect 5488 119 5582 223
rect 5734 60 5780 229
rect 0 -60 5936 60
<< obsm1 >>
rect 49 523 95 628
rect 1164 632 1558 678
rect 1164 615 1210 632
rect 654 569 1210 615
rect 1512 624 1558 632
rect 1773 624 2170 659
rect 1512 613 2170 624
rect 1512 578 1819 613
rect 1357 532 1414 567
rect 49 477 1013 523
rect 1357 486 1809 532
rect 1879 499 1999 567
rect 2102 531 2170 613
rect 2422 626 2490 671
rect 2864 632 3142 678
rect 2864 626 2910 632
rect 49 156 95 477
rect 520 421 566 477
rect 945 291 1013 477
rect 1763 279 1809 486
rect 1302 233 1809 279
rect 1942 456 1999 499
rect 1942 409 2258 456
rect 654 187 722 219
rect 1302 198 1370 233
rect 1942 198 2010 409
rect 2317 392 2363 603
rect 2422 580 2910 626
rect 2982 485 3050 556
rect 3096 540 3142 632
rect 3340 608 3598 662
rect 3340 540 3386 608
rect 3096 493 3386 540
rect 2570 438 3050 485
rect 2993 408 3050 438
rect 3434 408 3502 562
rect 3649 421 3695 578
rect 2317 345 2934 392
rect 2993 361 3502 408
rect 3562 375 3695 421
rect 3853 486 3899 578
rect 4201 486 4247 567
rect 3853 440 4247 486
rect 654 152 1250 187
rect 1522 152 1863 187
rect 2133 152 2179 194
rect 654 141 2179 152
rect 1204 106 1568 141
rect 1817 106 2179 141
rect 2357 136 2403 345
rect 2462 252 2995 299
rect 2949 152 2995 252
rect 3206 198 3274 361
rect 3562 244 3608 375
rect 3853 244 3899 440
rect 4661 439 4707 676
rect 4306 393 4707 439
rect 4614 361 4707 393
rect 3430 198 3608 244
rect 3654 198 3954 244
rect 4298 290 4555 337
rect 4614 315 5421 361
rect 3562 152 3608 198
rect 4298 152 4344 290
rect 2949 106 3362 152
rect 3562 106 4344 152
rect 4614 161 4660 315
<< labels >>
rlabel metal1 s 682 354 886 430 6 D
port 1 nsew default input
rlabel metal1 s 141 119 206 430 6 SE
port 2 nsew default input
rlabel metal1 s 4015 242 4246 318 6 SETN
port 3 nsew default input
rlabel metal1 s 365 119 430 430 6 SI
port 4 nsew default input
rlabel metal1 s 1242 354 1558 430 6 CLK
port 5 nsew clock input
rlabel metal1 s 5488 458 5582 676 6 Q
port 6 nsew default output
rlabel metal1 s 5062 458 5128 676 6 Q
port 6 nsew default output
rlabel metal1 s 5062 411 5582 458 6 Q
port 6 nsew default output
rlabel metal1 s 5488 269 5582 411 6 Q
port 6 nsew default output
rlabel metal1 s 5062 223 5582 269 6 Q
port 6 nsew default output
rlabel metal1 s 5488 161 5582 223 6 Q
port 6 nsew default output
rlabel metal1 s 5062 161 5108 223 6 Q
port 6 nsew default output
rlabel metal1 s 5488 119 5582 161 6 Q
port 6 nsew default output
rlabel metal1 s 0 724 5936 844 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 672 5760 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 672 5322 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 672 4911 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 672 4503 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 672 4054 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 672 3243 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2702 672 2770 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1620 672 1688 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 672 1118 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 672 320 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 670 5760 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 670 5322 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 670 4911 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 670 4503 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 670 4054 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 670 3243 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1620 670 1688 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 670 1118 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 672 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 661 5760 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 661 5322 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 661 4911 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 661 4503 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 661 4054 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 661 3243 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1050 661 1118 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 661 320 670 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 586 5760 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 586 5322 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 586 4911 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 586 4503 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 586 4054 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3197 586 3243 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 586 320 661 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 569 5760 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 569 5322 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 569 4911 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 569 4503 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 569 4054 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 586 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 532 5760 569 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 532 5322 569 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 532 4911 569 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 532 4503 569 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3986 532 4054 569 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5714 506 5760 532 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 5276 506 5322 532 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4865 506 4911 532 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4457 506 4503 532 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 273 229 319 232 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5734 204 5780 229 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4838 204 4884 229 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 204 319 229 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5734 183 5780 204 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4838 183 4884 204 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4390 183 4436 204 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 204 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5734 150 5780 183 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4838 150 4884 183 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4390 150 4436 183 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2770 150 2838 183 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 150 319 183 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5734 95 5780 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5275 95 5343 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4838 95 4884 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4390 95 4436 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2770 95 2838 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 95 319 150 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5734 60 5780 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 5275 60 5343 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4838 60 4884 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4390 60 4436 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2770 60 2838 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1614 60 1682 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1090 60 1158 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 95 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5936 60 8 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5936 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 310126
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 298366
<< end >>
