magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 568 894
<< polysilicon >>
rect -31 754 88 826
rect 193 754 312 826
rect -31 -74 88 -1
rect 193 -74 312 -1
use pmos_5p04310590878177_256x8m81  pmos_5p04310590878177_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 874
<< properties >>
string GDS_END 1066946
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1066504
<< end >>
