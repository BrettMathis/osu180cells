magic
tech gf180mcuB
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -143 448 143 453
rect -143 420 -138 448
rect -110 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 110 448
rect 138 420 143 448
rect -143 386 143 420
rect -143 358 -138 386
rect -110 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 110 386
rect 138 358 143 386
rect -143 324 143 358
rect -143 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 143 324
rect -143 262 143 296
rect -143 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 143 262
rect -143 200 143 234
rect -143 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 143 200
rect -143 138 143 172
rect -143 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 143 138
rect -143 76 143 110
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -110 143 -76
rect -143 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 143 -110
rect -143 -172 143 -138
rect -143 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 143 -172
rect -143 -234 143 -200
rect -143 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 143 -234
rect -143 -296 143 -262
rect -143 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 143 -296
rect -143 -358 143 -324
rect -143 -386 -138 -358
rect -110 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 110 -358
rect 138 -386 143 -358
rect -143 -420 143 -386
rect -143 -448 -138 -420
rect -110 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 110 -420
rect 138 -448 143 -420
rect -143 -453 143 -448
<< via2 >>
rect -138 420 -110 448
rect -76 420 -48 448
rect -14 420 14 448
rect 48 420 76 448
rect 110 420 138 448
rect -138 358 -110 386
rect -76 358 -48 386
rect -14 358 14 386
rect 48 358 76 386
rect 110 358 138 386
rect -138 296 -110 324
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect 110 296 138 324
rect -138 234 -110 262
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect 110 234 138 262
rect -138 172 -110 200
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect 110 172 138 200
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect -138 -200 -110 -172
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect 110 -200 138 -172
rect -138 -262 -110 -234
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect 110 -262 138 -234
rect -138 -324 -110 -296
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect 110 -324 138 -296
rect -138 -386 -110 -358
rect -76 -386 -48 -358
rect -14 -386 14 -358
rect 48 -386 76 -358
rect 110 -386 138 -358
rect -138 -448 -110 -420
rect -76 -448 -48 -420
rect -14 -448 14 -420
rect 48 -448 76 -420
rect 110 -448 138 -420
<< metal3 >>
rect -143 448 143 453
rect -143 420 -138 448
rect -110 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 110 448
rect 138 420 143 448
rect -143 386 143 420
rect -143 358 -138 386
rect -110 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 110 386
rect 138 358 143 386
rect -143 324 143 358
rect -143 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 143 324
rect -143 262 143 296
rect -143 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 143 262
rect -143 200 143 234
rect -143 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 143 200
rect -143 138 143 172
rect -143 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 143 138
rect -143 76 143 110
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -110 143 -76
rect -143 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 143 -110
rect -143 -172 143 -138
rect -143 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 143 -172
rect -143 -234 143 -200
rect -143 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 143 -234
rect -143 -296 143 -262
rect -143 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 143 -296
rect -143 -358 143 -324
rect -143 -386 -138 -358
rect -110 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 110 -358
rect 138 -386 143 -358
rect -143 -420 143 -386
rect -143 -448 -138 -420
rect -110 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 110 -420
rect 138 -448 143 -420
rect -143 -453 143 -448
<< properties >>
string GDS_END 2281524
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2276592
<< end >>
