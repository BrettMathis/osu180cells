magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -183 117 183 136
rect -183 -117 -164 117
rect 164 -117 183 117
rect -183 -136 183 -117
<< psubdiffcont >>
rect -164 -117 164 117
<< metal1 >>
rect -175 117 175 128
rect -175 -117 -164 117
rect 164 -117 175 117
rect -175 -128 175 -117
<< properties >>
string GDS_END 383080
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 382116
<< end >>
