magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -81 169 81 174
rect -81 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 81 169
rect -81 107 81 141
rect -81 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 81 107
rect -81 45 81 79
rect -81 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 81 45
rect -81 -17 81 17
rect -81 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 81 -17
rect -81 -79 81 -45
rect -81 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 81 -79
rect -81 -141 81 -107
rect -81 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 81 -141
rect -81 -174 81 -169
<< via2 >>
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
<< metal3 >>
rect -81 169 81 174
rect -81 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 81 169
rect -81 107 81 141
rect -81 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 81 107
rect -81 45 81 79
rect -81 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 81 45
rect -81 -17 81 17
rect -81 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 81 -17
rect -81 -79 81 -45
rect -81 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 81 -79
rect -81 -141 81 -107
rect -81 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 81 -141
rect -81 -174 81 -169
<< properties >>
string GDS_END 670932
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 669648
<< end >>
