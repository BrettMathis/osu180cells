magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 6944 844
rect 49 506 95 724
rect 477 600 523 724
rect 925 600 971 724
rect 1373 600 1419 724
rect 1821 600 1867 724
rect 2269 506 2315 724
rect 2513 600 2559 676
rect 2717 646 2763 724
rect 2941 600 2987 676
rect 3165 646 3211 724
rect 3389 600 3435 676
rect 3613 646 3659 724
rect 3837 600 3883 676
rect 4061 646 4107 724
rect 4285 600 4331 676
rect 4509 646 4555 724
rect 4733 600 4779 676
rect 4957 646 5003 724
rect 5181 600 5227 676
rect 5405 646 5451 724
rect 5629 600 5675 676
rect 5853 646 5899 724
rect 6077 600 6123 676
rect 6301 646 6347 724
rect 6525 600 6571 676
rect 126 348 1980 430
rect 2513 454 6571 600
rect 6749 506 6795 724
rect 4446 302 4626 454
rect 49 60 95 232
rect 497 60 543 192
rect 945 60 991 192
rect 1393 60 1439 192
rect 1841 60 1887 192
rect 2289 60 2335 192
rect 2513 173 6591 302
rect 2513 135 2565 173
rect 2961 135 3007 173
rect 3409 135 3455 173
rect 3857 135 3903 173
rect 4305 135 4351 173
rect 4753 135 4799 173
rect 5201 135 5247 173
rect 5649 135 5695 173
rect 6097 135 6143 173
rect 6545 135 6591 173
rect 2726 60 2794 127
rect 3174 60 3242 127
rect 3622 60 3690 127
rect 4070 60 4138 127
rect 4518 60 4586 127
rect 4966 60 5034 127
rect 5414 60 5482 127
rect 5862 60 5930 127
rect 6310 60 6378 127
rect 6769 60 6815 232
rect 0 -60 6944 60
<< obsm1 >>
rect 273 552 319 676
rect 701 552 747 676
rect 1149 552 1195 676
rect 1597 552 1643 676
rect 2045 552 2136 676
rect 273 506 2136 552
rect 2045 394 2136 506
rect 2045 348 4314 394
rect 2045 284 2136 348
rect 4736 348 6720 394
rect 273 238 2136 284
rect 273 135 319 238
rect 721 135 767 238
rect 1169 135 1215 238
rect 1617 135 1663 238
rect 2065 135 2136 238
<< labels >>
rlabel metal1 s 126 348 1980 430 6 I
port 1 nsew default input
rlabel metal1 s 6525 600 6571 676 6 Z
port 2 nsew default output
rlabel metal1 s 6077 600 6123 676 6 Z
port 2 nsew default output
rlabel metal1 s 5629 600 5675 676 6 Z
port 2 nsew default output
rlabel metal1 s 5181 600 5227 676 6 Z
port 2 nsew default output
rlabel metal1 s 4733 600 4779 676 6 Z
port 2 nsew default output
rlabel metal1 s 4285 600 4331 676 6 Z
port 2 nsew default output
rlabel metal1 s 3837 600 3883 676 6 Z
port 2 nsew default output
rlabel metal1 s 3389 600 3435 676 6 Z
port 2 nsew default output
rlabel metal1 s 2941 600 2987 676 6 Z
port 2 nsew default output
rlabel metal1 s 2513 600 2559 676 6 Z
port 2 nsew default output
rlabel metal1 s 2513 454 6571 600 6 Z
port 2 nsew default output
rlabel metal1 s 4446 302 4626 454 6 Z
port 2 nsew default output
rlabel metal1 s 2513 173 6591 302 6 Z
port 2 nsew default output
rlabel metal1 s 6545 135 6591 173 6 Z
port 2 nsew default output
rlabel metal1 s 6097 135 6143 173 6 Z
port 2 nsew default output
rlabel metal1 s 5649 135 5695 173 6 Z
port 2 nsew default output
rlabel metal1 s 5201 135 5247 173 6 Z
port 2 nsew default output
rlabel metal1 s 4753 135 4799 173 6 Z
port 2 nsew default output
rlabel metal1 s 4305 135 4351 173 6 Z
port 2 nsew default output
rlabel metal1 s 3857 135 3903 173 6 Z
port 2 nsew default output
rlabel metal1 s 3409 135 3455 173 6 Z
port 2 nsew default output
rlabel metal1 s 2961 135 3007 173 6 Z
port 2 nsew default output
rlabel metal1 s 2513 135 2565 173 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 6944 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 646 6795 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6301 646 6347 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5853 646 5899 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 646 5451 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 646 5003 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 646 4555 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 646 4107 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 646 3659 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 646 3211 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 646 2763 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 646 2315 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 646 1867 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 600 6795 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 600 2315 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 600 1867 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 600 1419 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 600 971 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 600 523 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 600 95 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 506 6795 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 506 2315 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6769 192 6815 232 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 192 95 232 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6769 127 6815 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 127 2335 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 127 1887 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 127 1439 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 127 991 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 127 543 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6769 60 6815 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6310 60 6378 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5862 60 5930 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5414 60 5482 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4966 60 5034 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4518 60 4586 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6944 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6944 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1359712
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1345148
<< end >>
