magic
tech gf180mcuC
timestamp 1669390400
<< properties >>
string GDS_END 500810
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 500550
<< end >>
