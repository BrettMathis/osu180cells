magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 896 844
rect 49 506 95 724
rect 273 536 319 678
rect 497 597 543 724
rect 682 536 767 678
rect 273 472 767 536
rect 82 352 603 424
rect 682 305 767 472
rect 273 258 767 305
rect 49 60 95 232
rect 273 106 319 258
rect 497 60 543 211
rect 682 106 767 258
rect 0 -60 896 60
<< labels >>
rlabel metal1 s 82 352 603 424 6 I
port 1 nsew default input
rlabel metal1 s 682 536 767 678 6 ZN
port 2 nsew default output
rlabel metal1 s 273 536 319 678 6 ZN
port 2 nsew default output
rlabel metal1 s 273 472 767 536 6 ZN
port 2 nsew default output
rlabel metal1 s 682 305 767 472 6 ZN
port 2 nsew default output
rlabel metal1 s 273 258 767 305 6 ZN
port 2 nsew default output
rlabel metal1 s 682 106 767 258 6 ZN
port 2 nsew default output
rlabel metal1 s 273 106 319 258 6 ZN
port 2 nsew default output
rlabel metal1 s 0 724 896 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 497 597 543 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 597 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 597 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 211 95 232 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 211 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 896 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 472800
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 469932
<< end >>
