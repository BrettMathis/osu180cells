magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 5014 1094
<< pwell >>
rect -86 -86 5014 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 215 836 333
rect 940 215 1060 333
rect 1164 215 1284 333
rect 1332 215 1452 333
rect 1532 215 1652 333
rect 1940 215 2060 333
rect 2108 215 2228 333
rect 2332 215 2452 333
rect 2556 215 2676 333
rect 3041 175 3161 333
rect 3209 175 3329 333
rect 3433 175 3553 333
rect 3601 175 3721 333
rect 3969 69 4089 333
rect 4193 69 4313 333
rect 4417 69 4537 333
rect 4641 69 4761 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 716 573 816 773
rect 920 573 1020 773
rect 1124 573 1224 773
rect 1332 573 1432 773
rect 1612 690 1712 890
rect 1960 690 2060 890
rect 2252 573 2352 773
rect 2456 573 2556 773
rect 2660 573 2760 773
rect 3025 575 3125 851
rect 3229 575 3329 851
rect 3433 575 3533 851
rect 3637 575 3737 851
rect 3989 573 4089 939
rect 4193 573 4293 939
rect 4397 573 4497 939
rect 4601 573 4701 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 274 716 333
rect 628 228 641 274
rect 687 228 716 274
rect 628 215 716 228
rect 836 320 940 333
rect 836 274 865 320
rect 911 274 940 320
rect 836 215 940 274
rect 1060 320 1164 333
rect 1060 274 1089 320
rect 1135 274 1164 320
rect 1060 215 1164 274
rect 1284 215 1332 333
rect 1452 215 1532 333
rect 1652 274 1940 333
rect 1652 228 1681 274
rect 1727 228 1940 274
rect 1652 215 1940 228
rect 2060 215 2108 333
rect 2228 320 2332 333
rect 2228 274 2257 320
rect 2303 274 2332 320
rect 2228 215 2332 274
rect 2452 320 2556 333
rect 2452 274 2481 320
rect 2527 274 2556 320
rect 2452 215 2556 274
rect 2676 320 2764 333
rect 2676 274 2705 320
rect 2751 274 2764 320
rect 2676 215 2764 274
rect 2953 308 3041 333
rect 2953 262 2966 308
rect 3012 262 3041 308
rect 2953 175 3041 262
rect 3161 175 3209 333
rect 3329 234 3433 333
rect 3329 188 3358 234
rect 3404 188 3433 234
rect 3329 175 3433 188
rect 3553 175 3601 333
rect 3721 320 3809 333
rect 3721 274 3750 320
rect 3796 274 3809 320
rect 3721 175 3809 274
rect 3881 222 3969 333
rect 3881 82 3894 222
rect 3940 82 3969 222
rect 3881 69 3969 82
rect 4089 320 4193 333
rect 4089 180 4118 320
rect 4164 180 4193 320
rect 4089 69 4193 180
rect 4313 222 4417 333
rect 4313 82 4342 222
rect 4388 82 4417 222
rect 4313 69 4417 82
rect 4537 314 4641 333
rect 4537 174 4566 314
rect 4612 174 4641 314
rect 4537 69 4641 174
rect 4761 222 4849 333
rect 4761 82 4790 222
rect 4836 82 4849 222
rect 4761 69 4849 82
<< mvpdiff >>
rect 1480 955 1552 968
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 1480 909 1493 955
rect 1539 909 1552 955
rect 2120 955 2192 968
rect 1480 896 1552 909
rect 1492 890 1552 896
rect 2120 909 2133 955
rect 2179 909 2192 955
rect 2120 890 2192 909
rect 1492 773 1612 890
rect 448 586 477 726
rect 523 586 536 726
rect 448 573 536 586
rect 628 760 716 773
rect 628 714 641 760
rect 687 714 716 760
rect 628 573 716 714
rect 816 726 920 773
rect 816 586 845 726
rect 891 586 920 726
rect 816 573 920 586
rect 1020 726 1124 773
rect 1020 586 1049 726
rect 1095 586 1124 726
rect 1020 573 1124 586
rect 1224 727 1332 773
rect 1224 681 1257 727
rect 1303 681 1332 727
rect 1224 573 1332 681
rect 1432 690 1612 773
rect 1712 749 1800 890
rect 1712 703 1741 749
rect 1787 703 1800 749
rect 1712 690 1800 703
rect 1872 749 1960 890
rect 1872 703 1885 749
rect 1931 703 1960 749
rect 1872 690 1960 703
rect 2060 773 2192 890
rect 3901 926 3989 939
rect 2937 838 3025 851
rect 2937 792 2950 838
rect 2996 792 3025 838
rect 2060 690 2252 773
rect 1432 573 1512 690
rect 2172 573 2252 690
rect 2352 726 2456 773
rect 2352 586 2381 726
rect 2427 586 2456 726
rect 2352 573 2456 586
rect 2556 726 2660 773
rect 2556 586 2585 726
rect 2631 586 2660 726
rect 2556 573 2660 586
rect 2760 632 2848 773
rect 2760 586 2789 632
rect 2835 586 2848 632
rect 2760 573 2848 586
rect 2937 575 3025 792
rect 3125 634 3229 851
rect 3125 588 3154 634
rect 3200 588 3229 634
rect 3125 575 3229 588
rect 3329 838 3433 851
rect 3329 792 3358 838
rect 3404 792 3433 838
rect 3329 575 3433 792
rect 3533 634 3637 851
rect 3533 588 3562 634
rect 3608 588 3637 634
rect 3533 575 3637 588
rect 3737 838 3825 851
rect 3737 698 3766 838
rect 3812 698 3825 838
rect 3737 575 3825 698
rect 3901 786 3914 926
rect 3960 786 3989 926
rect 3901 573 3989 786
rect 4089 726 4193 939
rect 4089 586 4118 726
rect 4164 586 4193 726
rect 4089 573 4193 586
rect 4293 926 4397 939
rect 4293 786 4322 926
rect 4368 786 4397 926
rect 4293 573 4397 786
rect 4497 726 4601 939
rect 4497 586 4526 726
rect 4572 586 4601 726
rect 4497 573 4601 586
rect 4701 926 4789 939
rect 4701 786 4730 926
rect 4776 786 4789 926
rect 4701 573 4789 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 228 687 274
rect 865 274 911 320
rect 1089 274 1135 320
rect 1681 228 1727 274
rect 2257 274 2303 320
rect 2481 274 2527 320
rect 2705 274 2751 320
rect 2966 262 3012 308
rect 3358 188 3404 234
rect 3750 274 3796 320
rect 3894 82 3940 222
rect 4118 180 4164 320
rect 4342 82 4388 222
rect 4566 174 4612 314
rect 4790 82 4836 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 1493 909 1539 955
rect 2133 909 2179 955
rect 477 586 523 726
rect 641 714 687 760
rect 845 586 891 726
rect 1049 586 1095 726
rect 1257 681 1303 727
rect 1741 703 1787 749
rect 1885 703 1931 749
rect 2950 792 2996 838
rect 2381 586 2427 726
rect 2585 586 2631 726
rect 2789 586 2835 632
rect 3154 588 3200 634
rect 3358 792 3404 838
rect 3562 588 3608 634
rect 3766 698 3812 838
rect 3914 786 3960 926
rect 4118 586 4164 726
rect 4322 786 4368 926
rect 4526 586 4572 726
rect 4730 786 4776 926
<< polysilicon >>
rect 348 909 1020 949
rect 144 849 244 893
rect 348 849 448 909
rect 716 773 816 817
rect 920 773 1020 909
rect 1612 890 1712 934
rect 1960 890 2060 934
rect 1124 852 1224 865
rect 1124 806 1137 852
rect 1183 806 1224 852
rect 1124 773 1224 806
rect 1332 773 1432 817
rect 2252 913 3125 953
rect 3989 939 4089 983
rect 4193 939 4293 983
rect 4397 939 4497 983
rect 4601 939 4701 983
rect 2252 773 2352 913
rect 2456 852 2556 865
rect 2456 806 2469 852
rect 2515 806 2556 852
rect 3025 851 3125 913
rect 3229 851 3329 895
rect 3433 851 3533 895
rect 3637 851 3737 895
rect 2456 773 2556 806
rect 2660 773 2760 817
rect 1612 646 1712 690
rect 144 516 244 573
rect 144 470 157 516
rect 203 470 244 516
rect 144 377 244 470
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 716 523 816 573
rect 920 529 1020 573
rect 1124 529 1224 573
rect 716 477 729 523
rect 775 477 816 523
rect 716 377 816 477
rect 1124 465 1164 529
rect 940 425 1164 465
rect 1332 480 1432 573
rect 1332 434 1373 480
rect 1419 434 1432 480
rect 407 366 468 377
rect 348 333 468 366
rect 716 333 836 377
rect 940 333 1060 425
rect 1212 412 1284 425
rect 1212 377 1225 412
rect 1164 366 1225 377
rect 1271 366 1284 412
rect 1164 333 1284 366
rect 1332 377 1432 434
rect 1612 377 1652 646
rect 1960 572 2060 690
rect 1960 526 1973 572
rect 2019 526 2060 572
rect 1960 377 2060 526
rect 2252 513 2352 573
rect 1332 333 1452 377
rect 1532 333 1652 377
rect 1940 333 2060 377
rect 2108 473 2352 513
rect 2456 513 2556 573
rect 2660 529 2760 573
rect 3025 542 3125 575
rect 3025 531 3054 542
rect 2456 473 2596 513
rect 2108 333 2228 473
rect 2556 377 2596 473
rect 2720 437 2760 529
rect 3041 496 3054 531
rect 3100 496 3125 542
rect 2720 397 2893 437
rect 2332 333 2452 377
rect 2556 333 2676 377
rect 124 131 244 175
rect 348 115 468 175
rect 716 171 836 215
rect 940 171 1060 215
rect 1164 115 1284 215
rect 1332 171 1452 215
rect 348 75 1284 115
rect 1532 75 1652 215
rect 1940 171 2060 215
rect 2108 171 2228 215
rect 2332 182 2452 215
rect 2332 136 2345 182
rect 2391 136 2452 182
rect 2556 171 2676 215
rect 2824 190 2893 397
rect 3041 377 3125 496
rect 3229 412 3329 575
rect 3229 377 3270 412
rect 3041 333 3161 377
rect 3209 366 3270 377
rect 3316 366 3329 412
rect 3209 333 3329 366
rect 3433 542 3533 575
rect 3433 496 3446 542
rect 3492 496 3533 542
rect 3433 377 3533 496
rect 3637 542 3737 575
rect 3637 496 3654 542
rect 3700 496 3737 542
rect 3637 483 3737 496
rect 3637 377 3721 483
rect 3989 465 4089 573
rect 4193 465 4293 573
rect 4397 465 4497 573
rect 4601 465 4701 573
rect 3989 447 4701 465
rect 3989 401 4002 447
rect 4048 401 4221 447
rect 4267 401 4430 447
rect 4476 401 4701 447
rect 3989 393 4701 401
rect 3989 377 4089 393
rect 3433 333 3553 377
rect 3601 333 3721 377
rect 3969 333 4089 377
rect 4193 333 4313 393
rect 4417 333 4537 393
rect 4641 377 4701 393
rect 4641 333 4761 377
rect 2821 182 2893 190
rect 2332 123 2452 136
rect 2821 136 2834 182
rect 2880 136 2893 182
rect 2821 123 2893 136
rect 3041 131 3161 175
rect 3209 131 3329 175
rect 3433 75 3553 175
rect 3601 131 3721 175
rect 1532 35 3553 75
rect 3969 25 4089 69
rect 4193 25 4313 69
rect 4417 25 4537 69
rect 4641 25 4761 69
<< polycontact >>
rect 1137 806 1183 852
rect 2469 806 2515 852
rect 157 470 203 516
rect 361 366 407 412
rect 729 477 775 523
rect 1373 434 1419 480
rect 1225 366 1271 412
rect 1973 526 2019 572
rect 3054 496 3100 542
rect 2345 136 2391 182
rect 3270 366 3316 412
rect 3446 496 3492 542
rect 3654 496 3700 542
rect 4002 401 4048 447
rect 4221 401 4267 447
rect 4430 401 4476 447
rect 2834 136 2880 182
<< metal1 >>
rect 0 955 4928 1098
rect 0 918 1493 955
rect 273 836 319 918
rect 69 739 115 750
rect 641 760 687 918
rect 1539 918 2133 955
rect 1493 898 1539 909
rect 2179 926 4928 955
rect 2179 918 3914 926
rect 2133 898 2179 909
rect 273 685 319 696
rect 477 726 523 737
rect 115 599 407 634
rect 69 588 407 599
rect 142 516 314 542
rect 142 470 157 516
rect 203 470 314 516
rect 142 459 314 470
rect 361 412 407 588
rect 49 366 361 401
rect 49 355 407 366
rect 641 703 687 714
rect 733 806 1137 852
rect 1183 806 2469 852
rect 2515 806 2526 852
rect 2939 838 3007 918
rect 733 657 779 806
rect 2939 792 2950 838
rect 2996 792 3007 838
rect 3347 838 3415 918
rect 3347 792 3358 838
rect 3404 792 3415 838
rect 3766 838 3812 918
rect 1257 749 1787 760
rect 523 611 779 657
rect 845 726 911 737
rect 523 586 543 611
rect 49 320 95 355
rect 49 263 95 274
rect 477 320 543 586
rect 891 586 911 726
rect 611 523 778 542
rect 611 477 729 523
rect 775 477 778 523
rect 611 466 778 477
rect 477 274 497 320
rect 845 320 911 586
rect 477 263 543 274
rect 641 274 687 285
rect 273 234 319 245
rect 273 90 319 188
rect 845 274 865 320
rect 845 263 911 274
rect 1049 726 1095 737
rect 1257 727 1741 749
rect 1303 703 1741 727
rect 1303 681 1787 703
rect 1885 749 2427 760
rect 1931 726 2427 749
rect 1931 714 2381 726
rect 1931 703 2303 714
rect 1885 692 2303 703
rect 1257 670 1787 681
rect 1049 583 1095 586
rect 1049 572 2019 583
rect 1049 537 1973 572
rect 1049 320 1135 537
rect 1973 515 2019 526
rect 1373 480 1419 491
rect 2257 469 2303 692
rect 2381 575 2427 586
rect 2585 726 3700 746
rect 2631 700 3700 726
rect 1419 434 2303 469
rect 1373 423 2303 434
rect 1225 412 1271 423
rect 1271 366 2211 377
rect 1225 331 2211 366
rect 1049 274 1089 320
rect 1049 263 1135 274
rect 1681 274 1727 285
rect 641 90 687 228
rect 1681 90 1727 228
rect 2165 182 2211 331
rect 2257 320 2303 423
rect 2585 331 2631 586
rect 2789 632 2835 643
rect 2789 331 2835 586
rect 3154 634 3200 645
rect 3054 542 3106 553
rect 3100 496 3106 542
rect 3054 354 3106 496
rect 2257 263 2303 274
rect 2481 320 2631 331
rect 2527 274 2631 320
rect 2481 263 2631 274
rect 2705 320 2835 331
rect 2751 308 2835 320
rect 3154 308 3200 588
rect 3390 542 3442 654
rect 3562 634 3608 645
rect 3390 496 3446 542
rect 3492 496 3503 542
rect 3562 423 3608 588
rect 3654 542 3700 700
rect 3960 918 4322 926
rect 3914 775 3960 786
rect 4368 918 4730 926
rect 4322 775 4368 786
rect 4776 918 4928 926
rect 4730 775 4776 786
rect 3766 687 3812 698
rect 4118 726 4164 737
rect 4526 726 4612 737
rect 4164 586 4526 621
rect 4572 586 4612 726
rect 4118 575 4612 586
rect 3654 485 3700 496
rect 4002 447 4487 458
rect 3562 412 4002 423
rect 3259 366 3270 412
rect 3316 401 4002 412
rect 4048 401 4221 447
rect 4267 401 4430 447
rect 4476 401 4487 447
rect 3316 366 4048 401
rect 2751 274 2966 308
rect 2705 262 2966 274
rect 3012 262 3200 308
rect 3750 355 4048 366
rect 3750 320 3796 355
rect 4533 331 4612 575
rect 3750 263 3796 274
rect 4118 320 4612 331
rect 3358 234 3404 245
rect 2165 136 2345 182
rect 2391 136 2834 182
rect 2880 136 2891 182
rect 3358 90 3404 188
rect 3894 222 3940 233
rect 0 82 3894 90
rect 4164 314 4612 320
rect 4164 279 4566 314
rect 4118 169 4164 180
rect 4342 222 4388 233
rect 3940 82 4342 90
rect 4510 174 4566 279
rect 4510 163 4612 174
rect 4790 222 4836 233
rect 4388 82 4790 90
rect 4836 82 4928 90
rect 0 -90 4928 82
<< labels >>
flabel metal1 s 142 459 314 542 0 FreeSans 200 0 0 0 CLKN
port 4 nsew clock input
flabel metal1 s 611 466 778 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4526 621 4612 737 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3390 542 3442 654 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 3054 354 3106 553 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 4928 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1681 245 1727 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3390 496 3503 542 1 RN
port 2 nsew default input
rlabel metal1 s 4118 621 4164 737 1 Q
port 5 nsew default output
rlabel metal1 s 4118 575 4612 621 1 Q
port 5 nsew default output
rlabel metal1 s 4533 331 4612 575 1 Q
port 5 nsew default output
rlabel metal1 s 4118 279 4612 331 1 Q
port 5 nsew default output
rlabel metal1 s 4510 169 4612 279 1 Q
port 5 nsew default output
rlabel metal1 s 4118 169 4164 279 1 Q
port 5 nsew default output
rlabel metal1 s 4510 163 4612 169 1 Q
port 5 nsew default output
rlabel metal1 s 4730 898 4776 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4322 898 4368 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3914 898 3960 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3766 898 3812 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3347 898 3415 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2939 898 3007 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2133 898 2179 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1493 898 1539 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 898 687 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 898 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4730 792 4776 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4322 792 4368 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3914 792 3960 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3766 792 3812 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3347 792 3415 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2939 792 3007 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 792 687 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 792 319 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4730 775 4776 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4322 775 4368 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3914 775 3960 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3766 775 3812 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 775 687 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3766 703 3812 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 703 687 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 703 319 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3766 687 3812 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 687 319 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 687 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 641 245 687 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3358 233 3404 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1681 233 1727 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4790 90 4836 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4342 90 4388 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3894 90 3940 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3358 90 3404 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1681 90 1727 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4928 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4928 1008
string GDS_END 541612
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 530856
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
