magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 -74 88 -1
rect 193 -74 312 -1
rect 417 -74 536 -1
rect 641 -74 760 -1
rect 865 -74 984 -1
use nmos_5p04310590878189_256x8m81  nmos_5p04310590878189_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 1104 2040
<< properties >>
string GDS_END 663898
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 663456
<< end >>
