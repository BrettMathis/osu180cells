magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -19 248 19 253
rect -19 -248 -14 248
rect 14 -248 19 248
rect -19 -253 19 -248
<< via2 >>
rect -14 -248 14 248
<< metal3 >>
rect -19 248 19 253
rect -19 -248 -14 248
rect 14 -248 19 248
rect -19 -253 19 -248
<< properties >>
string GDS_END 516010
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 515238
<< end >>
