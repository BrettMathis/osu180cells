magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 4775 50 5611 150
<< metal3 >>
rect 3339 1150 4353 1350
rect 3339 850 29240 1150
rect 3339 650 4353 850
rect 3339 -250 5045 450
use M2_M14310590878181_256x8m81  M2_M14310590878181_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 1000
box -162 -348 162 348
use M2_M14310590878181_256x8m81  M2_M14310590878181_256x8m81_1
timestamp 1669390400
transform 1 0 4883 0 1 100
box -162 -348 162 348
use M3_M24310590878182_256x8m81  M3_M24310590878182_256x8m81_0
timestamp 1669390400
transform 1 0 4883 0 1 100
box -162 -348 162 348
use M3_M24310590878182_256x8m81  M3_M24310590878182_256x8m81_1
timestamp 1669390400
transform 1 0 3783 0 1 1000
box -162 -348 162 348
<< properties >>
string GDS_END 1921008
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1920580
string path 25.225 0.500 16.695 0.500 
<< end >>
