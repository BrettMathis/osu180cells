magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 1720 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 850 190 910 360
rect 1020 190 1080 360
rect 1240 190 1300 360
rect 1410 190 1470 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 530 700 590 1040
rect 850 700 910 1040
rect 1020 700 1080 1040
rect 1240 700 1300 1040
rect 1410 700 1470 1040
<< ndiff >>
rect 90 278 190 360
rect 90 232 112 278
rect 158 232 190 278
rect 90 190 190 232
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 530 360
rect 590 298 690 360
rect 590 252 622 298
rect 668 252 690 298
rect 590 190 690 252
rect 750 263 850 360
rect 750 217 772 263
rect 818 217 850 263
rect 750 190 850 217
rect 910 338 1020 360
rect 910 292 942 338
rect 988 292 1020 338
rect 910 190 1020 292
rect 1080 263 1240 360
rect 1080 217 1112 263
rect 1158 217 1240 263
rect 1080 190 1240 217
rect 1300 298 1410 360
rect 1300 252 1332 298
rect 1378 252 1410 298
rect 1300 190 1410 252
rect 1470 298 1620 360
rect 1470 252 1552 298
rect 1598 252 1620 298
rect 1470 190 1620 252
<< pdiff >>
rect 90 1012 190 1040
rect 90 778 112 1012
rect 158 778 190 1012
rect 90 700 190 778
rect 250 987 360 1040
rect 250 753 282 987
rect 328 753 360 987
rect 250 700 360 753
rect 420 987 530 1040
rect 420 753 452 987
rect 498 753 530 987
rect 420 700 530 753
rect 590 987 690 1040
rect 590 753 622 987
rect 668 753 690 987
rect 590 700 690 753
rect 750 987 850 1040
rect 750 753 772 987
rect 818 753 850 987
rect 750 700 850 753
rect 910 700 1020 1040
rect 1080 987 1240 1040
rect 1080 753 1137 987
rect 1183 753 1240 987
rect 1080 700 1240 753
rect 1300 993 1410 1040
rect 1300 947 1332 993
rect 1378 947 1410 993
rect 1300 700 1410 947
rect 1470 987 1620 1040
rect 1470 753 1527 987
rect 1573 753 1620 987
rect 1470 700 1620 753
<< ndiffc >>
rect 112 232 158 278
rect 282 252 328 298
rect 622 252 668 298
rect 772 217 818 263
rect 942 292 988 338
rect 1112 217 1158 263
rect 1332 252 1378 298
rect 1552 252 1598 298
<< pdiffc >>
rect 112 778 158 1012
rect 282 753 328 987
rect 452 753 498 987
rect 622 753 668 987
rect 772 753 818 987
rect 1137 753 1183 987
rect 1332 947 1378 993
rect 1527 753 1573 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1340 98 1430 120
rect 1340 52 1362 98
rect 1408 52 1430 98
rect 1340 30 1430 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
rect 1290 1178 1380 1200
rect 1290 1132 1312 1178
rect 1358 1132 1380 1178
rect 1290 1110 1380 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1362 52 1408 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
rect 1312 1132 1358 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 850 1040 910 1090
rect 1020 1040 1080 1090
rect 1240 1040 1300 1090
rect 1410 1040 1470 1090
rect 190 670 250 700
rect 190 643 310 670
rect 190 597 237 643
rect 283 597 310 643
rect 190 570 310 597
rect 190 360 250 570
rect 360 520 420 700
rect 300 493 420 520
rect 530 510 590 700
rect 850 520 910 700
rect 300 447 327 493
rect 373 447 420 493
rect 300 420 420 447
rect 360 360 420 420
rect 470 483 590 510
rect 470 437 497 483
rect 543 437 590 483
rect 470 410 590 437
rect 780 493 910 520
rect 780 447 807 493
rect 853 447 910 493
rect 780 420 910 447
rect 530 360 590 410
rect 850 360 910 420
rect 1020 480 1080 700
rect 1240 680 1300 700
rect 1240 653 1360 680
rect 1240 607 1287 653
rect 1333 607 1360 653
rect 1240 580 1360 607
rect 1020 453 1120 480
rect 1020 407 1047 453
rect 1093 407 1120 453
rect 1020 380 1120 407
rect 1020 360 1080 380
rect 1240 360 1300 580
rect 1410 520 1470 700
rect 1350 493 1470 520
rect 1350 447 1377 493
rect 1423 447 1470 493
rect 1350 420 1470 447
rect 1410 360 1470 420
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 850 140 910 190
rect 1020 140 1080 190
rect 1240 140 1300 190
rect 1410 140 1470 190
<< polycontact >>
rect 237 597 283 643
rect 327 447 373 493
rect 497 437 543 483
rect 807 447 853 493
rect 1287 607 1333 653
rect 1047 407 1093 453
rect 1377 447 1423 493
<< metal1 >>
rect 0 1178 1720 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1312 1178
rect 1358 1176 1720 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 1126 1132 1312 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1314 1132
rect 1366 1124 1720 1176
rect 0 1110 1720 1124
rect 110 1012 160 1040
rect 110 778 112 1012
rect 158 778 160 1012
rect 110 760 160 778
rect 280 987 330 1110
rect 80 756 180 760
rect 80 704 104 756
rect 156 704 180 756
rect 80 700 180 704
rect 280 753 282 987
rect 328 753 330 987
rect 280 700 330 753
rect 450 987 500 1040
rect 450 753 452 987
rect 498 753 500 987
rect 110 278 160 700
rect 450 650 500 753
rect 620 987 670 1110
rect 620 753 622 987
rect 668 753 670 987
rect 620 700 670 753
rect 770 987 820 1110
rect 770 753 772 987
rect 818 753 820 987
rect 770 700 820 753
rect 1110 987 1210 1040
rect 1110 753 1137 987
rect 1183 753 1210 987
rect 1330 993 1380 1110
rect 1330 947 1332 993
rect 1378 947 1380 993
rect 1330 900 1380 947
rect 1500 987 1600 1040
rect 1110 700 1210 753
rect 1500 753 1527 987
rect 1573 753 1600 987
rect 1500 700 1600 753
rect 210 646 700 650
rect 210 643 624 646
rect 210 597 237 643
rect 283 597 624 643
rect 210 594 624 597
rect 676 594 700 646
rect 1110 600 1160 700
rect 1260 656 1360 660
rect 1260 604 1284 656
rect 1336 604 1360 656
rect 1550 640 1600 700
rect 1550 630 1620 640
rect 1260 600 1360 604
rect 1540 626 1640 630
rect 210 590 700 594
rect 300 496 400 500
rect 300 444 324 496
rect 376 444 400 496
rect 300 440 400 444
rect 470 483 570 490
rect 470 437 497 483
rect 543 437 570 483
rect 470 430 570 437
rect 490 370 550 430
rect 470 366 570 370
rect 110 232 112 278
rect 158 232 160 278
rect 110 190 160 232
rect 280 298 330 360
rect 470 314 494 366
rect 546 314 570 366
rect 470 310 570 314
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 620 298 670 590
rect 940 550 1210 600
rect 1540 574 1564 626
rect 1616 574 1640 626
rect 1540 570 1640 574
rect 1550 560 1620 570
rect 780 496 880 500
rect 780 444 804 496
rect 856 444 880 496
rect 780 440 880 444
rect 620 252 622 298
rect 668 252 670 298
rect 940 338 990 550
rect 1150 500 1350 550
rect 1300 493 1450 500
rect 1040 456 1100 480
rect 1040 404 1044 456
rect 1096 404 1100 456
rect 1300 447 1377 493
rect 1423 447 1450 493
rect 1300 440 1450 447
rect 1040 380 1100 404
rect 940 292 942 338
rect 988 292 990 338
rect 620 190 670 252
rect 770 263 820 290
rect 940 270 990 292
rect 1330 298 1380 360
rect 770 217 772 263
rect 818 220 820 263
rect 1110 263 1160 290
rect 1110 220 1112 263
rect 818 217 1112 220
rect 1158 217 1160 263
rect 770 170 1160 217
rect 1330 252 1332 298
rect 1378 252 1380 298
rect 1330 120 1380 252
rect 1550 298 1600 560
rect 1550 252 1552 298
rect 1598 252 1600 298
rect 1550 190 1600 252
rect 0 106 1720 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1364 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1362 98
rect 1416 54 1720 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1362 54
rect 1408 52 1720 54
rect 0 0 1720 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 1314 1132 1358 1176
rect 1358 1132 1366 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 104 704 156 756
rect 624 594 676 646
rect 1284 653 1336 656
rect 1284 607 1287 653
rect 1287 607 1333 653
rect 1333 607 1336 653
rect 1284 604 1336 607
rect 324 493 376 496
rect 324 447 327 493
rect 327 447 373 493
rect 373 447 376 493
rect 324 444 376 447
rect 494 314 546 366
rect 1564 574 1616 626
rect 804 493 856 496
rect 804 447 807 493
rect 807 447 853 493
rect 853 447 856 493
rect 804 444 856 447
rect 1044 453 1096 456
rect 1044 407 1047 453
rect 1047 407 1093 453
rect 1093 407 1096 453
rect 1044 404 1096 407
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1364 98 1416 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1364 54 1408 98
rect 1408 54 1416 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 80 756 180 770
rect 80 704 104 756
rect 156 704 180 756
rect 80 690 180 704
rect 600 650 700 660
rect 1260 656 1360 670
rect 1260 650 1284 656
rect 600 646 1284 650
rect 600 594 624 646
rect 676 604 1284 646
rect 1336 604 1360 656
rect 676 594 1360 604
rect 600 590 1360 594
rect 1540 626 1640 640
rect 600 580 700 590
rect 1540 574 1564 626
rect 1616 574 1640 626
rect 1540 560 1640 574
rect 300 500 400 510
rect 780 500 880 510
rect 300 496 880 500
rect 300 444 324 496
rect 376 444 804 496
rect 856 444 880 496
rect 1040 470 1100 480
rect 300 440 880 444
rect 300 430 400 440
rect 780 430 880 440
rect 1030 456 1110 470
rect 1030 404 1044 456
rect 1096 404 1110 456
rect 1030 390 1110 404
rect 480 370 560 380
rect 1030 370 1100 390
rect 470 366 1100 370
rect 470 314 494 366
rect 546 314 1100 366
rect 470 310 1100 314
rect 480 300 560 310
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1350 110 1430 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1340 106 1440 110
rect 1340 54 1364 106
rect 1416 54 1440 106
rect 1340 50 1440 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1350 40 1430 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 300 430 400 510 4 A
port 1 nsew signal input
rlabel metal2 s 1540 560 1640 640 4 S
port 2 nsew signal output
rlabel metal2 s 80 690 180 770 4 CO
port 3 nsew signal output
rlabel metal2 s 480 300 560 380 4 B
port 4 nsew signal input
rlabel metal2 s 300 440 880 500 1 A
port 1 nsew signal input
rlabel metal2 s 780 430 880 510 1 A
port 1 nsew signal input
rlabel metal1 s 300 440 400 500 1 A
port 1 nsew signal input
rlabel metal1 s 780 440 880 500 1 A
port 1 nsew signal input
rlabel metal2 s 470 310 1100 370 1 B
port 4 nsew signal input
rlabel metal2 s 1030 310 1100 470 1 B
port 4 nsew signal input
rlabel metal2 s 1040 310 1100 480 1 B
port 4 nsew signal input
rlabel metal2 s 1030 390 1110 470 1 B
port 4 nsew signal input
rlabel metal1 s 490 310 550 490 1 B
port 4 nsew signal input
rlabel metal1 s 470 310 570 370 1 B
port 4 nsew signal input
rlabel metal1 s 470 430 570 490 1 B
port 4 nsew signal input
rlabel metal1 s 1040 380 1100 480 1 B
port 4 nsew signal input
rlabel metal1 s 110 190 160 1040 1 CO
port 3 nsew signal output
rlabel metal1 s 80 700 180 760 1 CO
port 3 nsew signal output
rlabel metal1 s 1550 190 1600 1040 1 S
port 2 nsew signal output
rlabel metal1 s 1500 700 1600 1040 1 S
port 2 nsew signal output
rlabel metal1 s 1550 560 1620 640 1 S
port 2 nsew signal output
rlabel metal1 s 1540 570 1640 630 1 S
port 2 nsew signal output
rlabel metal2 s 90 1120 190 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 280 700 330 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 620 700 670 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 770 700 820 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1330 900 1380 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 1110 1720 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1350 40 1430 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1340 50 1440 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 280 0 330 360 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1330 0 1380 360 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 0 0 1720 120 1 VSS
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1720 1230
string GDS_END 40702
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 26130
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
