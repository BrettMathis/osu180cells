magic
tech gf180mcuC
timestamp 1669390400
<< properties >>
string GDS_END 7231850
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7230886
<< end >>
