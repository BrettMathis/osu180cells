magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 552 1220
<< mvpmos >>
rect 0 0 120 1100
rect 224 0 344 1100
<< mvpdiff >>
rect -88 1087 0 1100
rect -88 837 -75 1087
rect -29 837 0 1087
rect -88 780 0 837
rect -88 734 -75 780
rect -29 734 0 780
rect -88 677 0 734
rect -88 631 -75 677
rect -29 631 0 677
rect -88 574 0 631
rect -88 528 -75 574
rect -29 528 0 574
rect -88 471 0 528
rect -88 425 -75 471
rect -29 425 0 471
rect -88 368 0 425
rect -88 322 -75 368
rect -29 322 0 368
rect -88 265 0 322
rect -88 219 -75 265
rect -29 219 0 265
rect -88 162 0 219
rect -88 116 -75 162
rect -29 116 0 162
rect -88 59 0 116
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1087 224 1100
rect 120 837 149 1087
rect 195 837 224 1087
rect 120 780 224 837
rect 120 734 149 780
rect 195 734 224 780
rect 120 677 224 734
rect 120 631 149 677
rect 195 631 224 677
rect 120 574 224 631
rect 120 528 149 574
rect 195 528 224 574
rect 120 471 224 528
rect 120 425 149 471
rect 195 425 224 471
rect 120 368 224 425
rect 120 322 149 368
rect 195 322 224 368
rect 120 265 224 322
rect 120 219 149 265
rect 195 219 224 265
rect 120 162 224 219
rect 120 116 149 162
rect 195 116 224 162
rect 120 59 224 116
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 1087 432 1100
rect 344 837 373 1087
rect 419 837 432 1087
rect 344 780 432 837
rect 344 734 373 780
rect 419 734 432 780
rect 344 677 432 734
rect 344 631 373 677
rect 419 631 432 677
rect 344 574 432 631
rect 344 528 373 574
rect 419 528 432 574
rect 344 471 432 528
rect 344 425 373 471
rect 419 425 432 471
rect 344 368 432 425
rect 344 322 373 368
rect 419 322 432 368
rect 344 265 432 322
rect 344 219 373 265
rect 419 219 432 265
rect 344 162 432 219
rect 344 116 373 162
rect 419 116 432 162
rect 344 59 432 116
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 837 -29 1087
rect -75 734 -29 780
rect -75 631 -29 677
rect -75 528 -29 574
rect -75 425 -29 471
rect -75 322 -29 368
rect -75 219 -29 265
rect -75 116 -29 162
rect -75 13 -29 59
rect 149 837 195 1087
rect 149 734 195 780
rect 149 631 195 677
rect 149 528 195 574
rect 149 425 195 471
rect 149 322 195 368
rect 149 219 195 265
rect 149 116 195 162
rect 149 13 195 59
rect 373 837 419 1087
rect 373 734 419 780
rect 373 631 419 677
rect 373 528 419 574
rect 373 425 419 471
rect 373 322 419 368
rect 373 219 419 265
rect 373 116 419 162
rect 373 13 419 59
<< polysilicon >>
rect 0 1100 120 1144
rect 224 1100 344 1144
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 1087 -29 1100
rect -75 780 -29 837
rect -75 677 -29 734
rect -75 574 -29 631
rect -75 471 -29 528
rect -75 368 -29 425
rect -75 265 -29 322
rect -75 162 -29 219
rect -75 59 -29 116
rect -75 0 -29 13
rect 149 1087 195 1100
rect 149 780 195 837
rect 149 677 195 734
rect 149 574 195 631
rect 149 471 195 528
rect 149 368 195 425
rect 149 265 195 322
rect 149 162 195 219
rect 149 59 195 116
rect 149 0 195 13
rect 373 1087 419 1100
rect 373 780 419 837
rect 373 677 419 734
rect 373 574 419 631
rect 373 471 419 528
rect 373 368 419 425
rect 373 265 419 322
rect 373 162 419 219
rect 373 59 419 116
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 550 -52 550 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 550 396 550 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 550 172 550 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 76968
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 73514
<< end >>
