magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -42 16923 642 16942
rect -42 -23 -23 16923
rect 623 -23 642 16923
rect -42 -42 642 -23
<< psubdiffcont >>
rect -23 -23 623 16923
<< metal1 >>
rect -34 16923 634 16934
rect -34 -23 -23 16923
rect 623 -23 634 16923
rect -34 -34 634 -23
<< properties >>
string GDS_END 2188768
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2112412
<< end >>
