magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44892 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13291 44892 13323 44924 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13097 44878 13323 44892
tri 13323 44878 13337 44892 sw
rect 13097 44847 13337 44878
tri 13337 44847 13368 44878 sw
rect 13097 44846 13368 44847
tri 13368 44846 13369 44847 sw
rect 13097 44844 13369 44846
tri 13097 44831 13110 44844 ne
rect 13110 44833 13369 44844
tri 13369 44833 13382 44846 sw
rect 70802 44844 71000 44902
rect 13110 44831 13382 44833
tri 13110 44785 13155 44831 ne
rect 13155 44824 13382 44831
rect 13155 44785 13254 44824
tri 13155 44769 13172 44785 ne
rect 13172 44778 13254 44785
rect 13300 44801 13382 44824
tri 13382 44801 13414 44833 sw
rect 13300 44778 13414 44801
rect 13172 44769 13414 44778
tri 13172 44756 13185 44769 ne
rect 13185 44756 13414 44769
tri 13414 44756 13459 44801 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
tri 13185 44724 13217 44756 ne
rect 13217 44746 13459 44756
tri 13459 44746 13469 44756 sw
rect 13217 44724 13469 44746
tri 13217 44714 13227 44724 ne
rect 13227 44714 13469 44724
tri 13469 44714 13501 44746 sw
rect 70802 44740 71000 44798
tri 13227 44696 13245 44714 ne
rect 13245 44701 13501 44714
tri 13501 44701 13514 44714 sw
rect 13245 44696 13514 44701
tri 13514 44696 13519 44701 sw
tri 13245 44651 13290 44696 ne
rect 13290 44692 13519 44696
rect 13290 44651 13386 44692
tri 13290 44637 13304 44651 ne
rect 13304 44646 13386 44651
rect 13432 44651 13519 44692
tri 13519 44651 13565 44696 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13432 44646 13565 44651
rect 13304 44637 13565 44646
tri 13304 44624 13317 44637 ne
rect 13317 44624 13565 44637
tri 13565 44624 13591 44651 sw
rect 70802 44636 71000 44694
tri 13317 44592 13349 44624 ne
rect 13349 44614 13591 44624
tri 13591 44614 13601 44624 sw
rect 13349 44592 13601 44614
tri 13349 44573 13368 44592 ne
rect 13368 44582 13601 44592
tri 13601 44582 13633 44614 sw
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
rect 13368 44573 13633 44582
tri 13633 44573 13643 44582 sw
tri 13368 44527 13413 44573 ne
rect 13413 44569 13643 44573
tri 13643 44569 13646 44573 sw
rect 13413 44560 13646 44569
rect 13413 44527 13518 44560
tri 13413 44505 13436 44527 ne
rect 13436 44514 13518 44527
rect 13564 44537 13646 44560
tri 13646 44537 13678 44569 sw
rect 13564 44514 13678 44537
rect 13436 44505 13678 44514
tri 13436 44492 13449 44505 ne
rect 13449 44492 13678 44505
tri 13678 44492 13723 44537 sw
rect 70802 44532 71000 44590
tri 13449 44460 13481 44492 ne
rect 13481 44482 13723 44492
tri 13723 44482 13733 44492 sw
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 13481 44460 13733 44482
tri 13481 44450 13491 44460 ne
rect 13491 44450 13733 44460
tri 13733 44450 13765 44482 sw
tri 13491 44405 13536 44450 ne
rect 13536 44437 13765 44450
tri 13765 44437 13778 44450 sw
rect 13536 44428 13778 44437
rect 13536 44405 13650 44428
tri 13536 44376 13565 44405 ne
rect 13565 44382 13650 44405
rect 13696 44405 13778 44428
tri 13778 44405 13810 44437 sw
rect 70802 44428 71000 44486
rect 13696 44382 13810 44405
rect 13565 44376 13810 44382
tri 13565 44360 13581 44376 ne
rect 13581 44360 13810 44376
tri 13810 44360 13855 44405 sw
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13581 44328 13613 44360 ne
rect 13613 44350 13855 44360
tri 13855 44350 13865 44360 sw
rect 13613 44328 13865 44350
tri 13613 44298 13643 44328 ne
rect 13643 44318 13865 44328
tri 13865 44318 13897 44350 sw
rect 70802 44324 71000 44382
rect 13643 44298 13897 44318
tri 13897 44298 13917 44318 sw
tri 13643 44253 13688 44298 ne
rect 13688 44296 13917 44298
rect 13688 44253 13782 44296
tri 13688 44241 13700 44253 ne
rect 13700 44250 13782 44253
rect 13828 44286 13917 44296
tri 13917 44286 13929 44298 sw
rect 13828 44273 13929 44286
tri 13929 44273 13942 44286 sw
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13828 44250 13942 44273
rect 13700 44241 13942 44250
tri 13700 44228 13713 44241 ne
rect 13713 44228 13942 44241
tri 13942 44228 13987 44273 sw
tri 13713 44196 13745 44228 ne
rect 13745 44218 13987 44228
tri 13987 44218 13997 44228 sw
rect 70802 44220 71000 44278
rect 13745 44196 13997 44218
tri 13745 44186 13755 44196 ne
rect 13755 44186 13997 44196
tri 13997 44186 14029 44218 sw
tri 13755 44141 13800 44186 ne
rect 13800 44173 14029 44186
tri 14029 44173 14042 44186 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 13800 44164 14042 44173
rect 13800 44141 13914 44164
tri 13800 44109 13832 44141 ne
rect 13832 44118 13914 44141
rect 13960 44141 14042 44164
tri 14042 44141 14074 44173 sw
rect 13960 44118 14074 44141
rect 13832 44109 14074 44118
tri 13832 44096 13845 44109 ne
rect 13845 44096 14074 44109
tri 14074 44096 14119 44141 sw
rect 70802 44116 71000 44174
tri 13845 44064 13877 44096 ne
rect 13877 44086 14119 44096
tri 14119 44086 14129 44096 sw
rect 13877 44064 14129 44086
tri 13877 44024 13917 44064 ne
rect 13917 44054 14129 44064
tri 14129 44054 14161 44086 sw
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 13917 44041 14161 44054
tri 14161 44041 14174 44054 sw
rect 13917 44032 14174 44041
rect 13917 44024 14046 44032
tri 13917 44011 13929 44024 ne
rect 13929 44011 14046 44024
tri 13929 43966 13975 44011 ne
rect 13975 43986 14046 44011
rect 14092 44024 14174 44032
tri 14174 44024 14191 44041 sw
rect 14092 44011 14191 44024
tri 14191 44011 14204 44024 sw
rect 70802 44012 71000 44070
rect 14092 43986 14204 44011
rect 13975 43966 14204 43986
tri 14204 43966 14249 44011 sw
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13975 43964 13977 43966 ne
rect 13977 43964 14249 43966
tri 14249 43964 14251 43966 sw
tri 13977 43932 14009 43964 ne
rect 14009 43932 14251 43964
tri 14009 43922 14019 43932 ne
rect 14019 43922 14251 43932
tri 14251 43922 14293 43964 sw
tri 14019 43877 14064 43922 ne
rect 14064 43909 14293 43922
tri 14293 43909 14306 43922 sw
rect 14064 43900 14306 43909
rect 14064 43877 14178 43900
tri 14064 43845 14096 43877 ne
rect 14096 43854 14178 43877
rect 14224 43877 14306 43900
tri 14306 43877 14338 43909 sw
rect 70802 43908 71000 43966
rect 14224 43854 14338 43877
rect 14096 43845 14338 43854
tri 14096 43832 14109 43845 ne
rect 14109 43832 14338 43845
tri 14338 43832 14383 43877 sw
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
tri 14109 43800 14141 43832 ne
rect 14141 43822 14383 43832
tri 14383 43822 14393 43832 sw
rect 14141 43800 14393 43822
tri 14141 43755 14186 43800 ne
rect 14186 43790 14393 43800
tri 14393 43790 14425 43822 sw
rect 70802 43804 71000 43862
rect 14186 43777 14425 43790
tri 14425 43777 14438 43790 sw
rect 14186 43768 14438 43777
rect 14186 43755 14310 43768
tri 14186 43749 14191 43755 ne
rect 14191 43749 14310 43755
tri 14191 43713 14228 43749 ne
rect 14228 43722 14310 43749
rect 14356 43749 14438 43768
tri 14438 43749 14466 43777 sw
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43745 14466 43749
tri 14466 43745 14470 43749 sw
rect 14356 43722 14470 43745
rect 14228 43713 14470 43722
tri 14228 43700 14241 43713 ne
rect 14241 43700 14470 43713
tri 14470 43700 14515 43745 sw
rect 70802 43700 71000 43758
tri 14241 43668 14273 43700 ne
rect 14273 43690 14515 43700
tri 14515 43690 14525 43700 sw
rect 14273 43668 14525 43690
tri 14273 43658 14283 43668 ne
rect 14283 43658 14525 43668
tri 14525 43658 14557 43690 sw
tri 14283 43647 14294 43658 ne
rect 14294 43647 14557 43658
tri 14294 43601 14339 43647 ne
rect 14339 43645 14557 43647
tri 14557 43645 14570 43658 sw
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14339 43636 14570 43645
rect 14339 43601 14442 43636
tri 14339 43581 14360 43601 ne
rect 14360 43590 14442 43601
rect 14488 43601 14570 43636
tri 14570 43601 14614 43645 sw
rect 14488 43590 14614 43601
rect 14360 43581 14614 43590
tri 14360 43568 14373 43581 ne
rect 14373 43568 14614 43581
tri 14614 43568 14647 43601 sw
rect 70802 43596 71000 43654
tri 14373 43536 14405 43568 ne
rect 14405 43558 14647 43568
tri 14647 43558 14657 43568 sw
rect 14405 43536 14657 43558
tri 14405 43491 14450 43536 ne
rect 14450 43526 14657 43536
tri 14657 43526 14689 43558 sw
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14450 43513 14689 43526
tri 14689 43513 14702 43526 sw
rect 14450 43504 14702 43513
rect 14450 43491 14574 43504
tri 14450 43475 14466 43491 ne
rect 14466 43475 14574 43491
tri 14466 43449 14492 43475 ne
rect 14492 43458 14574 43475
rect 14620 43475 14702 43504
tri 14702 43475 14740 43513 sw
rect 70802 43492 71000 43550
rect 14620 43458 14740 43475
rect 14492 43449 14740 43458
tri 14492 43436 14505 43449 ne
rect 14505 43436 14740 43449
tri 14740 43436 14779 43475 sw
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14505 43404 14537 43436 ne
rect 14537 43426 14779 43436
tri 14779 43426 14789 43436 sw
rect 14537 43404 14789 43426
tri 14537 43394 14547 43404 ne
rect 14547 43394 14789 43404
tri 14789 43394 14821 43426 sw
tri 14547 43349 14592 43394 ne
rect 14592 43381 14821 43394
tri 14821 43381 14834 43394 sw
rect 70802 43388 71000 43446
rect 14592 43372 14834 43381
rect 14592 43349 14706 43372
tri 14592 43317 14624 43349 ne
rect 14624 43326 14706 43349
rect 14752 43349 14834 43372
tri 14834 43349 14866 43381 sw
rect 14752 43326 14866 43349
rect 14624 43317 14866 43326
tri 14624 43304 14637 43317 ne
rect 14637 43304 14866 43317
tri 14866 43304 14911 43349 sw
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
tri 14637 43272 14669 43304 ne
rect 14669 43294 14911 43304
tri 14911 43294 14921 43304 sw
rect 14669 43272 14921 43294
tri 14669 43237 14704 43272 ne
rect 14704 43262 14921 43272
tri 14921 43262 14953 43294 sw
rect 70802 43284 71000 43342
rect 14704 43249 14953 43262
tri 14953 43249 14966 43262 sw
rect 14704 43240 14966 43249
rect 14704 43237 14838 43240
tri 14704 43201 14740 43237 ne
rect 14740 43201 14838 43237
tri 14740 43185 14756 43201 ne
rect 14756 43194 14838 43201
rect 14884 43237 14966 43240
tri 14966 43237 14979 43249 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43201 14979 43237
tri 14979 43201 15015 43237 sw
rect 14884 43194 15015 43201
rect 14756 43191 15015 43194
tri 15015 43191 15024 43201 sw
rect 14756 43185 15024 43191
tri 14756 43172 14769 43185 ne
rect 14769 43172 15024 43185
tri 15024 43172 15043 43191 sw
rect 70802 43180 71000 43238
tri 14769 43140 14801 43172 ne
rect 14801 43162 15043 43172
tri 15043 43162 15053 43172 sw
rect 14801 43140 15053 43162
tri 14801 43130 14811 43140 ne
rect 14811 43130 15053 43140
tri 15053 43130 15085 43162 sw
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14811 43085 14856 43130 ne
rect 14856 43117 15085 43130
tri 15085 43117 15098 43130 sw
rect 14856 43108 15098 43117
rect 14856 43085 14970 43108
tri 14856 43053 14888 43085 ne
rect 14888 43062 14970 43085
rect 15016 43085 15098 43108
tri 15098 43085 15130 43117 sw
rect 15016 43062 15130 43085
rect 14888 43053 15130 43062
tri 14888 43040 14901 43053 ne
rect 14901 43040 15130 43053
tri 15130 43040 15175 43085 sw
rect 70802 43076 71000 43134
tri 14901 43008 14933 43040 ne
rect 14933 43030 15175 43040
tri 15175 43030 15185 43040 sw
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
rect 14933 43008 15185 43030
tri 14933 42963 14978 43008 ne
rect 14978 42998 15185 43008
tri 15185 42998 15217 43030 sw
rect 14978 42985 15217 42998
tri 15217 42985 15230 42998 sw
rect 14978 42976 15230 42985
rect 14978 42963 15102 42976
tri 14978 42926 15015 42963 ne
rect 15015 42930 15102 42963
rect 15148 42971 15230 42976
tri 15230 42971 15244 42985 sw
rect 70802 42972 71000 43030
rect 15148 42930 15244 42971
rect 15015 42926 15244 42930
tri 15244 42926 15289 42971 sw
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15015 42917 15024 42926 ne
rect 15024 42917 15289 42926
tri 15024 42908 15033 42917 ne
rect 15033 42908 15289 42917
tri 15289 42908 15307 42926 sw
tri 15033 42872 15069 42908 ne
rect 15069 42898 15307 42908
tri 15307 42898 15317 42908 sw
rect 15069 42872 15317 42898
tri 15069 42866 15075 42872 ne
rect 15075 42866 15317 42872
tri 15317 42866 15349 42898 sw
rect 70802 42868 71000 42926
tri 15075 42821 15120 42866 ne
rect 15120 42844 15349 42866
rect 15120 42821 15234 42844
tri 15120 42789 15152 42821 ne
rect 15152 42798 15234 42821
rect 15280 42827 15349 42844
tri 15349 42827 15389 42866 sw
rect 15280 42821 15389 42827
tri 15389 42821 15394 42827 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42798 15394 42821
rect 15152 42789 15394 42798
tri 15152 42776 15165 42789 ne
rect 15165 42776 15394 42789
tri 15394 42776 15439 42821 sw
tri 15165 42744 15197 42776 ne
rect 15197 42766 15439 42776
tri 15439 42766 15449 42776 sw
rect 15197 42744 15449 42766
tri 15197 42699 15242 42744 ne
rect 15242 42734 15449 42744
tri 15449 42734 15481 42766 sw
rect 70802 42764 71000 42822
rect 15242 42721 15481 42734
tri 15481 42721 15494 42734 sw
rect 15242 42712 15494 42721
rect 15242 42699 15366 42712
tri 15242 42657 15284 42699 ne
rect 15284 42666 15366 42699
rect 15412 42697 15494 42712
tri 15494 42697 15518 42721 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 15412 42666 15518 42697
rect 15284 42657 15518 42666
tri 15284 42652 15289 42657 ne
rect 15289 42652 15518 42657
tri 15518 42652 15563 42697 sw
rect 70802 42660 71000 42718
tri 15289 42644 15297 42652 ne
rect 15297 42644 15563 42652
tri 15563 42644 15571 42652 sw
tri 15297 42612 15329 42644 ne
rect 15329 42634 15571 42644
tri 15571 42634 15581 42644 sw
rect 15329 42612 15581 42634
tri 15329 42602 15339 42612 ne
rect 15339 42602 15581 42612
tri 15581 42602 15613 42634 sw
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15339 42557 15384 42602 ne
rect 15384 42589 15613 42602
tri 15613 42589 15626 42602 sw
rect 15384 42580 15626 42589
rect 15384 42557 15498 42580
tri 15384 42552 15389 42557 ne
rect 15389 42552 15498 42557
tri 15389 42512 15429 42552 ne
rect 15429 42534 15498 42552
rect 15544 42557 15626 42580
tri 15626 42557 15658 42589 sw
rect 15544 42534 15658 42557
rect 15429 42512 15658 42534
tri 15658 42512 15703 42557 sw
rect 70802 42556 71000 42614
tri 15429 42480 15461 42512 ne
rect 15461 42507 15703 42512
tri 15703 42507 15708 42512 sw
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15461 42480 15708 42507
tri 15461 42435 15506 42480 ne
rect 15506 42470 15708 42480
tri 15708 42470 15745 42507 sw
rect 15506 42457 15745 42470
tri 15745 42457 15758 42470 sw
rect 15506 42448 15758 42457
rect 15506 42435 15630 42448
tri 15506 42393 15548 42435 ne
rect 15548 42402 15630 42435
rect 15676 42425 15758 42448
tri 15758 42425 15790 42457 sw
rect 70802 42452 71000 42510
rect 15676 42402 15790 42425
rect 15548 42393 15790 42402
tri 15548 42377 15563 42393 ne
rect 15563 42380 15790 42393
tri 15790 42380 15835 42425 sw
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 15563 42377 15835 42380
tri 15835 42377 15838 42380 sw
tri 15563 42348 15593 42377 ne
rect 15593 42370 15838 42377
tri 15838 42370 15845 42377 sw
rect 15593 42348 15845 42370
tri 15593 42338 15603 42348 ne
rect 15603 42338 15845 42348
tri 15845 42338 15877 42370 sw
rect 70802 42348 71000 42406
tri 15603 42293 15648 42338 ne
rect 15648 42325 15877 42338
tri 15877 42325 15890 42338 sw
rect 15648 42316 15890 42325
rect 15648 42293 15762 42316
tri 15648 42261 15680 42293 ne
rect 15680 42270 15762 42293
rect 15808 42293 15890 42316
tri 15890 42293 15922 42325 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42270 15922 42293
rect 15680 42261 15922 42270
tri 15680 42248 15693 42261 ne
rect 15693 42248 15922 42261
tri 15922 42248 15967 42293 sw
tri 15693 42216 15725 42248 ne
rect 15725 42238 15967 42248
tri 15967 42238 15977 42248 sw
rect 70802 42244 71000 42302
rect 15725 42216 15977 42238
tri 15725 42187 15753 42216 ne
rect 15753 42206 15977 42216
tri 15977 42206 16009 42238 sw
rect 15753 42193 16009 42206
tri 16009 42193 16022 42206 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 15753 42187 16022 42193
tri 16022 42187 16028 42193 sw
tri 15753 42142 15799 42187 ne
rect 15799 42184 16028 42187
rect 15799 42142 15894 42184
tri 15799 42129 15812 42142 ne
rect 15812 42138 15894 42142
rect 15940 42142 16028 42184
tri 16028 42142 16073 42187 sw
rect 15940 42138 16073 42142
rect 15812 42129 16073 42138
tri 15812 42103 15838 42129 ne
rect 15838 42116 16073 42129
tri 16073 42116 16099 42142 sw
rect 70802 42140 71000 42198
rect 15838 42103 16099 42116
tri 16099 42103 16112 42116 sw
tri 15838 42084 15857 42103 ne
rect 15857 42084 16112 42103
tri 15857 42074 15867 42084 ne
rect 15867 42074 16112 42084
tri 16112 42074 16141 42103 sw
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15867 42029 15912 42074 ne
rect 15912 42061 16141 42074
tri 16141 42061 16154 42074 sw
rect 15912 42052 16154 42061
rect 15912 42029 16026 42052
tri 15912 41997 15944 42029 ne
rect 15944 42006 16026 42029
rect 16072 42029 16154 42052
tri 16154 42029 16186 42061 sw
rect 70802 42036 71000 42094
rect 16072 42006 16186 42029
rect 15944 41997 16186 42006
tri 15944 41984 15957 41997 ne
rect 15957 41984 16186 41997
tri 16186 41984 16231 42029 sw
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15957 41952 15989 41984 ne
rect 15989 41974 16231 41984
tri 16231 41974 16241 41984 sw
rect 15989 41952 16241 41974
tri 15989 41907 16034 41952 ne
rect 16034 41942 16241 41952
tri 16241 41942 16273 41974 sw
rect 16034 41929 16273 41942
tri 16273 41929 16286 41942 sw
rect 70802 41932 71000 41990
rect 16034 41920 16286 41929
rect 16034 41907 16158 41920
tri 16034 41865 16076 41907 ne
rect 16076 41874 16158 41907
rect 16204 41897 16286 41920
tri 16286 41897 16318 41929 sw
rect 16204 41874 16318 41897
rect 16076 41865 16318 41874
tri 16076 41829 16112 41865 ne
rect 16112 41852 16318 41865
tri 16318 41852 16363 41897 sw
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16112 41842 16363 41852
tri 16363 41842 16373 41852 sw
rect 16112 41829 16373 41842
tri 16373 41829 16387 41842 sw
tri 16112 41820 16121 41829 ne
rect 16121 41820 16387 41829
tri 16121 41810 16131 41820 ne
rect 16131 41810 16387 41820
tri 16387 41810 16405 41829 sw
rect 70802 41828 71000 41886
tri 16131 41777 16163 41810 ne
rect 16163 41797 16405 41810
tri 16405 41797 16418 41810 sw
rect 16163 41788 16418 41797
rect 16163 41777 16290 41788
tri 16163 41733 16208 41777 ne
rect 16208 41742 16290 41777
rect 16336 41777 16418 41788
tri 16418 41777 16438 41797 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16438 41777
rect 16208 41733 16438 41742
tri 16208 41720 16221 41733 ne
rect 16221 41732 16438 41733
tri 16438 41732 16483 41777 sw
rect 16221 41720 16483 41732
tri 16483 41720 16495 41732 sw
rect 70802 41724 71000 41782
tri 16221 41688 16253 41720 ne
rect 16253 41710 16495 41720
tri 16495 41710 16505 41720 sw
rect 16253 41688 16505 41710
tri 16253 41643 16298 41688 ne
rect 16298 41678 16505 41688
tri 16505 41678 16537 41710 sw
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16298 41665 16537 41678
tri 16537 41665 16550 41678 sw
rect 16298 41656 16550 41665
rect 16298 41643 16422 41656
tri 16298 41601 16340 41643 ne
rect 16340 41610 16422 41643
rect 16468 41633 16550 41656
tri 16550 41633 16582 41665 sw
rect 16468 41610 16582 41633
rect 16340 41601 16582 41610
tri 16340 41556 16385 41601 ne
rect 16385 41588 16582 41601
tri 16582 41588 16627 41633 sw
rect 70802 41620 71000 41678
rect 16385 41578 16627 41588
tri 16627 41578 16637 41588 sw
rect 16385 41556 16637 41578
tri 16385 41554 16387 41556 ne
rect 16387 41554 16637 41556
tri 16637 41554 16661 41578 sw
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16387 41546 16395 41554 ne
rect 16395 41546 16661 41554
tri 16661 41546 16669 41554 sw
tri 16395 41501 16440 41546 ne
rect 16440 41533 16669 41546
tri 16669 41533 16682 41546 sw
rect 16440 41524 16682 41533
rect 16440 41501 16554 41524
tri 16440 41458 16483 41501 ne
rect 16483 41478 16554 41501
rect 16600 41501 16682 41524
tri 16682 41501 16714 41533 sw
rect 70802 41516 71000 41574
rect 16600 41478 16714 41501
rect 16483 41458 16714 41478
tri 16483 41456 16485 41458 ne
rect 16485 41456 16714 41458
tri 16714 41456 16759 41501 sw
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
tri 16485 41413 16528 41456 ne
rect 16528 41446 16759 41456
tri 16759 41446 16769 41456 sw
rect 16528 41414 16769 41446
tri 16769 41414 16801 41446 sw
rect 16528 41413 16801 41414
tri 16801 41413 16803 41414 sw
tri 16528 41367 16573 41413 ne
rect 16573 41392 16803 41413
rect 16573 41367 16686 41392
tri 16573 41337 16604 41367 ne
rect 16604 41346 16686 41367
rect 16732 41367 16803 41392
tri 16803 41367 16848 41413 sw
rect 70802 41412 71000 41470
rect 16732 41346 16848 41367
rect 16604 41337 16848 41346
tri 16604 41292 16649 41337 ne
rect 16649 41324 16848 41337
tri 16848 41324 16891 41367 sw
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16649 41314 16891 41324
tri 16891 41314 16901 41324 sw
rect 16649 41292 16901 41314
tri 16649 41280 16661 41292 ne
rect 16661 41282 16901 41292
tri 16901 41282 16933 41314 sw
rect 70802 41308 71000 41366
rect 16661 41280 16933 41282
tri 16933 41280 16935 41282 sw
tri 16661 41235 16706 41280 ne
rect 16706 41269 16935 41280
tri 16935 41269 16946 41280 sw
rect 16706 41260 16946 41269
rect 16706 41235 16818 41260
tri 16706 41205 16736 41235 ne
rect 16736 41214 16818 41235
rect 16864 41237 16946 41260
tri 16946 41237 16978 41269 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 16864 41214 16978 41237
rect 16736 41205 16978 41214
tri 16736 41192 16749 41205 ne
rect 16749 41192 16978 41205
tri 16978 41192 17023 41237 sw
rect 70802 41204 71000 41262
tri 16749 41160 16781 41192 ne
rect 16781 41182 17023 41192
tri 17023 41182 17033 41192 sw
rect 16781 41160 17033 41182
tri 16781 41150 16791 41160 ne
rect 16791 41150 17033 41160
tri 17033 41150 17065 41182 sw
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16791 41105 16836 41150 ne
rect 16836 41137 17065 41150
tri 17065 41137 17078 41150 sw
rect 16836 41128 17078 41137
rect 16836 41105 16950 41128
tri 16836 41093 16848 41105 ne
rect 16848 41093 16950 41105
tri 16848 41060 16881 41093 ne
rect 16881 41082 16950 41093
rect 16996 41105 17078 41128
tri 17078 41105 17110 41137 sw
rect 16996 41082 17110 41105
rect 16881 41060 17110 41082
tri 17110 41060 17155 41105 sw
rect 70802 41100 71000 41158
tri 16881 41028 16913 41060 ne
rect 16913 41050 17155 41060
tri 17155 41050 17165 41060 sw
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 16913 41028 17165 41050
tri 16913 41005 16935 41028 ne
rect 16935 41018 17165 41028
tri 17165 41018 17197 41050 sw
rect 16935 41005 17197 41018
tri 17197 41005 17210 41018 sw
tri 16935 40960 16981 41005 ne
rect 16981 41003 17210 41005
tri 17210 41003 17213 41005 sw
rect 16981 40996 17213 41003
rect 16981 40960 17082 40996
tri 16981 40941 17000 40960 ne
rect 17000 40950 17082 40960
rect 17128 40973 17213 40996
tri 17213 40973 17242 41003 sw
rect 70802 40996 71000 41054
rect 17128 40950 17242 40973
rect 17000 40941 17242 40950
tri 17000 40928 17013 40941 ne
rect 17013 40928 17242 40941
tri 17242 40928 17287 40973 sw
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 17013 40896 17045 40928 ne
rect 17045 40918 17287 40928
tri 17287 40918 17297 40928 sw
rect 17045 40896 17297 40918
tri 17045 40886 17055 40896 ne
rect 17055 40886 17297 40896
tri 17297 40886 17329 40918 sw
rect 70802 40892 71000 40950
tri 17055 40841 17100 40886 ne
rect 17100 40873 17329 40886
tri 17329 40873 17342 40886 sw
rect 17100 40864 17342 40873
rect 17100 40841 17214 40864
tri 17100 40809 17132 40841 ne
rect 17132 40818 17214 40841
rect 17260 40841 17342 40864
tri 17342 40841 17374 40873 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17374 40841
rect 17132 40809 17374 40818
tri 17132 40796 17145 40809 ne
rect 17145 40796 17374 40809
tri 17374 40796 17419 40841 sw
tri 17145 40764 17177 40796 ne
rect 17177 40786 17419 40796
tri 17419 40786 17429 40796 sw
rect 70802 40788 71000 40846
rect 17177 40764 17429 40786
tri 17177 40731 17210 40764 ne
rect 17210 40754 17429 40764
tri 17429 40754 17461 40786 sw
rect 17210 40741 17461 40754
tri 17461 40741 17474 40754 sw
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17210 40732 17474 40741
rect 17210 40731 17346 40732
tri 17210 40728 17213 40731 ne
rect 17213 40728 17346 40731
tri 17213 40683 17258 40728 ne
rect 17258 40686 17346 40728
rect 17392 40731 17474 40732
tri 17474 40731 17484 40741 sw
rect 17392 40728 17484 40731
tri 17484 40728 17487 40731 sw
rect 17392 40686 17487 40728
rect 17258 40683 17487 40686
tri 17487 40683 17532 40728 sw
rect 70802 40684 71000 40742
tri 17258 40677 17264 40683 ne
rect 17264 40677 17532 40683
tri 17264 40664 17277 40677 ne
rect 17277 40664 17532 40677
tri 17532 40664 17551 40683 sw
tri 17277 40632 17309 40664 ne
rect 17309 40654 17551 40664
tri 17551 40654 17561 40664 sw
rect 17309 40632 17561 40654
tri 17309 40622 17319 40632 ne
rect 17319 40622 17561 40632
tri 17561 40622 17593 40654 sw
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17319 40577 17364 40622 ne
rect 17364 40609 17593 40622
tri 17593 40609 17606 40622 sw
rect 17364 40600 17606 40609
rect 17364 40577 17478 40600
tri 17364 40545 17396 40577 ne
rect 17396 40554 17478 40577
rect 17524 40577 17606 40600
tri 17606 40577 17638 40609 sw
rect 70802 40580 71000 40638
rect 17524 40554 17638 40577
rect 17396 40545 17638 40554
tri 17396 40532 17409 40545 ne
rect 17409 40532 17638 40545
tri 17638 40532 17683 40577 sw
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17409 40500 17441 40532 ne
rect 17441 40522 17683 40532
tri 17683 40522 17693 40532 sw
rect 17441 40500 17693 40522
tri 17441 40457 17484 40500 ne
rect 17484 40490 17693 40500
tri 17693 40490 17725 40522 sw
rect 17484 40477 17725 40490
tri 17725 40477 17738 40490 sw
rect 17484 40468 17738 40477
rect 17484 40457 17610 40468
tri 17484 40413 17528 40457 ne
rect 17528 40422 17610 40457
rect 17656 40457 17738 40468
tri 17738 40457 17759 40477 sw
rect 70802 40476 71000 40534
rect 17656 40445 17759 40457
tri 17759 40445 17770 40457 sw
rect 17656 40422 17770 40445
rect 17528 40413 17770 40422
tri 17528 40400 17541 40413 ne
rect 17541 40400 17770 40413
tri 17770 40400 17815 40445 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
tri 17541 40368 17573 40400 ne
rect 17573 40390 17815 40400
tri 17815 40390 17825 40400 sw
rect 17573 40368 17825 40390
tri 17573 40363 17577 40368 ne
rect 17577 40363 17825 40368
tri 17577 40358 17583 40363 ne
rect 17583 40358 17825 40363
tri 17825 40358 17857 40390 sw
rect 70802 40372 71000 40430
tri 17583 40318 17623 40358 ne
rect 17623 40345 17857 40358
tri 17857 40345 17870 40358 sw
rect 17623 40336 17870 40345
rect 17623 40318 17742 40336
tri 17623 40281 17660 40318 ne
rect 17660 40290 17742 40318
rect 17788 40318 17870 40336
tri 17870 40318 17897 40345 sw
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40290 17897 40318
rect 17660 40281 17897 40290
tri 17660 40268 17673 40281 ne
rect 17673 40273 17897 40281
tri 17897 40273 17942 40318 sw
rect 17673 40268 17942 40273
tri 17942 40268 17947 40273 sw
rect 70802 40268 71000 40326
tri 17673 40236 17705 40268 ne
rect 17705 40258 17947 40268
tri 17947 40258 17957 40268 sw
rect 17705 40236 17957 40258
tri 17705 40191 17750 40236 ne
rect 17750 40226 17957 40236
tri 17957 40226 17989 40258 sw
rect 17750 40213 17989 40226
tri 17989 40213 18002 40226 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17750 40204 18002 40213
rect 17750 40191 17874 40204
tri 17750 40182 17759 40191 ne
rect 17759 40182 17874 40191
tri 17759 40149 17792 40182 ne
rect 17792 40158 17874 40182
rect 17920 40182 18002 40204
tri 18002 40182 18033 40213 sw
rect 17920 40181 18033 40182
tri 18033 40181 18034 40182 sw
rect 17920 40158 18034 40181
rect 17792 40149 18034 40158
tri 17792 40136 17805 40149 ne
rect 17805 40136 18034 40149
tri 18034 40136 18079 40181 sw
rect 70802 40164 71000 40222
tri 17805 40104 17837 40136 ne
rect 17837 40126 18079 40136
tri 18079 40126 18089 40136 sw
rect 17837 40104 18089 40126
tri 17837 40094 17847 40104 ne
rect 17847 40094 18089 40104
tri 18089 40094 18121 40126 sw
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17847 40049 17892 40094 ne
rect 17892 40081 18121 40094
tri 18121 40081 18134 40094 sw
rect 17892 40072 18134 40081
rect 17892 40049 18006 40072
tri 17892 40004 17937 40049 ne
rect 17937 40026 18006 40049
rect 18052 40049 18134 40072
tri 18134 40049 18166 40081 sw
rect 70802 40060 71000 40118
rect 18052 40026 18166 40049
rect 17937 40004 18166 40026
tri 18166 40004 18211 40049 sw
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
tri 17937 39999 17942 40004 ne
rect 17942 39999 18211 40004
tri 17942 39953 17987 39999 ne
rect 17987 39994 18211 39999
tri 18211 39994 18221 40004 sw
rect 17987 39962 18221 39994
tri 18221 39962 18253 39994 sw
rect 17987 39953 18253 39962
tri 18253 39953 18262 39962 sw
rect 70802 39956 71000 40014
tri 17987 39908 18033 39953 ne
rect 18033 39940 18262 39953
rect 18033 39908 18138 39940
tri 18033 39885 18056 39908 ne
rect 18056 39894 18138 39908
rect 18184 39908 18262 39940
tri 18262 39908 18307 39953 sw
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39894 18307 39908
rect 18056 39885 18307 39894
tri 18056 39872 18069 39885 ne
rect 18069 39872 18307 39885
tri 18307 39872 18343 39908 sw
tri 18069 39840 18101 39872 ne
rect 18101 39862 18343 39872
tri 18343 39862 18353 39872 sw
rect 18101 39840 18353 39862
tri 18101 39830 18111 39840 ne
rect 18111 39830 18353 39840
tri 18353 39830 18385 39862 sw
rect 70802 39852 71000 39910
tri 18111 39785 18156 39830 ne
rect 18156 39817 18385 39830
tri 18385 39817 18398 39830 sw
rect 18156 39808 18398 39817
rect 18156 39785 18270 39808
tri 18156 39753 18188 39785 ne
rect 18188 39762 18270 39785
rect 18316 39785 18398 39808
tri 18398 39785 18430 39817 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39762 18430 39785
rect 18188 39753 18430 39762
tri 18188 39740 18201 39753 ne
rect 18201 39740 18430 39753
tri 18430 39740 18475 39785 sw
rect 70802 39748 71000 39806
tri 18201 39708 18233 39740 ne
rect 18233 39730 18475 39740
tri 18475 39730 18485 39740 sw
rect 18233 39708 18485 39730
tri 18233 39663 18278 39708 ne
rect 18278 39698 18485 39708
tri 18485 39698 18517 39730 sw
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18278 39685 18517 39698
tri 18517 39685 18530 39698 sw
rect 18278 39679 18530 39685
tri 18530 39679 18537 39685 sw
rect 18278 39676 18537 39679
rect 18278 39663 18402 39676
tri 18278 39634 18307 39663 ne
rect 18307 39633 18402 39663
tri 18307 39608 18333 39633 ne
rect 18333 39630 18402 39633
rect 18448 39633 18537 39676
tri 18537 39633 18582 39679 sw
rect 70802 39644 71000 39702
rect 18448 39630 18582 39633
rect 18333 39608 18582 39630
tri 18582 39608 18607 39633 sw
tri 18333 39576 18365 39608 ne
rect 18365 39598 18607 39608
tri 18607 39598 18617 39608 sw
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
rect 18365 39576 18617 39598
tri 18365 39566 18375 39576 ne
rect 18375 39566 18617 39576
tri 18617 39566 18649 39598 sw
tri 18375 39521 18420 39566 ne
rect 18420 39544 18649 39566
rect 18420 39521 18534 39544
tri 18420 39489 18452 39521 ne
rect 18452 39498 18534 39521
rect 18580 39543 18649 39544
tri 18649 39543 18672 39566 sw
rect 18580 39521 18672 39543
tri 18672 39521 18694 39543 sw
rect 70802 39540 71000 39598
rect 18580 39498 18694 39521
rect 18452 39489 18694 39498
tri 18452 39476 18465 39489 ne
rect 18465 39476 18694 39489
tri 18694 39476 18739 39521 sw
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18465 39444 18497 39476 ne
rect 18497 39466 18739 39476
tri 18739 39466 18749 39476 sw
rect 18497 39444 18749 39466
tri 18497 39399 18542 39444 ne
rect 18542 39434 18749 39444
tri 18749 39434 18781 39466 sw
rect 70802 39436 71000 39494
rect 18542 39421 18781 39434
tri 18781 39421 18794 39434 sw
rect 18542 39412 18794 39421
rect 18542 39399 18666 39412
tri 18542 39359 18582 39399 ne
rect 18582 39366 18666 39399
rect 18712 39404 18794 39412
tri 18794 39404 18811 39421 sw
rect 18712 39366 18811 39404
rect 18582 39359 18811 39366
tri 18811 39359 18856 39404 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
tri 18582 39357 18584 39359 ne
rect 18584 39357 18856 39359
tri 18584 39344 18597 39357 ne
rect 18597 39344 18856 39357
tri 18856 39344 18871 39359 sw
tri 18597 39312 18629 39344 ne
rect 18629 39334 18871 39344
tri 18871 39334 18881 39344 sw
rect 18629 39312 18881 39334
tri 18629 39302 18639 39312 ne
rect 18639 39302 18881 39312
tri 18881 39302 18913 39334 sw
rect 70802 39332 71000 39390
tri 18639 39269 18672 39302 ne
rect 18672 39289 18913 39302
tri 18913 39289 18926 39302 sw
rect 18672 39280 18926 39289
rect 18672 39269 18798 39280
tri 18672 39224 18717 39269 ne
rect 18717 39234 18798 39269
rect 18844 39269 18926 39280
tri 18926 39269 18946 39289 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 18844 39234 18946 39269
rect 18717 39224 18946 39234
tri 18946 39224 18991 39269 sw
rect 70802 39228 71000 39286
tri 18717 39212 18729 39224 ne
rect 18729 39212 18991 39224
tri 18991 39212 19003 39224 sw
tri 18729 39180 18761 39212 ne
rect 18761 39202 19003 39212
tri 19003 39202 19013 39212 sw
rect 18761 39180 19013 39202
tri 18761 39135 18806 39180 ne
rect 18806 39170 19013 39180
tri 19013 39170 19045 39202 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18806 39157 19045 39170
tri 19045 39157 19058 39170 sw
rect 18806 39148 19058 39157
rect 18806 39135 18930 39148
tri 18806 39093 18848 39135 ne
rect 18848 39102 18930 39135
rect 18976 39130 19058 39148
tri 19058 39130 19085 39157 sw
rect 18976 39102 19085 39130
rect 18848 39093 19085 39102
tri 18848 39085 18856 39093 ne
rect 18856 39085 19085 39093
tri 19085 39085 19131 39130 sw
rect 70802 39124 71000 39182
tri 18856 39080 18861 39085 ne
rect 18861 39080 19131 39085
tri 19131 39080 19135 39085 sw
tri 18861 39048 18893 39080 ne
rect 18893 39070 19135 39080
tri 19135 39070 19145 39080 sw
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
rect 18893 39048 19145 39070
tri 18893 39038 18903 39048 ne
rect 18903 39038 19145 39048
tri 19145 39038 19177 39070 sw
tri 18903 38993 18948 39038 ne
rect 18948 39025 19177 39038
tri 19177 39025 19190 39038 sw
rect 18948 39016 19190 39025
rect 18948 38993 19062 39016
tri 18948 38961 18980 38993 ne
rect 18980 38970 19062 38993
rect 19108 38993 19190 39016
tri 19190 38993 19222 39025 sw
rect 70802 39020 71000 39078
rect 19108 38970 19222 38993
rect 18980 38961 19222 38970
tri 18980 38948 18993 38961 ne
rect 18993 38948 19222 38961
tri 19222 38948 19267 38993 sw
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
tri 18993 38916 19025 38948 ne
rect 19025 38938 19267 38948
tri 19267 38938 19277 38948 sw
rect 19025 38916 19277 38938
tri 19025 38904 19037 38916 ne
rect 19037 38906 19277 38916
tri 19277 38906 19309 38938 sw
rect 70802 38916 71000 38974
rect 19037 38904 19309 38906
tri 19037 38859 19082 38904 ne
rect 19082 38893 19309 38904
tri 19309 38893 19322 38906 sw
rect 19082 38884 19322 38893
rect 19082 38859 19194 38884
tri 19082 38829 19112 38859 ne
rect 19112 38838 19194 38859
rect 19240 38859 19322 38884
tri 19322 38859 19356 38893 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19356 38859
rect 19112 38829 19356 38838
tri 19112 38810 19131 38829 ne
rect 19131 38816 19356 38829
tri 19356 38816 19399 38859 sw
rect 19131 38814 19399 38816
tri 19399 38814 19401 38816 sw
rect 19131 38810 19401 38814
tri 19401 38810 19405 38814 sw
rect 70802 38812 71000 38870
tri 19131 38784 19157 38810 ne
rect 19157 38806 19405 38810
tri 19405 38806 19409 38810 sw
rect 19157 38784 19409 38806
tri 19157 38774 19167 38784 ne
rect 19167 38774 19409 38784
tri 19409 38774 19441 38806 sw
tri 19167 38729 19212 38774 ne
rect 19212 38761 19441 38774
tri 19441 38761 19454 38774 sw
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
rect 19212 38752 19454 38761
rect 19212 38729 19326 38752
tri 19212 38697 19244 38729 ne
rect 19244 38706 19326 38729
rect 19372 38729 19454 38752
tri 19454 38729 19486 38761 sw
rect 19372 38706 19486 38729
rect 19244 38697 19486 38706
tri 19244 38684 19257 38697 ne
rect 19257 38684 19486 38697
tri 19486 38684 19531 38729 sw
rect 70802 38708 71000 38766
tri 19257 38652 19289 38684 ne
rect 19289 38674 19531 38684
tri 19531 38674 19541 38684 sw
rect 19289 38652 19541 38674
tri 19289 38607 19334 38652 ne
rect 19334 38642 19541 38652
tri 19541 38642 19573 38674 sw
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
rect 19334 38629 19573 38642
tri 19573 38629 19586 38642 sw
rect 19334 38620 19586 38629
rect 19334 38607 19458 38620
tri 19334 38585 19356 38607 ne
rect 19356 38585 19458 38607
tri 19356 38539 19401 38585 ne
rect 19401 38574 19458 38585
rect 19504 38597 19586 38620
tri 19586 38597 19618 38629 sw
rect 70802 38604 71000 38662
rect 19504 38574 19618 38597
rect 19401 38552 19618 38574
tri 19618 38552 19663 38597 sw
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 19401 38542 19663 38552
tri 19663 38542 19673 38552 sw
rect 19401 38539 19673 38542
tri 19401 38536 19405 38539 ne
rect 19405 38536 19673 38539
tri 19673 38536 19679 38542 sw
tri 19405 38510 19431 38536 ne
rect 19431 38510 19679 38536
tri 19679 38510 19705 38536 sw
tri 19431 38494 19447 38510 ne
rect 19447 38497 19705 38510
tri 19705 38497 19718 38510 sw
rect 70802 38500 71000 38558
rect 19447 38494 19718 38497
tri 19718 38494 19721 38497 sw
tri 19447 38449 19492 38494 ne
rect 19492 38488 19721 38494
rect 19492 38449 19590 38488
tri 19492 38433 19508 38449 ne
rect 19508 38442 19590 38449
rect 19636 38449 19721 38488
tri 19721 38449 19766 38494 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19766 38449
rect 19508 38433 19766 38442
tri 19508 38420 19521 38433 ne
rect 19521 38420 19766 38433
tri 19766 38420 19795 38449 sw
tri 19521 38388 19553 38420 ne
rect 19553 38410 19795 38420
tri 19795 38410 19805 38420 sw
rect 19553 38388 19805 38410
tri 19553 38343 19598 38388 ne
rect 19598 38378 19805 38388
tri 19805 38378 19837 38410 sw
rect 70802 38396 71000 38454
rect 19598 38365 19837 38378
tri 19837 38365 19850 38378 sw
rect 19598 38356 19850 38365
rect 19598 38343 19722 38356
tri 19598 38301 19640 38343 ne
rect 19640 38310 19722 38343
rect 19768 38333 19850 38356
tri 19850 38333 19882 38365 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38310 19882 38333
rect 19640 38301 19882 38310
tri 19640 38261 19679 38301 ne
rect 19679 38288 19882 38301
tri 19882 38288 19927 38333 sw
rect 70802 38292 71000 38350
rect 19679 38278 19927 38288
tri 19927 38278 19937 38288 sw
rect 19679 38261 19937 38278
tri 19937 38261 19954 38278 sw
tri 19679 38256 19685 38261 ne
rect 19685 38256 19954 38261
tri 19685 38246 19695 38256 ne
rect 19695 38246 19954 38256
tri 19954 38246 19969 38261 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
tri 19695 38201 19740 38246 ne
rect 19740 38233 19969 38246
tri 19969 38233 19982 38246 sw
rect 19740 38224 19982 38233
rect 19740 38201 19854 38224
tri 19740 38175 19766 38201 ne
rect 19766 38178 19854 38201
rect 19900 38201 19982 38224
tri 19982 38201 20014 38233 sw
rect 19900 38178 20014 38201
rect 19766 38175 20014 38178
tri 19766 38156 19785 38175 ne
rect 19785 38156 20014 38175
tri 20014 38156 20059 38201 sw
rect 70802 38188 71000 38246
tri 19785 38124 19817 38156 ne
rect 19817 38146 20059 38156
tri 20059 38146 20069 38156 sw
rect 19817 38124 20069 38146
tri 19817 38079 19862 38124 ne
rect 19862 38114 20069 38124
tri 20069 38114 20101 38146 sw
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19862 38092 20101 38114
rect 19862 38079 19986 38092
tri 19862 38037 19904 38079 ne
rect 19904 38046 19986 38079
rect 20032 38084 20101 38092
tri 20101 38084 20131 38114 sw
rect 70802 38084 71000 38142
rect 20032 38069 20131 38084
tri 20131 38069 20146 38084 sw
rect 20032 38046 20146 38069
rect 19904 38037 20146 38046
tri 19904 37992 19949 38037 ne
rect 19949 38024 20146 38037
tri 20146 38024 20191 38069 sw
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 19949 38014 20191 38024
tri 20191 38014 20201 38024 sw
rect 19949 37992 20201 38014
tri 19949 37987 19954 37992 ne
rect 19954 37987 20201 37992
tri 20201 37987 20228 38014 sw
tri 19954 37982 19959 37987 ne
rect 19959 37982 20228 37987
tri 20228 37982 20233 37987 sw
tri 19959 37937 20004 37982 ne
rect 20004 37969 20233 37982
tri 20233 37969 20246 37982 sw
rect 70802 37980 71000 38038
rect 20004 37960 20246 37969
rect 20004 37937 20118 37960
tri 20004 37905 20036 37937 ne
rect 20036 37914 20118 37937
rect 20164 37937 20246 37960
tri 20246 37937 20278 37969 sw
rect 20164 37914 20278 37937
rect 20036 37905 20278 37914
tri 20036 37892 20049 37905 ne
rect 20049 37892 20278 37905
tri 20278 37892 20323 37937 sw
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
tri 20049 37860 20081 37892 ne
rect 20081 37882 20323 37892
tri 20323 37882 20333 37892 sw
rect 20081 37860 20333 37882
tri 20081 37850 20091 37860 ne
rect 20091 37850 20333 37860
tri 20333 37850 20365 37882 sw
rect 70802 37876 71000 37934
tri 20091 37810 20131 37850 ne
rect 20131 37837 20365 37850
tri 20365 37837 20378 37850 sw
rect 20131 37828 20378 37837
rect 20131 37810 20250 37828
tri 20131 37765 20176 37810 ne
rect 20176 37782 20250 37810
rect 20296 37810 20378 37828
tri 20378 37810 20405 37837 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20296 37782 20405 37810
rect 20176 37765 20405 37782
tri 20405 37765 20451 37810 sw
rect 70802 37772 71000 37830
tri 20176 37760 20181 37765 ne
rect 20181 37760 20451 37765
tri 20451 37760 20455 37765 sw
tri 20181 37728 20213 37760 ne
rect 20213 37750 20455 37760
tri 20455 37750 20465 37760 sw
rect 20213 37728 20465 37750
tri 20213 37713 20228 37728 ne
rect 20228 37718 20465 37728
tri 20465 37718 20497 37750 sw
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 20228 37713 20497 37718
tri 20497 37713 20503 37718 sw
tri 20228 37667 20273 37713 ne
rect 20273 37705 20503 37713
tri 20503 37705 20510 37713 sw
rect 20273 37696 20510 37705
rect 20273 37667 20382 37696
tri 20273 37641 20300 37667 ne
rect 20300 37650 20382 37667
rect 20428 37673 20510 37696
tri 20510 37673 20542 37705 sw
rect 20428 37650 20542 37673
rect 20300 37641 20542 37650
tri 20300 37628 20313 37641 ne
rect 20313 37628 20542 37641
tri 20542 37628 20587 37673 sw
rect 70802 37668 71000 37726
tri 20313 37596 20345 37628 ne
rect 20345 37618 20587 37628
tri 20587 37618 20597 37628 sw
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
rect 20345 37596 20597 37618
tri 20345 37586 20355 37596 ne
rect 20355 37586 20597 37596
tri 20597 37586 20629 37618 sw
tri 20355 37541 20400 37586 ne
rect 20400 37573 20629 37586
tri 20629 37573 20642 37586 sw
rect 20400 37564 20642 37573
rect 20400 37541 20514 37564
tri 20400 37509 20432 37541 ne
rect 20432 37518 20514 37541
rect 20560 37541 20642 37564
tri 20642 37541 20674 37573 sw
rect 70802 37564 71000 37622
rect 20560 37518 20674 37541
rect 20432 37509 20674 37518
tri 20432 37496 20445 37509 ne
rect 20445 37496 20674 37509
tri 20674 37496 20719 37541 sw
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
tri 20445 37464 20477 37496 ne
rect 20477 37486 20719 37496
tri 20719 37486 20729 37496 sw
rect 20477 37464 20729 37486
tri 20477 37445 20496 37464 ne
rect 20496 37454 20729 37464
tri 20729 37454 20761 37486 sw
rect 70802 37460 71000 37518
rect 20496 37445 20761 37454
tri 20496 37438 20503 37445 ne
rect 20503 37441 20761 37445
tri 20761 37441 20774 37454 sw
rect 20503 37438 20774 37441
tri 20774 37438 20777 37441 sw
tri 20503 37400 20541 37438 ne
rect 20541 37432 20777 37438
rect 20541 37400 20646 37432
tri 20541 37377 20564 37400 ne
rect 20564 37386 20646 37400
rect 20692 37400 20777 37432
tri 20777 37400 20815 37438 sw
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37386 20815 37400
rect 20564 37377 20815 37386
tri 20564 37364 20577 37377 ne
rect 20577 37364 20815 37377
tri 20815 37364 20851 37400 sw
tri 20577 37332 20609 37364 ne
rect 20609 37355 20851 37364
tri 20851 37355 20861 37364 sw
rect 20609 37332 20861 37355
rect 70802 37356 71000 37414
tri 20609 37322 20619 37332 ne
rect 20619 37322 20861 37332
tri 20861 37322 20893 37354 sw
tri 20619 37277 20664 37322 ne
rect 20664 37309 20893 37322
tri 20893 37309 20906 37322 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 20664 37300 20906 37309
rect 20664 37277 20778 37300
tri 20664 37245 20696 37277 ne
rect 20696 37254 20778 37277
rect 20824 37277 20906 37300
tri 20906 37277 20938 37309 sw
rect 20824 37254 20938 37277
rect 20696 37245 20938 37254
tri 20696 37232 20709 37245 ne
rect 20709 37232 20938 37245
tri 20938 37232 20983 37277 sw
rect 70802 37252 71000 37310
tri 20709 37200 20741 37232 ne
rect 20741 37222 20983 37232
tri 20983 37222 20993 37232 sw
rect 20741 37200 20993 37222
tri 20741 37164 20777 37200 ne
rect 20777 37190 20993 37200
tri 20993 37190 21025 37222 sw
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20777 37177 21025 37190
tri 21025 37177 21038 37190 sw
rect 20777 37168 21038 37177
rect 20777 37164 20910 37168
tri 20777 37119 20822 37164 ne
rect 20822 37122 20910 37164
rect 20956 37164 21038 37168
tri 21038 37164 21051 37177 sw
rect 20956 37145 21051 37164
tri 21051 37145 21070 37164 sw
rect 70802 37148 71000 37206
rect 20956 37122 21070 37145
rect 20822 37119 21070 37122
tri 20822 37113 20828 37119 ne
rect 20828 37113 21070 37119
tri 20828 37100 20841 37113 ne
rect 20841 37100 21070 37113
tri 21070 37100 21115 37145 sw
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20841 37068 20873 37100 ne
rect 20873 37090 21115 37100
tri 21115 37090 21125 37100 sw
rect 20873 37068 21125 37090
tri 20873 37058 20883 37068 ne
rect 20883 37058 21125 37068
tri 21125 37058 21157 37090 sw
tri 20883 37035 20906 37058 ne
rect 20906 37045 21157 37058
tri 21157 37045 21170 37058 sw
rect 20906 37036 21170 37045
rect 20906 37035 21042 37036
tri 20906 36990 20951 37035 ne
rect 20951 36990 21042 37035
rect 21088 37035 21170 37036
tri 21170 37035 21180 37045 sw
rect 70802 37044 71000 37102
rect 21088 36990 21180 37035
tri 21180 36990 21225 37035 sw
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
tri 20951 36981 20960 36990 ne
rect 20960 36981 21225 36990
tri 20960 36968 20973 36981 ne
rect 20973 36968 21225 36981
tri 21225 36968 21247 36990 sw
tri 20973 36936 21005 36968 ne
rect 21005 36958 21247 36968
tri 21247 36958 21257 36968 sw
rect 21005 36936 21257 36958
tri 21005 36891 21050 36936 ne
rect 21050 36926 21257 36936
tri 21257 36926 21289 36958 sw
rect 70802 36940 71000 36998
rect 21050 36913 21289 36926
tri 21289 36913 21302 36926 sw
rect 21050 36904 21302 36913
rect 21050 36891 21174 36904
tri 21050 36889 21051 36891 ne
rect 21051 36889 21174 36891
tri 21051 36849 21092 36889 ne
rect 21092 36858 21174 36889
rect 21220 36889 21302 36904
tri 21302 36889 21326 36913 sw
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36881 21326 36889
tri 21326 36881 21334 36889 sw
rect 21220 36858 21334 36881
rect 21092 36849 21334 36858
tri 21092 36836 21105 36849 ne
rect 21105 36836 21334 36849
tri 21334 36836 21379 36881 sw
rect 70802 36836 71000 36894
tri 21105 36804 21137 36836 ne
rect 21137 36826 21379 36836
tri 21379 36826 21389 36836 sw
rect 21137 36804 21389 36826
tri 21137 36794 21147 36804 ne
rect 21147 36794 21389 36804
tri 21389 36794 21421 36826 sw
tri 21147 36749 21192 36794 ne
rect 21192 36781 21421 36794
tri 21421 36781 21434 36794 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21192 36772 21434 36781
rect 21192 36749 21306 36772
tri 21192 36715 21225 36749 ne
rect 21225 36726 21306 36749
rect 21352 36749 21434 36772
tri 21434 36749 21466 36781 sw
rect 21352 36726 21466 36749
rect 21225 36715 21466 36726
tri 21225 36704 21237 36715 ne
rect 21237 36704 21466 36715
tri 21466 36704 21511 36749 sw
rect 70802 36732 71000 36790
tri 21237 36670 21271 36704 ne
rect 21271 36694 21511 36704
tri 21511 36694 21521 36704 sw
rect 21271 36670 21521 36694
tri 21271 36625 21316 36670 ne
rect 21316 36662 21521 36670
tri 21521 36662 21553 36694 sw
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21316 36640 21553 36662
rect 21316 36625 21438 36640
tri 21316 36615 21326 36625 ne
rect 21326 36615 21438 36625
tri 21326 36585 21356 36615 ne
rect 21356 36594 21438 36615
rect 21484 36625 21553 36640
tri 21553 36625 21590 36662 sw
rect 70802 36628 71000 36686
rect 21484 36615 21590 36625
tri 21590 36615 21600 36625 sw
rect 21484 36594 21600 36615
rect 21356 36585 21600 36594
tri 21356 36572 21369 36585 ne
rect 21369 36572 21600 36585
tri 21600 36572 21643 36615 sw
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21369 36540 21401 36572 ne
rect 21401 36562 21643 36572
tri 21643 36562 21653 36572 sw
rect 21401 36540 21653 36562
tri 21401 36530 21411 36540 ne
rect 21411 36530 21653 36540
tri 21653 36530 21685 36562 sw
tri 21411 36485 21456 36530 ne
rect 21456 36517 21685 36530
tri 21685 36517 21698 36530 sw
rect 70802 36524 71000 36582
rect 21456 36508 21698 36517
rect 21456 36485 21570 36508
tri 21456 36453 21488 36485 ne
rect 21488 36462 21570 36485
rect 21616 36485 21698 36508
tri 21698 36485 21730 36517 sw
rect 21616 36462 21730 36485
rect 21488 36453 21730 36462
tri 21488 36440 21501 36453 ne
rect 21501 36440 21730 36453
tri 21730 36440 21775 36485 sw
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
tri 21501 36408 21533 36440 ne
rect 21533 36430 21775 36440
tri 21775 36430 21785 36440 sw
rect 21533 36408 21785 36430
tri 21533 36363 21578 36408 ne
rect 21578 36398 21785 36408
tri 21785 36398 21817 36430 sw
rect 70802 36420 71000 36478
rect 21578 36385 21817 36398
tri 21817 36385 21830 36398 sw
rect 21578 36376 21830 36385
rect 21578 36363 21702 36376
tri 21578 36351 21590 36363 ne
rect 21590 36351 21702 36363
tri 21590 36341 21600 36351 ne
rect 21600 36341 21702 36351
tri 21600 36308 21633 36341 ne
rect 21633 36330 21702 36341
rect 21748 36341 21830 36376
tri 21830 36341 21875 36385 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21875 36341
rect 21633 36308 21875 36330
tri 21875 36308 21907 36341 sw
rect 70802 36316 71000 36374
tri 21633 36276 21665 36308 ne
rect 21665 36305 21907 36308
tri 21907 36305 21910 36308 sw
rect 21665 36276 21910 36305
tri 21665 36266 21675 36276 ne
rect 21675 36266 21910 36276
tri 21910 36266 21949 36305 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21675 36221 21720 36266 ne
rect 21720 36253 21949 36266
tri 21949 36253 21962 36266 sw
rect 21720 36244 21962 36253
rect 21720 36221 21834 36244
tri 21720 36189 21752 36221 ne
rect 21752 36198 21834 36221
rect 21880 36221 21962 36244
tri 21962 36221 21994 36253 sw
rect 21880 36198 21994 36221
rect 21752 36189 21994 36198
tri 21752 36176 21765 36189 ne
rect 21765 36176 21994 36189
tri 21994 36176 22039 36221 sw
rect 70802 36212 71000 36270
tri 21765 36144 21797 36176 ne
rect 21797 36166 22039 36176
tri 22039 36166 22049 36176 sw
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
rect 21797 36144 22049 36166
tri 21797 36099 21842 36144 ne
rect 21842 36134 22049 36144
tri 22049 36134 22081 36166 sw
rect 21842 36121 22081 36134
tri 22081 36121 22094 36134 sw
rect 21842 36112 22094 36121
rect 21842 36099 21966 36112
tri 21842 36066 21875 36099 ne
rect 21875 36066 21966 36099
rect 22012 36111 22094 36112
tri 22094 36111 22104 36121 sw
rect 22012 36066 22104 36111
tri 22104 36066 22149 36111 sw
rect 70802 36108 71000 36166
tri 21875 36057 21884 36066 ne
rect 21884 36057 22149 36066
tri 21884 36044 21897 36057 ne
rect 21897 36044 22149 36057
tri 22149 36044 22171 36066 sw
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21897 36012 21929 36044 ne
rect 21929 36034 22171 36044
tri 22171 36034 22181 36044 sw
rect 21929 36012 22181 36034
tri 21929 36002 21939 36012 ne
rect 21939 36002 22181 36012
tri 22181 36002 22213 36034 sw
rect 70802 36004 71000 36062
tri 21939 35986 21955 36002 ne
rect 21955 35989 22213 36002
tri 22213 35989 22226 36002 sw
rect 21955 35986 22226 35989
tri 22226 35986 22229 35989 sw
tri 21955 35941 22000 35986 ne
rect 22000 35980 22229 35986
rect 22000 35941 22098 35980
tri 22000 35925 22016 35941 ne
rect 22016 35934 22098 35941
rect 22144 35941 22229 35980
tri 22229 35941 22275 35986 sw
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35934 22275 35941
rect 22016 35925 22275 35934
tri 22016 35912 22029 35925 ne
rect 22029 35912 22275 35925
tri 22275 35912 22303 35941 sw
tri 22029 35880 22061 35912 ne
rect 22061 35902 22303 35912
tri 22303 35902 22313 35912 sw
rect 22061 35880 22313 35902
tri 22061 35835 22106 35880 ne
rect 22106 35870 22313 35880
tri 22313 35870 22345 35902 sw
rect 70802 35900 71000 35958
rect 22106 35857 22345 35870
tri 22345 35857 22358 35870 sw
rect 22106 35848 22358 35857
rect 22106 35835 22230 35848
tri 22106 35793 22148 35835 ne
rect 22148 35802 22230 35835
rect 22276 35837 22358 35848
tri 22358 35837 22378 35857 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 22276 35802 22378 35837
rect 22148 35793 22378 35802
tri 22148 35792 22149 35793 ne
rect 22149 35792 22378 35793
tri 22378 35792 22423 35837 sw
rect 70802 35796 71000 35854
tri 22149 35780 22161 35792 ne
rect 22161 35780 22423 35792
tri 22423 35780 22435 35792 sw
tri 22161 35748 22193 35780 ne
rect 22193 35770 22435 35780
tri 22435 35770 22445 35780 sw
rect 22193 35748 22445 35770
tri 22193 35738 22203 35748 ne
rect 22203 35738 22445 35748
tri 22445 35738 22477 35770 sw
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22203 35693 22248 35738 ne
rect 22248 35725 22477 35738
tri 22477 35725 22490 35738 sw
rect 22248 35716 22490 35725
rect 22248 35693 22362 35716
tri 22248 35661 22280 35693 ne
rect 22280 35670 22362 35693
rect 22408 35693 22490 35716
tri 22490 35693 22522 35725 sw
rect 22408 35670 22522 35693
rect 22280 35661 22522 35670
tri 22280 35648 22293 35661 ne
rect 22293 35648 22522 35661
tri 22522 35648 22567 35693 sw
rect 70802 35692 71000 35750
tri 22293 35616 22325 35648 ne
rect 22325 35638 22567 35648
tri 22567 35638 22577 35648 sw
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 22325 35616 22577 35638
tri 22325 35576 22365 35616 ne
rect 22365 35606 22577 35616
tri 22577 35606 22609 35638 sw
rect 22365 35593 22609 35606
tri 22609 35593 22622 35606 sw
rect 22365 35584 22622 35593
rect 22365 35576 22494 35584
tri 22365 35531 22410 35576 ne
rect 22410 35538 22494 35576
rect 22540 35576 22622 35584
tri 22622 35576 22639 35593 sw
rect 70802 35588 71000 35646
rect 22540 35538 22639 35576
rect 22410 35531 22639 35538
tri 22639 35531 22685 35576 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
tri 22410 35529 22412 35531 ne
rect 22412 35529 22685 35531
tri 22412 35517 22423 35529 ne
rect 22423 35517 22685 35529
tri 22685 35517 22698 35531 sw
tri 22423 35516 22425 35517 ne
rect 22425 35516 22698 35517
tri 22698 35516 22699 35517 sw
tri 22425 35484 22457 35516 ne
rect 22457 35506 22699 35516
tri 22699 35506 22709 35516 sw
rect 22457 35484 22709 35506
tri 22457 35474 22467 35484 ne
rect 22467 35474 22709 35484
tri 22709 35474 22741 35506 sw
rect 70802 35484 71000 35542
tri 22467 35429 22512 35474 ne
rect 22512 35461 22741 35474
tri 22741 35461 22754 35474 sw
rect 22512 35452 22754 35461
rect 22512 35429 22626 35452
tri 22512 35397 22544 35429 ne
rect 22544 35406 22626 35429
rect 22672 35429 22754 35452
tri 22754 35429 22786 35461 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22786 35429
rect 22544 35397 22786 35406
tri 22544 35384 22557 35397 ne
rect 22557 35384 22786 35397
tri 22786 35384 22831 35429 sw
tri 22557 35352 22589 35384 ne
rect 22589 35374 22831 35384
tri 22831 35374 22841 35384 sw
rect 70802 35380 71000 35438
rect 22589 35352 22841 35374
tri 22589 35307 22634 35352 ne
rect 22634 35342 22841 35352
tri 22841 35342 22873 35374 sw
rect 22634 35329 22873 35342
tri 22873 35329 22886 35342 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22634 35320 22886 35329
rect 22634 35307 22758 35320
tri 22634 35301 22639 35307 ne
rect 22639 35301 22758 35307
tri 22639 35256 22685 35301 ne
rect 22685 35274 22758 35301
rect 22804 35297 22886 35320
tri 22886 35297 22918 35329 sw
rect 22804 35274 22918 35297
rect 22685 35256 22918 35274
tri 22685 35243 22698 35256 ne
rect 22698 35252 22918 35256
tri 22918 35252 22963 35297 sw
rect 70802 35276 71000 35334
rect 22698 35243 22963 35252
tri 22963 35243 22972 35252 sw
tri 22698 35211 22730 35243 ne
rect 22730 35242 22972 35243
tri 22972 35242 22973 35243 sw
rect 22730 35211 22973 35242
tri 22730 35210 22731 35211 ne
rect 22731 35210 22973 35211
tri 22973 35210 23005 35242 sw
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22731 35165 22776 35210 ne
rect 22776 35188 23005 35210
rect 22776 35165 22890 35188
tri 22776 35133 22808 35165 ne
rect 22808 35142 22890 35165
rect 22936 35166 23005 35188
tri 23005 35166 23049 35210 sw
rect 70802 35172 71000 35230
rect 22936 35165 23049 35166
tri 23049 35165 23050 35166 sw
rect 22936 35142 23050 35165
rect 22808 35133 23050 35142
tri 22808 35120 22821 35133 ne
rect 22821 35120 23050 35133
tri 23050 35120 23095 35165 sw
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22821 35088 22853 35120 ne
rect 22853 35110 23095 35120
tri 23095 35110 23105 35120 sw
rect 22853 35088 23105 35110
tri 22853 35043 22898 35088 ne
rect 22898 35078 23105 35088
tri 23105 35078 23137 35110 sw
rect 22898 35065 23137 35078
tri 23137 35065 23150 35078 sw
rect 70802 35068 71000 35126
rect 22898 35056 23150 35065
rect 22898 35043 23022 35056
tri 22898 35001 22940 35043 ne
rect 22940 35010 23022 35043
rect 23068 35033 23150 35056
tri 23150 35033 23182 35065 sw
rect 23068 35010 23182 35033
rect 22940 35001 23182 35010
tri 22940 34969 22972 35001 ne
rect 22972 34988 23182 35001
tri 23182 34988 23227 35033 sw
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 22972 34978 23227 34988
tri 23227 34978 23237 34988 sw
rect 22972 34969 23237 34978
tri 23237 34969 23247 34978 sw
tri 22972 34956 22985 34969 ne
rect 22985 34956 23247 34969
tri 22985 34946 22995 34956 ne
rect 22995 34946 23247 34956
tri 23247 34946 23269 34969 sw
rect 70802 34964 71000 35022
tri 22995 34901 23040 34946 ne
rect 23040 34933 23269 34946
tri 23269 34933 23282 34946 sw
rect 23040 34924 23282 34933
rect 23040 34901 23154 34924
tri 23040 34891 23049 34901 ne
rect 23049 34891 23154 34901
tri 23049 34856 23085 34891 ne
rect 23085 34878 23154 34891
rect 23200 34901 23282 34924
tri 23282 34901 23314 34933 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23314 34901
rect 23085 34856 23314 34878
tri 23314 34856 23359 34901 sw
rect 70802 34860 71000 34918
tri 23085 34824 23117 34856 ne
rect 23117 34846 23359 34856
tri 23359 34846 23369 34856 sw
rect 23117 34824 23369 34846
tri 23117 34779 23162 34824 ne
rect 23162 34814 23369 34824
tri 23369 34814 23401 34846 sw
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23162 34801 23401 34814
tri 23401 34801 23414 34814 sw
rect 23162 34792 23414 34801
rect 23162 34779 23286 34792
tri 23162 34737 23204 34779 ne
rect 23204 34746 23286 34779
rect 23332 34769 23414 34792
tri 23414 34769 23446 34801 sw
rect 23332 34746 23446 34769
rect 23204 34737 23446 34746
tri 23204 34694 23247 34737 ne
rect 23247 34724 23446 34737
tri 23446 34724 23491 34769 sw
rect 70802 34756 71000 34814
rect 23247 34714 23491 34724
tri 23491 34714 23501 34724 sw
rect 23247 34694 23501 34714
tri 23501 34694 23521 34714 sw
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23247 34692 23249 34694 ne
rect 23249 34692 23521 34694
tri 23249 34682 23259 34692 ne
rect 23259 34682 23521 34692
tri 23521 34682 23533 34694 sw
tri 23259 34637 23304 34682 ne
rect 23304 34669 23533 34682
tri 23533 34669 23546 34682 sw
rect 23304 34660 23546 34669
rect 23304 34637 23418 34660
tri 23304 34605 23336 34637 ne
rect 23336 34614 23418 34637
rect 23464 34637 23546 34660
tri 23546 34637 23578 34669 sw
rect 70802 34652 71000 34710
rect 23464 34614 23578 34637
rect 23336 34605 23578 34614
tri 23336 34592 23349 34605 ne
rect 23349 34592 23578 34605
tri 23578 34592 23623 34637 sw
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
tri 23349 34560 23381 34592 ne
rect 23381 34582 23623 34592
tri 23623 34582 23633 34592 sw
rect 23381 34560 23633 34582
tri 23381 34527 23414 34560 ne
rect 23414 34550 23633 34560
tri 23633 34550 23665 34582 sw
rect 23414 34537 23665 34550
tri 23665 34537 23678 34550 sw
rect 70802 34548 71000 34606
rect 23414 34528 23678 34537
rect 23414 34527 23550 34528
tri 23414 34481 23459 34527 ne
rect 23459 34482 23550 34527
rect 23596 34527 23678 34528
tri 23678 34527 23689 34537 sw
rect 23596 34482 23689 34527
rect 23459 34481 23689 34482
tri 23689 34481 23734 34527 sw
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
tri 23459 34473 23468 34481 ne
rect 23468 34473 23734 34481
tri 23468 34428 23513 34473 ne
rect 23513 34460 23734 34473
tri 23734 34460 23755 34481 sw
rect 23513 34450 23755 34460
tri 23755 34450 23765 34460 sw
rect 23513 34428 23765 34450
tri 23513 34420 23521 34428 ne
rect 23521 34420 23765 34428
tri 23765 34420 23795 34450 sw
rect 70802 34444 71000 34502
tri 23521 34418 23523 34420 ne
rect 23523 34418 23795 34420
tri 23795 34418 23797 34420 sw
tri 23523 34373 23568 34418 ne
rect 23568 34405 23797 34418
tri 23797 34405 23810 34418 sw
rect 23568 34396 23810 34405
rect 23568 34373 23682 34396
tri 23568 34341 23600 34373 ne
rect 23600 34350 23682 34373
rect 23728 34373 23810 34396
tri 23810 34373 23842 34405 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23728 34350 23842 34373
rect 23600 34341 23842 34350
tri 23600 34328 23613 34341 ne
rect 23613 34328 23842 34341
tri 23842 34328 23887 34373 sw
rect 70802 34340 71000 34398
tri 23613 34296 23645 34328 ne
rect 23645 34318 23887 34328
tri 23887 34318 23897 34328 sw
rect 23645 34296 23897 34318
tri 23645 34286 23655 34296 ne
rect 23655 34286 23897 34296
tri 23897 34286 23929 34318 sw
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23655 34241 23700 34286 ne
rect 23700 34273 23929 34286
tri 23929 34273 23942 34286 sw
rect 23700 34264 23942 34273
rect 23700 34241 23814 34264
tri 23700 34209 23732 34241 ne
rect 23732 34218 23814 34241
rect 23860 34241 23942 34264
tri 23942 34241 23974 34273 sw
rect 23860 34218 23974 34241
rect 23732 34209 23974 34218
tri 23732 34196 23745 34209 ne
rect 23745 34196 23974 34209
tri 23974 34196 24019 34241 sw
rect 70802 34236 71000 34294
tri 23745 34164 23777 34196 ne
rect 23777 34186 24019 34196
tri 24019 34186 24029 34196 sw
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23777 34164 24029 34186
tri 23777 34162 23779 34164 ne
rect 23779 34162 24029 34164
tri 23779 34145 23795 34162 ne
rect 23795 34154 24029 34162
tri 24029 34154 24061 34186 sw
rect 23795 34145 24061 34154
tri 24061 34145 24070 34154 sw
tri 23795 34117 23824 34145 ne
rect 23824 34141 24070 34145
tri 24070 34141 24074 34145 sw
rect 23824 34132 24074 34141
rect 23824 34117 23946 34132
tri 23824 34077 23864 34117 ne
rect 23864 34086 23946 34117
rect 23992 34117 24074 34132
tri 24074 34117 24099 34141 sw
rect 70802 34132 71000 34190
rect 23992 34086 24099 34117
rect 23864 34077 24099 34086
tri 23864 34064 23877 34077 ne
rect 23877 34071 24099 34077
tri 24099 34071 24144 34117 sw
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 23877 34064 24144 34071
tri 24144 34064 24151 34071 sw
tri 23877 34032 23909 34064 ne
rect 23909 34054 24151 34064
tri 24151 34054 24161 34064 sw
rect 23909 34032 24161 34054
tri 23909 34022 23919 34032 ne
rect 23919 34022 24161 34032
tri 24161 34022 24193 34054 sw
rect 70802 34028 71000 34086
tri 23919 33977 23964 34022 ne
rect 23964 34009 24193 34022
tri 24193 34009 24206 34022 sw
rect 23964 34000 24206 34009
rect 23964 33977 24078 34000
tri 23964 33945 23996 33977 ne
rect 23996 33954 24078 33977
rect 24124 33977 24206 34000
tri 24206 33977 24238 34009 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33954 24238 33977
rect 23996 33945 24238 33954
tri 23996 33932 24009 33945 ne
rect 24009 33932 24238 33945
tri 24238 33932 24283 33977 sw
tri 24009 33900 24041 33932 ne
rect 24041 33922 24283 33932
tri 24283 33922 24293 33932 sw
rect 70802 33924 71000 33982
rect 24041 33900 24293 33922
tri 24041 33871 24070 33900 ne
rect 24070 33890 24293 33900
tri 24293 33890 24325 33922 sw
rect 24070 33877 24325 33890
tri 24325 33877 24338 33890 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 24070 33871 24338 33877
tri 24338 33871 24344 33877 sw
tri 24070 33826 24115 33871 ne
rect 24115 33868 24344 33871
rect 24115 33826 24210 33868
tri 24115 33800 24141 33826 ne
rect 24141 33822 24210 33826
rect 24256 33845 24344 33868
tri 24344 33845 24370 33871 sw
rect 24256 33822 24370 33845
rect 24141 33800 24370 33822
tri 24370 33800 24415 33845 sw
rect 70802 33820 71000 33878
tri 24141 33797 24144 33800 ne
rect 24144 33797 24415 33800
tri 24144 33758 24183 33797 ne
rect 24183 33790 24415 33797
tri 24415 33790 24425 33800 sw
rect 24183 33758 24425 33790
tri 24425 33758 24457 33790 sw
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24183 33752 24189 33758 ne
rect 24189 33752 24457 33758
tri 24457 33752 24463 33758 sw
tri 24189 33707 24234 33752 ne
rect 24234 33736 24463 33752
rect 24234 33707 24342 33736
tri 24234 33681 24260 33707 ne
rect 24260 33690 24342 33707
rect 24388 33707 24463 33736
tri 24463 33707 24509 33752 sw
rect 70802 33716 71000 33774
rect 24388 33690 24509 33707
rect 24260 33681 24509 33690
tri 24260 33668 24273 33681 ne
rect 24273 33668 24509 33681
tri 24509 33668 24547 33707 sw
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24273 33636 24305 33668 ne
rect 24305 33658 24547 33668
tri 24547 33658 24557 33668 sw
rect 24305 33636 24557 33658
tri 24305 33597 24344 33636 ne
rect 24344 33626 24557 33636
tri 24557 33626 24589 33658 sw
rect 24344 33613 24589 33626
tri 24589 33613 24602 33626 sw
rect 24344 33604 24602 33613
rect 24344 33597 24474 33604
tri 24344 33551 24389 33597 ne
rect 24389 33558 24474 33597
rect 24520 33597 24602 33604
tri 24602 33597 24619 33613 sw
rect 70802 33612 71000 33670
rect 24520 33581 24619 33597
tri 24619 33581 24634 33597 sw
rect 24520 33558 24634 33581
rect 24389 33551 24634 33558
tri 24389 33549 24392 33551 ne
rect 24392 33549 24634 33551
tri 24392 33536 24405 33549 ne
rect 24405 33536 24634 33549
tri 24634 33536 24679 33581 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
tri 24405 33504 24437 33536 ne
rect 24437 33526 24679 33536
tri 24679 33526 24689 33536 sw
rect 24437 33504 24689 33526
tri 24437 33494 24447 33504 ne
rect 24447 33494 24689 33504
tri 24689 33494 24721 33526 sw
rect 70802 33508 71000 33566
tri 24447 33449 24492 33494 ne
rect 24492 33481 24721 33494
tri 24721 33481 24734 33494 sw
rect 24492 33472 24734 33481
rect 24492 33449 24606 33472
tri 24492 33432 24509 33449 ne
rect 24509 33432 24606 33449
tri 24509 33404 24537 33432 ne
rect 24537 33426 24606 33432
rect 24652 33449 24734 33472
tri 24734 33449 24766 33481 sw
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33426 24766 33449
rect 24537 33404 24766 33426
tri 24766 33404 24811 33449 sw
rect 70802 33404 71000 33462
tri 24537 33372 24569 33404 ne
rect 24569 33394 24811 33404
tri 24811 33394 24821 33404 sw
rect 24569 33372 24821 33394
tri 24569 33327 24614 33372 ne
rect 24614 33362 24821 33372
tri 24821 33362 24853 33394 sw
rect 24614 33342 24853 33362
tri 24853 33342 24873 33362 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 24614 33340 24873 33342
rect 24614 33327 24738 33340
tri 24614 33322 24619 33327 ne
rect 24619 33322 24738 33327
tri 24619 33285 24656 33322 ne
rect 24656 33294 24738 33322
rect 24784 33322 24873 33340
tri 24873 33322 24893 33342 sw
rect 24784 33317 24893 33322
tri 24893 33317 24898 33322 sw
rect 24784 33294 24898 33317
rect 24656 33285 24898 33294
tri 24656 33272 24669 33285 ne
rect 24669 33272 24898 33285
tri 24898 33272 24943 33317 sw
rect 70802 33300 71000 33358
tri 24669 33240 24701 33272 ne
rect 24701 33262 24943 33272
tri 24943 33262 24953 33272 sw
rect 24701 33240 24953 33262
tri 24701 33230 24711 33240 ne
rect 24711 33230 24953 33240
tri 24953 33230 24985 33262 sw
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24711 33185 24756 33230 ne
rect 24756 33217 24985 33230
tri 24985 33217 24998 33230 sw
rect 24756 33208 24998 33217
rect 24756 33185 24870 33208
tri 24756 33153 24788 33185 ne
rect 24788 33162 24870 33185
rect 24916 33185 24998 33208
tri 24998 33185 25030 33217 sw
rect 70802 33196 71000 33254
rect 24916 33162 25030 33185
rect 24788 33153 25030 33162
tri 24788 33140 24801 33153 ne
rect 24801 33140 25030 33153
tri 25030 33140 25075 33185 sw
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24801 33108 24833 33140 ne
rect 24833 33130 25075 33140
tri 25075 33130 25085 33140 sw
rect 24833 33108 25085 33130
tri 24833 33067 24873 33108 ne
rect 24873 33098 25085 33108
tri 25085 33098 25117 33130 sw
rect 24873 33085 25117 33098
tri 25117 33085 25130 33098 sw
rect 70802 33092 71000 33150
rect 24873 33076 25130 33085
rect 24873 33067 25002 33076
tri 24873 33048 24893 33067 ne
rect 24893 33048 25002 33067
tri 24893 33022 24919 33048 ne
rect 24919 33030 25002 33048
rect 25048 33048 25130 33076
tri 25130 33048 25167 33085 sw
rect 25048 33030 25167 33048
rect 24919 33022 25167 33030
tri 25167 33022 25193 33048 sw
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
tri 24919 33021 24920 33022 ne
rect 24920 33021 25193 33022
tri 24920 33008 24933 33021 ne
rect 24933 33008 25193 33021
tri 25193 33008 25207 33022 sw
tri 24933 32976 24965 33008 ne
rect 24965 32998 25207 33008
tri 25207 32998 25217 33008 sw
rect 24965 32976 25217 32998
tri 24965 32966 24975 32976 ne
rect 24975 32966 25217 32976
tri 25217 32966 25249 32998 sw
rect 70802 32988 71000 33046
tri 24975 32921 25020 32966 ne
rect 25020 32953 25249 32966
tri 25249 32953 25262 32966 sw
rect 25020 32944 25262 32953
rect 25020 32921 25134 32944
tri 25020 32889 25052 32921 ne
rect 25052 32898 25134 32921
rect 25180 32921 25262 32944
tri 25262 32921 25294 32953 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32898 25294 32921
rect 25052 32889 25294 32898
tri 25052 32876 25065 32889 ne
rect 25065 32876 25294 32889
tri 25294 32876 25339 32921 sw
rect 70802 32884 71000 32942
tri 25065 32844 25097 32876 ne
rect 25097 32866 25339 32876
tri 25339 32866 25349 32876 sw
rect 25097 32844 25349 32866
tri 25097 32799 25142 32844 ne
rect 25142 32834 25349 32844
tri 25349 32834 25381 32866 sw
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 25142 32821 25381 32834
tri 25381 32821 25394 32834 sw
rect 25142 32819 25394 32821
tri 25394 32819 25397 32821 sw
rect 25142 32812 25397 32819
rect 25142 32799 25266 32812
tri 25142 32773 25167 32799 ne
rect 25167 32773 25266 32799
tri 25167 32757 25184 32773 ne
rect 25184 32766 25266 32773
rect 25312 32773 25397 32812
tri 25397 32773 25442 32819 sw
rect 70802 32780 71000 32838
rect 25312 32766 25442 32773
rect 25184 32757 25442 32766
tri 25184 32744 25197 32757 ne
rect 25197 32744 25442 32757
tri 25442 32744 25471 32773 sw
tri 25197 32712 25229 32744 ne
rect 25229 32734 25471 32744
tri 25471 32734 25481 32744 sw
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
rect 25229 32712 25481 32734
tri 25229 32703 25238 32712 ne
rect 25238 32703 25481 32712
tri 25238 32702 25239 32703 ne
rect 25239 32702 25481 32703
tri 25481 32702 25513 32734 sw
tri 25239 32657 25283 32702 ne
rect 25283 32689 25513 32702
tri 25513 32689 25526 32702 sw
rect 25283 32680 25526 32689
rect 25283 32657 25398 32680
tri 25283 32625 25316 32657 ne
rect 25316 32634 25398 32657
rect 25444 32657 25526 32680
tri 25526 32657 25558 32689 sw
rect 70802 32676 71000 32734
rect 25444 32634 25558 32657
rect 25316 32625 25558 32634
tri 25316 32612 25329 32625 ne
rect 25329 32612 25558 32625
tri 25558 32612 25603 32657 sw
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25329 32580 25361 32612 ne
rect 25361 32602 25603 32612
tri 25603 32602 25613 32612 sw
rect 25361 32580 25613 32602
tri 25361 32535 25406 32580 ne
rect 25406 32570 25613 32580
tri 25613 32570 25645 32602 sw
rect 70802 32572 71000 32630
rect 25406 32557 25645 32570
tri 25645 32557 25658 32570 sw
rect 25406 32548 25658 32557
rect 25406 32535 25530 32548
tri 25406 32499 25442 32535 ne
rect 25442 32502 25530 32535
rect 25576 32544 25658 32548
tri 25658 32544 25671 32557 sw
rect 25576 32502 25671 32544
rect 25442 32499 25671 32502
tri 25671 32499 25716 32544 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
tri 25442 32493 25448 32499 ne
rect 25448 32493 25716 32499
tri 25448 32480 25461 32493 ne
rect 25461 32480 25716 32493
tri 25716 32480 25735 32499 sw
tri 25461 32448 25493 32480 ne
rect 25493 32470 25735 32480
tri 25735 32470 25745 32480 sw
rect 25493 32448 25745 32470
tri 25493 32438 25503 32448 ne
rect 25503 32438 25745 32448
tri 25745 32438 25777 32470 sw
rect 70802 32468 71000 32526
tri 25503 32393 25548 32438 ne
rect 25548 32425 25777 32438
tri 25777 32425 25790 32438 sw
rect 25548 32416 25790 32425
rect 25548 32393 25662 32416
tri 25548 32348 25593 32393 ne
rect 25593 32370 25662 32393
rect 25708 32393 25790 32416
tri 25790 32393 25822 32425 sw
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 25708 32370 25822 32393
rect 25593 32348 25822 32370
tri 25822 32348 25867 32393 sw
rect 70802 32364 71000 32422
tri 25593 32338 25603 32348 ne
rect 25603 32338 25867 32348
tri 25867 32338 25877 32348 sw
tri 25603 32293 25648 32338 ne
rect 25648 32306 25877 32338
tri 25877 32306 25909 32338 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 25648 32293 25909 32306
tri 25909 32293 25922 32306 sw
tri 25648 32247 25693 32293 ne
rect 25693 32284 25923 32293
rect 25693 32247 25794 32284
tri 25693 32229 25712 32247 ne
rect 25712 32238 25794 32247
rect 25840 32247 25923 32284
tri 25923 32247 25968 32293 sw
rect 70802 32260 71000 32318
rect 25840 32238 25968 32247
rect 25712 32229 25968 32238
tri 25712 32225 25716 32229 ne
rect 25716 32225 25968 32229
tri 25968 32225 25991 32247 sw
tri 25716 32216 25725 32225 ne
rect 25725 32216 25991 32225
tri 25991 32216 25999 32225 sw
tri 25725 32184 25757 32216 ne
rect 25757 32206 25999 32216
tri 25999 32206 26009 32216 sw
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
rect 25757 32184 26009 32206
tri 25757 32174 25767 32184 ne
rect 25767 32174 26009 32184
tri 26009 32174 26041 32206 sw
tri 25767 32129 25812 32174 ne
rect 25812 32161 26041 32174
tri 26041 32161 26054 32174 sw
rect 25812 32152 26054 32161
rect 25812 32129 25926 32152
tri 25812 32097 25844 32129 ne
rect 25844 32106 25926 32129
rect 25972 32129 26054 32152
tri 26054 32129 26086 32161 sw
rect 70802 32156 71000 32214
rect 25972 32106 26086 32129
rect 25844 32097 26086 32106
tri 25844 32084 25857 32097 ne
rect 25857 32084 26086 32097
tri 26086 32084 26131 32129 sw
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
tri 25857 32052 25889 32084 ne
rect 25889 32074 26131 32084
tri 26131 32074 26141 32084 sw
rect 25889 32052 26141 32074
tri 25889 32007 25934 32052 ne
rect 25934 32042 26141 32052
tri 26141 32042 26173 32074 sw
rect 70802 32052 71000 32110
rect 25934 32029 26173 32042
tri 26173 32029 26186 32042 sw
rect 25934 32020 26186 32029
rect 25934 32007 26058 32020
tri 25934 31973 25968 32007 ne
rect 25968 31974 26058 32007
rect 26104 31997 26186 32020
tri 26186 31997 26218 32029 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31974 26218 31997
rect 25968 31973 26218 31974
tri 25968 31950 25991 31973 ne
rect 25991 31952 26218 31973
tri 26218 31952 26263 31997 sw
rect 25991 31950 26263 31952
tri 26263 31950 26265 31952 sw
tri 25991 31920 26021 31950 ne
rect 26021 31942 26265 31950
tri 26265 31942 26273 31950 sw
rect 70802 31948 71000 32006
rect 26021 31920 26273 31942
tri 26021 31910 26031 31920 ne
rect 26031 31910 26273 31920
tri 26273 31910 26305 31942 sw
tri 26031 31865 26076 31910 ne
rect 26076 31888 26305 31910
rect 26076 31865 26190 31888
tri 26076 31833 26108 31865 ne
rect 26108 31842 26190 31865
rect 26236 31883 26305 31888
tri 26305 31883 26333 31910 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26236 31865 26333 31883
tri 26333 31865 26350 31883 sw
rect 26236 31842 26350 31865
rect 26108 31833 26350 31842
tri 26108 31820 26121 31833 ne
rect 26121 31820 26350 31833
tri 26350 31820 26395 31865 sw
rect 70802 31844 71000 31902
tri 26121 31788 26153 31820 ne
rect 26153 31810 26395 31820
tri 26395 31810 26405 31820 sw
rect 26153 31788 26405 31810
tri 26153 31743 26198 31788 ne
rect 26198 31778 26405 31788
tri 26405 31778 26437 31810 sw
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26198 31765 26437 31778
tri 26437 31765 26450 31778 sw
rect 26198 31756 26450 31765
rect 26198 31743 26322 31756
tri 26198 31701 26240 31743 ne
rect 26240 31710 26322 31743
rect 26368 31733 26450 31756
tri 26450 31733 26482 31765 sw
rect 70802 31740 71000 31798
rect 26368 31710 26482 31733
rect 26240 31701 26482 31710
tri 26240 31676 26265 31701 ne
rect 26265 31688 26482 31701
tri 26482 31688 26527 31733 sw
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 26265 31678 26527 31688
tri 26527 31678 26537 31688 sw
rect 26265 31676 26537 31678
tri 26537 31676 26539 31678 sw
tri 26265 31656 26285 31676 ne
rect 26285 31656 26539 31676
tri 26285 31646 26295 31656 ne
rect 26295 31646 26539 31656
tri 26539 31646 26569 31676 sw
tri 26295 31608 26333 31646 ne
rect 26333 31633 26569 31646
tri 26569 31633 26582 31646 sw
rect 70802 31636 71000 31694
rect 26333 31624 26582 31633
rect 26333 31608 26454 31624
tri 26333 31563 26378 31608 ne
rect 26378 31578 26454 31608
rect 26500 31608 26582 31624
tri 26582 31608 26607 31633 sw
rect 26500 31578 26607 31608
rect 26378 31563 26607 31578
tri 26607 31563 26652 31608 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
tri 26378 31556 26385 31563 ne
rect 26385 31556 26652 31563
tri 26652 31556 26659 31563 sw
tri 26385 31524 26417 31556 ne
rect 26417 31546 26659 31556
tri 26659 31546 26669 31556 sw
rect 26417 31524 26669 31546
tri 26417 31479 26462 31524 ne
rect 26462 31514 26669 31524
tri 26669 31514 26701 31546 sw
rect 70802 31532 71000 31590
rect 26462 31501 26701 31514
tri 26701 31501 26714 31514 sw
rect 26462 31492 26714 31501
rect 26462 31479 26586 31492
tri 26462 31437 26504 31479 ne
rect 26504 31446 26586 31479
rect 26632 31469 26714 31492
tri 26714 31469 26746 31501 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31446 26746 31469
rect 26504 31437 26746 31446
tri 26504 31401 26539 31437 ne
rect 26539 31424 26746 31437
tri 26746 31424 26791 31469 sw
rect 70802 31428 71000 31486
rect 26539 31414 26791 31424
tri 26791 31414 26801 31424 sw
rect 26539 31401 26801 31414
tri 26801 31401 26814 31414 sw
tri 26539 31392 26549 31401 ne
rect 26549 31392 26814 31401
tri 26549 31382 26559 31392 ne
rect 26559 31382 26814 31392
tri 26814 31382 26833 31401 sw
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26559 31337 26604 31382 ne
rect 26604 31369 26833 31382
tri 26833 31369 26846 31382 sw
rect 26604 31360 26846 31369
rect 26604 31337 26718 31360
tri 26604 31305 26636 31337 ne
rect 26636 31314 26718 31337
rect 26764 31337 26846 31360
tri 26846 31337 26878 31369 sw
rect 26764 31314 26878 31337
rect 26636 31305 26878 31314
tri 26636 31292 26649 31305 ne
rect 26649 31292 26878 31305
tri 26878 31292 26923 31337 sw
rect 70802 31324 71000 31382
tri 26649 31260 26681 31292 ne
rect 26681 31282 26923 31292
tri 26923 31282 26933 31292 sw
rect 26681 31260 26933 31282
tri 26681 31243 26697 31260 ne
rect 26697 31250 26933 31260
tri 26933 31250 26965 31282 sw
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26697 31243 26965 31250
tri 26697 31198 26743 31243 ne
rect 26743 31237 26965 31243
tri 26965 31237 26978 31250 sw
rect 26743 31228 26978 31237
rect 26743 31198 26850 31228
tri 26743 31173 26768 31198 ne
rect 26768 31182 26850 31198
rect 26896 31198 26978 31228
tri 26978 31198 27017 31237 sw
rect 70802 31220 71000 31278
rect 26896 31182 27017 31198
rect 26768 31173 27017 31182
tri 26768 31128 26813 31173 ne
rect 26813 31160 27017 31173
tri 27017 31160 27055 31198 sw
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 26813 31153 27055 31160
tri 27055 31153 27062 31160 sw
rect 26813 31150 27062 31153
tri 27062 31150 27065 31153 sw
rect 26813 31128 27065 31150
tri 26813 31127 26814 31128 ne
rect 26814 31127 27065 31128
tri 27065 31127 27088 31150 sw
tri 26814 31118 26823 31127 ne
rect 26823 31118 27088 31127
tri 27088 31118 27097 31127 sw
tri 26823 31073 26868 31118 ne
rect 26868 31105 27097 31118
tri 27097 31105 27110 31118 sw
rect 70802 31116 71000 31174
rect 26868 31096 27110 31105
rect 26868 31073 26982 31096
tri 26868 31041 26900 31073 ne
rect 26900 31050 26982 31073
rect 27028 31073 27110 31096
tri 27110 31073 27142 31105 sw
rect 27028 31050 27142 31073
rect 26900 31041 27142 31050
tri 26900 31028 26913 31041 ne
rect 26913 31028 27142 31041
tri 27142 31028 27187 31073 sw
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
tri 26913 30996 26945 31028 ne
rect 26945 31018 27187 31028
tri 27187 31018 27197 31028 sw
rect 26945 30996 27197 31018
tri 26945 30951 26990 30996 ne
rect 26990 30986 27197 30996
tri 27197 30986 27229 31018 sw
rect 70802 31012 71000 31070
rect 26990 30973 27229 30986
tri 27229 30973 27242 30986 sw
rect 26990 30964 27242 30973
rect 26990 30951 27114 30964
tri 26990 30909 27032 30951 ne
rect 27032 30918 27114 30951
rect 27160 30941 27242 30964
tri 27242 30941 27274 30973 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27160 30918 27274 30941
rect 27032 30909 27274 30918
tri 27032 30864 27077 30909 ne
rect 27077 30896 27274 30909
tri 27274 30896 27319 30941 sw
rect 70802 30908 71000 30966
rect 27077 30886 27319 30896
tri 27319 30886 27329 30896 sw
rect 27077 30864 27329 30886
tri 27077 30853 27088 30864 ne
rect 27088 30854 27329 30864
tri 27329 30854 27361 30886 sw
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27088 30853 27361 30854
tri 27361 30853 27363 30854 sw
tri 27088 30833 27107 30853 ne
rect 27107 30841 27363 30853
tri 27363 30841 27374 30853 sw
rect 27107 30833 27374 30841
tri 27374 30833 27382 30841 sw
tri 27107 30788 27153 30833 ne
rect 27153 30832 27382 30833
rect 27153 30788 27246 30832
tri 27153 30777 27164 30788 ne
rect 27164 30786 27246 30788
rect 27292 30788 27382 30832
tri 27382 30788 27427 30833 sw
rect 70802 30804 71000 30862
rect 27292 30786 27427 30788
rect 27164 30777 27427 30786
tri 27164 30764 27177 30777 ne
rect 27177 30764 27427 30777
tri 27427 30764 27451 30788 sw
tri 27177 30732 27209 30764 ne
rect 27209 30754 27451 30764
tri 27451 30754 27461 30764 sw
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
rect 27209 30732 27461 30754
tri 27209 30722 27219 30732 ne
rect 27219 30722 27461 30732
tri 27461 30722 27493 30754 sw
tri 27219 30677 27264 30722 ne
rect 27264 30709 27493 30722
tri 27493 30709 27506 30722 sw
rect 27264 30700 27506 30709
rect 27264 30677 27378 30700
tri 27264 30645 27296 30677 ne
rect 27296 30654 27378 30677
rect 27424 30677 27506 30700
tri 27506 30677 27538 30709 sw
rect 70802 30700 71000 30758
rect 27424 30654 27538 30677
rect 27296 30645 27538 30654
tri 27296 30632 27309 30645 ne
rect 27309 30632 27538 30645
tri 27538 30632 27583 30677 sw
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27309 30600 27341 30632 ne
rect 27341 30622 27583 30632
tri 27583 30622 27593 30632 sw
rect 27341 30600 27593 30622
tri 27341 30578 27363 30600 ne
rect 27363 30590 27593 30600
tri 27593 30590 27625 30622 sw
rect 70802 30596 71000 30654
rect 27363 30578 27625 30590
tri 27625 30578 27637 30590 sw
tri 27363 30533 27408 30578 ne
rect 27408 30577 27637 30578
tri 27637 30577 27638 30578 sw
rect 27408 30568 27638 30577
rect 27408 30533 27510 30568
tri 27408 30514 27427 30533 ne
rect 27427 30522 27510 30533
rect 27556 30545 27638 30568
tri 27638 30545 27670 30577 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30522 27670 30545
rect 27427 30514 27670 30522
tri 27427 30500 27441 30514 ne
rect 27441 30500 27670 30514
tri 27670 30500 27715 30545 sw
tri 27441 30468 27473 30500 ne
rect 27473 30490 27715 30500
tri 27715 30490 27725 30500 sw
rect 70802 30492 71000 30550
rect 27473 30468 27725 30490
tri 27473 30458 27483 30468 ne
rect 27483 30458 27725 30468
tri 27725 30458 27757 30490 sw
tri 27483 30413 27528 30458 ne
rect 27528 30436 27757 30458
rect 27528 30413 27642 30436
tri 27528 30381 27560 30413 ne
rect 27560 30390 27642 30413
rect 27688 30423 27757 30436
tri 27757 30423 27792 30458 sw
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 27688 30413 27792 30423
tri 27792 30413 27802 30423 sw
rect 27688 30390 27802 30413
rect 27560 30381 27802 30390
tri 27560 30368 27573 30381 ne
rect 27573 30368 27802 30381
tri 27802 30368 27847 30413 sw
rect 70802 30388 71000 30446
tri 27573 30336 27605 30368 ne
rect 27605 30358 27847 30368
tri 27847 30358 27857 30368 sw
rect 27605 30336 27857 30358
tri 27605 30304 27637 30336 ne
rect 27637 30326 27857 30336
tri 27857 30326 27889 30358 sw
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
rect 27637 30313 27889 30326
tri 27889 30313 27902 30326 sw
rect 27637 30304 27902 30313
tri 27902 30304 27911 30313 sw
tri 27637 30259 27682 30304 ne
rect 27682 30259 27774 30304
tri 27682 30249 27692 30259 ne
rect 27692 30258 27774 30259
rect 27820 30281 27911 30304
tri 27911 30281 27934 30304 sw
rect 70802 30284 71000 30342
rect 27820 30258 27934 30281
rect 27692 30249 27934 30258
tri 27692 30236 27705 30249 ne
rect 27705 30236 27934 30249
tri 27934 30236 27979 30281 sw
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27705 30204 27737 30236 ne
rect 27737 30226 27979 30236
tri 27979 30226 27989 30236 sw
rect 27737 30204 27989 30226
tri 27737 30194 27747 30204 ne
rect 27747 30194 27989 30204
tri 27989 30194 28021 30226 sw
tri 27747 30149 27792 30194 ne
rect 27792 30181 28021 30194
tri 28021 30181 28034 30194 sw
rect 27792 30172 28034 30181
rect 27792 30149 27906 30172
tri 27792 30104 27837 30149 ne
rect 27837 30126 27906 30149
rect 27952 30149 28034 30172
tri 28034 30149 28066 30181 sw
rect 70802 30180 71000 30238
rect 27952 30126 28066 30149
rect 27837 30104 28066 30126
tri 28066 30104 28111 30149 sw
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
tri 27837 30072 27869 30104 ne
rect 27869 30072 28111 30104
tri 27869 30029 27911 30072 ne
rect 27911 30062 28111 30072
tri 28111 30062 28153 30104 sw
rect 70802 30076 71000 30134
rect 27911 30049 28153 30062
tri 28153 30049 28166 30062 sw
rect 27911 30040 28166 30049
rect 27911 30029 28038 30040
tri 27911 29985 27956 30029 ne
rect 27956 29994 28038 30029
rect 28084 30029 28166 30040
tri 28166 30029 28186 30049 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 30017 28186 30029
tri 28186 30017 28198 30029 sw
rect 28084 29994 28198 30017
rect 27956 29985 28198 29994
tri 27956 29972 27969 29985 ne
rect 27969 29972 28198 29985
tri 28198 29972 28243 30017 sw
rect 70802 29972 71000 30030
tri 27969 29940 28001 29972 ne
rect 28001 29962 28243 29972
tri 28243 29962 28253 29972 sw
rect 28001 29940 28253 29962
tri 28001 29930 28011 29940 ne
rect 28011 29930 28253 29940
tri 28253 29930 28285 29962 sw
tri 28011 29885 28056 29930 ne
rect 28056 29917 28285 29930
tri 28285 29917 28298 29930 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28056 29908 28298 29917
rect 28056 29885 28170 29908
tri 28056 29853 28088 29885 ne
rect 28088 29862 28170 29885
rect 28216 29885 28298 29908
tri 28298 29885 28330 29917 sw
rect 28216 29862 28330 29885
rect 28088 29853 28330 29862
tri 28088 29840 28101 29853 ne
rect 28101 29840 28330 29853
tri 28330 29840 28375 29885 sw
rect 70802 29868 71000 29926
tri 28101 29808 28133 29840 ne
rect 28133 29830 28375 29840
tri 28375 29830 28385 29840 sw
rect 28133 29808 28385 29830
tri 28133 29784 28157 29808 ne
rect 28157 29798 28385 29808
tri 28385 29798 28417 29830 sw
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28157 29785 28417 29798
tri 28417 29785 28430 29798 sw
rect 28157 29784 28430 29785
tri 28157 29755 28186 29784 ne
rect 28186 29776 28430 29784
rect 28186 29755 28302 29776
tri 28186 29739 28202 29755 ne
rect 28202 29739 28302 29755
tri 28202 29721 28220 29739 ne
rect 28220 29730 28302 29739
rect 28348 29755 28430 29776
tri 28430 29755 28460 29785 sw
rect 70802 29764 71000 29822
rect 28348 29739 28460 29755
tri 28460 29739 28476 29755 sw
rect 28348 29730 28476 29739
rect 28220 29721 28476 29730
tri 28220 29708 28233 29721 ne
rect 28233 29708 28476 29721
tri 28476 29708 28507 29739 sw
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28233 29676 28265 29708 ne
rect 28265 29698 28507 29708
tri 28507 29698 28517 29708 sw
rect 28265 29676 28517 29698
tri 28265 29666 28275 29676 ne
rect 28275 29666 28517 29676
tri 28517 29666 28549 29698 sw
tri 28275 29621 28320 29666 ne
rect 28320 29653 28549 29666
tri 28549 29653 28562 29666 sw
rect 70802 29660 71000 29718
rect 28320 29644 28562 29653
rect 28320 29621 28434 29644
tri 28320 29589 28352 29621 ne
rect 28352 29598 28434 29621
rect 28480 29621 28562 29644
tri 28562 29621 28594 29653 sw
rect 28480 29598 28594 29621
rect 28352 29589 28594 29598
tri 28352 29576 28365 29589 ne
rect 28365 29576 28594 29589
tri 28594 29576 28639 29621 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
tri 28365 29544 28397 29576 ne
rect 28397 29566 28639 29576
tri 28639 29566 28649 29576 sw
rect 28397 29544 28649 29566
tri 28397 29499 28442 29544 ne
rect 28442 29534 28649 29544
tri 28649 29534 28681 29566 sw
rect 70802 29556 71000 29614
rect 28442 29521 28681 29534
tri 28681 29521 28694 29534 sw
rect 28442 29512 28694 29521
rect 28442 29499 28566 29512
tri 28442 29481 28460 29499 ne
rect 28460 29481 28566 29499
tri 28460 29457 28484 29481 ne
rect 28484 29466 28566 29481
rect 28612 29481 28694 29512
tri 28694 29481 28735 29521 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28735 29481
rect 28484 29457 28735 29466
tri 28484 29444 28497 29457 ne
rect 28497 29444 28735 29457
tri 28735 29444 28771 29481 sw
rect 70802 29452 71000 29510
tri 28497 29412 28529 29444 ne
rect 28529 29434 28771 29444
tri 28771 29434 28781 29444 sw
rect 28529 29412 28781 29434
tri 28529 29402 28539 29412 ne
rect 28539 29402 28781 29412
tri 28781 29402 28813 29434 sw
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28539 29374 28567 29402 ne
rect 28567 29389 28813 29402
tri 28813 29389 28826 29402 sw
rect 28567 29380 28826 29389
rect 28567 29374 28698 29380
tri 28567 29329 28612 29374 ne
rect 28612 29334 28698 29374
rect 28744 29374 28826 29380
tri 28826 29374 28841 29389 sw
rect 28744 29334 28841 29374
rect 28612 29329 28841 29334
tri 28841 29329 28886 29374 sw
rect 70802 29348 71000 29406
tri 28612 29325 28616 29329 ne
rect 28616 29325 28886 29329
tri 28616 29312 28629 29325 ne
rect 28629 29312 28886 29325
tri 28886 29312 28903 29329 sw
tri 28629 29280 28661 29312 ne
rect 28661 29302 28903 29312
tri 28903 29302 28913 29312 sw
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
rect 28661 29280 28913 29302
tri 28661 29235 28706 29280 ne
rect 28706 29270 28913 29280
tri 28913 29270 28945 29302 sw
rect 28706 29257 28945 29270
tri 28945 29257 28958 29270 sw
rect 28706 29251 28958 29257
tri 28958 29251 28964 29257 sw
rect 28706 29248 28964 29251
rect 28706 29235 28830 29248
tri 28706 29206 28735 29235 ne
rect 28735 29206 28830 29235
tri 28735 29193 28748 29206 ne
rect 28748 29202 28830 29206
rect 28876 29206 28964 29248
tri 28964 29206 29009 29251 sw
rect 70802 29244 71000 29302
rect 28876 29202 29009 29206
rect 28748 29193 29009 29202
tri 28748 29180 28761 29193 ne
rect 28761 29180 29009 29193
tri 29009 29180 29035 29206 sw
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28761 29148 28793 29180 ne
rect 28793 29170 29035 29180
tri 29035 29170 29045 29180 sw
rect 28793 29148 29045 29170
tri 28793 29138 28803 29148 ne
rect 28803 29138 29045 29148
tri 29045 29138 29077 29170 sw
rect 70802 29140 71000 29198
tri 28803 29093 28848 29138 ne
rect 28848 29125 29077 29138
tri 29077 29125 29090 29138 sw
rect 28848 29116 29090 29125
rect 28848 29093 28962 29116
tri 28848 29055 28886 29093 ne
rect 28886 29070 28962 29093
rect 29008 29093 29090 29116
tri 29090 29093 29122 29125 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 29008 29070 29122 29093
rect 28886 29055 29122 29070
tri 28886 29048 28893 29055 ne
rect 28893 29048 29122 29055
tri 29122 29048 29167 29093 sw
tri 28893 29009 28931 29048 ne
rect 28931 29038 29167 29048
tri 29167 29038 29177 29048 sw
rect 28931 29009 29177 29038
tri 28931 28964 28977 29009 ne
rect 28977 29006 29177 29009
tri 29177 29006 29209 29038 sw
rect 70802 29036 71000 29094
rect 28977 28984 29209 29006
rect 28977 28964 29094 28984
tri 28977 28932 29009 28964 ne
rect 29009 28938 29094 28964
rect 29140 28964 29209 28984
tri 29209 28964 29251 29006 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29140 28938 29251 28964
rect 29009 28932 29251 28938
tri 29251 28932 29283 28964 sw
rect 70802 28932 71000 28990
tri 29009 28929 29012 28932 ne
rect 29012 28929 29283 28932
tri 29012 28916 29025 28929 ne
rect 29025 28916 29283 28929
tri 29283 28916 29299 28932 sw
tri 29025 28884 29057 28916 ne
rect 29057 28906 29299 28916
tri 29299 28906 29309 28916 sw
rect 29057 28884 29309 28906
tri 29057 28874 29067 28884 ne
rect 29067 28874 29309 28884
tri 29309 28874 29341 28906 sw
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29067 28829 29112 28874 ne
rect 29112 28861 29341 28874
tri 29341 28861 29354 28874 sw
rect 29112 28852 29354 28861
rect 29112 28829 29226 28852
tri 29112 28797 29144 28829 ne
rect 29144 28806 29226 28829
rect 29272 28829 29354 28852
tri 29354 28829 29386 28861 sw
rect 29272 28806 29386 28829
rect 29144 28797 29386 28806
tri 29144 28784 29157 28797 ne
rect 29157 28784 29386 28797
tri 29386 28784 29431 28829 sw
rect 70802 28828 71000 28886
tri 29157 28752 29189 28784 ne
rect 29189 28774 29431 28784
tri 29431 28774 29441 28784 sw
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29189 28752 29441 28774
tri 29189 28707 29234 28752 ne
rect 29234 28742 29441 28752
tri 29441 28742 29473 28774 sw
rect 29234 28729 29473 28742
tri 29473 28729 29486 28742 sw
rect 29234 28720 29486 28729
rect 29234 28707 29358 28720
tri 29234 28690 29251 28707 ne
rect 29251 28690 29358 28707
tri 29251 28657 29283 28690 ne
rect 29283 28674 29358 28690
rect 29404 28703 29486 28720
tri 29486 28703 29513 28729 sw
rect 70802 28724 71000 28782
rect 29404 28674 29513 28703
rect 29283 28657 29513 28674
tri 29513 28657 29558 28703 sw
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
tri 29283 28652 29289 28657 ne
rect 29289 28652 29558 28657
tri 29558 28652 29563 28657 sw
tri 29289 28620 29321 28652 ne
rect 29321 28645 29563 28652
tri 29563 28645 29571 28652 sw
rect 29321 28620 29571 28645
tri 29321 28610 29331 28620 ne
rect 29331 28610 29571 28620
tri 29571 28610 29605 28645 sw
rect 70802 28620 71000 28678
tri 29331 28565 29376 28610 ne
rect 29376 28597 29605 28610
tri 29605 28597 29618 28610 sw
rect 29376 28588 29618 28597
rect 29376 28565 29490 28588
tri 29376 28533 29408 28565 ne
rect 29408 28542 29490 28565
rect 29536 28565 29618 28588
tri 29618 28565 29650 28597 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29650 28565
rect 29408 28533 29650 28542
tri 29408 28520 29421 28533 ne
rect 29421 28520 29650 28533
tri 29650 28520 29695 28565 sw
tri 29421 28488 29453 28520 ne
rect 29453 28510 29695 28520
tri 29695 28510 29705 28520 sw
rect 70802 28516 71000 28574
rect 29453 28488 29705 28510
tri 29453 28443 29498 28488 ne
rect 29498 28478 29705 28488
tri 29705 28478 29737 28510 sw
rect 29498 28465 29737 28478
tri 29737 28465 29750 28478 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29498 28456 29750 28465
rect 29498 28443 29622 28456
tri 29498 28401 29540 28443 ne
rect 29540 28410 29622 28443
rect 29668 28433 29750 28456
tri 29750 28433 29782 28465 sw
rect 29668 28410 29782 28433
rect 29540 28401 29782 28410
tri 29540 28383 29558 28401 ne
rect 29558 28388 29782 28401
tri 29782 28388 29827 28433 sw
rect 70802 28412 71000 28470
rect 29558 28383 29827 28388
tri 29827 28383 29832 28388 sw
tri 29558 28356 29585 28383 ne
rect 29585 28378 29832 28383
tri 29832 28378 29837 28383 sw
rect 29585 28356 29837 28378
tri 29585 28346 29595 28356 ne
rect 29595 28346 29837 28356
tri 29837 28346 29869 28378 sw
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29595 28325 29616 28346 ne
rect 29616 28333 29869 28346
tri 29869 28333 29882 28346 sw
rect 29616 28325 29882 28333
tri 29882 28325 29890 28333 sw
tri 29616 28280 29661 28325 ne
rect 29661 28324 29890 28325
rect 29661 28280 29754 28324
tri 29661 28269 29672 28280 ne
rect 29672 28278 29754 28280
rect 29800 28280 29890 28324
tri 29890 28280 29935 28325 sw
rect 70802 28308 71000 28366
rect 29800 28278 29935 28280
rect 29672 28269 29935 28278
tri 29672 28256 29685 28269 ne
rect 29685 28256 29935 28269
tri 29935 28256 29959 28280 sw
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29685 28224 29717 28256 ne
rect 29717 28246 29959 28256
tri 29959 28246 29969 28256 sw
rect 29717 28224 29969 28246
tri 29717 28179 29762 28224 ne
rect 29762 28214 29969 28224
tri 29969 28214 30001 28246 sw
rect 29762 28201 30001 28214
tri 30001 28201 30014 28214 sw
rect 70802 28204 71000 28262
rect 29762 28192 30014 28201
rect 29762 28179 29886 28192
tri 29762 28137 29804 28179 ne
rect 29804 28146 29886 28179
rect 29932 28169 30014 28192
tri 30014 28169 30046 28201 sw
rect 29932 28146 30046 28169
rect 29804 28137 30046 28146
tri 29804 28109 29832 28137 ne
rect 29832 28124 30046 28137
tri 30046 28124 30091 28169 sw
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29832 28114 30091 28124
tri 30091 28114 30101 28124 sw
rect 29832 28109 30101 28114
tri 30101 28109 30107 28114 sw
tri 29832 28092 29849 28109 ne
rect 29849 28092 30107 28109
tri 29849 28082 29859 28092 ne
rect 29859 28082 30107 28092
tri 30107 28082 30133 28109 sw
rect 70802 28100 71000 28158
tri 29859 28037 29904 28082 ne
rect 29904 28069 30133 28082
tri 30133 28069 30146 28082 sw
rect 29904 28060 30146 28069
rect 29904 28037 30018 28060
tri 29904 28005 29936 28037 ne
rect 29936 28014 30018 28037
rect 30064 28037 30146 28060
tri 30146 28037 30178 28069 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30178 28037
rect 29936 28005 30178 28014
tri 29936 27992 29949 28005 ne
rect 29949 27992 30178 28005
tri 30178 27992 30223 28037 sw
rect 70802 27996 71000 28054
tri 29949 27960 29981 27992 ne
rect 29981 27982 30223 27992
tri 30223 27982 30233 27992 sw
rect 29981 27960 30233 27982
tri 29981 27915 30026 27960 ne
rect 30026 27950 30233 27960
tri 30233 27950 30265 27982 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30026 27937 30265 27950
tri 30265 27937 30278 27950 sw
rect 30026 27928 30278 27937
rect 30026 27915 30150 27928
tri 30026 27873 30068 27915 ne
rect 30068 27882 30150 27915
rect 30196 27915 30278 27928
tri 30278 27915 30300 27937 sw
rect 30196 27882 30300 27915
rect 30068 27873 30300 27882
tri 30068 27834 30107 27873 ne
rect 30107 27870 30300 27873
tri 30300 27870 30345 27915 sw
rect 70802 27892 71000 27950
rect 30107 27860 30345 27870
tri 30345 27860 30355 27870 sw
rect 30107 27850 30355 27860
tri 30355 27850 30365 27860 sw
rect 30107 27834 30365 27850
tri 30365 27834 30381 27850 sw
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30107 27828 30113 27834 ne
rect 30113 27828 30381 27834
tri 30113 27818 30123 27828 ne
rect 30123 27818 30381 27828
tri 30381 27818 30397 27834 sw
tri 30123 27773 30168 27818 ne
rect 30168 27805 30397 27818
tri 30397 27805 30410 27818 sw
rect 30168 27796 30410 27805
rect 30168 27773 30282 27796
tri 30168 27741 30200 27773 ne
rect 30200 27750 30282 27773
rect 30328 27773 30410 27796
tri 30410 27773 30442 27805 sw
rect 70802 27788 71000 27846
rect 30328 27750 30442 27773
rect 30200 27741 30442 27750
tri 30200 27728 30213 27741 ne
rect 30213 27728 30442 27741
tri 30442 27728 30487 27773 sw
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30213 27696 30245 27728 ne
rect 30245 27718 30487 27728
tri 30487 27718 30497 27728 sw
rect 30245 27696 30497 27718
tri 30245 27651 30290 27696 ne
rect 30290 27686 30497 27696
tri 30497 27686 30529 27718 sw
rect 30290 27673 30529 27686
tri 30529 27673 30542 27686 sw
rect 70802 27684 71000 27742
rect 30290 27664 30542 27673
rect 30290 27651 30414 27664
tri 30290 27641 30300 27651 ne
rect 30300 27641 30414 27651
tri 30300 27595 30345 27641 ne
rect 30345 27618 30414 27641
rect 30460 27641 30542 27664
tri 30542 27641 30574 27673 sw
rect 30460 27618 30574 27641
rect 30345 27596 30574 27618
tri 30574 27596 30619 27641 sw
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30345 27595 30619 27596
tri 30345 27560 30381 27595 ne
rect 30381 27586 30619 27595
tri 30619 27586 30629 27596 sw
rect 30381 27560 30629 27586
tri 30629 27560 30655 27586 sw
rect 70802 27580 71000 27638
tri 30381 27554 30387 27560 ne
rect 30387 27554 30655 27560
tri 30655 27554 30661 27560 sw
tri 30387 27550 30391 27554 ne
rect 30391 27550 30661 27554
tri 30661 27550 30665 27554 sw
tri 30391 27505 30436 27550 ne
rect 30436 27532 30665 27550
rect 30436 27505 30546 27532
tri 30436 27477 30464 27505 ne
rect 30464 27486 30546 27505
rect 30592 27505 30665 27532
tri 30665 27505 30710 27550 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30592 27486 30710 27505
rect 30464 27477 30710 27486
tri 30464 27464 30477 27477 ne
rect 30477 27464 30710 27477
tri 30710 27464 30751 27505 sw
rect 70802 27476 71000 27534
tri 30477 27432 30509 27464 ne
rect 30509 27454 30751 27464
tri 30751 27454 30761 27464 sw
rect 30509 27432 30761 27454
tri 30509 27387 30554 27432 ne
rect 30554 27422 30761 27432
tri 30761 27422 30793 27454 sw
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
rect 30554 27409 30793 27422
tri 30793 27409 30806 27422 sw
rect 30554 27400 30806 27409
rect 30554 27387 30678 27400
tri 30554 27345 30596 27387 ne
rect 30596 27354 30678 27387
rect 30724 27377 30806 27400
tri 30806 27377 30838 27409 sw
rect 30724 27354 30838 27377
rect 30596 27345 30838 27354
tri 30596 27300 30641 27345 ne
rect 30641 27332 30838 27345
tri 30838 27332 30883 27377 sw
rect 70802 27372 71000 27430
rect 30641 27322 30883 27332
tri 30883 27322 30893 27332 sw
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 30641 27300 30893 27322
tri 30641 27285 30655 27300 ne
rect 30655 27290 30893 27300
tri 30893 27290 30925 27322 sw
rect 30655 27285 30925 27290
tri 30925 27285 30930 27290 sw
tri 30655 27240 30701 27285 ne
rect 30701 27277 30930 27285
tri 30930 27277 30938 27285 sw
rect 30701 27268 30938 27277
rect 30701 27240 30810 27268
tri 30701 27231 30710 27240 ne
rect 30710 27231 30810 27240
tri 30710 27200 30741 27231 ne
rect 30741 27222 30810 27231
rect 30856 27245 30938 27268
tri 30938 27245 30970 27277 sw
rect 70802 27268 71000 27326
rect 30856 27222 30970 27245
rect 30741 27200 30970 27222
tri 30970 27200 31015 27245 sw
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30741 27168 30773 27200 ne
rect 30773 27190 31015 27200
tri 31015 27190 31025 27200 sw
rect 30773 27168 31025 27190
tri 30773 27158 30783 27168 ne
rect 30783 27158 31025 27168
tri 31025 27158 31057 27190 sw
rect 70802 27164 71000 27222
tri 30783 27113 30828 27158 ne
rect 30828 27140 31057 27158
tri 31057 27140 31075 27158 sw
rect 30828 27136 31075 27140
rect 30828 27113 30942 27136
tri 30828 27081 30860 27113 ne
rect 30860 27090 30942 27113
rect 30988 27113 31075 27136
tri 31075 27113 31102 27140 sw
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27090 31102 27113
rect 30860 27081 31102 27090
tri 30860 27068 30873 27081 ne
rect 30873 27068 31102 27081
tri 31102 27068 31147 27113 sw
tri 30873 27036 30905 27068 ne
rect 30905 27058 31147 27068
tri 31147 27058 31157 27068 sw
rect 70802 27060 71000 27118
rect 30905 27036 31157 27058
tri 30905 27011 30930 27036 ne
rect 30930 27026 31157 27036
tri 31157 27026 31189 27058 sw
rect 30930 27013 31189 27026
tri 31189 27013 31202 27026 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 30930 27011 31202 27013
tri 31202 27011 31204 27013 sw
tri 30930 26966 30975 27011 ne
rect 30975 27004 31204 27011
rect 30975 26966 31074 27004
tri 30975 26949 30992 26966 ne
rect 30992 26958 31074 26966
rect 31120 26981 31204 27004
tri 31204 26981 31234 27011 sw
rect 31120 26958 31234 26981
rect 30992 26949 31234 26958
tri 30992 26936 31005 26949 ne
rect 31005 26936 31234 26949
tri 31234 26936 31279 26981 sw
rect 70802 26956 71000 27014
tri 31005 26904 31037 26936 ne
rect 31037 26926 31279 26936
tri 31279 26926 31289 26936 sw
rect 31037 26904 31289 26926
tri 31037 26894 31047 26904 ne
rect 31047 26894 31289 26904
tri 31289 26894 31321 26926 sw
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31047 26866 31075 26894 ne
rect 31075 26881 31321 26894
tri 31321 26881 31334 26894 sw
rect 31075 26872 31334 26881
rect 31075 26866 31206 26872
tri 31075 26821 31120 26866 ne
rect 31120 26826 31206 26866
rect 31252 26866 31334 26872
tri 31334 26866 31349 26881 sw
rect 31252 26826 31349 26866
rect 31120 26821 31349 26826
tri 31349 26821 31395 26866 sw
rect 70802 26852 71000 26910
tri 31120 26817 31124 26821 ne
rect 31124 26817 31395 26821
tri 31124 26804 31137 26817 ne
rect 31137 26804 31395 26817
tri 31395 26804 31411 26821 sw
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
tri 31137 26772 31169 26804 ne
rect 31169 26794 31411 26804
tri 31411 26794 31421 26804 sw
rect 31169 26772 31421 26794
tri 31169 26737 31204 26772 ne
rect 31204 26762 31421 26772
tri 31421 26762 31453 26794 sw
rect 31204 26749 31453 26762
tri 31453 26749 31466 26762 sw
rect 31204 26740 31466 26749
rect 31204 26737 31338 26740
tri 31204 26691 31249 26737 ne
rect 31249 26694 31338 26737
rect 31384 26737 31466 26740
tri 31466 26737 31479 26749 sw
rect 70802 26748 71000 26806
rect 31384 26717 31479 26737
tri 31479 26717 31498 26737 sw
rect 31384 26694 31498 26717
rect 31249 26691 31498 26694
tri 31249 26685 31256 26691 ne
rect 31256 26685 31498 26691
tri 31256 26672 31269 26685 ne
rect 31269 26672 31498 26685
tri 31498 26672 31543 26717 sw
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
tri 31269 26640 31301 26672 ne
rect 31301 26662 31543 26672
tri 31543 26662 31553 26672 sw
rect 31301 26640 31553 26662
tri 31301 26630 31311 26640 ne
rect 31311 26630 31553 26640
tri 31553 26630 31585 26662 sw
rect 70802 26644 71000 26702
tri 31311 26585 31356 26630 ne
rect 31356 26617 31585 26630
tri 31585 26617 31598 26630 sw
rect 31356 26608 31598 26617
rect 31356 26585 31470 26608
tri 31356 26553 31388 26585 ne
rect 31388 26562 31470 26585
rect 31516 26585 31598 26608
tri 31598 26585 31630 26617 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26562 31630 26585
rect 31388 26553 31630 26562
tri 31388 26540 31401 26553 ne
rect 31401 26540 31630 26553
tri 31630 26540 31675 26585 sw
rect 70802 26540 71000 26598
tri 31401 26508 31433 26540 ne
rect 31433 26530 31675 26540
tri 31675 26530 31685 26540 sw
rect 31433 26508 31685 26530
tri 31433 26501 31440 26508 ne
rect 31440 26501 31685 26508
tri 31440 26462 31479 26501 ne
rect 31479 26498 31685 26501
tri 31685 26498 31717 26530 sw
rect 31479 26485 31717 26498
tri 31717 26485 31730 26498 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31479 26476 31730 26485
rect 31479 26462 31602 26476
tri 31479 26456 31485 26462 ne
rect 31485 26456 31602 26462
tri 31485 26421 31520 26456 ne
rect 31520 26430 31602 26456
rect 31648 26462 31730 26476
tri 31730 26462 31753 26485 sw
rect 31648 26456 31753 26462
tri 31753 26456 31759 26462 sw
rect 31648 26430 31759 26456
rect 31520 26421 31759 26430
tri 31520 26408 31533 26421 ne
rect 31533 26411 31759 26421
tri 31759 26411 31805 26456 sw
rect 70802 26436 71000 26494
rect 31533 26408 31805 26411
tri 31805 26408 31807 26411 sw
tri 31533 26376 31565 26408 ne
rect 31565 26398 31807 26408
tri 31807 26398 31817 26408 sw
rect 31565 26376 31817 26398
tri 31565 26366 31575 26376 ne
rect 31575 26366 31817 26376
tri 31817 26366 31849 26398 sw
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31575 26321 31620 26366 ne
rect 31620 26353 31849 26366
tri 31849 26353 31862 26366 sw
rect 31620 26344 31862 26353
rect 31620 26321 31734 26344
tri 31620 26289 31652 26321 ne
rect 31652 26298 31734 26321
rect 31780 26321 31862 26344
tri 31862 26321 31894 26353 sw
rect 70802 26332 71000 26390
rect 31780 26298 31894 26321
rect 31652 26289 31894 26298
tri 31652 26276 31665 26289 ne
rect 31665 26276 31894 26289
tri 31894 26276 31939 26321 sw
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31665 26244 31697 26276 ne
rect 31697 26266 31939 26276
tri 31939 26266 31949 26276 sw
rect 31697 26244 31949 26266
tri 31697 26199 31742 26244 ne
rect 31742 26234 31949 26244
tri 31949 26234 31981 26266 sw
rect 31742 26221 31981 26234
tri 31981 26221 31994 26234 sw
rect 70802 26228 71000 26286
rect 31742 26212 31994 26221
rect 31742 26199 31866 26212
tri 31742 26188 31753 26199 ne
rect 31753 26188 31866 26199
tri 31753 26144 31797 26188 ne
rect 31797 26166 31866 26188
rect 31912 26188 31994 26212
tri 31994 26188 32027 26221 sw
rect 31912 26166 32027 26188
rect 31797 26144 32027 26166
tri 32027 26144 32071 26188 sw
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
tri 31797 26136 31805 26144 ne
rect 31805 26136 32071 26144
tri 31805 26102 31839 26136 ne
rect 31839 26134 32071 26136
tri 32071 26134 32081 26144 sw
rect 31839 26102 32081 26134
tri 32081 26102 32113 26134 sw
rect 70802 26124 71000 26182
tri 31839 26091 31850 26102 ne
rect 31850 26091 32113 26102
tri 32113 26091 32124 26102 sw
tri 31850 26046 31895 26091 ne
rect 31895 26080 32124 26091
rect 31895 26046 31998 26080
tri 31895 26025 31916 26046 ne
rect 31916 26034 31998 26046
rect 32044 26046 32124 26080
tri 32124 26046 32169 26091 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26034 32169 26046
rect 31916 26025 32169 26034
tri 31916 26012 31929 26025 ne
rect 31929 26012 32169 26025
tri 32169 26012 32203 26046 sw
rect 70802 26020 71000 26078
tri 31929 25980 31961 26012 ne
rect 31961 26002 32203 26012
tri 32203 26002 32213 26012 sw
rect 31961 25980 32213 26002
tri 31961 25935 32006 25980 ne
rect 32006 25970 32213 25980
tri 32213 25970 32245 26002 sw
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32006 25957 32245 25970
tri 32245 25957 32258 25970 sw
rect 32006 25948 32258 25957
rect 32006 25935 32130 25948
tri 32006 25913 32027 25935 ne
rect 32027 25913 32130 25935
tri 32027 25893 32048 25913 ne
rect 32048 25902 32130 25913
rect 32176 25913 32258 25948
tri 32258 25913 32302 25957 sw
rect 70802 25916 71000 25974
rect 32176 25902 32302 25913
rect 32048 25893 32302 25902
tri 32048 25880 32061 25893 ne
rect 32061 25880 32302 25893
tri 32302 25880 32335 25913 sw
tri 32061 25848 32093 25880 ne
rect 32093 25870 32335 25880
tri 32335 25870 32345 25880 sw
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
rect 32093 25848 32345 25870
tri 32093 25838 32103 25848 ne
rect 32103 25838 32345 25848
tri 32345 25838 32377 25870 sw
tri 32103 25793 32148 25838 ne
rect 32148 25825 32377 25838
tri 32377 25825 32390 25838 sw
rect 32148 25816 32390 25825
rect 32148 25793 32262 25816
tri 32148 25771 32169 25793 ne
rect 32169 25771 32262 25793
tri 32169 25748 32193 25771 ne
rect 32193 25770 32262 25771
rect 32308 25793 32390 25816
tri 32390 25793 32422 25825 sw
rect 70802 25812 71000 25870
rect 32308 25770 32422 25793
rect 32193 25748 32422 25770
tri 32422 25748 32467 25793 sw
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
tri 32193 25716 32225 25748 ne
rect 32225 25738 32467 25748
tri 32467 25738 32477 25748 sw
rect 32225 25716 32477 25738
tri 32225 25671 32270 25716 ne
rect 32270 25706 32477 25716
tri 32477 25706 32509 25738 sw
rect 70802 25708 71000 25766
rect 32270 25684 32509 25706
rect 32270 25671 32394 25684
tri 32270 25639 32302 25671 ne
rect 32302 25639 32394 25671
tri 32302 25629 32312 25639 ne
rect 32312 25638 32394 25639
rect 32440 25681 32509 25684
tri 32509 25681 32534 25706 sw
rect 32440 25639 32534 25681
tri 32534 25639 32576 25681 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25638 32576 25639
rect 32312 25629 32576 25638
tri 32312 25616 32325 25629 ne
rect 32325 25616 32576 25629
tri 32576 25616 32599 25639 sw
tri 32325 25584 32357 25616 ne
rect 32357 25606 32599 25616
tri 32599 25606 32609 25616 sw
rect 32357 25584 32609 25606
tri 32357 25574 32367 25584 ne
rect 32367 25574 32609 25584
tri 32609 25574 32641 25606 sw
rect 70802 25604 71000 25662
tri 32367 25529 32412 25574 ne
rect 32412 25561 32641 25574
tri 32641 25561 32654 25574 sw
rect 32412 25552 32654 25561
rect 32412 25529 32526 25552
tri 32412 25497 32444 25529 ne
rect 32444 25506 32526 25529
rect 32572 25529 32654 25552
tri 32654 25529 32686 25561 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32572 25506 32686 25529
rect 32444 25497 32686 25506
tri 32444 25484 32457 25497 ne
rect 32457 25484 32686 25497
tri 32686 25484 32731 25529 sw
rect 70802 25500 71000 25558
tri 32457 25452 32489 25484 ne
rect 32489 25474 32731 25484
tri 32731 25474 32741 25484 sw
rect 32489 25452 32741 25474
tri 32489 25407 32534 25452 ne
rect 32534 25442 32741 25452
tri 32741 25442 32773 25474 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32534 25429 32773 25442
tri 32773 25429 32786 25442 sw
rect 32534 25420 32786 25429
rect 32534 25407 32658 25420
tri 32534 25365 32576 25407 ne
rect 32576 25374 32658 25407
rect 32704 25410 32786 25420
tri 32786 25410 32805 25429 sw
rect 32704 25374 32805 25410
rect 32576 25365 32805 25374
tri 32805 25365 32851 25410 sw
rect 70802 25396 71000 25454
tri 32576 25352 32589 25365 ne
rect 32589 25361 32851 25365
tri 32851 25361 32854 25365 sw
rect 32589 25352 32854 25361
tri 32854 25352 32863 25361 sw
tri 32589 25320 32621 25352 ne
rect 32621 25342 32863 25352
tri 32863 25342 32873 25352 sw
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 32621 25320 32873 25342
tri 32621 25310 32631 25320 ne
rect 32631 25310 32873 25320
tri 32873 25310 32905 25342 sw
tri 32631 25265 32676 25310 ne
rect 32676 25297 32905 25310
tri 32905 25297 32918 25310 sw
rect 32676 25288 32918 25297
rect 32676 25265 32790 25288
tri 32676 25233 32708 25265 ne
rect 32708 25242 32790 25265
rect 32836 25265 32918 25288
tri 32918 25265 32950 25297 sw
rect 70802 25292 71000 25350
rect 32836 25242 32950 25265
rect 32708 25233 32950 25242
tri 32708 25220 32721 25233 ne
rect 32721 25220 32950 25233
tri 32950 25220 32995 25265 sw
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
tri 32721 25188 32753 25220 ne
rect 32753 25210 32995 25220
tri 32995 25210 33005 25220 sw
rect 32753 25188 33005 25210
tri 32753 25143 32798 25188 ne
rect 32798 25178 33005 25188
tri 33005 25178 33037 25210 sw
rect 70802 25188 71000 25246
rect 32798 25165 33037 25178
tri 33037 25165 33050 25178 sw
rect 32798 25156 33050 25165
rect 32798 25143 32922 25156
tri 32798 25101 32840 25143 ne
rect 32840 25110 32922 25143
rect 32968 25135 33050 25156
tri 33050 25135 33080 25165 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25110 33080 25135
rect 32840 25101 33080 25110
tri 32840 25090 32851 25101 ne
rect 32851 25090 33080 25101
tri 33080 25090 33125 25135 sw
tri 32851 25088 32853 25090 ne
rect 32853 25088 33125 25090
tri 33125 25088 33127 25090 sw
tri 32853 25056 32885 25088 ne
rect 32885 25078 33127 25088
tri 33127 25078 33137 25088 sw
rect 70802 25084 71000 25142
rect 32885 25056 33137 25078
tri 32885 25046 32895 25056 ne
rect 32895 25046 33137 25056
tri 33137 25046 33169 25078 sw
tri 32895 25042 32899 25046 ne
rect 32899 25042 33169 25046
tri 32899 24997 32944 25042 ne
rect 32944 25033 33169 25042
tri 33169 25033 33182 25046 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 32944 25024 33182 25033
rect 32944 24997 33054 25024
tri 32944 24969 32972 24997 ne
rect 32972 24978 33054 24997
rect 33100 24997 33182 25024
tri 33182 24997 33219 25033 sw
rect 33100 24978 33219 24997
rect 32972 24969 33219 24978
tri 32972 24956 32985 24969 ne
rect 32985 24956 33219 24969
tri 33219 24956 33259 24997 sw
rect 70802 24980 71000 25038
tri 32985 24924 33017 24956 ne
rect 33017 24951 33259 24956
tri 33259 24951 33264 24956 sw
rect 33017 24946 33264 24951
tri 33264 24946 33269 24951 sw
rect 33017 24924 33269 24946
tri 33017 24879 33062 24924 ne
rect 33062 24914 33269 24924
tri 33269 24914 33301 24946 sw
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
rect 33062 24901 33301 24914
tri 33301 24901 33314 24914 sw
rect 33062 24892 33314 24901
rect 33062 24879 33186 24892
tri 33062 24837 33104 24879 ne
rect 33104 24846 33186 24879
rect 33232 24869 33314 24892
tri 33314 24869 33346 24901 sw
rect 70802 24876 71000 24934
rect 33232 24846 33346 24869
rect 33104 24837 33346 24846
tri 33104 24816 33125 24837 ne
rect 33125 24824 33346 24837
tri 33346 24824 33391 24869 sw
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33125 24816 33391 24824
tri 33391 24816 33399 24824 sw
tri 33125 24792 33149 24816 ne
rect 33149 24814 33399 24816
tri 33399 24814 33401 24816 sw
rect 33149 24792 33401 24814
tri 33149 24782 33159 24792 ne
rect 33159 24782 33401 24792
tri 33401 24782 33433 24814 sw
tri 33159 24737 33204 24782 ne
rect 33204 24769 33433 24782
tri 33433 24769 33446 24782 sw
rect 70802 24772 71000 24830
rect 33204 24760 33446 24769
rect 33204 24737 33318 24760
tri 33204 24692 33249 24737 ne
rect 33249 24714 33318 24737
rect 33364 24737 33446 24760
tri 33446 24737 33478 24769 sw
rect 33364 24714 33478 24737
rect 33249 24692 33478 24714
tri 33478 24692 33523 24737 sw
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
tri 33249 24677 33264 24692 ne
rect 33264 24682 33523 24692
tri 33523 24682 33533 24692 sw
rect 33264 24677 33533 24682
tri 33264 24632 33309 24677 ne
rect 33309 24650 33533 24677
tri 33533 24650 33565 24682 sw
rect 70802 24668 71000 24726
rect 33309 24637 33565 24650
tri 33565 24637 33578 24650 sw
rect 33309 24632 33578 24637
tri 33578 24632 33583 24637 sw
tri 33309 24587 33354 24632 ne
rect 33354 24628 33583 24632
rect 33354 24587 33450 24628
tri 33354 24573 33368 24587 ne
rect 33368 24582 33450 24587
rect 33496 24587 33583 24628
tri 33583 24587 33629 24632 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33629 24587
rect 33368 24573 33629 24582
tri 33368 24541 33399 24573 ne
rect 33399 24560 33629 24573
tri 33629 24560 33655 24587 sw
rect 70802 24564 71000 24622
rect 33399 24550 33655 24560
tri 33655 24550 33665 24560 sw
rect 33399 24541 33665 24550
tri 33665 24541 33674 24550 sw
tri 33399 24528 33413 24541 ne
rect 33413 24528 33674 24541
tri 33413 24518 33423 24528 ne
rect 33423 24518 33674 24528
tri 33674 24518 33697 24541 sw
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33423 24473 33468 24518 ne
rect 33468 24505 33697 24518
tri 33697 24505 33710 24518 sw
rect 33468 24496 33710 24505
rect 33468 24473 33582 24496
tri 33468 24441 33500 24473 ne
rect 33500 24450 33582 24473
rect 33628 24473 33710 24496
tri 33710 24473 33742 24505 sw
rect 33628 24450 33742 24473
rect 33500 24441 33742 24450
tri 33500 24428 33513 24441 ne
rect 33513 24428 33742 24441
tri 33742 24428 33787 24473 sw
rect 70802 24460 71000 24518
tri 33513 24396 33545 24428 ne
rect 33545 24418 33787 24428
tri 33787 24418 33797 24428 sw
rect 33545 24396 33797 24418
tri 33545 24351 33590 24396 ne
rect 33590 24386 33797 24396
tri 33797 24386 33829 24418 sw
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
rect 33590 24373 33829 24386
tri 33829 24373 33842 24386 sw
rect 33590 24364 33842 24373
rect 33590 24351 33714 24364
tri 33590 24312 33629 24351 ne
rect 33629 24318 33714 24351
rect 33760 24341 33842 24364
tri 33842 24341 33874 24373 sw
rect 70802 24356 71000 24414
rect 33760 24318 33874 24341
rect 33629 24312 33874 24318
tri 33629 24267 33674 24312 ne
rect 33674 24296 33874 24312
tri 33874 24296 33919 24341 sw
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 33674 24286 33919 24296
tri 33919 24286 33929 24296 sw
rect 33674 24267 33929 24286
tri 33929 24267 33948 24286 sw
tri 33674 24264 33677 24267 ne
rect 33677 24264 33948 24267
tri 33677 24254 33687 24264 ne
rect 33687 24254 33948 24264
tri 33948 24254 33961 24267 sw
tri 33687 24209 33732 24254 ne
rect 33732 24232 33961 24254
rect 33732 24209 33846 24232
tri 33732 24177 33764 24209 ne
rect 33764 24186 33846 24209
rect 33892 24222 33961 24232
tri 33961 24222 33993 24254 sw
rect 70802 24252 71000 24310
rect 33892 24209 33993 24222
tri 33993 24209 34006 24222 sw
rect 33892 24186 34006 24209
rect 33764 24177 34006 24186
tri 33764 24164 33777 24177 ne
rect 33777 24164 34006 24177
tri 34006 24164 34051 24209 sw
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
tri 33777 24132 33809 24164 ne
rect 33809 24154 34051 24164
tri 34051 24154 34061 24164 sw
rect 33809 24132 34061 24154
tri 33809 24087 33854 24132 ne
rect 33854 24122 34061 24132
tri 34061 24122 34093 24154 sw
rect 70802 24148 71000 24206
rect 33854 24109 34093 24122
tri 34093 24109 34106 24122 sw
rect 33854 24100 34106 24109
rect 33854 24087 33978 24100
tri 33854 24045 33896 24087 ne
rect 33896 24054 33978 24087
rect 34024 24077 34106 24100
tri 34106 24077 34138 24109 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 34024 24054 34138 24077
rect 33896 24045 34138 24054
tri 33896 24000 33941 24045 ne
rect 33941 24032 34138 24045
tri 34138 24032 34183 24077 sw
rect 70802 24044 71000 24102
rect 33941 24022 34183 24032
tri 34183 24022 34193 24032 sw
rect 33941 24000 34193 24022
tri 33941 23993 33948 24000 ne
rect 33948 23993 34193 24000
tri 34193 23993 34223 24022 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33948 23990 33951 23993 ne
rect 33951 23990 34223 23993
tri 34223 23990 34225 23993 sw
tri 33951 23947 33993 23990 ne
rect 33993 23977 34225 23990
tri 34225 23977 34238 23990 sw
rect 33993 23968 34238 23977
rect 33993 23947 34110 23968
tri 33993 23902 34039 23947 ne
rect 34039 23922 34110 23947
rect 34156 23947 34238 23968
tri 34238 23947 34268 23977 sw
rect 34156 23922 34268 23947
rect 34039 23902 34268 23922
tri 34268 23902 34313 23947 sw
rect 70802 23940 71000 23998
tri 34039 23900 34041 23902 ne
rect 34041 23900 34313 23902
tri 34313 23900 34315 23902 sw
tri 34041 23868 34073 23900 ne
rect 34073 23868 34315 23900
tri 34073 23858 34083 23868 ne
rect 34083 23858 34315 23868
tri 34315 23858 34357 23900 sw
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34083 23813 34128 23858 ne
rect 34128 23845 34357 23858
tri 34357 23845 34370 23858 sw
rect 34128 23836 34370 23845
rect 34128 23813 34242 23836
tri 34128 23781 34160 23813 ne
rect 34160 23790 34242 23813
rect 34288 23813 34370 23836
tri 34370 23813 34402 23845 sw
rect 70802 23836 71000 23894
rect 34288 23790 34402 23813
rect 34160 23781 34402 23790
tri 34160 23768 34173 23781 ne
rect 34173 23768 34402 23781
tri 34402 23768 34447 23813 sw
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34173 23736 34205 23768 ne
rect 34205 23758 34447 23768
tri 34447 23758 34457 23768 sw
rect 34205 23736 34457 23758
tri 34205 23718 34223 23736 ne
rect 34223 23726 34457 23736
tri 34457 23726 34489 23758 sw
rect 70802 23732 71000 23790
rect 34223 23718 34489 23726
tri 34489 23718 34497 23726 sw
tri 34223 23673 34268 23718 ne
rect 34268 23713 34497 23718
tri 34497 23713 34502 23718 sw
rect 34268 23704 34502 23713
rect 34268 23673 34374 23704
tri 34268 23649 34292 23673 ne
rect 34292 23658 34374 23673
rect 34420 23681 34502 23704
tri 34502 23681 34534 23713 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34534 23681
rect 34292 23649 34534 23658
tri 34292 23636 34305 23649 ne
rect 34305 23636 34534 23649
tri 34534 23636 34579 23681 sw
tri 34305 23604 34337 23636 ne
rect 34337 23626 34579 23636
tri 34579 23626 34589 23636 sw
rect 70802 23628 71000 23686
rect 34337 23604 34589 23626
tri 34337 23594 34347 23604 ne
rect 34347 23594 34589 23604
tri 34589 23594 34621 23626 sw
tri 34347 23583 34358 23594 ne
rect 34358 23583 34621 23594
tri 34358 23537 34403 23583 ne
rect 34403 23581 34621 23583
tri 34621 23581 34634 23594 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34403 23572 34634 23581
rect 34403 23537 34506 23572
tri 34403 23517 34424 23537 ne
rect 34424 23526 34506 23537
rect 34552 23537 34634 23572
tri 34634 23537 34678 23581 sw
rect 34552 23526 34678 23537
rect 34424 23517 34678 23526
tri 34424 23504 34437 23517 ne
rect 34437 23504 34678 23517
tri 34678 23504 34711 23537 sw
rect 70802 23524 71000 23582
tri 34437 23472 34469 23504 ne
rect 34469 23494 34711 23504
tri 34711 23494 34721 23504 sw
rect 34469 23472 34721 23494
tri 34469 23444 34497 23472 ne
rect 34497 23462 34721 23472
tri 34721 23462 34753 23494 sw
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34497 23449 34753 23462
tri 34753 23449 34766 23462 sw
rect 34497 23444 34766 23449
tri 34766 23444 34771 23449 sw
tri 34497 23399 34542 23444 ne
rect 34542 23440 34771 23444
rect 34542 23399 34638 23440
tri 34542 23385 34556 23399 ne
rect 34556 23394 34638 23399
rect 34684 23417 34771 23440
tri 34771 23417 34798 23444 sw
rect 70802 23420 71000 23478
rect 34684 23394 34798 23417
rect 34556 23385 34798 23394
tri 34556 23372 34569 23385 ne
rect 34569 23372 34798 23385
tri 34798 23372 34843 23417 sw
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34569 23340 34601 23372 ne
rect 34601 23362 34843 23372
tri 34843 23362 34853 23372 sw
rect 34601 23340 34853 23362
tri 34601 23330 34611 23340 ne
rect 34611 23330 34853 23340
tri 34853 23330 34885 23362 sw
tri 34611 23285 34656 23330 ne
rect 34656 23317 34885 23330
tri 34885 23317 34898 23330 sw
rect 34656 23308 34898 23317
rect 34656 23285 34770 23308
tri 34656 23253 34688 23285 ne
rect 34688 23262 34770 23285
rect 34816 23285 34898 23308
tri 34898 23285 34930 23317 sw
rect 70802 23316 71000 23374
rect 34816 23262 34930 23285
rect 34688 23253 34930 23262
tri 34688 23240 34701 23253 ne
rect 34701 23240 34930 23253
tri 34930 23240 34975 23285 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
tri 34701 23208 34733 23240 ne
rect 34733 23230 34975 23240
tri 34975 23230 34985 23240 sw
rect 34733 23208 34985 23230
tri 34733 23173 34768 23208 ne
rect 34768 23198 34985 23208
tri 34985 23198 35017 23230 sw
rect 70802 23212 71000 23270
rect 34768 23185 35017 23198
tri 35017 23185 35030 23198 sw
rect 34768 23176 35030 23185
rect 34768 23173 34902 23176
tri 34768 23169 34771 23173 ne
rect 34771 23169 34902 23173
tri 34771 23124 34817 23169 ne
rect 34817 23130 34902 23169
rect 34948 23173 35030 23176
tri 35030 23173 35043 23185 sw
rect 34948 23169 35043 23173
tri 35043 23169 35046 23173 sw
rect 34948 23130 35046 23169
rect 34817 23127 35046 23130
tri 35046 23127 35088 23169 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34817 23124 35088 23127
tri 34817 23121 34820 23124 ne
rect 34820 23121 35088 23124
tri 34820 23108 34833 23121 ne
rect 34833 23108 35088 23121
tri 35088 23108 35107 23127 sw
rect 70802 23108 71000 23166
tri 34833 23076 34865 23108 ne
rect 34865 23098 35107 23108
tri 35107 23098 35117 23108 sw
rect 34865 23076 35117 23098
tri 34865 23066 34875 23076 ne
rect 34875 23066 35117 23076
tri 35117 23066 35149 23098 sw
tri 34875 23021 34920 23066 ne
rect 34920 23053 35149 23066
tri 35149 23053 35162 23066 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 34920 23044 35162 23053
rect 34920 23021 35034 23044
tri 34920 22989 34952 23021 ne
rect 34952 22998 35034 23021
rect 35080 23021 35162 23044
tri 35162 23021 35194 23053 sw
rect 35080 22998 35194 23021
rect 34952 22989 35194 22998
tri 34952 22976 34965 22989 ne
rect 34965 22976 35194 22989
tri 35194 22976 35239 23021 sw
rect 70802 23004 71000 23062
tri 34965 22944 34997 22976 ne
rect 34997 22966 35239 22976
tri 35239 22966 35249 22976 sw
rect 34997 22944 35249 22966
tri 34997 22899 35042 22944 ne
rect 35042 22934 35249 22944
tri 35249 22934 35281 22966 sw
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
rect 35042 22921 35281 22934
tri 35281 22921 35294 22934 sw
rect 35042 22912 35294 22921
rect 35042 22899 35166 22912
tri 35042 22895 35046 22899 ne
rect 35046 22895 35166 22899
tri 35046 22853 35088 22895 ne
rect 35088 22866 35166 22895
rect 35212 22895 35294 22912
tri 35294 22895 35320 22921 sw
rect 70802 22900 71000 22958
rect 35212 22889 35320 22895
tri 35320 22889 35326 22895 sw
rect 35212 22866 35326 22889
rect 35088 22853 35326 22866
tri 35088 22844 35097 22853 ne
rect 35097 22844 35326 22853
tri 35326 22844 35371 22889 sw
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35097 22808 35133 22844 ne
rect 35133 22834 35371 22844
tri 35371 22834 35381 22844 sw
rect 35133 22808 35381 22834
tri 35133 22802 35139 22808 ne
rect 35139 22802 35381 22808
tri 35381 22802 35413 22834 sw
tri 35139 22757 35184 22802 ne
rect 35184 22780 35413 22802
rect 35184 22757 35298 22780
tri 35184 22725 35216 22757 ne
rect 35216 22734 35298 22757
rect 35344 22763 35413 22780
tri 35413 22763 35453 22802 sw
rect 70802 22796 71000 22854
rect 35344 22757 35453 22763
tri 35453 22757 35458 22763 sw
rect 35344 22734 35458 22757
rect 35216 22725 35458 22734
tri 35216 22712 35229 22725 ne
rect 35229 22712 35458 22725
tri 35458 22712 35503 22757 sw
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
tri 35229 22680 35261 22712 ne
rect 35261 22702 35503 22712
tri 35503 22702 35513 22712 sw
rect 35261 22680 35513 22702
tri 35261 22635 35306 22680 ne
rect 35306 22670 35513 22680
tri 35513 22670 35545 22702 sw
rect 70802 22692 71000 22750
rect 35306 22657 35545 22670
tri 35545 22657 35558 22670 sw
rect 35306 22648 35558 22657
rect 35306 22635 35430 22648
tri 35306 22621 35320 22635 ne
rect 35320 22621 35430 22635
tri 35320 22593 35348 22621 ne
rect 35348 22602 35430 22621
rect 35476 22621 35558 22648
tri 35558 22621 35595 22657 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22602 35595 22621
rect 35348 22593 35595 22602
tri 35348 22580 35361 22593 ne
rect 35361 22580 35595 22593
tri 35595 22580 35635 22621 sw
rect 70802 22588 71000 22646
tri 35361 22548 35393 22580 ne
rect 35393 22570 35635 22580
tri 35635 22570 35645 22580 sw
rect 35393 22548 35645 22570
tri 35393 22538 35403 22548 ne
rect 35403 22538 35645 22548
tri 35645 22538 35677 22570 sw
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35403 22493 35448 22538 ne
rect 35448 22525 35677 22538
tri 35677 22525 35690 22538 sw
rect 35448 22516 35690 22525
rect 35448 22493 35562 22516
tri 35448 22488 35453 22493 ne
rect 35453 22488 35562 22493
tri 35453 22448 35493 22488 ne
rect 35493 22470 35562 22488
rect 35608 22493 35690 22516
tri 35690 22493 35722 22525 sw
rect 35608 22470 35722 22493
rect 35493 22448 35722 22470
tri 35722 22448 35767 22493 sw
rect 70802 22484 71000 22542
tri 35493 22416 35525 22448 ne
rect 35525 22443 35767 22448
tri 35767 22443 35772 22448 sw
rect 35525 22416 35772 22443
tri 35525 22371 35570 22416 ne
rect 35570 22406 35772 22416
tri 35772 22406 35809 22443 sw
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
rect 35570 22393 35809 22406
tri 35809 22393 35822 22406 sw
rect 35570 22391 35822 22393
tri 35822 22391 35824 22393 sw
rect 35570 22384 35824 22391
rect 35570 22371 35694 22384
tri 35570 22346 35595 22371 ne
rect 35595 22346 35694 22371
tri 35595 22329 35612 22346 ne
rect 35612 22338 35694 22346
rect 35740 22346 35824 22384
tri 35824 22346 35869 22391 sw
rect 70802 22380 71000 22438
rect 35740 22338 35869 22346
rect 35612 22329 35869 22338
tri 35612 22316 35625 22329 ne
rect 35625 22316 35869 22329
tri 35869 22316 35899 22346 sw
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35625 22284 35657 22316 ne
rect 35657 22306 35899 22316
tri 35899 22306 35909 22316 sw
rect 35657 22284 35909 22306
tri 35657 22274 35667 22284 ne
rect 35667 22274 35909 22284
tri 35909 22274 35941 22306 sw
rect 70802 22276 71000 22334
tri 35667 22229 35712 22274 ne
rect 35712 22261 35941 22274
tri 35941 22261 35954 22274 sw
rect 35712 22252 35954 22261
rect 35712 22229 35826 22252
tri 35712 22197 35744 22229 ne
rect 35744 22206 35826 22229
rect 35872 22229 35954 22252
tri 35954 22229 35986 22261 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 35986 22229
rect 35744 22197 35986 22206
tri 35744 22184 35757 22197 ne
rect 35757 22184 35986 22197
tri 35986 22184 36031 22229 sw
tri 35757 22152 35789 22184 ne
rect 35789 22174 36031 22184
tri 36031 22174 36041 22184 sw
rect 35789 22152 36041 22174
tri 35789 22123 35817 22152 ne
rect 35817 22142 36041 22152
tri 36041 22142 36073 22174 sw
rect 70802 22172 71000 22230
rect 35817 22129 36073 22142
tri 36073 22129 36086 22142 sw
rect 35817 22123 36086 22129
tri 36086 22123 36092 22129 sw
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
tri 35817 22078 35863 22123 ne
rect 35863 22120 36092 22123
rect 35863 22078 35958 22120
tri 35863 22072 35869 22078 ne
rect 35869 22074 35958 22078
rect 36004 22078 36092 22120
tri 36092 22078 36137 22123 sw
rect 36004 22074 36137 22078
rect 35869 22072 36137 22074
tri 36137 22072 36143 22078 sw
tri 35869 22065 35876 22072 ne
rect 35876 22065 36143 22072
tri 35876 22052 35889 22065 ne
rect 35889 22052 36143 22065
tri 36143 22052 36163 22072 sw
rect 70802 22068 71000 22126
tri 35889 22020 35921 22052 ne
rect 35921 22042 36163 22052
tri 36163 22042 36173 22052 sw
rect 35921 22020 36173 22042
tri 35921 22010 35931 22020 ne
rect 35931 22010 36173 22020
tri 36173 22010 36205 22042 sw
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35931 21965 35976 22010 ne
rect 35976 21997 36205 22010
tri 36205 21997 36218 22010 sw
rect 35976 21988 36218 21997
rect 35976 21965 36090 21988
tri 35976 21933 36008 21965 ne
rect 36008 21942 36090 21965
rect 36136 21965 36218 21988
tri 36218 21965 36250 21997 sw
rect 36136 21942 36250 21965
rect 36008 21933 36250 21942
tri 36008 21920 36021 21933 ne
rect 36021 21920 36250 21933
tri 36250 21920 36295 21965 sw
rect 70802 21964 71000 22022
tri 36021 21888 36053 21920 ne
rect 36053 21910 36295 21920
tri 36295 21910 36305 21920 sw
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36053 21888 36305 21910
tri 36053 21843 36098 21888 ne
rect 36098 21878 36305 21888
tri 36305 21878 36337 21910 sw
rect 36098 21865 36337 21878
tri 36337 21865 36350 21878 sw
rect 36098 21856 36350 21865
rect 36098 21843 36222 21856
tri 36098 21801 36140 21843 ne
rect 36140 21810 36222 21843
rect 36268 21843 36350 21856
tri 36350 21843 36373 21865 sw
rect 70802 21860 71000 21918
rect 36268 21810 36373 21843
rect 36140 21801 36373 21810
tri 36140 21797 36143 21801 ne
rect 36143 21797 36373 21801
tri 36373 21797 36418 21843 sw
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
tri 36143 21788 36153 21797 ne
rect 36153 21788 36418 21797
tri 36418 21788 36427 21797 sw
tri 36153 21756 36185 21788 ne
rect 36185 21778 36427 21788
tri 36427 21778 36437 21788 sw
rect 36185 21756 36437 21778
tri 36185 21746 36195 21756 ne
rect 36195 21746 36437 21756
tri 36437 21746 36469 21778 sw
rect 70802 21756 71000 21814
tri 36195 21713 36227 21746 ne
rect 36227 21733 36469 21746
tri 36469 21733 36482 21746 sw
rect 36227 21724 36482 21733
rect 36227 21713 36354 21724
tri 36227 21669 36272 21713 ne
rect 36272 21678 36354 21713
rect 36400 21713 36482 21724
tri 36482 21713 36502 21733 sw
rect 36400 21678 36502 21713
rect 36272 21669 36502 21678
tri 36272 21656 36285 21669 ne
rect 36285 21668 36502 21669
tri 36502 21668 36547 21713 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36285 21656 36547 21668
tri 36547 21656 36559 21668 sw
tri 36285 21624 36317 21656 ne
rect 36317 21646 36559 21656
tri 36559 21646 36569 21656 sw
rect 70802 21652 71000 21710
rect 36317 21624 36569 21646
tri 36317 21579 36362 21624 ne
rect 36362 21614 36569 21624
tri 36569 21614 36601 21646 sw
rect 36362 21601 36601 21614
tri 36601 21601 36614 21614 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36362 21592 36614 21601
rect 36362 21579 36486 21592
tri 36362 21537 36404 21579 ne
rect 36404 21546 36486 21579
rect 36532 21569 36614 21592
tri 36614 21569 36646 21601 sw
rect 36532 21546 36646 21569
rect 36404 21537 36646 21546
tri 36404 21523 36418 21537 ne
rect 36418 21524 36646 21537
tri 36646 21524 36691 21569 sw
rect 70802 21548 71000 21606
rect 36418 21523 36691 21524
tri 36691 21523 36692 21524 sw
tri 36418 21492 36449 21523 ne
rect 36449 21514 36692 21523
tri 36692 21514 36701 21523 sw
rect 36449 21492 36701 21514
tri 36449 21482 36459 21492 ne
rect 36459 21482 36701 21492
tri 36701 21482 36733 21514 sw
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36459 21437 36504 21482 ne
rect 36504 21469 36733 21482
tri 36733 21469 36746 21482 sw
rect 36504 21460 36746 21469
rect 36504 21437 36618 21460
tri 36504 21394 36547 21437 ne
rect 36547 21414 36618 21437
rect 36664 21437 36746 21460
tri 36746 21437 36778 21469 sw
rect 70802 21444 71000 21502
rect 36664 21414 36778 21437
rect 36547 21394 36778 21414
tri 36547 21392 36549 21394 ne
rect 36549 21392 36778 21394
tri 36778 21392 36823 21437 sw
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36549 21349 36592 21392 ne
rect 36592 21382 36823 21392
tri 36823 21382 36833 21392 sw
rect 36592 21350 36833 21382
tri 36833 21350 36865 21382 sw
rect 36592 21349 36865 21350
tri 36865 21349 36867 21350 sw
tri 36592 21303 36637 21349 ne
rect 36637 21328 36867 21349
rect 36637 21303 36750 21328
tri 36637 21273 36668 21303 ne
rect 36668 21282 36750 21303
rect 36796 21303 36867 21328
tri 36867 21303 36912 21349 sw
rect 70802 21340 71000 21398
rect 36796 21282 36912 21303
rect 36668 21273 36912 21282
tri 36668 21249 36692 21273 ne
rect 36692 21260 36912 21273
tri 36912 21260 36955 21303 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36692 21250 36955 21260
tri 36955 21250 36965 21260 sw
rect 36692 21249 36965 21250
tri 36965 21249 36967 21250 sw
tri 36692 21228 36713 21249 ne
rect 36713 21228 36967 21249
tri 36713 21218 36723 21228 ne
rect 36723 21218 36967 21228
tri 36967 21218 36997 21249 sw
rect 70802 21236 71000 21294
tri 36723 21173 36768 21218 ne
rect 36768 21205 36997 21218
tri 36997 21205 37010 21218 sw
rect 36768 21196 37010 21205
rect 36768 21173 36882 21196
tri 36768 21141 36800 21173 ne
rect 36800 21150 36882 21173
rect 36928 21173 37010 21196
tri 37010 21173 37042 21205 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21150 37042 21173
rect 36800 21141 37042 21150
tri 36800 21128 36813 21141 ne
rect 36813 21128 37042 21141
tri 37042 21128 37087 21173 sw
rect 70802 21132 71000 21190
tri 36813 21096 36845 21128 ne
rect 36845 21118 37087 21128
tri 37087 21118 37097 21128 sw
rect 36845 21096 37097 21118
tri 36845 21051 36890 21096 ne
rect 36890 21086 37097 21096
tri 37097 21086 37129 21118 sw
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 36890 21073 37129 21086
tri 37129 21073 37142 21086 sw
rect 36890 21064 37142 21073
rect 36890 21051 37014 21064
tri 36890 21029 36912 21051 ne
rect 36912 21029 37014 21051
tri 36912 20984 36957 21029 ne
rect 36957 21018 37014 21029
rect 37060 21041 37142 21064
tri 37142 21041 37174 21073 sw
rect 37060 21018 37174 21041
rect 36957 20996 37174 21018
tri 37174 20996 37219 21041 sw
rect 70802 21028 71000 21086
rect 36957 20986 37219 20996
tri 37219 20986 37229 20996 sw
rect 36957 20984 37229 20986
tri 36957 20974 36967 20984 ne
rect 36967 20974 37229 20984
tri 37229 20974 37241 20986 sw
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 36967 20964 36977 20974 ne
rect 36977 20964 37241 20974
tri 36977 20954 36987 20964 ne
rect 36987 20954 37241 20964
tri 37241 20954 37261 20974 sw
tri 36987 20909 37032 20954 ne
rect 37032 20939 37261 20954
tri 37261 20939 37277 20954 sw
rect 37032 20932 37277 20939
rect 37032 20909 37146 20932
tri 37032 20877 37064 20909 ne
rect 37064 20886 37146 20909
rect 37192 20909 37277 20932
tri 37277 20909 37306 20939 sw
rect 70802 20924 71000 20982
rect 37192 20886 37306 20909
rect 37064 20877 37306 20886
tri 37064 20864 37077 20877 ne
rect 37077 20864 37306 20877
tri 37306 20864 37351 20909 sw
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
tri 37077 20832 37109 20864 ne
rect 37109 20854 37351 20864
tri 37351 20854 37361 20864 sw
rect 37109 20832 37361 20854
tri 37109 20787 37154 20832 ne
rect 37154 20822 37361 20832
tri 37361 20822 37393 20854 sw
rect 37154 20809 37393 20822
tri 37393 20809 37406 20822 sw
rect 70802 20820 71000 20878
rect 37154 20800 37406 20809
rect 37154 20787 37278 20800
tri 37154 20745 37196 20787 ne
rect 37196 20754 37278 20787
rect 37324 20777 37406 20800
tri 37406 20777 37438 20809 sw
rect 37324 20754 37438 20777
rect 37196 20745 37438 20754
tri 37196 20700 37241 20745 ne
rect 37241 20732 37438 20745
tri 37438 20732 37483 20777 sw
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 37241 20722 37483 20732
tri 37483 20722 37493 20732 sw
rect 37241 20700 37493 20722
tri 37493 20700 37515 20722 sw
rect 70802 20716 71000 20774
tri 37241 20690 37251 20700 ne
rect 37251 20690 37515 20700
tri 37515 20690 37525 20700 sw
tri 37251 20664 37277 20690 ne
rect 37277 20677 37525 20690
tri 37525 20677 37538 20690 sw
rect 37277 20668 37538 20677
rect 37277 20664 37410 20668
tri 37277 20619 37322 20664 ne
rect 37322 20622 37410 20664
rect 37456 20664 37538 20668
tri 37538 20664 37551 20677 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37456 20622 37551 20664
rect 37322 20619 37551 20622
tri 37551 20619 37596 20664 sw
tri 37322 20613 37328 20619 ne
rect 37328 20613 37596 20619
tri 37328 20600 37341 20613 ne
rect 37341 20600 37596 20613
tri 37596 20600 37615 20619 sw
rect 70802 20612 71000 20670
tri 37341 20568 37373 20600 ne
rect 37373 20590 37615 20600
tri 37615 20590 37625 20600 sw
rect 37373 20568 37625 20590
tri 37373 20523 37418 20568 ne
rect 37418 20558 37625 20568
tri 37625 20558 37657 20590 sw
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37418 20545 37657 20558
tri 37657 20545 37670 20558 sw
rect 37418 20536 37670 20545
rect 37418 20523 37542 20536
tri 37418 20481 37460 20523 ne
rect 37460 20490 37542 20523
rect 37588 20513 37670 20536
tri 37670 20513 37702 20545 sw
rect 37588 20490 37702 20513
rect 37460 20481 37702 20490
tri 37460 20436 37505 20481 ne
rect 37505 20468 37702 20481
tri 37702 20468 37747 20513 sw
rect 70802 20508 71000 20566
rect 37505 20458 37747 20468
tri 37747 20458 37757 20468 sw
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 37505 20436 37757 20458
tri 37505 20425 37515 20436 ne
rect 37515 20426 37757 20436
tri 37757 20426 37789 20458 sw
rect 37515 20425 37789 20426
tri 37789 20425 37790 20426 sw
tri 37515 20380 37561 20425 ne
rect 37561 20413 37790 20425
tri 37790 20413 37802 20425 sw
rect 37561 20404 37802 20413
rect 37561 20380 37674 20404
tri 37561 20349 37592 20380 ne
rect 37592 20358 37674 20380
rect 37720 20381 37802 20404
tri 37802 20381 37834 20413 sw
rect 70802 20404 71000 20462
rect 37720 20358 37834 20381
rect 37592 20349 37834 20358
tri 37592 20336 37605 20349 ne
rect 37605 20336 37834 20349
tri 37834 20336 37879 20381 sw
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37605 20304 37637 20336 ne
rect 37637 20326 37879 20336
tri 37879 20326 37889 20336 sw
rect 37637 20304 37889 20326
tri 37637 20299 37641 20304 ne
rect 37641 20299 37889 20304
tri 37641 20294 37647 20299 ne
rect 37647 20294 37889 20299
tri 37889 20294 37921 20326 sw
rect 70802 20300 71000 20358
tri 37647 20254 37687 20294 ne
rect 37687 20281 37921 20294
tri 37921 20281 37934 20294 sw
rect 37687 20272 37934 20281
rect 37687 20254 37806 20272
tri 37687 20217 37724 20254 ne
rect 37724 20226 37806 20254
rect 37852 20254 37934 20272
tri 37934 20254 37961 20281 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37961 20254
rect 37724 20217 37961 20226
tri 37724 20204 37737 20217 ne
rect 37737 20209 37961 20217
tri 37961 20209 38006 20254 sw
rect 37737 20204 38006 20209
tri 38006 20204 38011 20209 sw
tri 37737 20172 37769 20204 ne
rect 37769 20194 38011 20204
tri 38011 20194 38021 20204 sw
rect 70802 20196 71000 20254
rect 37769 20172 38021 20194
tri 37769 20151 37790 20172 ne
rect 37790 20162 38021 20172
tri 38021 20162 38053 20194 sw
rect 37790 20151 38053 20162
tri 38053 20151 38064 20162 sw
tri 37790 20106 37835 20151 ne
rect 37835 20149 38064 20151
tri 38064 20149 38066 20151 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 37835 20140 38066 20149
rect 37835 20106 37938 20140
tri 37835 20085 37856 20106 ne
rect 37856 20094 37938 20106
rect 37984 20117 38066 20140
tri 38066 20117 38098 20149 sw
rect 37984 20094 38098 20117
rect 37856 20085 38098 20094
tri 37856 20072 37869 20085 ne
rect 37869 20072 38098 20085
tri 38098 20072 38143 20117 sw
rect 70802 20092 71000 20150
tri 37869 20040 37901 20072 ne
rect 37901 20062 38143 20072
tri 38143 20062 38153 20072 sw
rect 37901 20040 38153 20062
tri 37901 20030 37911 20040 ne
rect 37911 20030 38153 20040
tri 38153 20030 38185 20062 sw
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37911 19985 37956 20030 ne
rect 37956 20017 38185 20030
tri 38185 20017 38198 20030 sw
rect 37956 20008 38198 20017
rect 37956 19985 38070 20008
tri 37956 19940 38001 19985 ne
rect 38001 19962 38070 19985
rect 38116 19985 38198 20008
tri 38198 19985 38230 20017 sw
rect 70802 19988 71000 20046
rect 38116 19962 38230 19985
rect 38001 19940 38230 19962
tri 38230 19940 38275 19985 sw
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
tri 38001 19935 38006 19940 ne
rect 38006 19935 38275 19940
tri 38006 19889 38051 19935 ne
rect 38051 19930 38275 19935
tri 38275 19930 38285 19940 sw
rect 38051 19898 38285 19930
tri 38285 19898 38317 19930 sw
rect 38051 19889 38317 19898
tri 38317 19889 38326 19898 sw
tri 38051 19877 38064 19889 ne
rect 38064 19877 38326 19889
tri 38326 19877 38339 19889 sw
rect 70802 19884 71000 19942
tri 38064 19831 38109 19877 ne
rect 38109 19876 38339 19877
rect 38109 19831 38202 19876
tri 38109 19821 38120 19831 ne
rect 38120 19830 38202 19831
rect 38248 19844 38339 19876
tri 38339 19844 38371 19877 sw
rect 38248 19830 38371 19844
rect 38120 19821 38371 19830
tri 38120 19808 38133 19821 ne
rect 38133 19808 38371 19821
tri 38371 19808 38407 19844 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
tri 38133 19776 38165 19808 ne
rect 38165 19798 38407 19808
tri 38407 19798 38417 19808 sw
rect 38165 19776 38417 19798
tri 38165 19766 38175 19776 ne
rect 38175 19766 38417 19776
tri 38417 19766 38449 19798 sw
rect 70802 19780 71000 19838
tri 38175 19721 38220 19766 ne
rect 38220 19753 38449 19766
tri 38449 19753 38462 19766 sw
rect 38220 19744 38462 19753
rect 38220 19721 38334 19744
tri 38220 19689 38252 19721 ne
rect 38252 19698 38334 19721
rect 38380 19721 38462 19744
tri 38462 19721 38494 19753 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19698 38494 19721
rect 38252 19689 38494 19698
tri 38252 19676 38265 19689 ne
rect 38265 19676 38494 19689
tri 38494 19676 38539 19721 sw
rect 70802 19676 71000 19734
tri 38265 19644 38297 19676 ne
rect 38297 19666 38539 19676
tri 38539 19666 38549 19676 sw
rect 38297 19644 38549 19666
tri 38297 19602 38339 19644 ne
rect 38339 19634 38549 19644
tri 38549 19634 38581 19666 sw
rect 38339 19621 38581 19634
tri 38581 19621 38594 19634 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38339 19612 38594 19621
rect 38339 19602 38466 19612
tri 38339 19570 38371 19602 ne
rect 38371 19570 38466 19602
tri 38371 19544 38397 19570 ne
rect 38397 19566 38466 19570
rect 38512 19602 38594 19612
tri 38594 19602 38613 19621 sw
rect 38512 19589 38613 19602
tri 38613 19589 38626 19602 sw
rect 38512 19566 38626 19589
rect 38397 19544 38626 19566
tri 38626 19544 38671 19589 sw
rect 70802 19572 71000 19630
tri 38397 19512 38429 19544 ne
rect 38429 19534 38671 19544
tri 38671 19534 38681 19544 sw
rect 38429 19512 38681 19534
tri 38429 19502 38439 19512 ne
rect 38439 19502 38681 19512
tri 38681 19502 38713 19534 sw
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38439 19457 38484 19502 ne
rect 38484 19480 38713 19502
rect 38484 19457 38598 19480
tri 38484 19425 38516 19457 ne
rect 38516 19434 38598 19457
rect 38644 19479 38713 19480
tri 38713 19479 38736 19502 sw
rect 38644 19457 38736 19479
tri 38736 19457 38758 19479 sw
rect 70802 19468 71000 19526
rect 38644 19434 38758 19457
rect 38516 19425 38758 19434
tri 38516 19412 38529 19425 ne
rect 38529 19412 38758 19425
tri 38758 19412 38803 19457 sw
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38529 19380 38561 19412 ne
rect 38561 19402 38803 19412
tri 38803 19402 38813 19412 sw
rect 38561 19380 38813 19402
tri 38561 19335 38606 19380 ne
rect 38606 19370 38813 19380
tri 38813 19370 38845 19402 sw
rect 38606 19357 38845 19370
tri 38845 19357 38858 19370 sw
rect 70802 19364 71000 19422
rect 38606 19348 38858 19357
rect 38606 19335 38730 19348
tri 38606 19328 38613 19335 ne
rect 38613 19328 38730 19335
tri 38613 19293 38648 19328 ne
rect 38648 19302 38730 19328
rect 38776 19328 38858 19348
tri 38858 19328 38887 19357 sw
rect 38776 19325 38887 19328
tri 38887 19325 38890 19328 sw
rect 38776 19302 38890 19325
rect 38648 19293 38890 19302
tri 38648 19280 38661 19293 ne
rect 38661 19280 38890 19293
tri 38890 19280 38935 19325 sw
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
tri 38661 19248 38693 19280 ne
rect 38693 19270 38935 19280
tri 38935 19270 38945 19280 sw
rect 38693 19248 38945 19270
tri 38693 19238 38703 19248 ne
rect 38703 19238 38945 19248
tri 38945 19238 38977 19270 sw
rect 70802 19260 71000 19318
tri 38703 19205 38736 19238 ne
rect 38736 19225 38977 19238
tri 38977 19225 38990 19238 sw
rect 38736 19216 38990 19225
rect 38736 19205 38862 19216
tri 38736 19160 38781 19205 ne
rect 38781 19170 38862 19205
rect 38908 19205 38990 19216
tri 38990 19205 39010 19225 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19170 39010 19205
rect 38781 19160 39010 19170
tri 39010 19160 39055 19205 sw
tri 38781 19148 38793 19160 ne
rect 38793 19148 39055 19160
tri 39055 19148 39067 19160 sw
rect 70802 19156 71000 19214
tri 38793 19116 38825 19148 ne
rect 38825 19138 39067 19148
tri 39067 19138 39077 19148 sw
rect 38825 19116 39077 19138
tri 38825 19071 38870 19116 ne
rect 38870 19106 39077 19116
tri 39077 19106 39109 19138 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 38870 19093 39109 19106
tri 39109 19093 39122 19106 sw
rect 38870 19084 39122 19093
rect 38870 19071 38994 19084
tri 38870 19053 38887 19071 ne
rect 38887 19053 38994 19071
tri 38887 19029 38912 19053 ne
rect 38912 19038 38994 19053
rect 39040 19053 39122 19084
tri 39122 19053 39162 19093 sw
rect 39040 19038 39162 19053
rect 38912 19029 39162 19038
tri 38912 19016 38925 19029 ne
rect 38925 19016 39162 19029
tri 39162 19016 39199 19053 sw
rect 70802 19052 71000 19110
tri 38925 18984 38957 19016 ne
rect 38957 19006 39199 19016
tri 39199 19006 39209 19016 sw
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38957 18984 39209 19006
tri 38957 18974 38967 18984 ne
rect 38967 18974 39209 18984
tri 39209 18974 39241 19006 sw
tri 38967 18929 39012 18974 ne
rect 39012 18961 39241 18974
tri 39241 18961 39254 18974 sw
rect 39012 18952 39254 18961
rect 39012 18929 39126 18952
tri 39012 18897 39044 18929 ne
rect 39044 18906 39126 18929
rect 39172 18929 39254 18952
tri 39254 18929 39286 18961 sw
rect 70802 18948 71000 19006
rect 39172 18906 39286 18929
rect 39044 18897 39286 18906
tri 39044 18884 39057 18897 ne
rect 39057 18884 39286 18897
tri 39286 18884 39331 18929 sw
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39057 18852 39089 18884 ne
rect 39089 18874 39331 18884
tri 39331 18874 39341 18884 sw
rect 39089 18852 39341 18874
tri 39089 18840 39101 18852 ne
rect 39101 18842 39341 18852
tri 39341 18842 39373 18874 sw
rect 70802 18844 71000 18902
rect 39101 18840 39373 18842
tri 39101 18795 39146 18840 ne
rect 39146 18829 39373 18840
tri 39373 18829 39386 18842 sw
rect 39146 18820 39386 18829
rect 39146 18795 39258 18820
tri 39146 18779 39162 18795 ne
rect 39162 18779 39258 18795
tri 39162 18765 39176 18779 ne
rect 39176 18774 39258 18779
rect 39304 18795 39386 18820
tri 39386 18795 39420 18829 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18779 39420 18795
tri 39420 18779 39436 18795 sw
rect 39304 18774 39436 18779
rect 39176 18765 39436 18774
tri 39176 18752 39189 18765 ne
rect 39189 18752 39436 18765
tri 39436 18752 39463 18779 sw
tri 39189 18720 39221 18752 ne
rect 39221 18750 39463 18752
tri 39463 18750 39465 18752 sw
rect 39221 18742 39465 18750
tri 39465 18742 39473 18750 sw
rect 39221 18720 39473 18742
tri 39221 18710 39231 18720 ne
rect 39231 18710 39473 18720
tri 39473 18710 39505 18742 sw
rect 70802 18740 71000 18798
tri 39231 18665 39276 18710 ne
rect 39276 18697 39505 18710
tri 39505 18697 39518 18710 sw
rect 39276 18688 39518 18697
rect 39276 18665 39390 18688
tri 39276 18633 39308 18665 ne
rect 39308 18642 39390 18665
rect 39436 18665 39518 18688
tri 39518 18665 39550 18697 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39436 18642 39550 18665
rect 39308 18633 39550 18642
tri 39308 18620 39321 18633 ne
rect 39321 18620 39550 18633
tri 39550 18620 39595 18665 sw
rect 70802 18636 71000 18694
tri 39321 18588 39353 18620 ne
rect 39353 18610 39595 18620
tri 39595 18610 39605 18620 sw
rect 39353 18588 39605 18610
tri 39353 18543 39398 18588 ne
rect 39398 18578 39605 18588
tri 39605 18578 39637 18610 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39398 18565 39637 18578
tri 39637 18565 39650 18578 sw
rect 39398 18556 39650 18565
rect 39398 18543 39522 18556
tri 39398 18505 39436 18543 ne
rect 39436 18510 39522 18543
rect 39568 18550 39650 18556
tri 39650 18550 39665 18565 sw
rect 39568 18510 39665 18550
rect 39436 18505 39665 18510
tri 39665 18505 39711 18550 sw
rect 70802 18532 71000 18590
tri 39436 18488 39453 18505 ne
rect 39453 18488 39711 18505
tri 39711 18488 39727 18505 sw
tri 39453 18475 39465 18488 ne
rect 39465 18478 39727 18488
tri 39727 18478 39737 18488 sw
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39465 18475 39737 18478
tri 39465 18446 39495 18475 ne
rect 39495 18446 39737 18475
tri 39737 18446 39769 18478 sw
tri 39495 18430 39511 18446 ne
rect 39511 18433 39769 18446
tri 39769 18433 39782 18446 sw
rect 39511 18430 39782 18433
tri 39782 18430 39785 18433 sw
tri 39511 18385 39556 18430 ne
rect 39556 18424 39785 18430
rect 39556 18385 39654 18424
tri 39556 18369 39572 18385 ne
rect 39572 18378 39654 18385
rect 39700 18385 39785 18424
tri 39785 18385 39830 18430 sw
rect 70802 18428 71000 18486
rect 39700 18378 39830 18385
rect 39572 18369 39830 18378
tri 39572 18356 39585 18369 ne
rect 39585 18356 39830 18369
tri 39830 18356 39859 18385 sw
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
tri 39585 18324 39617 18356 ne
rect 39617 18346 39859 18356
tri 39859 18346 39869 18356 sw
rect 39617 18324 39869 18346
tri 39617 18279 39662 18324 ne
rect 39662 18314 39869 18324
tri 39869 18314 39901 18346 sw
rect 70802 18324 71000 18382
rect 39662 18301 39901 18314
tri 39901 18301 39914 18314 sw
rect 39662 18292 39914 18301
rect 39662 18279 39786 18292
tri 39662 18237 39704 18279 ne
rect 39704 18246 39786 18279
rect 39832 18275 39914 18292
tri 39914 18275 39940 18301 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18246 39940 18275
rect 39704 18237 39940 18246
tri 39704 18230 39711 18237 ne
rect 39711 18230 39940 18237
tri 39940 18230 39985 18275 sw
tri 39711 18224 39717 18230 ne
rect 39717 18224 39985 18230
tri 39985 18224 39991 18230 sw
tri 39717 18192 39749 18224 ne
rect 39749 18214 39991 18224
tri 39991 18214 40001 18224 sw
rect 70802 18220 71000 18278
rect 39749 18192 40001 18214
tri 39749 18182 39759 18192 ne
rect 39759 18182 40001 18192
tri 40001 18182 40033 18214 sw
tri 39759 18137 39804 18182 ne
rect 39804 18169 40033 18182
tri 40033 18169 40046 18182 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39804 18160 40046 18169
rect 39804 18137 39918 18160
tri 39804 18111 39830 18137 ne
rect 39830 18114 39918 18137
rect 39964 18137 40046 18160
tri 40046 18137 40078 18169 sw
rect 39964 18114 40078 18137
rect 39830 18111 40078 18114
tri 39830 18092 39849 18111 ne
rect 39849 18092 40078 18111
tri 40078 18092 40123 18137 sw
rect 70802 18116 71000 18174
tri 39849 18060 39881 18092 ne
rect 39881 18082 40123 18092
tri 40123 18082 40133 18092 sw
rect 39881 18060 40133 18082
tri 39881 18015 39926 18060 ne
rect 39926 18050 40133 18060
tri 40133 18050 40165 18082 sw
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
rect 39926 18028 40165 18050
rect 39926 18015 40050 18028
tri 39926 17973 39968 18015 ne
rect 39968 17982 40050 18015
rect 40096 18020 40165 18028
tri 40165 18020 40195 18050 sw
rect 40096 18005 40195 18020
tri 40195 18005 40210 18020 sw
rect 70802 18012 71000 18070
rect 40096 17982 40210 18005
rect 39968 17973 40210 17982
tri 39968 17956 39985 17973 ne
rect 39985 17960 40210 17973
tri 40210 17960 40255 18005 sw
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 39985 17956 40255 17960
tri 40255 17956 40259 17960 sw
tri 39985 17928 40013 17956 ne
rect 40013 17950 40259 17956
tri 40259 17950 40265 17956 sw
rect 40013 17928 40265 17950
tri 40013 17918 40023 17928 ne
rect 40023 17918 40265 17928
tri 40265 17918 40297 17950 sw
tri 40023 17873 40068 17918 ne
rect 40068 17905 40297 17918
tri 40297 17905 40310 17918 sw
rect 70802 17908 71000 17966
rect 40068 17896 40310 17905
rect 40068 17873 40182 17896
tri 40068 17841 40100 17873 ne
rect 40100 17850 40182 17873
rect 40228 17873 40310 17896
tri 40310 17873 40342 17905 sw
rect 40228 17850 40342 17873
rect 40100 17841 40342 17850
tri 40100 17828 40113 17841 ne
rect 40113 17828 40342 17841
tri 40342 17828 40387 17873 sw
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
tri 40113 17796 40145 17828 ne
rect 40145 17818 40387 17828
tri 40387 17818 40397 17828 sw
rect 40145 17796 40397 17818
tri 40145 17751 40190 17796 ne
rect 40190 17786 40397 17796
tri 40397 17786 40429 17818 sw
rect 70802 17804 71000 17862
rect 40190 17773 40429 17786
tri 40429 17773 40442 17786 sw
rect 40190 17764 40442 17773
rect 40190 17751 40314 17764
tri 40190 17746 40195 17751 ne
rect 40195 17746 40314 17751
tri 40195 17701 40240 17746 ne
rect 40240 17718 40314 17746
rect 40360 17746 40442 17764
tri 40442 17746 40469 17773 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17718 40469 17746
rect 40240 17701 40469 17718
tri 40469 17701 40515 17746 sw
tri 40240 17681 40259 17701 ne
rect 40259 17696 40515 17701
tri 40515 17696 40519 17701 sw
rect 70802 17700 71000 17758
rect 40259 17681 40519 17696
tri 40519 17681 40534 17696 sw
tri 40259 17664 40277 17681 ne
rect 40277 17664 40534 17681
tri 40277 17654 40287 17664 ne
rect 40287 17654 40534 17664
tri 40534 17654 40561 17681 sw
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40287 17609 40332 17654 ne
rect 40332 17641 40561 17654
tri 40561 17641 40574 17654 sw
rect 40332 17632 40574 17641
rect 40332 17609 40446 17632
tri 40332 17577 40364 17609 ne
rect 40364 17586 40446 17609
rect 40492 17609 40574 17632
tri 40574 17609 40606 17641 sw
rect 40492 17586 40606 17609
rect 40364 17577 40606 17586
tri 40364 17564 40377 17577 ne
rect 40377 17564 40606 17577
tri 40606 17564 40651 17609 sw
rect 70802 17596 71000 17654
tri 40377 17532 40409 17564 ne
rect 40409 17554 40651 17564
tri 40651 17554 40661 17564 sw
rect 40409 17532 40661 17554
tri 40409 17487 40454 17532 ne
rect 40454 17522 40661 17532
tri 40661 17522 40693 17554 sw
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40454 17509 40693 17522
tri 40693 17509 40706 17522 sw
rect 40454 17500 40706 17509
rect 40454 17487 40578 17500
tri 40454 17445 40496 17487 ne
rect 40496 17454 40578 17487
rect 40624 17477 40706 17500
tri 40706 17477 40738 17509 sw
rect 70802 17492 71000 17550
rect 40624 17454 40738 17477
rect 40496 17445 40738 17454
tri 40496 17407 40534 17445 ne
rect 40534 17432 40738 17445
tri 40738 17432 40783 17477 sw
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 40534 17422 40783 17432
tri 40783 17422 40793 17432 sw
rect 40534 17407 40793 17422
tri 40793 17407 40808 17422 sw
tri 40534 17400 40541 17407 ne
rect 40541 17400 40808 17407
tri 40541 17390 40551 17400 ne
rect 40551 17390 40808 17400
tri 40808 17390 40825 17407 sw
tri 40551 17381 40560 17390 ne
rect 40560 17381 40825 17390
tri 40560 17336 40605 17381 ne
rect 40605 17377 40825 17381
tri 40825 17377 40838 17390 sw
rect 70802 17388 71000 17446
rect 40605 17368 40838 17377
rect 40605 17336 40710 17368
tri 40605 17313 40628 17336 ne
rect 40628 17322 40710 17336
rect 40756 17336 40838 17368
tri 40838 17336 40879 17377 sw
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40879 17336
rect 40628 17313 40879 17322
tri 40628 17300 40641 17313 ne
rect 40641 17300 40879 17313
tri 40879 17300 40915 17336 sw
tri 40641 17268 40673 17300 ne
rect 40673 17291 40915 17300
tri 40915 17291 40925 17300 sw
rect 40673 17268 40925 17291
tri 40673 17223 40718 17268 ne
rect 40718 17258 40925 17268
tri 40925 17258 40957 17290 sw
rect 70802 17284 71000 17342
rect 40718 17245 40957 17258
tri 40957 17245 40970 17258 sw
rect 40718 17236 40970 17245
rect 40718 17223 40842 17236
tri 40718 17181 40760 17223 ne
rect 40760 17190 40842 17223
rect 40888 17213 40970 17236
tri 40970 17213 41002 17245 sw
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 40888 17190 41002 17213
rect 40760 17181 41002 17190
tri 40760 17136 40805 17181 ne
rect 40805 17168 41002 17181
tri 41002 17168 41047 17213 sw
rect 70802 17180 71000 17238
rect 40805 17158 41047 17168
tri 41047 17158 41057 17168 sw
rect 40805 17136 41057 17158
tri 40805 17133 40808 17136 ne
rect 40808 17133 41057 17136
tri 41057 17133 41083 17158 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40808 17126 40815 17133 ne
rect 40815 17126 41083 17133
tri 41083 17126 41089 17133 sw
tri 40815 17081 40860 17126 ne
rect 40860 17113 41089 17126
tri 41089 17113 41102 17126 sw
rect 40860 17104 41102 17113
rect 40860 17081 40974 17104
tri 40860 17049 40892 17081 ne
rect 40892 17058 40974 17081
rect 41020 17081 41102 17104
tri 41102 17081 41134 17113 sw
rect 41020 17058 41134 17081
rect 40892 17049 41134 17058
tri 40892 17036 40905 17049 ne
rect 40905 17036 41134 17049
tri 41134 17036 41179 17081 sw
rect 70802 17076 71000 17134
tri 40905 17004 40937 17036 ne
rect 40937 17026 41179 17036
tri 41179 17026 41189 17036 sw
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40937 17004 41189 17026
tri 40937 16971 40970 17004 ne
rect 40970 16994 41189 17004
tri 41189 16994 41221 17026 sw
rect 40970 16981 41221 16994
tri 41221 16981 41234 16994 sw
rect 40970 16972 41234 16981
rect 40970 16971 41106 16972
tri 40970 16926 41015 16971 ne
rect 41015 16926 41106 16971
rect 41152 16971 41234 16972
tri 41234 16971 41244 16981 sw
rect 70802 16972 71000 17030
rect 41152 16926 41244 16971
tri 41244 16926 41289 16971 sw
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41015 16917 41024 16926 ne
rect 41024 16917 41289 16926
tri 41024 16872 41069 16917 ne
rect 41069 16904 41289 16917
tri 41289 16904 41311 16926 sw
rect 41069 16894 41311 16904
tri 41311 16894 41321 16904 sw
rect 41069 16872 41321 16894
tri 41069 16858 41083 16872 ne
rect 41083 16862 41321 16872
tri 41321 16862 41353 16894 sw
rect 70802 16868 71000 16926
rect 41083 16858 41353 16862
tri 41353 16858 41357 16862 sw
tri 41083 16813 41128 16858 ne
rect 41128 16849 41357 16858
tri 41357 16849 41366 16858 sw
rect 41128 16840 41366 16849
rect 41128 16813 41238 16840
tri 41128 16785 41156 16813 ne
rect 41156 16794 41238 16813
rect 41284 16817 41366 16840
tri 41366 16817 41398 16849 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41398 16817
rect 41156 16785 41398 16794
tri 41156 16772 41169 16785 ne
rect 41169 16772 41398 16785
tri 41398 16772 41443 16817 sw
tri 41169 16740 41201 16772 ne
rect 41201 16762 41443 16772
tri 41443 16762 41453 16772 sw
rect 70802 16764 71000 16822
rect 41201 16740 41453 16762
tri 41201 16730 41211 16740 ne
rect 41211 16730 41453 16740
tri 41453 16730 41485 16762 sw
tri 41211 16685 41256 16730 ne
rect 41256 16717 41485 16730
tri 41485 16717 41498 16730 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41256 16708 41498 16717
rect 41256 16685 41370 16708
tri 41256 16651 41289 16685 ne
rect 41289 16662 41370 16685
rect 41416 16685 41498 16708
tri 41498 16685 41530 16717 sw
rect 41416 16662 41530 16685
rect 41289 16651 41530 16662
tri 41289 16640 41301 16651 ne
rect 41301 16640 41530 16651
tri 41530 16640 41575 16685 sw
rect 70802 16660 71000 16718
tri 41301 16606 41335 16640 ne
rect 41335 16630 41575 16640
tri 41575 16630 41585 16640 sw
rect 41335 16606 41585 16630
tri 41335 16584 41357 16606 ne
rect 41357 16598 41585 16606
tri 41585 16598 41617 16630 sw
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41357 16584 41617 16598
tri 41617 16584 41631 16598 sw
tri 41357 16539 41402 16584 ne
rect 41402 16576 41631 16584
rect 41402 16539 41502 16576
tri 41402 16521 41420 16539 ne
rect 41420 16530 41502 16539
rect 41548 16561 41631 16576
tri 41631 16561 41654 16584 sw
rect 41548 16553 41654 16561
tri 41654 16553 41662 16561 sw
rect 70802 16556 71000 16614
rect 41548 16530 41662 16553
rect 41420 16521 41662 16530
tri 41420 16508 41433 16521 ne
rect 41433 16508 41662 16521
tri 41662 16508 41707 16553 sw
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41433 16476 41465 16508 ne
rect 41465 16498 41707 16508
tri 41707 16498 41717 16508 sw
rect 41465 16476 41717 16498
tri 41465 16466 41475 16476 ne
rect 41475 16466 41717 16476
tri 41717 16466 41749 16498 sw
tri 41475 16421 41520 16466 ne
rect 41520 16453 41749 16466
tri 41749 16453 41762 16466 sw
rect 41520 16444 41762 16453
rect 41520 16421 41634 16444
tri 41520 16389 41552 16421 ne
rect 41552 16398 41634 16421
rect 41680 16421 41762 16444
tri 41762 16421 41794 16453 sw
rect 70802 16452 71000 16510
rect 41680 16398 41794 16421
rect 41552 16389 41794 16398
tri 41552 16376 41565 16389 ne
rect 41565 16376 41794 16389
tri 41794 16376 41839 16421 sw
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
tri 41565 16344 41597 16376 ne
rect 41597 16366 41839 16376
tri 41839 16366 41849 16376 sw
rect 41597 16344 41849 16366
tri 41597 16309 41631 16344 ne
rect 41631 16334 41849 16344
tri 41849 16334 41881 16366 sw
rect 70802 16348 71000 16406
rect 41631 16321 41881 16334
tri 41881 16321 41894 16334 sw
rect 41631 16312 41894 16321
rect 41631 16309 41766 16312
tri 41631 16287 41654 16309 ne
rect 41654 16287 41766 16309
tri 41654 16244 41697 16287 ne
rect 41697 16266 41766 16287
rect 41812 16309 41894 16312
tri 41894 16309 41906 16321 sw
rect 41812 16289 41906 16309
tri 41906 16289 41926 16309 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16266 41926 16289
rect 41697 16244 41926 16266
tri 41926 16244 41971 16289 sw
rect 70802 16244 71000 16302
tri 41697 16212 41729 16244 ne
rect 41729 16241 41971 16244
tri 41971 16241 41974 16244 sw
rect 41729 16212 41974 16241
tri 41729 16202 41739 16212 ne
rect 41739 16202 41974 16212
tri 41974 16202 42013 16241 sw
tri 41739 16157 41784 16202 ne
rect 41784 16189 42013 16202
tri 42013 16189 42026 16202 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41784 16180 42026 16189
rect 41784 16157 41898 16180
tri 41784 16125 41816 16157 ne
rect 41816 16134 41898 16157
rect 41944 16157 42026 16180
tri 42026 16157 42058 16189 sw
rect 41944 16134 42058 16157
rect 41816 16125 42058 16134
tri 41816 16112 41829 16125 ne
rect 41829 16112 42058 16125
tri 42058 16112 42103 16157 sw
rect 70802 16140 71000 16198
tri 41829 16080 41861 16112 ne
rect 41861 16102 42103 16112
tri 42103 16102 42113 16112 sw
rect 41861 16080 42113 16102
tri 41861 16035 41906 16080 ne
rect 41906 16070 42113 16080
tri 42113 16070 42145 16102 sw
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
rect 41906 16057 42145 16070
tri 42145 16057 42158 16070 sw
rect 41906 16048 42158 16057
rect 41906 16035 42030 16048
tri 41906 15993 41948 16035 ne
rect 41948 16002 42030 16035
rect 42076 16035 42158 16048
tri 42158 16035 42180 16057 sw
rect 70802 16036 71000 16094
rect 42076 16025 42180 16035
tri 42180 16025 42190 16035 sw
rect 42076 16002 42190 16025
rect 41948 15993 42190 16002
tri 41948 15980 41961 15993 ne
rect 41961 15980 42190 15993
tri 42190 15980 42235 16025 sw
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41961 15948 41993 15980 ne
rect 41993 15970 42235 15980
tri 42235 15970 42245 15980 sw
rect 41993 15948 42245 15970
tri 41993 15938 42003 15948 ne
rect 42003 15938 42245 15948
tri 42245 15938 42277 15970 sw
tri 42003 15922 42019 15938 ne
rect 42019 15925 42277 15938
tri 42277 15925 42290 15938 sw
rect 70802 15932 71000 15990
rect 42019 15922 42290 15925
tri 42290 15922 42293 15925 sw
tri 42019 15877 42064 15922 ne
rect 42064 15916 42293 15922
rect 42064 15877 42162 15916
tri 42064 15861 42080 15877 ne
rect 42080 15870 42162 15877
rect 42208 15877 42293 15916
tri 42293 15877 42339 15922 sw
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15870 42339 15877
rect 42080 15861 42339 15870
tri 42080 15848 42093 15861 ne
rect 42093 15848 42339 15861
tri 42339 15848 42367 15877 sw
tri 42093 15816 42125 15848 ne
rect 42125 15838 42367 15848
tri 42367 15838 42377 15848 sw
rect 42125 15816 42377 15838
tri 42125 15771 42170 15816 ne
rect 42170 15806 42377 15816
tri 42377 15806 42409 15838 sw
rect 70802 15828 71000 15886
rect 42170 15793 42409 15806
tri 42409 15793 42422 15806 sw
rect 42170 15784 42422 15793
rect 42170 15771 42294 15784
tri 42170 15761 42180 15771 ne
rect 42180 15761 42294 15771
tri 42180 15729 42212 15761 ne
rect 42212 15738 42294 15761
rect 42340 15761 42422 15784
tri 42422 15761 42455 15793 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15738 42455 15761
rect 42212 15729 42455 15738
tri 42212 15716 42225 15729 ne
rect 42225 15716 42455 15729
tri 42455 15716 42499 15761 sw
rect 70802 15724 71000 15782
tri 42225 15684 42257 15716 ne
rect 42257 15706 42499 15716
tri 42499 15706 42509 15716 sw
rect 42257 15684 42509 15706
tri 42257 15674 42267 15684 ne
rect 42267 15674 42509 15684
tri 42509 15674 42541 15706 sw
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42267 15629 42312 15674 ne
rect 42312 15661 42541 15674
tri 42541 15661 42554 15674 sw
rect 42312 15652 42554 15661
rect 42312 15629 42426 15652
tri 42312 15597 42344 15629 ne
rect 42344 15606 42426 15629
rect 42472 15629 42554 15652
tri 42554 15629 42586 15661 sw
rect 42472 15606 42586 15629
rect 42344 15597 42586 15606
tri 42344 15584 42357 15597 ne
rect 42357 15584 42586 15597
tri 42586 15584 42631 15629 sw
rect 70802 15620 71000 15678
tri 42357 15552 42389 15584 ne
rect 42389 15574 42631 15584
tri 42631 15574 42641 15584 sw
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42389 15552 42641 15574
tri 42389 15512 42429 15552 ne
rect 42429 15542 42641 15552
tri 42641 15542 42673 15574 sw
rect 42429 15529 42673 15542
tri 42673 15529 42686 15542 sw
rect 42429 15520 42686 15529
rect 42429 15512 42558 15520
tri 42429 15486 42455 15512 ne
rect 42455 15486 42558 15512
tri 42455 15465 42476 15486 ne
rect 42476 15474 42558 15486
rect 42604 15512 42686 15520
tri 42686 15512 42703 15529 sw
rect 70802 15516 71000 15574
rect 42604 15486 42703 15512
tri 42703 15486 42729 15512 sw
rect 42604 15474 42729 15486
rect 42476 15467 42729 15474
tri 42729 15467 42749 15486 sw
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 42476 15465 42749 15467
tri 42476 15452 42489 15465 ne
rect 42489 15452 42749 15465
tri 42749 15452 42763 15467 sw
tri 42489 15420 42521 15452 ne
rect 42521 15442 42763 15452
tri 42763 15442 42773 15452 sw
rect 42521 15420 42773 15442
tri 42521 15410 42531 15420 ne
rect 42531 15410 42773 15420
tri 42773 15410 42805 15442 sw
rect 70802 15412 71000 15470
tri 42531 15365 42576 15410 ne
rect 42576 15397 42805 15410
tri 42805 15397 42818 15410 sw
rect 42576 15388 42818 15397
rect 42576 15365 42690 15388
tri 42576 15333 42608 15365 ne
rect 42608 15342 42690 15365
rect 42736 15365 42818 15388
tri 42818 15365 42850 15397 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42850 15365
rect 42608 15333 42850 15342
tri 42608 15320 42621 15333 ne
rect 42621 15320 42850 15333
tri 42850 15320 42895 15365 sw
tri 42621 15288 42653 15320 ne
rect 42653 15310 42895 15320
tri 42895 15310 42905 15320 sw
rect 42653 15288 42905 15310
tri 42653 15243 42698 15288 ne
rect 42698 15278 42905 15288
tri 42905 15278 42937 15310 sw
rect 70802 15308 71000 15366
rect 42698 15265 42937 15278
tri 42937 15265 42950 15278 sw
rect 42698 15257 42950 15265
tri 42950 15257 42958 15265 sw
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 42698 15256 42958 15257
rect 42698 15243 42822 15256
tri 42698 15212 42729 15243 ne
rect 42729 15212 42822 15243
tri 42729 15192 42749 15212 ne
rect 42749 15210 42822 15212
rect 42868 15212 42958 15256
tri 42958 15212 43003 15257 sw
rect 42868 15210 43003 15212
rect 42749 15192 43003 15210
tri 42749 15188 42753 15192 ne
rect 42753 15188 43003 15192
tri 43003 15188 43027 15212 sw
rect 70802 15204 71000 15262
tri 42753 15147 42794 15188 ne
rect 42794 15178 43027 15188
tri 43027 15178 43037 15188 sw
rect 42794 15147 43037 15178
tri 42794 15146 42795 15147 ne
rect 42795 15146 43037 15147
tri 43037 15146 43069 15178 sw
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42795 15101 42840 15146 ne
rect 42840 15124 43069 15146
rect 42840 15101 42954 15124
tri 42840 15069 42872 15101 ne
rect 42872 15078 42954 15101
rect 43000 15102 43069 15124
tri 43069 15102 43113 15146 sw
rect 43000 15101 43113 15102
tri 43113 15101 43114 15102 sw
rect 43000 15078 43114 15101
rect 42872 15069 43114 15078
tri 42872 15056 42885 15069 ne
rect 42885 15056 43114 15069
tri 43114 15056 43159 15101 sw
rect 70802 15100 71000 15158
tri 42885 15024 42917 15056 ne
rect 42917 15046 43159 15056
tri 43159 15046 43169 15056 sw
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
rect 42917 15024 43169 15046
tri 42917 14979 42962 15024 ne
rect 42962 15014 43169 15024
tri 43169 15014 43201 15046 sw
rect 42962 15001 43201 15014
tri 43201 15001 43214 15014 sw
rect 42962 14992 43214 15001
rect 42962 14979 43086 14992
tri 42962 14937 43003 14979 ne
rect 43003 14946 43086 14979
rect 43132 14983 43214 14992
tri 43214 14983 43233 15001 sw
rect 70802 14996 71000 15054
rect 43132 14946 43233 14983
rect 43003 14937 43233 14946
tri 43233 14937 43278 14983 sw
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
tri 43004 14924 43017 14937 ne
rect 43017 14924 43278 14937
tri 43278 14924 43291 14937 sw
tri 43017 14892 43049 14924 ne
rect 43049 14914 43291 14924
tri 43291 14914 43301 14924 sw
rect 43049 14892 43301 14914
tri 43049 14882 43059 14892 ne
rect 43059 14882 43301 14892
tri 43301 14882 43333 14914 sw
rect 70802 14892 71000 14950
tri 43059 14837 43104 14882 ne
rect 43104 14869 43333 14882
tri 43333 14869 43346 14882 sw
rect 43104 14860 43346 14869
rect 43104 14837 43218 14860
tri 43104 14827 43113 14837 ne
rect 43113 14827 43218 14837
tri 43113 14792 43149 14827 ne
rect 43149 14814 43218 14827
rect 43264 14837 43346 14860
tri 43346 14837 43378 14869 sw
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14814 43378 14837
rect 43149 14792 43378 14814
tri 43378 14792 43423 14837 sw
tri 43149 14760 43181 14792 ne
rect 43181 14782 43423 14792
tri 43423 14782 43433 14792 sw
rect 70802 14788 71000 14846
rect 43181 14760 43433 14782
tri 43181 14715 43226 14760 ne
rect 43226 14750 43433 14760
tri 43433 14750 43465 14782 sw
rect 43226 14737 43465 14750
tri 43465 14737 43478 14750 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 43226 14728 43478 14737
rect 43226 14715 43350 14728
tri 43226 14673 43268 14715 ne
rect 43268 14682 43350 14715
rect 43396 14708 43478 14728
tri 43478 14708 43507 14737 sw
rect 43396 14682 43507 14708
rect 43268 14673 43507 14682
tri 43268 14663 43278 14673 ne
rect 43278 14663 43507 14673
tri 43507 14663 43552 14708 sw
rect 70802 14684 71000 14742
tri 43278 14660 43281 14663 ne
rect 43281 14660 43552 14663
tri 43552 14660 43555 14663 sw
tri 43281 14628 43313 14660 ne
rect 43313 14650 43555 14660
tri 43555 14650 43565 14660 sw
rect 43313 14628 43565 14650
tri 43313 14618 43323 14628 ne
rect 43323 14618 43565 14628
tri 43565 14618 43597 14650 sw
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43323 14573 43368 14618 ne
rect 43368 14605 43597 14618
tri 43597 14605 43610 14618 sw
rect 43368 14596 43610 14605
rect 43368 14573 43482 14596
tri 43368 14541 43400 14573 ne
rect 43400 14550 43482 14573
rect 43528 14573 43610 14596
tri 43610 14573 43642 14605 sw
rect 70802 14580 71000 14638
rect 43528 14550 43642 14573
rect 43400 14541 43642 14550
tri 43400 14528 43413 14541 ne
rect 43413 14528 43642 14541
tri 43642 14528 43687 14573 sw
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43413 14496 43445 14528 ne
rect 43445 14518 43687 14528
tri 43687 14518 43697 14528 sw
rect 43445 14496 43697 14518
tri 43445 14463 43478 14496 ne
rect 43478 14486 43697 14496
tri 43697 14486 43729 14518 sw
rect 43478 14473 43729 14486
tri 43729 14473 43742 14486 sw
rect 70802 14476 71000 14534
rect 43478 14464 43742 14473
rect 43478 14463 43614 14464
tri 43478 14417 43523 14463 ne
rect 43523 14418 43614 14463
rect 43660 14463 43742 14464
tri 43742 14463 43753 14473 sw
rect 43660 14418 43753 14463
rect 43523 14417 43753 14418
tri 43753 14417 43798 14463 sw
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
tri 43523 14409 43532 14417 ne
rect 43532 14409 43798 14417
tri 43532 14389 43552 14409 ne
rect 43552 14396 43798 14409
tri 43798 14396 43819 14417 sw
rect 43552 14389 43819 14396
tri 43819 14389 43827 14396 sw
tri 43552 14364 43577 14389 ne
rect 43577 14386 43827 14389
tri 43827 14386 43829 14389 sw
rect 43577 14364 43829 14386
tri 43577 14354 43587 14364 ne
rect 43587 14354 43829 14364
tri 43829 14354 43861 14386 sw
rect 70802 14372 71000 14430
tri 43587 14309 43632 14354 ne
rect 43632 14341 43861 14354
tri 43861 14341 43874 14354 sw
rect 43632 14332 43874 14341
rect 43632 14309 43746 14332
tri 43632 14277 43664 14309 ne
rect 43664 14286 43746 14309
rect 43792 14309 43874 14332
tri 43874 14309 43906 14341 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14286 43906 14309
rect 43664 14277 43906 14286
tri 43664 14264 43677 14277 ne
rect 43677 14264 43906 14277
tri 43906 14264 43951 14309 sw
rect 70802 14268 71000 14326
tri 43677 14232 43709 14264 ne
rect 43709 14254 43951 14264
tri 43951 14254 43961 14264 sw
rect 43709 14232 43961 14254
tri 43709 14187 43754 14232 ne
rect 43754 14222 43961 14232
tri 43961 14222 43993 14254 sw
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
rect 43754 14209 43993 14222
tri 43993 14209 44006 14222 sw
rect 43754 14200 44006 14209
rect 43754 14187 43878 14200
tri 43754 14145 43796 14187 ne
rect 43796 14154 43878 14187
rect 43924 14177 44006 14200
tri 44006 14177 44038 14209 sw
rect 43924 14154 44038 14177
rect 43796 14145 44038 14154
tri 43796 14114 43827 14145 ne
rect 43827 14132 44038 14145
tri 44038 14132 44083 14177 sw
rect 70802 14164 71000 14222
rect 43827 14122 44083 14132
tri 44083 14122 44093 14132 sw
rect 43827 14114 44093 14122
tri 44093 14114 44101 14122 sw
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43827 14100 43841 14114 ne
rect 43841 14100 44101 14114
tri 43841 14098 43843 14100 ne
rect 43843 14098 44101 14100
tri 43843 14090 43851 14098 ne
rect 43851 14090 44101 14098
tri 44101 14090 44125 14114 sw
tri 43851 14053 43888 14090 ne
rect 43888 14077 44125 14090
tri 44125 14077 44138 14090 sw
rect 43888 14068 44138 14077
rect 43888 14053 44010 14068
tri 43888 14013 43928 14053 ne
rect 43928 14022 44010 14053
rect 44056 14053 44138 14068
tri 44138 14053 44163 14077 sw
rect 70802 14060 71000 14118
rect 44056 14022 44163 14053
rect 43928 14013 44163 14022
tri 43928 14000 43941 14013 ne
rect 43941 14007 44163 14013
tri 44163 14007 44208 14053 sw
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 43941 14000 44208 14007
tri 44208 14000 44215 14007 sw
tri 43941 13968 43973 14000 ne
rect 43973 13990 44215 14000
tri 44215 13990 44225 14000 sw
rect 43973 13968 44225 13990
tri 43973 13923 44018 13968 ne
rect 44018 13958 44225 13968
tri 44225 13958 44257 13990 sw
rect 44018 13945 44257 13958
tri 44257 13945 44270 13958 sw
rect 70802 13956 71000 14014
rect 44018 13936 44270 13945
rect 44018 13923 44142 13936
tri 44018 13881 44060 13923 ne
rect 44060 13890 44142 13923
rect 44188 13913 44270 13936
tri 44270 13913 44302 13945 sw
rect 44188 13890 44302 13913
rect 44060 13881 44302 13890
tri 44060 13840 44101 13881 ne
rect 44101 13868 44302 13881
tri 44302 13868 44347 13913 sw
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 44101 13858 44347 13868
tri 44347 13858 44357 13868 sw
rect 44101 13840 44357 13858
tri 44357 13840 44375 13858 sw
rect 70802 13852 71000 13910
tri 44101 13836 44105 13840 ne
rect 44105 13836 44375 13840
tri 44105 13826 44115 13836 ne
rect 44115 13826 44375 13836
tri 44375 13826 44389 13840 sw
tri 44115 13781 44160 13826 ne
rect 44160 13813 44389 13826
tri 44389 13813 44402 13826 sw
rect 44160 13804 44402 13813
rect 44160 13781 44274 13804
tri 44160 13736 44205 13781 ne
rect 44205 13758 44274 13781
rect 44320 13781 44402 13804
tri 44402 13781 44434 13813 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44320 13758 44434 13781
rect 44205 13736 44434 13758
tri 44434 13736 44479 13781 sw
rect 70802 13748 71000 13806
tri 44205 13733 44208 13736 ne
rect 44208 13733 44479 13736
tri 44208 13688 44253 13733 ne
rect 44253 13726 44479 13733
tri 44479 13726 44489 13736 sw
rect 44253 13694 44489 13726
tri 44489 13694 44521 13726 sw
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44253 13688 44521 13694
tri 44521 13688 44527 13694 sw
tri 44253 13643 44298 13688 ne
rect 44298 13672 44527 13688
rect 44298 13643 44406 13672
tri 44298 13617 44324 13643 ne
rect 44324 13626 44406 13643
rect 44452 13643 44527 13672
tri 44527 13643 44573 13688 sw
rect 70802 13644 71000 13702
rect 44452 13626 44573 13643
rect 44324 13617 44573 13626
tri 44324 13572 44369 13617 ne
rect 44369 13604 44573 13617
tri 44573 13604 44611 13643 sw
rect 44369 13594 44611 13604
tri 44611 13594 44621 13604 sw
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44369 13572 44621 13594
tri 44369 13565 44375 13572 ne
rect 44375 13565 44621 13572
tri 44621 13565 44650 13594 sw
tri 44375 13562 44379 13565 ne
rect 44379 13562 44650 13565
tri 44650 13562 44653 13565 sw
tri 44379 13517 44424 13562 ne
rect 44424 13549 44653 13562
tri 44653 13549 44666 13562 sw
rect 44424 13540 44666 13549
rect 44424 13517 44538 13540
tri 44424 13485 44456 13517 ne
rect 44456 13494 44538 13517
rect 44584 13517 44666 13540
tri 44666 13517 44698 13549 sw
rect 70802 13540 71000 13598
rect 44584 13494 44698 13517
rect 44456 13485 44698 13494
tri 44456 13472 44469 13485 ne
rect 44469 13472 44698 13485
tri 44698 13472 44743 13517 sw
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44469 13440 44501 13472 ne
rect 44501 13462 44743 13472
tri 44743 13462 44753 13472 sw
rect 44501 13440 44753 13462
tri 44501 13430 44511 13440 ne
rect 44511 13430 44753 13440
tri 44753 13430 44785 13462 sw
rect 70802 13436 71000 13494
tri 44511 13385 44556 13430 ne
rect 44556 13417 44785 13430
tri 44785 13417 44798 13430 sw
rect 44556 13413 44798 13417
tri 44798 13413 44802 13417 sw
rect 44556 13408 44802 13413
rect 44556 13385 44670 13408
tri 44556 13368 44573 13385 ne
rect 44573 13368 44670 13385
tri 44573 13340 44601 13368 ne
rect 44601 13362 44670 13368
rect 44716 13368 44802 13408
tri 44802 13368 44847 13413 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13362 44847 13368
rect 44601 13340 44847 13362
tri 44847 13340 44875 13368 sw
tri 44601 13308 44633 13340 ne
rect 44633 13336 44875 13340
tri 44875 13336 44879 13340 sw
rect 44633 13308 44879 13336
tri 44633 13291 44650 13308 ne
rect 44650 13291 44879 13308
tri 44879 13291 44924 13336 sw
rect 70802 13291 71000 13390
tri 44650 13278 44663 13291 ne
rect 44663 13278 71000 13291
tri 44663 13233 44708 13278 ne
rect 44708 13269 71000 13278
rect 44708 13256 45088 13269
rect 44708 13233 44850 13256
tri 44708 13201 44740 13233 ne
rect 44740 13210 44850 13233
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44740 13201 71000 13210
tri 44740 13188 44753 13201 ne
rect 44753 13188 71000 13201
tri 44753 13156 44785 13188 ne
rect 44785 13165 71000 13188
rect 44785 13156 45088 13165
tri 44785 13111 44830 13156 ne
rect 44830 13119 45088 13156
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44830 13111 71000 13119
tri 44830 13110 44831 13111 ne
rect 44831 13110 71000 13111
tri 44831 13097 44844 13110 ne
rect 44844 13097 71000 13110
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 13914 44118 13960 44164
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 14970 43062 15016 43108
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 15366 42666 15412 42712
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 15894 42138 15940 42184
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 16422 41610 16468 41656
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 16818 41214 16864 41260
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 17346 40686 17392 40732
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 17874 40158 17920 40204
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 18798 39234 18844 39280
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 18930 39102 18976 39148
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 19854 38178 19900 38224
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 20778 37254 20824 37300
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 20910 37122 20956 37168
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 21306 36726 21352 36772
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 21834 36198 21880 36244
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 22230 35802 22276 35848
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 22758 35274 22804 35320
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 24210 33822 24256 33868
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 24738 33294 24784 33340
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 25662 32370 25708 32416
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 25794 32238 25840 32284
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 26190 31842 26236 31888
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 26718 31314 26764 31360
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 27642 30390 27688 30436
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 28170 29862 28216 29908
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 28698 29334 28744 29380
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 29226 28806 29272 28852
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 29622 28410 29668 28456
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 30150 27882 30196 27928
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 31074 26958 31120 27004
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 31206 26826 31252 26872
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 31602 26430 31648 26476
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 32526 25506 32572 25552
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 32658 25374 32704 25420
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 33054 24978 33100 25024
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 34110 23922 34156 23968
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 34506 23526 34552 23572
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 35034 22998 35080 23044
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 36486 21546 36532 21592
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 37542 20490 37588 20536
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 37938 20094 37984 20140
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 38466 19566 38512 19612
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 38994 19038 39040 19084
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 39390 18642 39436 18688
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 39522 18510 39568 18556
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 39918 18114 39964 18160
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 40446 17586 40492 17632
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 40842 17190 40888 17236
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 40974 17058 41020 17104
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 41370 16662 41416 16708
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 41898 16134 41944 16180
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 43350 14682 43396 14728
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 45022 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 70813 44844 71000 44902
rect 13243 44824 13311 44835
rect 13243 44778 13254 44824
rect 13300 44778 13311 44824
rect 13243 44767 13311 44778
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 70813 44740 71000 44798
rect 13375 44692 13443 44703
rect 13375 44646 13386 44692
rect 13432 44646 13443 44692
rect 13375 44635 13443 44646
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 70813 44636 71000 44694
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
rect 13507 44560 13575 44571
rect 13507 44514 13518 44560
rect 13564 44514 13575 44560
rect 13507 44503 13575 44514
rect 70813 44532 71000 44590
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 13639 44428 13707 44439
rect 13639 44382 13650 44428
rect 13696 44382 13707 44428
rect 13639 44371 13707 44382
rect 70813 44428 71000 44486
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 70813 44324 71000 44382
rect 13771 44296 13839 44307
rect 13771 44250 13782 44296
rect 13828 44250 13839 44296
rect 13771 44239 13839 44250
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 70813 44220 71000 44278
rect 13903 44164 13971 44175
rect 13903 44118 13914 44164
rect 13960 44118 13971 44164
rect 13903 44107 13971 44118
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 70813 44116 71000 44174
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 14035 44032 14103 44043
rect 14035 43986 14046 44032
rect 14092 43986 14103 44032
rect 14035 43975 14103 43986
rect 70813 44012 71000 44070
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
rect 14167 43900 14235 43911
rect 14167 43854 14178 43900
rect 14224 43854 14235 43900
rect 14167 43843 14235 43854
rect 70813 43908 71000 43966
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 70813 43804 71000 43862
rect 14299 43768 14367 43779
rect 14299 43722 14310 43768
rect 14356 43722 14367 43768
rect 14299 43711 14367 43722
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 70813 43700 71000 43758
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14431 43636 14499 43647
rect 14431 43590 14442 43636
rect 14488 43590 14499 43636
rect 14431 43579 14499 43590
rect 70813 43596 71000 43654
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14563 43504 14631 43515
rect 14563 43458 14574 43504
rect 14620 43458 14631 43504
rect 14563 43447 14631 43458
rect 70813 43492 71000 43550
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
rect 70813 43388 71000 43446
rect 14695 43372 14763 43383
rect 14695 43326 14706 43372
rect 14752 43326 14763 43372
rect 14695 43315 14763 43326
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 70813 43284 71000 43342
rect 14827 43240 14895 43251
rect 14827 43194 14838 43240
rect 14884 43194 14895 43240
rect 14827 43183 14895 43194
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 70813 43180 71000 43238
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
rect 14959 43108 15027 43119
rect 14959 43062 14970 43108
rect 15016 43062 15027 43108
rect 14959 43051 15027 43062
rect 70813 43076 71000 43134
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
rect 15091 42976 15159 42987
rect 15091 42930 15102 42976
rect 15148 42930 15159 42976
rect 15091 42919 15159 42930
rect 70813 42972 71000 43030
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
rect 70813 42868 71000 42926
rect 15223 42844 15291 42855
rect 15223 42798 15234 42844
rect 15280 42798 15291 42844
rect 15223 42787 15291 42798
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 70813 42764 71000 42822
rect 15355 42712 15423 42723
rect 15355 42666 15366 42712
rect 15412 42666 15423 42712
rect 15355 42655 15423 42666
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 70813 42660 71000 42718
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
rect 15487 42580 15555 42591
rect 15487 42534 15498 42580
rect 15544 42534 15555 42580
rect 15487 42523 15555 42534
rect 70813 42556 71000 42614
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15619 42448 15687 42459
rect 15619 42402 15630 42448
rect 15676 42402 15687 42448
rect 15619 42391 15687 42402
rect 70813 42452 71000 42510
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 70813 42348 71000 42406
rect 15751 42316 15819 42327
rect 15751 42270 15762 42316
rect 15808 42270 15819 42316
rect 15751 42259 15819 42270
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 70813 42244 71000 42302
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 15883 42184 15951 42195
rect 15883 42138 15894 42184
rect 15940 42138 15951 42184
rect 15883 42127 15951 42138
rect 70813 42140 71000 42198
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
rect 16015 42052 16083 42063
rect 16015 42006 16026 42052
rect 16072 42006 16083 42052
rect 16015 41995 16083 42006
rect 70813 42036 71000 42094
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
rect 70813 41932 71000 41990
rect 16147 41920 16215 41931
rect 16147 41874 16158 41920
rect 16204 41874 16215 41920
rect 16147 41863 16215 41874
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 70813 41828 71000 41886
rect 16279 41788 16347 41799
rect 16279 41742 16290 41788
rect 16336 41742 16347 41788
rect 16279 41731 16347 41742
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 70813 41724 71000 41782
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16411 41656 16479 41667
rect 16411 41610 16422 41656
rect 16468 41610 16479 41656
rect 16411 41599 16479 41610
rect 70813 41620 71000 41678
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
rect 16543 41524 16611 41535
rect 16543 41478 16554 41524
rect 16600 41478 16611 41524
rect 16543 41467 16611 41478
rect 70813 41516 71000 41574
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 70813 41412 71000 41470
rect 16675 41392 16743 41403
rect 16675 41346 16686 41392
rect 16732 41346 16743 41392
rect 16675 41335 16743 41346
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 70813 41308 71000 41366
rect 16807 41260 16875 41271
rect 16807 41214 16818 41260
rect 16864 41214 16875 41260
rect 16807 41203 16875 41214
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 70813 41204 71000 41262
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 16939 41128 17007 41139
rect 16939 41082 16950 41128
rect 16996 41082 17007 41128
rect 16939 41071 17007 41082
rect 70813 41100 71000 41158
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 17071 40996 17139 41007
rect 17071 40950 17082 40996
rect 17128 40950 17139 40996
rect 17071 40939 17139 40950
rect 70813 40996 71000 41054
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 70813 40892 71000 40950
rect 17203 40864 17271 40875
rect 17203 40818 17214 40864
rect 17260 40818 17271 40864
rect 17203 40807 17271 40818
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 70813 40788 71000 40846
rect 17335 40732 17403 40743
rect 17335 40686 17346 40732
rect 17392 40686 17403 40732
rect 17335 40675 17403 40686
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 70813 40684 71000 40742
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
rect 17467 40600 17535 40611
rect 17467 40554 17478 40600
rect 17524 40554 17535 40600
rect 17467 40543 17535 40554
rect 70813 40580 71000 40638
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
rect 17599 40468 17667 40479
rect 17599 40422 17610 40468
rect 17656 40422 17667 40468
rect 17599 40411 17667 40422
rect 70813 40476 71000 40534
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 70813 40372 71000 40430
rect 17731 40336 17799 40347
rect 17731 40290 17742 40336
rect 17788 40290 17799 40336
rect 17731 40279 17799 40290
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 70813 40268 71000 40326
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17863 40204 17931 40215
rect 17863 40158 17874 40204
rect 17920 40158 17931 40204
rect 17863 40147 17931 40158
rect 70813 40164 71000 40222
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
rect 17995 40072 18063 40083
rect 17995 40026 18006 40072
rect 18052 40026 18063 40072
rect 17995 40015 18063 40026
rect 70813 40060 71000 40118
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 70813 39956 71000 40014
rect 18127 39940 18195 39951
rect 18127 39894 18138 39940
rect 18184 39894 18195 39940
rect 18127 39883 18195 39894
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 70813 39852 71000 39910
rect 18259 39808 18327 39819
rect 18259 39762 18270 39808
rect 18316 39762 18327 39808
rect 18259 39751 18327 39762
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 70813 39748 71000 39806
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18391 39676 18459 39687
rect 18391 39630 18402 39676
rect 18448 39630 18459 39676
rect 18391 39619 18459 39630
rect 70813 39644 71000 39702
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
rect 18523 39544 18591 39555
rect 18523 39498 18534 39544
rect 18580 39498 18591 39544
rect 18523 39487 18591 39498
rect 70813 39540 71000 39598
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
rect 70813 39436 71000 39494
rect 18655 39412 18723 39423
rect 18655 39366 18666 39412
rect 18712 39366 18723 39412
rect 18655 39355 18723 39366
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 70813 39332 71000 39390
rect 18787 39280 18855 39291
rect 18787 39234 18798 39280
rect 18844 39234 18855 39280
rect 18787 39223 18855 39234
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 70813 39228 71000 39286
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18919 39148 18987 39159
rect 18919 39102 18930 39148
rect 18976 39102 18987 39148
rect 18919 39091 18987 39102
rect 70813 39124 71000 39182
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
rect 19051 39016 19119 39027
rect 19051 38970 19062 39016
rect 19108 38970 19119 39016
rect 19051 38959 19119 38970
rect 70813 39020 71000 39078
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 70813 38916 71000 38974
rect 19183 38884 19251 38895
rect 19183 38838 19194 38884
rect 19240 38838 19251 38884
rect 19183 38827 19251 38838
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 70813 38812 71000 38870
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
rect 19315 38752 19383 38763
rect 19315 38706 19326 38752
rect 19372 38706 19383 38752
rect 19315 38695 19383 38706
rect 70813 38708 71000 38766
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
rect 19447 38620 19515 38631
rect 19447 38574 19458 38620
rect 19504 38574 19515 38620
rect 19447 38563 19515 38574
rect 70813 38604 71000 38662
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 70813 38500 71000 38558
rect 19579 38488 19647 38499
rect 19579 38442 19590 38488
rect 19636 38442 19647 38488
rect 19579 38431 19647 38442
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 70813 38396 71000 38454
rect 19711 38356 19779 38367
rect 19711 38310 19722 38356
rect 19768 38310 19779 38356
rect 19711 38299 19779 38310
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 70813 38292 71000 38350
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19843 38224 19911 38235
rect 19843 38178 19854 38224
rect 19900 38178 19911 38224
rect 19843 38167 19911 38178
rect 70813 38188 71000 38246
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19975 38092 20043 38103
rect 19975 38046 19986 38092
rect 20032 38046 20043 38092
rect 19975 38035 20043 38046
rect 70813 38084 71000 38142
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 70813 37980 71000 38038
rect 20107 37960 20175 37971
rect 20107 37914 20118 37960
rect 20164 37914 20175 37960
rect 20107 37903 20175 37914
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 70813 37876 71000 37934
rect 20239 37828 20307 37839
rect 20239 37782 20250 37828
rect 20296 37782 20307 37828
rect 20239 37771 20307 37782
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 70813 37772 71000 37830
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 20371 37696 20439 37707
rect 20371 37650 20382 37696
rect 20428 37650 20439 37696
rect 20371 37639 20439 37650
rect 70813 37668 71000 37726
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
rect 20503 37564 20571 37575
rect 20503 37518 20514 37564
rect 20560 37518 20571 37564
rect 20503 37507 20571 37518
rect 70813 37564 71000 37622
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 70813 37460 71000 37518
rect 20635 37432 20703 37443
rect 20635 37386 20646 37432
rect 20692 37386 20703 37432
rect 20635 37375 20703 37386
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 70813 37356 71000 37414
rect 20767 37300 20835 37311
rect 20767 37254 20778 37300
rect 20824 37254 20835 37300
rect 20767 37243 20835 37254
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 70813 37252 71000 37310
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20899 37168 20967 37179
rect 20899 37122 20910 37168
rect 20956 37122 20967 37168
rect 20899 37111 20967 37122
rect 70813 37148 71000 37206
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
rect 21031 37036 21099 37047
rect 21031 36990 21042 37036
rect 21088 36990 21099 37036
rect 21031 36979 21099 36990
rect 70813 37044 71000 37102
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 70813 36940 71000 36998
rect 21163 36904 21231 36915
rect 21163 36858 21174 36904
rect 21220 36858 21231 36904
rect 21163 36847 21231 36858
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 70813 36836 71000 36894
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21295 36772 21363 36783
rect 21295 36726 21306 36772
rect 21352 36726 21363 36772
rect 21295 36715 21363 36726
rect 70813 36732 71000 36790
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21427 36640 21495 36651
rect 21427 36594 21438 36640
rect 21484 36594 21495 36640
rect 21427 36583 21495 36594
rect 70813 36628 71000 36686
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
rect 70813 36524 71000 36582
rect 21559 36508 21627 36519
rect 21559 36462 21570 36508
rect 21616 36462 21627 36508
rect 21559 36451 21627 36462
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 70813 36420 71000 36478
rect 21691 36376 21759 36387
rect 21691 36330 21702 36376
rect 21748 36330 21759 36376
rect 21691 36319 21759 36330
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 70813 36316 71000 36374
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 21823 36244 21891 36255
rect 21823 36198 21834 36244
rect 21880 36198 21891 36244
rect 21823 36187 21891 36198
rect 70813 36212 71000 36270
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
rect 21955 36112 22023 36123
rect 21955 36066 21966 36112
rect 22012 36066 22023 36112
rect 21955 36055 22023 36066
rect 70813 36108 71000 36166
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 70813 36004 71000 36062
rect 22087 35980 22155 35991
rect 22087 35934 22098 35980
rect 22144 35934 22155 35980
rect 22087 35923 22155 35934
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 70813 35900 71000 35958
rect 22219 35848 22287 35859
rect 22219 35802 22230 35848
rect 22276 35802 22287 35848
rect 22219 35791 22287 35802
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 70813 35796 71000 35854
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
rect 22351 35716 22419 35727
rect 22351 35670 22362 35716
rect 22408 35670 22419 35716
rect 22351 35659 22419 35670
rect 70813 35692 71000 35750
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 22483 35584 22551 35595
rect 22483 35538 22494 35584
rect 22540 35538 22551 35584
rect 22483 35527 22551 35538
rect 70813 35588 71000 35646
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 70813 35484 71000 35542
rect 22615 35452 22683 35463
rect 22615 35406 22626 35452
rect 22672 35406 22683 35452
rect 22615 35395 22683 35406
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 70813 35380 71000 35438
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22747 35320 22815 35331
rect 22747 35274 22758 35320
rect 22804 35274 22815 35320
rect 22747 35263 22815 35274
rect 70813 35276 71000 35334
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
rect 22879 35188 22947 35199
rect 22879 35142 22890 35188
rect 22936 35142 22947 35188
rect 22879 35131 22947 35142
rect 70813 35172 71000 35230
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 70813 35068 71000 35126
rect 23011 35056 23079 35067
rect 23011 35010 23022 35056
rect 23068 35010 23079 35056
rect 23011 34999 23079 35010
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 70813 34964 71000 35022
rect 23143 34924 23211 34935
rect 23143 34878 23154 34924
rect 23200 34878 23211 34924
rect 23143 34867 23211 34878
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 70813 34860 71000 34918
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23275 34792 23343 34803
rect 23275 34746 23286 34792
rect 23332 34746 23343 34792
rect 23275 34735 23343 34746
rect 70813 34756 71000 34814
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
rect 23407 34660 23475 34671
rect 23407 34614 23418 34660
rect 23464 34614 23475 34660
rect 23407 34603 23475 34614
rect 70813 34652 71000 34710
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 70813 34548 71000 34606
rect 23539 34528 23607 34539
rect 23539 34482 23550 34528
rect 23596 34482 23607 34528
rect 23539 34471 23607 34482
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 70813 34444 71000 34502
rect 23671 34396 23739 34407
rect 23671 34350 23682 34396
rect 23728 34350 23739 34396
rect 23671 34339 23739 34350
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 70813 34340 71000 34398
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
rect 23803 34264 23871 34275
rect 23803 34218 23814 34264
rect 23860 34218 23871 34264
rect 23803 34207 23871 34218
rect 70813 34236 71000 34294
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23935 34132 24003 34143
rect 23935 34086 23946 34132
rect 23992 34086 24003 34132
rect 23935 34075 24003 34086
rect 70813 34132 71000 34190
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 70813 34028 71000 34086
rect 24067 34000 24135 34011
rect 24067 33954 24078 34000
rect 24124 33954 24135 34000
rect 24067 33943 24135 33954
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 70813 33924 71000 33982
rect 24199 33868 24267 33879
rect 24199 33822 24210 33868
rect 24256 33822 24267 33868
rect 24199 33811 24267 33822
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 70813 33820 71000 33878
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
rect 24331 33736 24399 33747
rect 24331 33690 24342 33736
rect 24388 33690 24399 33736
rect 24331 33679 24399 33690
rect 70813 33716 71000 33774
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 24463 33604 24531 33615
rect 24463 33558 24474 33604
rect 24520 33558 24531 33604
rect 24463 33547 24531 33558
rect 70813 33612 71000 33670
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 70813 33508 71000 33566
rect 24595 33472 24663 33483
rect 24595 33426 24606 33472
rect 24652 33426 24663 33472
rect 24595 33415 24663 33426
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 70813 33404 71000 33462
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 24727 33340 24795 33351
rect 24727 33294 24738 33340
rect 24784 33294 24795 33340
rect 24727 33283 24795 33294
rect 70813 33300 71000 33358
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
rect 24859 33208 24927 33219
rect 24859 33162 24870 33208
rect 24916 33162 24927 33208
rect 24859 33151 24927 33162
rect 70813 33196 71000 33254
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 70813 33092 71000 33150
rect 24991 33076 25059 33087
rect 24991 33030 25002 33076
rect 25048 33030 25059 33076
rect 24991 33019 25059 33030
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 70813 32988 71000 33046
rect 25123 32944 25191 32955
rect 25123 32898 25134 32944
rect 25180 32898 25191 32944
rect 25123 32887 25191 32898
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 70813 32884 71000 32942
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 25255 32812 25323 32823
rect 25255 32766 25266 32812
rect 25312 32766 25323 32812
rect 25255 32755 25323 32766
rect 70813 32780 71000 32838
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
rect 25387 32680 25455 32691
rect 25387 32634 25398 32680
rect 25444 32634 25455 32680
rect 25387 32623 25455 32634
rect 70813 32676 71000 32734
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
rect 70813 32572 71000 32630
rect 25519 32548 25587 32559
rect 25519 32502 25530 32548
rect 25576 32502 25587 32548
rect 25519 32491 25587 32502
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 70813 32468 71000 32526
rect 25651 32416 25719 32427
rect 25651 32370 25662 32416
rect 25708 32370 25719 32416
rect 25651 32359 25719 32370
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 70813 32364 71000 32422
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 25783 32284 25851 32295
rect 25783 32238 25794 32284
rect 25840 32238 25851 32284
rect 25783 32227 25851 32238
rect 70813 32260 71000 32318
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
rect 25915 32152 25983 32163
rect 25915 32106 25926 32152
rect 25972 32106 25983 32152
rect 25915 32095 25983 32106
rect 70813 32156 71000 32214
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 70813 32052 71000 32110
rect 26047 32020 26115 32031
rect 26047 31974 26058 32020
rect 26104 31974 26115 32020
rect 26047 31963 26115 31974
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 70813 31948 71000 32006
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26179 31888 26247 31899
rect 26179 31842 26190 31888
rect 26236 31842 26247 31888
rect 26179 31831 26247 31842
rect 70813 31844 71000 31902
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26311 31756 26379 31767
rect 26311 31710 26322 31756
rect 26368 31710 26379 31756
rect 26311 31699 26379 31710
rect 70813 31740 71000 31798
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 70813 31636 71000 31694
rect 26443 31624 26511 31635
rect 26443 31578 26454 31624
rect 26500 31578 26511 31624
rect 26443 31567 26511 31578
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 70813 31532 71000 31590
rect 26575 31492 26643 31503
rect 26575 31446 26586 31492
rect 26632 31446 26643 31492
rect 26575 31435 26643 31446
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 70813 31428 71000 31486
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 26707 31360 26775 31371
rect 26707 31314 26718 31360
rect 26764 31314 26775 31360
rect 26707 31303 26775 31314
rect 70813 31324 71000 31382
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26839 31228 26907 31239
rect 26839 31182 26850 31228
rect 26896 31182 26907 31228
rect 26839 31171 26907 31182
rect 70813 31220 71000 31278
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 70813 31116 71000 31174
rect 26971 31096 27039 31107
rect 26971 31050 26982 31096
rect 27028 31050 27039 31096
rect 26971 31039 27039 31050
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 70813 31012 71000 31070
rect 27103 30964 27171 30975
rect 27103 30918 27114 30964
rect 27160 30918 27171 30964
rect 27103 30907 27171 30918
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 70813 30908 71000 30966
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27235 30832 27303 30843
rect 27235 30786 27246 30832
rect 27292 30786 27303 30832
rect 27235 30775 27303 30786
rect 70813 30804 71000 30862
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
rect 27367 30700 27435 30711
rect 27367 30654 27378 30700
rect 27424 30654 27435 30700
rect 27367 30643 27435 30654
rect 70813 30700 71000 30758
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 70813 30596 71000 30654
rect 27499 30568 27567 30579
rect 27499 30522 27510 30568
rect 27556 30522 27567 30568
rect 27499 30511 27567 30522
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 70813 30492 71000 30550
rect 27631 30436 27699 30447
rect 27631 30390 27642 30436
rect 27688 30390 27699 30436
rect 27631 30379 27699 30390
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 70813 30388 71000 30446
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
rect 27763 30304 27831 30315
rect 27763 30258 27774 30304
rect 27820 30258 27831 30304
rect 27763 30247 27831 30258
rect 70813 30284 71000 30342
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
rect 27895 30172 27963 30183
rect 27895 30126 27906 30172
rect 27952 30126 27963 30172
rect 27895 30115 27963 30126
rect 70813 30180 71000 30238
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 70813 30076 71000 30134
rect 28027 30040 28095 30051
rect 28027 29994 28038 30040
rect 28084 29994 28095 30040
rect 28027 29983 28095 29994
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 70813 29972 71000 30030
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28159 29908 28227 29919
rect 28159 29862 28170 29908
rect 28216 29862 28227 29908
rect 28159 29851 28227 29862
rect 70813 29868 71000 29926
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28291 29776 28359 29787
rect 28291 29730 28302 29776
rect 28348 29730 28359 29776
rect 28291 29719 28359 29730
rect 70813 29764 71000 29822
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 70813 29660 71000 29718
rect 28423 29644 28491 29655
rect 28423 29598 28434 29644
rect 28480 29598 28491 29644
rect 28423 29587 28491 29598
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 70813 29556 71000 29614
rect 28555 29512 28623 29523
rect 28555 29466 28566 29512
rect 28612 29466 28623 29512
rect 28555 29455 28623 29466
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 70813 29452 71000 29510
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
rect 28687 29380 28755 29391
rect 28687 29334 28698 29380
rect 28744 29334 28755 29380
rect 28687 29323 28755 29334
rect 70813 29348 71000 29406
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
rect 28819 29248 28887 29259
rect 28819 29202 28830 29248
rect 28876 29202 28887 29248
rect 28819 29191 28887 29202
rect 70813 29244 71000 29302
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 70813 29140 71000 29198
rect 28951 29116 29019 29127
rect 28951 29070 28962 29116
rect 29008 29070 29019 29116
rect 28951 29059 29019 29070
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 70813 29036 71000 29094
rect 29083 28984 29151 28995
rect 29083 28938 29094 28984
rect 29140 28938 29151 28984
rect 29083 28927 29151 28938
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 70813 28932 71000 28990
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
rect 29215 28852 29283 28863
rect 29215 28806 29226 28852
rect 29272 28806 29283 28852
rect 29215 28795 29283 28806
rect 70813 28828 71000 28886
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29347 28720 29415 28731
rect 29347 28674 29358 28720
rect 29404 28674 29415 28720
rect 29347 28663 29415 28674
rect 70813 28724 71000 28782
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 70813 28620 71000 28678
rect 29479 28588 29547 28599
rect 29479 28542 29490 28588
rect 29536 28542 29547 28588
rect 29479 28531 29547 28542
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 70813 28516 71000 28574
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29611 28456 29679 28467
rect 29611 28410 29622 28456
rect 29668 28410 29679 28456
rect 29611 28399 29679 28410
rect 70813 28412 71000 28470
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
rect 29743 28324 29811 28335
rect 29743 28278 29754 28324
rect 29800 28278 29811 28324
rect 29743 28267 29811 28278
rect 70813 28308 71000 28366
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 70813 28204 71000 28262
rect 29875 28192 29943 28203
rect 29875 28146 29886 28192
rect 29932 28146 29943 28192
rect 29875 28135 29943 28146
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 70813 28100 71000 28158
rect 30007 28060 30075 28071
rect 30007 28014 30018 28060
rect 30064 28014 30075 28060
rect 30007 28003 30075 28014
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 70813 27996 71000 28054
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30139 27928 30207 27939
rect 30139 27882 30150 27928
rect 30196 27882 30207 27928
rect 30139 27871 30207 27882
rect 70813 27892 71000 27950
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
rect 30271 27796 30339 27807
rect 30271 27750 30282 27796
rect 30328 27750 30339 27796
rect 30271 27739 30339 27750
rect 70813 27788 71000 27846
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 70813 27684 71000 27742
rect 30403 27664 30471 27675
rect 30403 27618 30414 27664
rect 30460 27618 30471 27664
rect 30403 27607 30471 27618
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 70813 27580 71000 27638
rect 30535 27532 30603 27543
rect 30535 27486 30546 27532
rect 30592 27486 30603 27532
rect 30535 27475 30603 27486
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 70813 27476 71000 27534
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
rect 30667 27400 30735 27411
rect 30667 27354 30678 27400
rect 30724 27354 30735 27400
rect 30667 27343 30735 27354
rect 70813 27372 71000 27430
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 30799 27268 30867 27279
rect 30799 27222 30810 27268
rect 30856 27222 30867 27268
rect 30799 27211 30867 27222
rect 70813 27268 71000 27326
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
rect 70813 27164 71000 27222
rect 30931 27136 30999 27147
rect 30931 27090 30942 27136
rect 30988 27090 30999 27136
rect 30931 27079 30999 27090
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 70813 27060 71000 27118
rect 31063 27004 31131 27015
rect 31063 26958 31074 27004
rect 31120 26958 31131 27004
rect 31063 26947 31131 26958
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 70813 26956 71000 27014
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
rect 31195 26872 31263 26883
rect 31195 26826 31206 26872
rect 31252 26826 31263 26872
rect 31195 26815 31263 26826
rect 70813 26852 71000 26910
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31327 26740 31395 26751
rect 31327 26694 31338 26740
rect 31384 26694 31395 26740
rect 31327 26683 31395 26694
rect 70813 26748 71000 26806
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 70813 26644 71000 26702
rect 31459 26608 31527 26619
rect 31459 26562 31470 26608
rect 31516 26562 31527 26608
rect 31459 26551 31527 26562
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 70813 26540 71000 26598
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31591 26476 31659 26487
rect 31591 26430 31602 26476
rect 31648 26430 31659 26476
rect 31591 26419 31659 26430
rect 70813 26436 71000 26494
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
rect 31723 26344 31791 26355
rect 31723 26298 31734 26344
rect 31780 26298 31791 26344
rect 31723 26287 31791 26298
rect 70813 26332 71000 26390
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
rect 70813 26228 71000 26286
rect 31855 26212 31923 26223
rect 31855 26166 31866 26212
rect 31912 26166 31923 26212
rect 31855 26155 31923 26166
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 70813 26124 71000 26182
rect 31987 26080 32055 26091
rect 31987 26034 31998 26080
rect 32044 26034 32055 26080
rect 31987 26023 32055 26034
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 70813 26020 71000 26078
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32119 25948 32187 25959
rect 32119 25902 32130 25948
rect 32176 25902 32187 25948
rect 32119 25891 32187 25902
rect 70813 25916 71000 25974
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
rect 32251 25816 32319 25827
rect 32251 25770 32262 25816
rect 32308 25770 32319 25816
rect 32251 25759 32319 25770
rect 70813 25812 71000 25870
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 70813 25708 71000 25766
rect 32383 25684 32451 25695
rect 32383 25638 32394 25684
rect 32440 25638 32451 25684
rect 32383 25627 32451 25638
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 70813 25604 71000 25662
rect 32515 25552 32583 25563
rect 32515 25506 32526 25552
rect 32572 25506 32583 25552
rect 32515 25495 32583 25506
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 70813 25500 71000 25558
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32647 25420 32715 25431
rect 32647 25374 32658 25420
rect 32704 25374 32715 25420
rect 32647 25363 32715 25374
rect 70813 25396 71000 25454
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 32779 25288 32847 25299
rect 32779 25242 32790 25288
rect 32836 25242 32847 25288
rect 32779 25231 32847 25242
rect 70813 25292 71000 25350
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 70813 25188 71000 25246
rect 32911 25156 32979 25167
rect 32911 25110 32922 25156
rect 32968 25110 32979 25156
rect 32911 25099 32979 25110
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 70813 25084 71000 25142
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 33043 25024 33111 25035
rect 33043 24978 33054 25024
rect 33100 24978 33111 25024
rect 33043 24967 33111 24978
rect 70813 24980 71000 25038
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
rect 33175 24892 33243 24903
rect 33175 24846 33186 24892
rect 33232 24846 33243 24892
rect 33175 24835 33243 24846
rect 70813 24876 71000 24934
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 70813 24772 71000 24830
rect 33307 24760 33375 24771
rect 33307 24714 33318 24760
rect 33364 24714 33375 24760
rect 33307 24703 33375 24714
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 70813 24668 71000 24726
rect 33439 24628 33507 24639
rect 33439 24582 33450 24628
rect 33496 24582 33507 24628
rect 33439 24571 33507 24582
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 70813 24564 71000 24622
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
rect 33571 24496 33639 24507
rect 33571 24450 33582 24496
rect 33628 24450 33639 24496
rect 33571 24439 33639 24450
rect 70813 24460 71000 24518
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
rect 33703 24364 33771 24375
rect 33703 24318 33714 24364
rect 33760 24318 33771 24364
rect 33703 24307 33771 24318
rect 70813 24356 71000 24414
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 70813 24252 71000 24310
rect 33835 24232 33903 24243
rect 33835 24186 33846 24232
rect 33892 24186 33903 24232
rect 33835 24175 33903 24186
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 70813 24148 71000 24206
rect 33967 24100 34035 24111
rect 33967 24054 33978 24100
rect 34024 24054 34035 24100
rect 33967 24043 34035 24054
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 70813 24044 71000 24102
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
rect 34099 23968 34167 23979
rect 34099 23922 34110 23968
rect 34156 23922 34167 23968
rect 34099 23911 34167 23922
rect 70813 23940 71000 23998
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
rect 34231 23836 34299 23847
rect 34231 23790 34242 23836
rect 34288 23790 34299 23836
rect 34231 23779 34299 23790
rect 70813 23836 71000 23894
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 70813 23732 71000 23790
rect 34363 23704 34431 23715
rect 34363 23658 34374 23704
rect 34420 23658 34431 23704
rect 34363 23647 34431 23658
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 70813 23628 71000 23686
rect 34495 23572 34563 23583
rect 34495 23526 34506 23572
rect 34552 23526 34563 23572
rect 34495 23515 34563 23526
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 70813 23524 71000 23582
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34627 23440 34695 23451
rect 34627 23394 34638 23440
rect 34684 23394 34695 23440
rect 34627 23383 34695 23394
rect 70813 23420 71000 23478
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
rect 34759 23308 34827 23319
rect 34759 23262 34770 23308
rect 34816 23262 34827 23308
rect 34759 23251 34827 23262
rect 70813 23316 71000 23374
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 70813 23212 71000 23270
rect 34891 23176 34959 23187
rect 34891 23130 34902 23176
rect 34948 23130 34959 23176
rect 34891 23119 34959 23130
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 70813 23108 71000 23166
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 35023 23044 35091 23055
rect 35023 22998 35034 23044
rect 35080 22998 35091 23044
rect 35023 22987 35091 22998
rect 70813 23004 71000 23062
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
rect 35155 22912 35223 22923
rect 35155 22866 35166 22912
rect 35212 22866 35223 22912
rect 35155 22855 35223 22866
rect 70813 22900 71000 22958
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 70813 22796 71000 22854
rect 35287 22780 35355 22791
rect 35287 22734 35298 22780
rect 35344 22734 35355 22780
rect 35287 22723 35355 22734
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 70813 22692 71000 22750
rect 35419 22648 35487 22659
rect 35419 22602 35430 22648
rect 35476 22602 35487 22648
rect 35419 22591 35487 22602
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 70813 22588 71000 22646
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
rect 35551 22516 35619 22527
rect 35551 22470 35562 22516
rect 35608 22470 35619 22516
rect 35551 22459 35619 22470
rect 70813 22484 71000 22542
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
rect 35683 22384 35751 22395
rect 35683 22338 35694 22384
rect 35740 22338 35751 22384
rect 35683 22327 35751 22338
rect 70813 22380 71000 22438
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
rect 70813 22276 71000 22334
rect 35815 22252 35883 22263
rect 35815 22206 35826 22252
rect 35872 22206 35883 22252
rect 35815 22195 35883 22206
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 70813 22172 71000 22230
rect 35947 22120 36015 22131
rect 35947 22074 35958 22120
rect 36004 22074 36015 22120
rect 35947 22063 36015 22074
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 70813 22068 71000 22126
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
rect 36079 21988 36147 21999
rect 36079 21942 36090 21988
rect 36136 21942 36147 21988
rect 36079 21931 36147 21942
rect 70813 21964 71000 22022
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36211 21856 36279 21867
rect 36211 21810 36222 21856
rect 36268 21810 36279 21856
rect 36211 21799 36279 21810
rect 70813 21860 71000 21918
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 70813 21756 71000 21814
rect 36343 21724 36411 21735
rect 36343 21678 36354 21724
rect 36400 21678 36411 21724
rect 36343 21667 36411 21678
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 70813 21652 71000 21710
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36475 21592 36543 21603
rect 36475 21546 36486 21592
rect 36532 21546 36543 21592
rect 36475 21535 36543 21546
rect 70813 21548 71000 21606
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
rect 36607 21460 36675 21471
rect 36607 21414 36618 21460
rect 36664 21414 36675 21460
rect 36607 21403 36675 21414
rect 70813 21444 71000 21502
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
rect 70813 21340 71000 21398
rect 36739 21328 36807 21339
rect 36739 21282 36750 21328
rect 36796 21282 36807 21328
rect 36739 21271 36807 21282
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 70813 21236 71000 21294
rect 36871 21196 36939 21207
rect 36871 21150 36882 21196
rect 36928 21150 36939 21196
rect 36871 21139 36939 21150
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 70813 21132 71000 21190
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 37003 21064 37071 21075
rect 37003 21018 37014 21064
rect 37060 21018 37071 21064
rect 37003 21007 37071 21018
rect 70813 21028 71000 21086
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
rect 37135 20932 37203 20943
rect 37135 20886 37146 20932
rect 37192 20886 37203 20932
rect 37135 20875 37203 20886
rect 70813 20924 71000 20982
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 70813 20820 71000 20878
rect 37267 20800 37335 20811
rect 37267 20754 37278 20800
rect 37324 20754 37335 20800
rect 37267 20743 37335 20754
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 70813 20716 71000 20774
rect 37399 20668 37467 20679
rect 37399 20622 37410 20668
rect 37456 20622 37467 20668
rect 37399 20611 37467 20622
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 70813 20612 71000 20670
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37531 20536 37599 20547
rect 37531 20490 37542 20536
rect 37588 20490 37599 20536
rect 37531 20479 37599 20490
rect 70813 20508 71000 20566
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 37663 20404 37731 20415
rect 37663 20358 37674 20404
rect 37720 20358 37731 20404
rect 37663 20347 37731 20358
rect 70813 20404 71000 20462
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
rect 70813 20300 71000 20358
rect 37795 20272 37863 20283
rect 37795 20226 37806 20272
rect 37852 20226 37863 20272
rect 37795 20215 37863 20226
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 70813 20196 71000 20254
rect 37927 20140 37995 20151
rect 37927 20094 37938 20140
rect 37984 20094 37995 20140
rect 37927 20083 37995 20094
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 70813 20092 71000 20150
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
rect 38059 20008 38127 20019
rect 38059 19962 38070 20008
rect 38116 19962 38127 20008
rect 38059 19951 38127 19962
rect 70813 19988 71000 20046
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 38191 19876 38259 19887
rect 38191 19830 38202 19876
rect 38248 19830 38259 19876
rect 38191 19819 38259 19830
rect 70813 19884 71000 19942
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 70813 19780 71000 19838
rect 38323 19744 38391 19755
rect 38323 19698 38334 19744
rect 38380 19698 38391 19744
rect 38323 19687 38391 19698
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 70813 19676 71000 19734
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38455 19612 38523 19623
rect 38455 19566 38466 19612
rect 38512 19566 38523 19612
rect 38455 19555 38523 19566
rect 70813 19572 71000 19630
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
rect 38587 19480 38655 19491
rect 38587 19434 38598 19480
rect 38644 19434 38655 19480
rect 38587 19423 38655 19434
rect 70813 19468 71000 19526
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 70813 19364 71000 19422
rect 38719 19348 38787 19359
rect 38719 19302 38730 19348
rect 38776 19302 38787 19348
rect 38719 19291 38787 19302
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 70813 19260 71000 19318
rect 38851 19216 38919 19227
rect 38851 19170 38862 19216
rect 38908 19170 38919 19216
rect 38851 19159 38919 19170
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 70813 19156 71000 19214
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 38983 19084 39051 19095
rect 38983 19038 38994 19084
rect 39040 19038 39051 19084
rect 38983 19027 39051 19038
rect 70813 19052 71000 19110
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 39115 18952 39183 18963
rect 39115 18906 39126 18952
rect 39172 18906 39183 18952
rect 39115 18895 39183 18906
rect 70813 18948 71000 19006
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 70813 18844 71000 18902
rect 39247 18820 39315 18831
rect 39247 18774 39258 18820
rect 39304 18774 39315 18820
rect 39247 18763 39315 18774
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 70813 18740 71000 18798
rect 39379 18688 39447 18699
rect 39379 18642 39390 18688
rect 39436 18642 39447 18688
rect 39379 18631 39447 18642
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 70813 18636 71000 18694
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39511 18556 39579 18567
rect 39511 18510 39522 18556
rect 39568 18510 39579 18556
rect 39511 18499 39579 18510
rect 70813 18532 71000 18590
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39643 18424 39711 18435
rect 39643 18378 39654 18424
rect 39700 18378 39711 18424
rect 39643 18367 39711 18378
rect 70813 18428 71000 18486
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 70813 18324 71000 18382
rect 39775 18292 39843 18303
rect 39775 18246 39786 18292
rect 39832 18246 39843 18292
rect 39775 18235 39843 18246
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 70813 18220 71000 18278
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39907 18160 39975 18171
rect 39907 18114 39918 18160
rect 39964 18114 39975 18160
rect 39907 18103 39975 18114
rect 70813 18116 71000 18174
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
rect 40039 18028 40107 18039
rect 40039 17982 40050 18028
rect 40096 17982 40107 18028
rect 40039 17971 40107 17982
rect 70813 18012 71000 18070
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 70813 17908 71000 17966
rect 40171 17896 40239 17907
rect 40171 17850 40182 17896
rect 40228 17850 40239 17896
rect 40171 17839 40239 17850
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 70813 17804 71000 17862
rect 40303 17764 40371 17775
rect 40303 17718 40314 17764
rect 40360 17718 40371 17764
rect 40303 17707 40371 17718
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 70813 17700 71000 17758
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
rect 40435 17632 40503 17643
rect 40435 17586 40446 17632
rect 40492 17586 40503 17632
rect 40435 17575 40503 17586
rect 70813 17596 71000 17654
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40567 17500 40635 17511
rect 40567 17454 40578 17500
rect 40624 17454 40635 17500
rect 40567 17443 40635 17454
rect 70813 17492 71000 17550
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 70813 17388 71000 17446
rect 40699 17368 40767 17379
rect 40699 17322 40710 17368
rect 40756 17322 40767 17368
rect 40699 17311 40767 17322
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 70813 17284 71000 17342
rect 40831 17236 40899 17247
rect 40831 17190 40842 17236
rect 40888 17190 40899 17236
rect 40831 17179 40899 17190
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 70813 17180 71000 17238
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
rect 40963 17104 41031 17115
rect 40963 17058 40974 17104
rect 41020 17058 41031 17104
rect 40963 17047 41031 17058
rect 70813 17076 71000 17134
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 41095 16972 41163 16983
rect 41095 16926 41106 16972
rect 41152 16926 41163 16972
rect 41095 16915 41163 16926
rect 70813 16972 71000 17030
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
rect 70813 16868 71000 16926
rect 41227 16840 41295 16851
rect 41227 16794 41238 16840
rect 41284 16794 41295 16840
rect 41227 16783 41295 16794
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 70813 16764 71000 16822
rect 41359 16708 41427 16719
rect 41359 16662 41370 16708
rect 41416 16662 41427 16708
rect 41359 16651 41427 16662
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 70813 16660 71000 16718
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41491 16576 41559 16587
rect 41491 16530 41502 16576
rect 41548 16530 41559 16576
rect 41491 16519 41559 16530
rect 70813 16556 71000 16614
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
rect 41623 16444 41691 16455
rect 41623 16398 41634 16444
rect 41680 16398 41691 16444
rect 41623 16387 41691 16398
rect 70813 16452 71000 16510
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 70813 16348 71000 16406
rect 41755 16312 41823 16323
rect 41755 16266 41766 16312
rect 41812 16266 41823 16312
rect 41755 16255 41823 16266
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 70813 16244 71000 16302
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41887 16180 41955 16191
rect 41887 16134 41898 16180
rect 41944 16134 41955 16180
rect 41887 16123 41955 16134
rect 70813 16140 71000 16198
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
rect 42019 16048 42087 16059
rect 42019 16002 42030 16048
rect 42076 16002 42087 16048
rect 42019 15991 42087 16002
rect 70813 16036 71000 16094
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 70813 15932 71000 15990
rect 42151 15916 42219 15927
rect 42151 15870 42162 15916
rect 42208 15870 42219 15916
rect 42151 15859 42219 15870
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 70813 15828 71000 15886
rect 42283 15784 42351 15795
rect 42283 15738 42294 15784
rect 42340 15738 42351 15784
rect 42283 15727 42351 15738
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 70813 15724 71000 15782
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42415 15652 42483 15663
rect 42415 15606 42426 15652
rect 42472 15606 42483 15652
rect 42415 15595 42483 15606
rect 70813 15620 71000 15678
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42547 15520 42615 15531
rect 42547 15474 42558 15520
rect 42604 15474 42615 15520
rect 42547 15463 42615 15474
rect 70813 15516 71000 15574
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 70813 15412 71000 15470
rect 42679 15388 42747 15399
rect 42679 15342 42690 15388
rect 42736 15342 42747 15388
rect 42679 15331 42747 15342
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 70813 15308 71000 15366
rect 42811 15256 42879 15267
rect 42811 15210 42822 15256
rect 42868 15210 42879 15256
rect 42811 15199 42879 15210
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 70813 15204 71000 15262
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
rect 42943 15124 43011 15135
rect 42943 15078 42954 15124
rect 43000 15078 43011 15124
rect 42943 15067 43011 15078
rect 70813 15100 71000 15158
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
rect 43075 14992 43143 15003
rect 43075 14946 43086 14992
rect 43132 14946 43143 14992
rect 43075 14935 43143 14946
rect 70813 14996 71000 15054
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 70813 14892 71000 14950
rect 43207 14860 43275 14871
rect 43207 14814 43218 14860
rect 43264 14814 43275 14860
rect 43207 14803 43275 14814
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 70813 14788 71000 14846
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 43339 14728 43407 14739
rect 43339 14682 43350 14728
rect 43396 14682 43407 14728
rect 43339 14671 43407 14682
rect 70813 14684 71000 14742
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
rect 43471 14596 43539 14607
rect 43471 14550 43482 14596
rect 43528 14550 43539 14596
rect 43471 14539 43539 14550
rect 70813 14580 71000 14638
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 70813 14476 71000 14534
rect 43603 14464 43671 14475
rect 43603 14418 43614 14464
rect 43660 14418 43671 14464
rect 43603 14407 43671 14418
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 70813 14372 71000 14430
rect 43735 14332 43803 14343
rect 43735 14286 43746 14332
rect 43792 14286 43803 14332
rect 43735 14275 43803 14286
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 70813 14268 71000 14326
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
rect 43867 14200 43935 14211
rect 43867 14154 43878 14200
rect 43924 14154 43935 14200
rect 43867 14143 43935 14154
rect 70813 14164 71000 14222
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 43999 14068 44067 14079
rect 43999 14022 44010 14068
rect 44056 14022 44067 14068
rect 43999 14011 44067 14022
rect 70813 14060 71000 14118
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 70813 13956 71000 14014
rect 44131 13936 44199 13947
rect 44131 13890 44142 13936
rect 44188 13890 44199 13936
rect 44131 13879 44199 13890
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 70813 13852 71000 13910
rect 44263 13804 44331 13815
rect 44263 13758 44274 13804
rect 44320 13758 44331 13804
rect 44263 13747 44331 13758
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 70813 13748 71000 13806
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44395 13672 44463 13683
rect 44395 13626 44406 13672
rect 44452 13626 44463 13672
rect 44395 13615 44463 13626
rect 70813 13644 71000 13702
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44527 13540 44595 13551
rect 44527 13494 44538 13540
rect 44584 13494 44595 13540
rect 44527 13483 44595 13494
rect 70813 13540 71000 13598
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 70813 13436 71000 13494
rect 44659 13408 44727 13419
rect 44659 13362 44670 13408
rect 44716 13362 44727 13408
rect 44659 13351 44727 13362
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 70813 13280 71000 13390
rect 45077 13269 71000 13280
rect 44839 13256 44907 13267
rect 44839 13210 44850 13256
rect 44896 13210 44907 13256
rect 44839 13199 44907 13210
rect 45077 13223 45088 13269
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 45077 13165 71000 13223
rect 45077 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 45077 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47111 17000 71000
rect 17200 48447 20200 71000
rect 20400 49773 23400 71000
rect 23600 50451 25000 71000
rect 25200 51120 26600 71000
rect 26800 52512 29800 71000
rect 30000 53791 33000 71000
rect 33200 55312 36200 71000
rect 36400 56464 39400 71000
rect 39600 57138 41000 71000
rect 41200 57810 42600 71000
rect 42800 59140 45800 71000
rect 46000 60508 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63320 55400 71000
rect 55600 63836 57000 71000
rect 57200 64540 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68200 68200 71000
tri 68200 68200 68693 68693 sw
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66800 68029 66884 68113 ne
rect 66884 68029 70613 68113
tri 66600 67829 66800 68029 sw
tri 66884 67829 67084 68029 ne
rect 67084 67829 70613 68029
rect 65200 67650 66800 67829
tri 66800 67650 66979 67829 sw
tri 67084 67650 67263 67829 ne
rect 67263 67650 70613 67829
rect 65200 67449 66979 67650
tri 65200 67366 65283 67449 ne
rect 65283 67366 66979 67449
tri 66979 67366 67263 67650 sw
tri 67263 67366 67547 67650 ne
rect 67547 67366 70613 67650
tri 65000 67166 65200 67366 sw
tri 65283 67166 65483 67366 ne
rect 65483 67264 67263 67366
tri 67263 67264 67365 67366 sw
tri 67547 67264 67649 67366 ne
rect 67649 67264 70613 67366
rect 65483 67166 67365 67264
rect 63600 66980 65200 67166
tri 65200 66980 65386 67166 sw
tri 65483 66980 65669 67166 ne
rect 65669 66980 67365 67166
tri 67365 66980 67649 67264 sw
tri 67649 66980 67933 67264 ne
rect 67933 66980 70613 67264
rect 63600 66906 65386 66980
tri 65386 66906 65460 66980 sw
tri 65669 66906 65743 66980 ne
rect 65743 66906 67649 66980
tri 67649 66906 67723 66980 sw
tri 67933 66906 68007 66980 ne
rect 68007 66916 70613 66980
rect 70669 66916 71000 68116
rect 68007 66906 71000 66916
rect 63600 66786 65460 66906
tri 63600 66694 63692 66786 ne
rect 63692 66694 65460 66786
tri 65460 66694 65672 66906 sw
tri 65743 66694 65955 66906 ne
rect 65955 66800 67723 66906
tri 67723 66800 67829 66906 sw
tri 68007 66800 68113 66906 ne
rect 68113 66800 71000 66906
rect 65955 66694 67829 66800
tri 67829 66694 67935 66800 sw
tri 63400 66494 63600 66694 sw
tri 63692 66494 63892 66694 ne
rect 63892 66494 65672 66694
rect 62000 66323 63600 66494
tri 63600 66323 63771 66494 sw
tri 63892 66323 64063 66494 ne
rect 64063 66411 65672 66494
tri 65672 66411 65955 66694 sw
tri 65955 66411 66238 66694 ne
rect 66238 66600 67935 66694
tri 67935 66600 68029 66694 sw
rect 66238 66411 71000 66600
rect 64063 66332 65955 66411
tri 65955 66332 66034 66411 sw
tri 66238 66332 66317 66411 ne
rect 66317 66332 71000 66411
rect 64063 66323 66034 66332
rect 62000 66114 63771 66323
tri 62000 66031 62083 66114 ne
rect 62083 66031 63771 66114
tri 63771 66031 64063 66323 sw
tri 64063 66031 64355 66323 ne
rect 64355 66049 66034 66323
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64355 66031 66317 66049
tri 66317 66031 66335 66049 sw
tri 66600 66031 66618 66049 ne
rect 66618 66031 71000 66049
tri 61800 65831 62000 66031 sw
tri 62083 65831 62283 66031 ne
rect 62283 65831 64063 66031
rect 60400 65760 62000 65831
tri 62000 65760 62071 65831 sw
tri 62283 65760 62354 65831 ne
rect 62354 65760 64063 65831
tri 64063 65760 64334 66031 sw
tri 64355 65760 64626 66031 ne
rect 64626 65766 66335 66031
tri 66335 65766 66600 66031 sw
tri 66618 65766 66883 66031 ne
rect 66883 65766 71000 66031
rect 64626 65760 66600 65766
tri 66600 65760 66606 65766 sw
tri 66883 65760 66889 65766 ne
rect 66889 65760 71000 65766
rect 60400 65649 62071 65760
tri 62071 65649 62182 65760 sw
tri 62354 65649 62465 65760 ne
rect 62465 65672 64334 65760
tri 64334 65672 64422 65760 sw
tri 64626 65672 64714 65760 ne
rect 64714 65672 66606 65760
rect 62465 65649 64422 65672
rect 60400 65451 62182 65649
tri 60400 65366 60485 65451 ne
rect 60485 65366 62182 65451
tri 62182 65366 62465 65649 sw
tri 62465 65380 62734 65649 ne
rect 62734 65380 64422 65649
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65663 66606 65672
tri 66606 65663 66703 65760 sw
tri 66889 65663 66986 65760 ne
rect 66986 65663 71000 65760
rect 65006 65380 66703 65663
tri 66703 65380 66986 65663 sw
tri 66986 65380 67269 65663 ne
rect 67269 65380 71000 65663
tri 62734 65366 62748 65380 ne
rect 62748 65366 64714 65380
tri 64714 65366 64728 65380 sw
tri 65006 65366 65020 65380 ne
rect 65020 65366 66986 65380
tri 66986 65366 67000 65380 sw
tri 67269 65366 67283 65380 ne
rect 67283 65366 71000 65380
tri 60200 65166 60400 65366 sw
tri 60485 65166 60685 65366 ne
rect 60685 65166 62465 65366
rect 58800 64984 60400 65166
tri 60400 64984 60582 65166 sw
tri 60685 64984 60867 65166 ne
rect 60867 65083 62465 65166
tri 62465 65083 62748 65366 sw
tri 62748 65083 63031 65366 ne
rect 63031 65292 64728 65366
tri 64728 65292 64802 65366 sw
tri 65020 65292 65094 65366 ne
rect 65094 65292 67000 65366
rect 63031 65083 64802 65292
rect 60867 64997 62748 65083
tri 62748 64997 62834 65083 sw
tri 63031 64997 63117 65083 ne
rect 63117 65000 64802 65083
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 67000 65292
tri 67000 65200 67166 65366 sw
tri 67283 65200 67449 65366 ne
rect 67449 65200 71000 65366
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60867 64984 62834 64997
rect 58800 64786 60582 64984
tri 58800 64699 58887 64786 ne
rect 58887 64699 60582 64786
tri 60582 64699 60867 64984 sw
tri 60867 64699 61152 64984 ne
rect 61152 64714 62834 64984
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61152 64699 63117 64714
tri 63117 64699 63132 64714 sw
tri 63400 64699 63415 64714 ne
rect 63415 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63415 64699 65386 64708
tri 65386 64699 65395 64708 sw
tri 65678 64699 65687 64708 ne
rect 65687 64699 71000 64708
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60867 64699
tri 60867 64540 61026 64699 sw
tri 61152 64540 61311 64699 ne
rect 61311 64540 63132 64699
tri 63132 64540 63291 64699 sw
tri 63415 64540 63574 64699 ne
rect 63574 64540 65395 64699
tri 65395 64540 65554 64699 sw
tri 65687 64540 65846 64699 ne
rect 65846 64540 71000 64699
rect 57200 64499 58759 64540
tri 58759 64499 58800 64540 sw
tri 59046 64499 59087 64540 ne
rect 59087 64499 61026 64540
rect 57200 64323 58800 64499
tri 58800 64323 58976 64499 sw
tri 59087 64323 59263 64499 ne
rect 59263 64445 61026 64499
tri 61026 64445 61121 64540 sw
tri 61311 64445 61406 64540 ne
rect 61406 64445 63291 64540
rect 59263 64323 61121 64445
rect 57200 64119 58976 64323
tri 57200 64036 57283 64119 ne
rect 57283 64036 58976 64119
tri 58976 64036 59263 64323 sw
tri 59263 64160 59426 64323 ne
rect 59426 64160 61121 64323
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63291 64445
tri 63291 64431 63400 64540 sw
tri 63574 64431 63683 64540 ne
rect 63683 64452 65554 64540
tri 65554 64452 65642 64540 sw
tri 65846 64452 65934 64540 ne
rect 65934 64452 71000 64540
rect 63683 64431 65642 64452
rect 61691 64160 63400 64431
tri 63400 64160 63671 64431 sw
tri 63683 64160 63954 64431 ne
rect 63954 64160 65642 64431
tri 65642 64160 65934 64452 sw
tri 65934 64160 66226 64452 ne
rect 66226 64160 71000 64452
tri 59426 64036 59550 64160 ne
rect 59550 64036 61406 64160
tri 61406 64036 61530 64160 sw
tri 61691 64036 61815 64160 ne
rect 61815 64036 63671 64160
tri 63671 64036 63795 64160 sw
tri 63954 64036 64078 64160 ne
rect 64078 64036 65934 64160
tri 65934 64036 66058 64160 sw
tri 66226 64036 66350 64160 ne
rect 66350 64036 71000 64160
tri 57000 63836 57200 64036 sw
tri 57283 63836 57483 64036 ne
rect 57483 63836 59263 64036
rect 55600 63656 57200 63836
tri 57200 63656 57380 63836 sw
tri 57483 63656 57663 63836 ne
rect 57663 63749 59263 63836
tri 59263 63749 59550 64036 sw
tri 59550 63749 59837 64036 ne
rect 59837 63780 61530 64036
tri 61530 63780 61786 64036 sw
tri 61815 63780 62071 64036 ne
rect 62071 63780 63795 64036
tri 63795 63780 64051 64036 sw
tri 64078 63780 64334 64036 ne
rect 64334 63780 66058 64036
tri 66058 63780 66314 64036 sw
tri 66350 63780 66606 64036 ne
rect 66606 63780 71000 64036
rect 59837 63749 61786 63780
rect 57663 63673 59550 63749
tri 59550 63673 59626 63749 sw
tri 59837 63673 59913 63749 ne
rect 59913 63673 61786 63749
rect 57663 63656 59626 63673
rect 55600 63456 57380 63656
tri 55600 63373 55683 63456 ne
rect 55683 63373 57380 63456
tri 57380 63373 57663 63656 sw
tri 57663 63373 57946 63656 ne
rect 57946 63386 59626 63656
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 64051 63780
tri 64051 63683 64148 63780 sw
tri 64334 63683 64431 63780 ne
rect 64431 63683 66314 63780
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 57946 63373 59913 63386
tri 59913 63373 59926 63386 sw
tri 60200 63373 60213 63386 ne
rect 60213 63373 62071 63386
tri 62071 63373 62193 63495 sw
tri 62356 63373 62478 63495 ne
rect 62478 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66314 63683
tri 66314 63600 66494 63780 sw
tri 66606 63600 66786 63780 ne
rect 66786 63600 71000 63780
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62478 63373 64431 63400
tri 64431 63373 64458 63400 sw
tri 64714 63373 64741 63400 ne
rect 64741 63373 71000 63400
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57663 63373
tri 57663 63320 57716 63373 sw
tri 57946 63320 57999 63373 ne
rect 57999 63320 59926 63373
tri 59926 63320 59979 63373 sw
tri 60213 63320 60266 63373 ne
rect 60266 63320 62193 63373
tri 62193 63320 62246 63373 sw
tri 62478 63320 62531 63373 ne
rect 62531 63320 64458 63373
tri 64458 63320 64511 63373 sw
tri 64741 63320 64794 63373 ne
rect 64794 63320 71000 63373
rect 54000 63173 55453 63320
tri 55453 63173 55600 63320 sw
tri 55736 63173 55883 63320 ne
rect 55883 63223 57716 63320
tri 57716 63223 57813 63320 sw
tri 57999 63223 58096 63320 ne
rect 58096 63223 59979 63320
rect 55883 63173 57813 63223
rect 54000 62990 55600 63173
tri 55600 62990 55783 63173 sw
tri 55883 62990 56066 63173 ne
rect 56066 62990 57813 63173
rect 54000 62793 55783 62990
tri 54000 62707 54086 62793 ne
rect 54086 62707 55783 62793
tri 55783 62707 56066 62990 sw
tri 56066 62940 56116 62990 ne
rect 56116 62940 57813 62990
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59979 63223
tri 59979 63099 60200 63320 sw
tri 60266 63099 60487 63320 ne
rect 60487 63225 62246 63320
tri 62246 63225 62341 63320 sw
tri 62531 63225 62626 63320 ne
rect 62626 63225 64511 63320
rect 60487 63099 62341 63225
rect 58379 62940 60200 63099
tri 60200 62940 60359 63099 sw
tri 60487 62940 60646 63099 ne
rect 60646 62940 62341 63099
tri 62341 62940 62626 63225 sw
tri 62626 62940 62911 63225 ne
rect 62911 63117 64511 63225
tri 64511 63117 64714 63320 sw
tri 64794 63117 64997 63320 ne
rect 64997 63117 71000 63320
rect 62911 62940 64714 63117
tri 64714 62940 64891 63117 sw
tri 64997 62940 65174 63117 ne
rect 65174 62940 71000 63117
tri 56116 62707 56349 62940 ne
rect 56349 62707 58096 62940
tri 58096 62707 58329 62940 sw
tri 58379 62707 58612 62940 ne
rect 58612 62707 60359 62940
tri 60359 62707 60592 62940 sw
tri 60646 62707 60879 62940 ne
rect 60879 62707 62626 62940
tri 62626 62707 62859 62940 sw
tri 62911 62707 63144 62940 ne
rect 63144 62707 64891 62940
tri 64891 62707 65124 62940 sw
tri 65174 62707 65407 62940 ne
rect 65407 62707 71000 62940
tri 53800 62507 54000 62707 sw
tri 54086 62507 54286 62707 ne
rect 54286 62507 56066 62707
rect 52400 62325 54000 62507
tri 54000 62325 54182 62507 sw
tri 54286 62325 54468 62507 ne
rect 54468 62424 56066 62507
tri 56066 62424 56349 62707 sw
tri 56349 62424 56632 62707 ne
rect 56632 62560 58329 62707
tri 58329 62560 58476 62707 sw
tri 58612 62560 58759 62707 ne
rect 58759 62560 60592 62707
tri 60592 62560 60739 62707 sw
tri 60879 62560 61026 62707 ne
rect 61026 62560 62859 62707
tri 62859 62560 63006 62707 sw
tri 63144 62560 63291 62707 ne
rect 63291 62560 65124 62707
tri 65124 62560 65271 62707 sw
tri 65407 62560 65554 62707 ne
rect 65554 62560 71000 62707
rect 56632 62424 58476 62560
rect 54468 62339 56349 62424
tri 56349 62339 56434 62424 sw
tri 56632 62339 56717 62424 ne
rect 56717 62339 58476 62424
rect 54468 62325 56434 62339
rect 52400 62127 54182 62325
tri 52400 62039 52488 62127 ne
rect 52488 62039 54182 62127
tri 54182 62039 54468 62325 sw
tri 54468 62039 54754 62325 ne
rect 54754 62056 56434 62325
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60739 62560
tri 60739 62467 60832 62560 sw
tri 61026 62467 61119 62560 ne
rect 61119 62467 63006 62560
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54754 62039 56717 62056
tri 56717 62039 56734 62056 sw
tri 57000 62039 57017 62056 ne
rect 57017 62039 58759 62056
tri 58759 62039 58997 62277 sw
tri 59042 62039 59280 62277 ne
rect 59280 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 63006 62467
tri 63006 62465 63101 62560 sw
tri 63291 62465 63386 62560 ne
rect 63386 62465 65271 62560
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62463 65271 62465
tri 65271 62463 65368 62560 sw
tri 65554 62463 65651 62560 ne
rect 65651 62463 71000 62560
rect 63671 62180 65368 62463
tri 65368 62180 65651 62463 sw
tri 65651 62180 65934 62463 ne
rect 65934 62180 71000 62463
rect 59280 62039 61119 62180
tri 61119 62039 61260 62180 sw
tri 61406 62039 61547 62180 ne
rect 61547 62039 63386 62180
tri 63386 62039 63527 62180 sw
tri 63671 62039 63812 62180 ne
rect 63812 62039 65651 62180
tri 65651 62039 65792 62180 sw
tri 65934 62039 66075 62180 ne
rect 66075 62039 71000 62180
tri 52200 61839 52400 62039 sw
tri 52488 61839 52688 62039 ne
rect 52688 62006 54468 62039
tri 54468 62006 54501 62039 sw
tri 54754 62006 54787 62039 ne
rect 54787 62006 56734 62039
rect 52688 61839 54501 62006
rect 50800 61663 52400 61839
tri 52400 61663 52576 61839 sw
tri 52688 61663 52864 61839 ne
rect 52864 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56734 62006
tri 56734 61773 57000 62039 sw
tri 57017 61773 57283 62039 ne
rect 57283 62003 58997 62039
tri 58997 62003 59033 62039 sw
tri 59280 62003 59316 62039 ne
rect 59316 62003 61260 62039
rect 57283 61773 59033 62003
rect 55073 61720 57000 61773
tri 57000 61720 57053 61773 sw
tri 57283 61720 57336 61773 ne
rect 57336 61720 59033 61773
tri 59033 61720 59316 62003 sw
tri 59316 61720 59599 62003 ne
rect 59599 61893 61260 62003
tri 61260 61893 61406 62039 sw
tri 61547 61893 61693 62039 ne
rect 61693 61893 63527 62039
rect 59599 61720 61406 61893
tri 61406 61720 61579 61893 sw
tri 61693 61720 61866 61893 ne
rect 61866 61800 63527 61893
tri 63527 61800 63766 62039 sw
tri 63812 61800 64051 62039 ne
rect 64051 62000 65792 62039
tri 65792 62000 65831 62039 sw
tri 66075 62000 66114 62039 ne
rect 66114 62000 71000 62039
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61866 61720 63766 61800
tri 63766 61720 63846 61800 sw
tri 64051 61720 64131 61800 ne
rect 64131 61720 71000 61800
rect 52864 61663 54787 61720
rect 50800 61459 52576 61663
tri 50800 61375 50884 61459 ne
rect 50884 61375 52576 61459
tri 52576 61375 52864 61663 sw
tri 52864 61375 53152 61663 ne
rect 53152 61661 54787 61663
tri 54787 61661 54846 61720 sw
tri 55073 61661 55132 61720 ne
rect 55132 61661 57053 61720
rect 53152 61375 54846 61661
tri 54846 61375 55132 61661 sw
tri 55132 61375 55418 61661 ne
rect 55418 61658 57053 61661
tri 57053 61658 57115 61720 sw
tri 57336 61658 57398 61720 ne
rect 57398 61658 59316 61720
tri 59316 61658 59378 61720 sw
tri 59599 61658 59661 61720 ne
rect 59661 61662 61579 61720
tri 61579 61662 61637 61720 sw
tri 61866 61662 61924 61720 ne
rect 61924 61662 63846 61720
rect 59661 61658 61637 61662
rect 55418 61375 57115 61658
tri 57115 61375 57398 61658 sw
tri 57398 61375 57681 61658 ne
rect 57681 61375 59378 61658
tri 59378 61375 59661 61658 sw
tri 59661 61375 59944 61658 ne
rect 59944 61375 61637 61658
tri 61637 61375 61924 61662 sw
tri 61924 61375 62211 61662 ne
rect 62211 61515 63846 61662
tri 63846 61515 64051 61720 sw
tri 64131 61515 64336 61720 ne
rect 64336 61515 71000 61720
rect 62211 61375 64051 61515
tri 64051 61375 64191 61515 sw
tri 64336 61375 64476 61515 ne
rect 64476 61375 71000 61515
tri 50600 61175 50800 61375 sw
tri 50884 61175 51084 61375 ne
rect 51084 61175 52864 61375
rect 49200 60992 50800 61175
tri 50800 60992 50983 61175 sw
tri 51084 60992 51267 61175 ne
rect 51267 61087 52864 61175
tri 52864 61087 53152 61375 sw
tri 53152 61087 53440 61375 ne
rect 53440 61340 55132 61375
tri 55132 61340 55167 61375 sw
tri 55418 61340 55453 61375 ne
rect 55453 61340 57398 61375
tri 57398 61340 57433 61375 sw
tri 57681 61340 57716 61375 ne
rect 57716 61340 59661 61375
tri 59661 61340 59696 61375 sw
tri 59944 61340 59979 61375 ne
rect 59979 61340 61924 61375
tri 61924 61340 61959 61375 sw
tri 62211 61340 62246 61375 ne
rect 62246 61340 64191 61375
tri 64191 61340 64226 61375 sw
tri 64476 61340 64511 61375 ne
rect 64511 61340 71000 61375
rect 53440 61087 55167 61340
rect 51267 61015 53152 61087
tri 53152 61015 53224 61087 sw
tri 53440 61015 53512 61087 ne
rect 53512 61054 55167 61087
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57433 61340
tri 57433 61243 57530 61340 sw
tri 57716 61243 57813 61340 ne
rect 57813 61243 59696 61340
tri 59696 61243 59793 61340 sw
tri 59979 61243 60076 61340 ne
rect 60076 61247 61959 61340
tri 61959 61247 62052 61340 sw
tri 62246 61247 62339 61340 ne
rect 62339 61247 64226 61340
rect 60076 61243 62052 61247
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51267 60992 53224 61015
rect 49200 60795 50983 60992
tri 49200 60708 49287 60795 ne
rect 49287 60708 50983 60795
tri 50983 60708 51267 60992 sw
tri 51267 60708 51551 60992 ne
rect 51551 60727 53224 60992
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60994 55453 61015
tri 55453 60994 55513 61054 sw
tri 55739 60994 55799 61054 ne
rect 55799 60994 57530 61054
rect 53800 60727 55513 60994
rect 51551 60708 53512 60727
tri 53512 60708 53531 60727 sw
tri 53800 60708 53819 60727 ne
rect 53819 60708 55513 60727
tri 55513 60708 55799 60994 sw
tri 55799 60708 56085 60994 ne
rect 56085 60960 57530 60994
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 60960 62052 61243
tri 62052 60960 62339 61247 sw
tri 62339 60960 62626 61247 ne
rect 62626 61245 64226 61247
tri 64226 61245 64321 61340 sw
tri 64511 61245 64606 61340 ne
rect 64606 61245 71000 61340
rect 62626 60960 64321 61245
tri 64321 60960 64606 61245 sw
tri 64606 60960 64891 61245 ne
rect 64891 60960 71000 61245
rect 56085 60708 57813 60960
tri 57813 60708 58065 60960 sw
tri 58096 60708 58348 60960 ne
rect 58348 60708 60076 60960
tri 60076 60708 60328 60960 sw
tri 60359 60708 60611 60960 ne
rect 60611 60708 62339 60960
tri 62339 60708 62591 60960 sw
tri 62626 60708 62878 60960 ne
rect 62878 60708 64606 60960
tri 64606 60708 64858 60960 sw
tri 64891 60708 65143 60960 ne
rect 65143 60708 71000 60960
tri 49000 60508 49200 60708 sw
tri 49287 60508 49487 60708 ne
rect 49487 60508 51267 60708
rect 46000 60417 49200 60508
tri 49200 60417 49292 60508 sw
tri 49487 60417 49578 60508 ne
rect 49578 60500 51267 60508
tri 51267 60500 51475 60708 sw
tri 51551 60500 51759 60708 ne
rect 51759 60500 53531 60708
tri 53531 60500 53739 60708 sw
tri 53819 60500 54027 60708 ne
rect 54027 60500 55799 60708
tri 55799 60500 56007 60708 sw
tri 56085 60500 56293 60708 ne
rect 56293 60677 58065 60708
tri 58065 60677 58096 60708 sw
tri 58348 60677 58379 60708 ne
rect 58379 60677 60328 60708
rect 56293 60500 58096 60677
tri 58096 60500 58273 60677 sw
tri 58379 60500 58556 60677 ne
rect 58556 60580 60328 60677
tri 60328 60580 60456 60708 sw
tri 60611 60580 60739 60708 ne
rect 60739 60580 62591 60708
tri 62591 60580 62719 60708 sw
tri 62878 60580 63006 60708 ne
rect 63006 60580 64858 60708
tri 64858 60580 64986 60708 sw
tri 65143 60580 65271 60708 ne
rect 65271 60580 71000 60708
rect 58556 60500 60456 60580
tri 60456 60500 60536 60580 sw
tri 60739 60500 60819 60580 ne
rect 60819 60500 62719 60580
tri 62719 60500 62799 60580 sw
tri 63006 60500 63086 60580 ne
rect 63086 60500 64986 60580
tri 64986 60500 65066 60580 sw
tri 65271 60500 65351 60580 ne
rect 65351 60500 71000 60580
rect 49578 60417 51475 60500
rect 46000 60130 49292 60417
tri 49292 60130 49578 60417 sw
tri 49578 60130 49865 60417 ne
rect 49865 60414 51475 60417
tri 51475 60414 51561 60500 sw
tri 51759 60414 51845 60500 ne
rect 51845 60439 53739 60500
tri 53739 60439 53800 60500 sw
tri 54027 60439 54088 60500 ne
rect 54088 60439 56007 60500
rect 51845 60418 53800 60439
tri 53800 60418 53821 60439 sw
tri 54088 60418 54109 60439 ne
rect 54109 60418 56007 60439
rect 51845 60414 53821 60418
rect 49865 60130 51561 60414
tri 51561 60130 51845 60414 sw
tri 51845 60130 52129 60414 ne
rect 52129 60130 53821 60414
tri 53821 60130 54109 60418 sw
tri 54109 60130 54397 60418 ne
rect 54397 60416 56007 60418
tri 56007 60416 56091 60500 sw
tri 56293 60416 56377 60500 ne
rect 56377 60416 58273 60500
rect 54397 60130 56091 60416
tri 56091 60130 56377 60416 sw
tri 56377 60130 56663 60416 ne
rect 56663 60413 58273 60416
tri 58273 60413 58360 60500 sw
tri 58556 60413 58643 60500 ne
rect 58643 60413 60536 60500
rect 56663 60130 58360 60413
tri 58360 60130 58643 60413 sw
tri 58643 60130 58926 60413 ne
rect 58926 60297 60536 60413
tri 60536 60297 60739 60500 sw
tri 60819 60297 61022 60500 ne
rect 61022 60487 62799 60500
tri 62799 60487 62812 60500 sw
tri 63086 60487 63099 60500 ne
rect 63099 60487 65066 60500
rect 61022 60297 62812 60487
rect 58926 60130 60739 60297
tri 60739 60130 60906 60297 sw
tri 61022 60130 61189 60297 ne
rect 61189 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 65066 60487
tri 65066 60400 65166 60500 sw
tri 65351 60400 65451 60500 ne
rect 65451 60400 71000 60500
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61189 60130 63099 60200
tri 63099 60130 63169 60200 sw
tri 63386 60130 63456 60200 ne
rect 63456 60130 71000 60200
rect 46000 59843 49578 60130
tri 49578 59843 49865 60130 sw
tri 49865 59843 50152 60130 ne
rect 50152 60120 51845 60130
tri 51845 60120 51855 60130 sw
tri 52129 60120 52139 60130 ne
rect 52139 60120 54109 60130
tri 54109 60120 54119 60130 sw
tri 54397 60120 54407 60130 ne
rect 54407 60120 56377 60130
tri 56377 60120 56387 60130 sw
tri 56663 60120 56673 60130 ne
rect 56673 60120 58643 60130
tri 58643 60120 58653 60130 sw
tri 58926 60120 58936 60130 ne
rect 58936 60120 60906 60130
tri 60906 60120 60916 60130 sw
tri 61189 60120 61199 60130 ne
rect 61199 60120 63169 60130
tri 63169 60120 63179 60130 sw
tri 63456 60120 63466 60130 ne
rect 63466 60120 71000 60130
rect 50152 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54119 60120
rect 50152 59843 51916 60059
rect 46000 59682 49865 59843
tri 49865 59682 50027 59843 sw
tri 50152 59682 50313 59843 ne
rect 50313 59775 51916 59843
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54119 60059
tri 54119 60028 54211 60120 sw
tri 54407 60028 54499 60120 ne
rect 54499 60028 56387 60120
rect 52484 59775 54211 60028
rect 50313 59682 52200 59775
rect 46000 59466 50027 59682
tri 46000 59340 46125 59466 ne
rect 46125 59395 50027 59466
tri 50027 59395 50313 59682 sw
tri 50313 59395 50600 59682 ne
rect 50600 59624 52200 59682
tri 52200 59624 52351 59775 sw
tri 52484 59624 52635 59775 ne
rect 52635 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56387 60028
tri 56387 60026 56481 60120 sw
tri 56673 60026 56767 60120 ne
rect 56767 60026 58653 60120
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 60023 58653 60026
tri 58653 60023 58750 60120 sw
tri 58936 60023 59033 60120 ne
rect 59033 60023 60916 60120
tri 60916 60023 61013 60120 sw
tri 61199 60023 61296 60120 ne
rect 61296 60023 63179 60120
rect 57053 59740 58750 60023
tri 58750 59740 59033 60023 sw
tri 59033 59740 59316 60023 ne
rect 59316 59740 61013 60023
tri 61013 59740 61296 60023 sw
tri 61296 59740 61579 60023 ne
rect 61579 59913 63179 60023
tri 63179 59913 63386 60120 sw
tri 63466 59913 63673 60120 ne
rect 63673 59913 70613 60120
rect 61579 59740 63386 59913
tri 63386 59740 63559 59913 sw
tri 63673 59740 63846 59913 ne
rect 63846 59740 70613 59913
rect 52635 59624 54499 59740
rect 50600 59395 52351 59624
rect 46125 59340 50313 59395
tri 50313 59340 50368 59395 sw
tri 50600 59340 50655 59395 ne
rect 50655 59340 52351 59395
tri 52351 59340 52635 59624 sw
tri 52635 59340 52919 59624 ne
rect 52919 59452 54499 59624
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 59033 59740
rect 55075 59452 56861 59646
rect 52919 59340 54787 59452
tri 54787 59340 54899 59452 sw
tri 55075 59340 55187 59452 ne
rect 55187 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 59033 59646
tri 59033 59643 59130 59740 sw
tri 59316 59643 59413 59740 ne
rect 59413 59643 61296 59740
tri 61296 59643 61393 59740 sw
tri 61579 59643 61676 59740 ne
rect 61676 59647 63559 59740
tri 63559 59647 63652 59740 sw
tri 63846 59647 63939 59740 ne
rect 63939 59647 70613 59740
rect 61676 59643 63652 59647
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59360 61393 59643
tri 61393 59360 61676 59643 sw
tri 61676 59360 61959 59643 ne
rect 61959 59360 63652 59643
tri 63652 59360 63939 59647 sw
tri 63939 59360 64226 59647 ne
rect 64226 59360 70613 59647
rect 55187 59340 57147 59360
tri 57147 59340 57167 59360 sw
tri 57433 59340 57453 59360 ne
rect 57453 59340 59413 59360
tri 59413 59340 59433 59360 sw
tri 59696 59340 59716 59360 ne
rect 59716 59340 61676 59360
tri 61676 59340 61696 59360 sw
tri 61959 59340 61979 59360 ne
rect 61979 59340 63939 59360
tri 63939 59340 63959 59360 sw
tri 64226 59340 64246 59360 ne
rect 64246 59340 70613 59360
tri 45800 59140 46000 59340 sw
tri 46125 59140 46325 59340 ne
rect 46325 59140 50368 59340
rect 42800 58910 46000 59140
tri 46000 58910 46230 59140 sw
tri 46325 58910 46556 59140 ne
rect 46556 59108 50368 59140
tri 50368 59108 50600 59340 sw
tri 50655 59108 50887 59340 ne
rect 50887 59194 52635 59340
tri 52635 59194 52781 59340 sw
tri 52919 59194 53065 59340 ne
rect 53065 59198 54899 59340
tri 54899 59198 55041 59340 sw
tri 55187 59198 55329 59340 ne
rect 55329 59198 57167 59340
rect 53065 59194 55041 59198
rect 50887 59108 52781 59194
rect 46556 58910 50600 59108
tri 50600 58910 50798 59108 sw
tri 50887 58910 51085 59108 ne
rect 51085 58910 52781 59108
tri 52781 58910 53065 59194 sw
tri 53065 58910 53349 59194 ne
rect 53349 58910 55041 59194
tri 55041 58910 55329 59198 sw
tri 55329 58910 55617 59198 ne
rect 55617 59074 57167 59198
tri 57167 59074 57433 59340 sw
tri 57453 59074 57719 59340 ne
rect 57719 59263 59433 59340
tri 59433 59263 59510 59340 sw
tri 59716 59263 59793 59340 ne
rect 59793 59263 61696 59340
tri 61696 59263 61773 59340 sw
tri 61979 59263 62056 59340 ne
rect 62056 59267 63959 59340
tri 63959 59267 64032 59340 sw
tri 64246 59267 64319 59340 ne
rect 64319 59267 70613 59340
rect 62056 59263 64032 59267
rect 57719 59074 59510 59263
rect 55617 58910 57433 59074
tri 57433 58910 57597 59074 sw
tri 57719 58910 57883 59074 ne
rect 57883 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 58980 64032 59263
tri 64032 58980 64319 59267 sw
tri 64319 58980 64606 59267 ne
rect 64606 58980 70613 59267
rect 57883 58910 59793 58980
tri 59793 58910 59863 58980 sw
tri 60076 58910 60146 58980 ne
rect 60146 58910 62056 58980
tri 62056 58910 62126 58980 sw
tri 62339 58910 62409 58980 ne
rect 62409 58910 64319 58980
tri 64319 58910 64389 58980 sw
tri 64606 58910 64676 58980 ne
rect 64676 58920 70613 58980
rect 70669 58920 71000 60120
rect 64676 58910 71000 58920
rect 42800 58854 46230 58910
tri 46230 58854 46287 58910 sw
tri 46556 58854 46612 58910 ne
rect 46612 58854 50798 58910
rect 42800 58528 46287 58854
tri 46287 58528 46612 58854 sw
tri 46612 58528 46937 58854 ne
rect 46937 58815 50798 58854
tri 50798 58815 50893 58910 sw
tri 51085 58815 51180 58910 ne
rect 51180 58815 53065 58910
rect 46937 58528 50893 58815
tri 50893 58528 51180 58815 sw
tri 51180 58528 51467 58815 ne
rect 51467 58812 53065 58815
tri 53065 58812 53163 58910 sw
tri 53349 58812 53447 58910 ne
rect 53447 58816 55329 58910
tri 55329 58816 55423 58910 sw
tri 55617 58816 55711 58910 ne
rect 55711 58816 57597 58910
rect 53447 58812 55423 58816
rect 51467 58528 53163 58812
tri 53163 58528 53447 58812 sw
tri 53447 58528 53731 58812 ne
rect 53731 58528 55423 58812
tri 55423 58528 55711 58816 sw
tri 55711 58528 55999 58816 ne
rect 55999 58814 57597 58816
tri 57597 58814 57693 58910 sw
tri 57883 58814 57979 58910 ne
rect 57979 58814 59863 58910
rect 55999 58528 57693 58814
tri 57693 58528 57979 58814 sw
tri 57979 58528 58265 58814 ne
rect 58265 58697 59863 58814
tri 59863 58697 60076 58910 sw
tri 60146 58697 60359 58910 ne
rect 60359 58883 62126 58910
tri 62126 58883 62153 58910 sw
tri 62409 58883 62436 58910 ne
rect 62436 58883 64389 58910
rect 60359 58697 62153 58883
rect 58265 58528 60076 58697
tri 60076 58528 60245 58697 sw
tri 60359 58528 60528 58697 ne
rect 60528 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64389 58883
tri 64389 58800 64499 58910 sw
tri 64676 58800 64786 58910 ne
rect 64786 58800 71000 58910
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60528 58528 62436 58600
tri 62436 58528 62508 58600 sw
tri 62719 58528 62791 58600 ne
rect 62791 58528 71000 58600
rect 42800 58335 46612 58528
tri 46612 58335 46805 58528 sw
tri 46937 58335 47130 58528 ne
rect 47130 58520 51180 58528
tri 51180 58520 51188 58528 sw
tri 51467 58520 51475 58528 ne
rect 51475 58520 53447 58528
tri 53447 58520 53455 58528 sw
tri 53731 58520 53739 58528 ne
rect 53739 58520 55711 58528
tri 55711 58520 55719 58528 sw
tri 55999 58520 56007 58528 ne
rect 56007 58520 57979 58528
tri 57979 58520 57987 58528 sw
tri 58265 58520 58273 58528 ne
rect 58273 58520 60245 58528
tri 60245 58520 60253 58528 sw
tri 60528 58520 60536 58528 ne
rect 60536 58520 62508 58528
tri 62508 58520 62516 58528 sw
tri 62791 58520 62799 58528 ne
rect 62799 58520 71000 58528
rect 47130 58335 51188 58520
rect 42800 58098 46805 58335
tri 42800 58010 42888 58098 ne
rect 42888 58010 46805 58098
tri 46805 58010 47130 58335 sw
tri 47130 58010 47456 58335 ne
rect 47456 58233 51188 58335
tri 51188 58233 51475 58520 sw
tri 51475 58233 51762 58520 ne
rect 51762 58424 53455 58520
tri 53455 58424 53551 58520 sw
tri 53739 58424 53835 58520 ne
rect 53835 58428 55719 58520
tri 55719 58428 55811 58520 sw
tri 56007 58428 56099 58520 ne
rect 56099 58428 57987 58520
rect 53835 58424 55811 58428
rect 51762 58233 53551 58424
rect 47456 58010 51475 58233
tri 51475 58010 51698 58233 sw
tri 51762 58010 51985 58233 ne
rect 51985 58140 53551 58233
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58426 57987 58428
tri 57987 58426 58081 58520 sw
tri 58273 58426 58367 58520 ne
rect 58367 58426 60253 58520
rect 56387 58140 58081 58426
tri 58081 58140 58367 58426 sw
tri 58367 58140 58653 58426 ne
rect 58653 58423 60253 58426
tri 60253 58423 60350 58520 sw
tri 60536 58423 60633 58520 ne
rect 60633 58423 62516 58520
rect 58653 58140 60350 58423
tri 60350 58140 60633 58423 sw
tri 60633 58140 60916 58423 ne
rect 60916 58317 62516 58423
tri 62516 58317 62719 58520 sw
tri 62799 58317 63002 58520 ne
rect 63002 58317 71000 58520
rect 60916 58140 62719 58317
tri 62719 58140 62896 58317 sw
tri 63002 58140 63179 58317 ne
rect 63179 58140 71000 58317
rect 51985 58010 53835 58140
tri 53835 58010 53965 58140 sw
tri 54119 58010 54249 58140 ne
rect 54249 58010 56099 58140
tri 56099 58010 56229 58140 sw
tri 56387 58010 56517 58140 ne
rect 56517 58010 58367 58140
tri 58367 58010 58497 58140 sw
tri 58653 58010 58783 58140 ne
rect 58783 58010 60633 58140
tri 60633 58010 60763 58140 sw
tri 60916 58010 61046 58140 ne
rect 61046 58010 62896 58140
tri 62896 58010 63026 58140 sw
tri 63179 58010 63309 58140 ne
rect 63309 58010 71000 58140
tri 42600 57810 42800 58010 sw
tri 42888 57810 43088 58010 ne
rect 43088 57810 47130 58010
rect 41200 57626 42800 57810
tri 42800 57626 42984 57810 sw
tri 43088 57626 43272 57810 ne
rect 43272 57685 47130 57810
tri 47130 57685 47456 58010 sw
tri 47456 57685 47781 58010 ne
rect 47781 57772 51698 58010
tri 51698 57772 51936 58010 sw
tri 51985 57772 52223 58010 ne
rect 52223 57856 53965 58010
tri 53965 57856 54119 58010 sw
tri 54249 57856 54403 58010 ne
rect 54403 57856 56229 58010
rect 52223 57772 54119 57856
rect 47781 57685 51936 57772
rect 43272 57663 47456 57685
tri 47456 57663 47477 57685 sw
tri 47781 57663 47802 57685 ne
rect 47802 57663 51936 57685
rect 43272 57626 47477 57663
rect 41200 57430 42984 57626
tri 41200 57338 41292 57430 ne
rect 41292 57338 42984 57430
tri 42984 57338 43272 57626 sw
tri 43272 57338 43560 57626 ne
rect 43560 57338 47477 57626
tri 47477 57338 47802 57663 sw
tri 47802 57486 47980 57663 ne
rect 47980 57486 51936 57663
tri 51936 57486 52223 57772 sw
tri 52223 57486 52509 57772 ne
rect 52509 57770 54119 57772
tri 54119 57770 54205 57856 sw
tri 54403 57770 54489 57856 ne
rect 54489 57770 56229 57856
rect 52509 57486 54205 57770
tri 54205 57486 54489 57770 sw
tri 54489 57486 54773 57770 ne
rect 54773 57760 56229 57770
tri 56229 57760 56479 58010 sw
tri 56517 57760 56767 58010 ne
rect 56767 57760 58497 58010
tri 58497 57760 58747 58010 sw
tri 58783 57760 59033 58010 ne
rect 59033 57760 60763 58010
tri 60763 57760 61013 58010 sw
tri 61046 57760 61296 58010 ne
rect 61296 57760 63026 58010
tri 63026 57760 63276 58010 sw
tri 63309 57760 63559 58010 ne
rect 63559 57760 71000 58010
rect 54773 57486 56479 57760
tri 56479 57486 56753 57760 sw
tri 56767 57486 57041 57760 ne
rect 57041 57486 58747 57760
tri 58747 57486 59021 57760 sw
tri 59033 57486 59307 57760 ne
rect 59307 57486 61013 57760
tri 61013 57486 61287 57760 sw
tri 61296 57486 61570 57760 ne
rect 61570 57486 63276 57760
tri 63276 57486 63550 57760 sw
tri 63559 57486 63833 57760 ne
rect 63833 57486 71000 57760
tri 47980 57338 48128 57486 ne
rect 48128 57338 52223 57486
tri 52223 57338 52370 57486 sw
tri 52509 57338 52657 57486 ne
rect 52657 57338 54489 57486
tri 54489 57338 54637 57486 sw
tri 54773 57338 54921 57486 ne
rect 54921 57472 56753 57486
tri 56753 57472 56767 57486 sw
tri 57041 57472 57055 57486 ne
rect 57055 57472 59021 57486
rect 54921 57338 56767 57472
tri 56767 57338 56901 57472 sw
tri 57055 57338 57189 57472 ne
rect 57189 57380 59021 57472
tri 59021 57380 59127 57486 sw
tri 59307 57380 59413 57486 ne
rect 59413 57380 61287 57486
tri 61287 57380 61393 57486 sw
tri 61570 57380 61676 57486 ne
rect 61676 57380 63550 57486
tri 63550 57380 63656 57486 sw
tri 63833 57380 63939 57486 ne
rect 63939 57380 71000 57486
rect 57189 57338 59127 57380
tri 59127 57338 59169 57380 sw
tri 59413 57338 59455 57380 ne
rect 59455 57338 61393 57380
tri 61393 57338 61435 57380 sw
tri 61676 57338 61718 57380 ne
rect 61718 57338 63656 57380
tri 63656 57338 63698 57380 sw
tri 63939 57338 63981 57380 ne
rect 63981 57338 71000 57380
tri 41000 57138 41200 57338 sw
tri 41292 57138 41492 57338 ne
rect 41492 57208 43272 57338
tri 43272 57208 43402 57338 sw
tri 43560 57208 43690 57338 ne
rect 43690 57245 47802 57338
tri 47802 57245 47895 57338 sw
tri 48128 57245 48220 57338 ne
rect 48220 57245 52370 57338
rect 43690 57208 47895 57245
rect 41492 57138 43402 57208
rect 39600 56920 41200 57138
tri 41200 56920 41418 57138 sw
tri 41492 56920 41710 57138 ne
rect 41710 56920 43402 57138
tri 43402 56920 43690 57208 sw
tri 43690 56920 43978 57208 ne
rect 43978 56920 47895 57208
tri 47895 56920 48220 57245 sw
tri 48220 56920 48546 57245 ne
rect 48546 57207 52370 57245
tri 52370 57207 52502 57338 sw
tri 52657 57207 52788 57338 ne
rect 52788 57207 54637 57338
rect 48546 56920 52502 57207
tri 52502 56920 52788 57207 sw
tri 52788 56920 53075 57207 ne
rect 53075 57204 54637 57207
tri 54637 57204 54771 57338 sw
tri 54921 57204 55055 57338 ne
rect 55055 57208 56901 57338
tri 56901 57208 57031 57338 sw
tri 57189 57208 57319 57338 ne
rect 57319 57208 59169 57338
rect 55055 57204 57031 57208
rect 53075 56920 54771 57204
tri 54771 56920 55055 57204 sw
tri 55055 56920 55339 57204 ne
rect 55339 56920 57031 57204
tri 57031 56920 57319 57208 sw
tri 57319 56920 57607 57208 ne
rect 57607 57094 59169 57208
tri 59169 57094 59413 57338 sw
tri 59455 57094 59699 57338 ne
rect 59699 57283 61435 57338
tri 61435 57283 61490 57338 sw
tri 61718 57283 61773 57338 ne
rect 61773 57283 63698 57338
rect 59699 57094 61490 57283
rect 57607 56920 59413 57094
tri 59413 56920 59587 57094 sw
tri 59699 56920 59873 57094 ne
rect 59873 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63698 57283
tri 63698 57200 63836 57338 sw
tri 63981 57200 64119 57338 ne
rect 64119 57200 71000 57338
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59873 56920 61773 57000
tri 61773 56920 61853 57000 sw
tri 62056 56920 62136 57000 ne
rect 62136 56920 71000 57000
rect 39600 56840 41418 56920
tri 41418 56840 41498 56920 sw
tri 41710 56840 41790 56920 ne
rect 41790 56840 43690 56920
tri 43690 56840 43770 56920 sw
tri 43978 56840 44058 56920 ne
rect 44058 56840 48220 56920
tri 48220 56840 48300 56920 sw
tri 48546 56840 48626 56920 ne
rect 48626 56840 52788 56920
tri 52788 56840 52868 56920 sw
tri 53075 56840 53155 56920 ne
rect 53155 56840 55055 56920
tri 55055 56840 55135 56920 sw
tri 55339 56840 55419 56920 ne
rect 55419 56840 57319 56920
tri 57319 56840 57399 56920 sw
tri 57607 56840 57687 56920 ne
rect 57687 56840 59587 56920
tri 59587 56840 59667 56920 sw
tri 59873 56840 59953 56920 ne
rect 59953 56840 61853 56920
tri 61853 56840 61933 56920 sw
tri 62136 56840 62216 56920 ne
rect 62216 56910 71000 56920
rect 62216 56840 70613 56910
rect 39600 56758 41498 56840
tri 39600 56664 39694 56758 ne
rect 39694 56664 41498 56758
tri 41498 56664 41674 56840 sw
tri 41790 56664 41966 56840 ne
rect 41966 56664 43770 56840
tri 43770 56664 43946 56840 sw
tri 44058 56664 44233 56840 ne
rect 44233 56664 48300 56840
tri 48300 56664 48476 56840 sw
tri 48626 56664 48801 56840 ne
rect 48801 56664 52868 56840
tri 52868 56664 53044 56840 sw
tri 53155 56664 53331 56840 ne
rect 53331 56664 55135 56840
tri 55135 56664 55311 56840 sw
tri 55419 56664 55595 56840 ne
rect 55595 56664 57399 56840
tri 57399 56664 57575 56840 sw
tri 57687 56664 57863 56840 ne
rect 57863 56664 59667 56840
tri 59667 56664 59843 56840 sw
tri 59953 56664 60129 56840 ne
rect 60129 56717 61933 56840
tri 61933 56717 62056 56840 sw
tri 62216 56717 62339 56840 ne
rect 62339 56717 70613 56840
rect 60129 56664 62056 56717
tri 62056 56664 62109 56717 sw
tri 62339 56664 62392 56717 ne
rect 62392 56664 70613 56717
tri 39400 56464 39600 56664 sw
tri 39694 56464 39894 56664 ne
rect 39894 56663 41674 56664
tri 41674 56663 41675 56664 sw
tri 41966 56663 41967 56664 ne
rect 41967 56663 43946 56664
rect 39894 56464 41675 56663
rect 36400 56371 39600 56464
tri 39600 56371 39693 56464 sw
tri 39894 56371 39987 56464 ne
rect 39987 56371 41675 56464
tri 41675 56371 41967 56663 sw
tri 41967 56460 42170 56663 ne
rect 42170 56460 43946 56663
tri 43946 56460 44150 56664 sw
tri 44233 56460 44438 56664 ne
rect 44438 56466 48476 56664
tri 48476 56466 48675 56664 sw
tri 48801 56466 49000 56664 ne
rect 49000 56540 53044 56664
tri 53044 56540 53168 56664 sw
tri 53331 56540 53455 56664 ne
rect 53455 56540 55311 56664
tri 55311 56540 55435 56664 sw
tri 55595 56540 55719 56664 ne
rect 55719 56540 57575 56664
tri 57575 56540 57699 56664 sw
tri 57863 56540 57987 56664 ne
rect 57987 56540 59843 56664
tri 59843 56540 59967 56664 sw
tri 60129 56540 60253 56664 ne
rect 60253 56540 62109 56664
tri 62109 56540 62233 56664 sw
tri 62392 56540 62516 56664 ne
rect 62516 56540 70613 56664
rect 49000 56466 53168 56540
rect 44438 56460 48675 56466
tri 48675 56460 48680 56466 sw
tri 49000 56460 49006 56466 ne
rect 49006 56460 53168 56466
tri 53168 56460 53248 56540 sw
tri 53455 56460 53535 56540 ne
rect 53535 56460 55435 56540
tri 55435 56460 55515 56540 sw
tri 55719 56460 55799 56540 ne
rect 55799 56460 57699 56540
tri 57699 56460 57779 56540 sw
tri 57987 56460 58067 56540 ne
rect 58067 56460 59967 56540
tri 59967 56460 60047 56540 sw
tri 60253 56460 60333 56540 ne
rect 60333 56460 62233 56540
tri 62233 56460 62313 56540 sw
tri 62516 56460 62596 56540 ne
rect 62596 56460 70613 56540
tri 42170 56371 42259 56460 ne
rect 42259 56371 44150 56460
tri 44150 56371 44239 56460 sw
tri 44438 56371 44526 56460 ne
rect 44526 56371 48680 56460
tri 48680 56371 48769 56460 sw
tri 49006 56371 49094 56460 ne
rect 49094 56371 53248 56460
tri 53248 56371 53337 56460 sw
tri 53535 56371 53624 56460 ne
rect 53624 56371 55515 56460
tri 55515 56371 55604 56460 sw
tri 55799 56371 55888 56460 ne
rect 55888 56371 57779 56460
tri 57779 56371 57868 56460 sw
tri 58067 56371 58156 56460 ne
rect 58156 56371 60047 56460
tri 60047 56371 60136 56460 sw
tri 60333 56371 60422 56460 ne
rect 60422 56371 62313 56460
tri 62313 56371 62402 56460 sw
tri 62596 56371 62685 56460 ne
rect 62685 56371 70613 56460
rect 36400 56078 39693 56371
tri 39693 56078 39987 56371 sw
tri 39987 56078 40280 56371 ne
rect 40280 56322 41967 56371
tri 41967 56322 42016 56371 sw
tri 42259 56322 42308 56371 ne
rect 42308 56322 44239 56371
rect 40280 56078 42016 56322
rect 36400 55994 39987 56078
tri 39987 55994 40071 56078 sw
tri 40280 55994 40364 56078 ne
rect 40364 56030 42016 56078
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56084 44239 56322
tri 44239 56084 44526 56371 sw
tri 44526 56084 44814 56371 ne
rect 44814 56140 48769 56371
tri 48769 56140 49000 56371 sw
tri 49094 56140 49325 56371 ne
rect 49325 56253 53337 56371
tri 53337 56253 53455 56371 sw
tri 53624 56253 53742 56371 ne
rect 53742 56253 55604 56371
rect 49325 56140 53455 56253
rect 44814 56084 49000 56140
rect 42600 56030 44526 56084
rect 40364 55994 42308 56030
rect 36400 55700 40071 55994
tri 40071 55700 40364 55994 sw
tri 40364 55700 40658 55994 ne
rect 40658 55738 42308 55994
tri 42308 55738 42600 56030 sw
tri 42600 55830 42800 56030 ne
rect 42800 55988 44526 56030
tri 44526 55988 44622 56084 sw
tri 44814 55988 44910 56084 ne
rect 44910 56025 49000 56084
tri 49000 56025 49115 56140 sw
tri 49325 56025 49440 56140 ne
rect 49440 56025 53455 56140
rect 44910 55988 49115 56025
rect 42800 55830 44622 55988
tri 42800 55738 42892 55830 ne
rect 42892 55738 44622 55830
rect 40658 55700 42600 55738
tri 42600 55700 42638 55738 sw
tri 42892 55700 42930 55738 ne
rect 42930 55700 44622 55738
tri 44622 55700 44910 55988 sw
tri 44910 55700 45198 55988 ne
rect 45198 55700 49115 55988
tri 49115 55700 49440 56025 sw
tri 49440 55700 49766 56025 ne
rect 49766 55987 53455 56025
tri 53455 55987 53722 56253 sw
tri 53742 55987 54008 56253 ne
rect 54008 56160 55604 56253
tri 55604 56160 55815 56371 sw
tri 55888 56160 56099 56371 ne
rect 56099 56160 57868 56371
tri 57868 56160 58079 56371 sw
tri 58156 56160 58367 56371 ne
rect 58367 56160 60136 56371
tri 60136 56160 60347 56371 sw
tri 60422 56160 60633 56371 ne
rect 60633 56160 62402 56371
tri 62402 56160 62613 56371 sw
tri 62685 56160 62896 56371 ne
rect 62896 56160 70613 56371
rect 54008 55987 55815 56160
rect 49766 55700 53722 55987
tri 53722 55700 54008 55987 sw
tri 54008 55700 54295 55987 ne
rect 54295 55876 55815 55987
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60347 56160
rect 56383 55876 58171 56068
rect 54295 55700 56099 55876
tri 56099 55700 56275 55876 sw
tri 56383 55700 56559 55876 ne
rect 56559 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60347 56068
tri 60347 56066 60441 56160 sw
tri 60633 56066 60727 56160 ne
rect 60727 56066 62613 56160
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 56063 62613 56066
tri 62613 56063 62710 56160 sw
tri 62896 56063 62993 56160 ne
rect 62993 56063 70613 56160
rect 61013 55780 62710 56063
tri 62710 55780 62993 56063 sw
tri 62993 55780 63276 56063 ne
rect 63276 55780 70613 56063
rect 56559 55700 58459 55780
tri 58459 55700 58539 55780 sw
tri 58747 55700 58827 55780 ne
rect 58827 55700 60727 55780
tri 60727 55700 60807 55780 sw
tri 61013 55700 61093 55780 ne
rect 61093 55700 62993 55780
tri 62993 55700 63073 55780 sw
tri 63276 55700 63356 55780 ne
rect 63356 55710 70613 55780
rect 70669 55710 71000 56910
rect 63356 55700 71000 55710
rect 36400 55617 40364 55700
tri 40364 55617 40447 55700 sw
tri 40658 55617 40741 55700 ne
rect 40741 55617 42638 55700
rect 36400 55422 40447 55617
tri 36400 55323 36498 55422 ne
rect 36498 55323 40447 55422
tri 40447 55323 40741 55617 sw
tri 40741 55323 41035 55617 ne
rect 41035 55615 42638 55617
tri 42638 55615 42723 55700 sw
tri 42930 55615 43015 55700 ne
rect 43015 55615 44910 55700
rect 41035 55538 42723 55615
tri 42723 55538 42800 55615 sw
tri 43015 55538 43092 55615 ne
rect 43092 55611 44910 55615
tri 44910 55611 44999 55700 sw
tri 45198 55611 45287 55700 ne
rect 45287 55649 49440 55700
tri 49440 55649 49492 55700 sw
tri 49766 55649 49817 55700 ne
rect 49817 55649 54008 55700
rect 45287 55611 49492 55649
rect 43092 55538 44999 55611
rect 41035 55323 42800 55538
tri 42800 55323 43015 55538 sw
tri 43092 55323 43307 55538 ne
rect 43307 55323 44999 55538
tri 44999 55323 45287 55611 sw
tri 45287 55323 45574 55611 ne
rect 45574 55323 49492 55611
tri 49492 55323 49817 55649 sw
tri 49817 55323 50142 55649 ne
rect 50142 55610 54008 55649
tri 54008 55610 54098 55700 sw
tri 54295 55610 54385 55700 ne
rect 54385 55610 56275 55700
rect 50142 55323 54098 55610
tri 54098 55323 54385 55610 sw
tri 54385 55323 54672 55610 ne
rect 54672 55607 56275 55610
tri 56275 55607 56368 55700 sw
tri 56559 55607 56652 55700 ne
rect 56652 55607 58539 55700
rect 54672 55323 56368 55607
tri 56368 55323 56652 55607 sw
tri 56652 55323 56936 55607 ne
rect 56936 55492 58539 55607
tri 58539 55492 58747 55700 sw
tri 58827 55492 59035 55700 ne
rect 59035 55686 60807 55700
tri 60807 55686 60821 55700 sw
tri 61093 55686 61107 55700 ne
rect 61107 55686 63073 55700
rect 59035 55492 60821 55686
rect 56936 55323 58747 55492
tri 58747 55323 58916 55492 sw
tri 59035 55323 59204 55492 ne
rect 59204 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 63073 55686
tri 63073 55600 63173 55700 sw
tri 63356 55600 63456 55700 ne
rect 63456 55600 71000 55700
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59204 55323 61107 55400
tri 61107 55323 61184 55400 sw
tri 61393 55323 61470 55400 ne
rect 61470 55323 71000 55400
tri 36200 55312 36211 55323 sw
tri 36498 55312 36510 55323 ne
rect 36510 55312 40741 55323
tri 40741 55312 40752 55323 sw
tri 41035 55312 41046 55323 ne
rect 41046 55312 43015 55323
tri 43015 55312 43026 55323 sw
tri 43307 55312 43318 55323 ne
rect 43318 55312 45287 55323
tri 45287 55312 45298 55323 sw
tri 45574 55312 45586 55323 ne
rect 45586 55312 49817 55323
tri 49817 55312 49828 55323 sw
tri 50142 55312 50154 55323 ne
rect 50154 55312 54385 55323
tri 54385 55312 54396 55323 sw
tri 54672 55312 54683 55323 ne
rect 54683 55312 56652 55323
tri 56652 55312 56663 55323 sw
tri 56936 55312 56947 55323 ne
rect 56947 55312 58916 55323
tri 58916 55312 58927 55323 sw
tri 59204 55312 59215 55323 ne
rect 59215 55312 61184 55323
tri 61184 55312 61195 55323 sw
tri 61470 55312 61481 55323 ne
rect 61481 55312 71000 55323
rect 33200 55123 36211 55312
tri 36211 55123 36400 55312 sw
tri 36510 55123 36698 55312 ne
rect 36698 55154 40752 55312
tri 40752 55154 40911 55312 sw
tri 41046 55154 41204 55312 ne
rect 41204 55154 43026 55312
rect 36698 55123 40911 55154
rect 33200 54825 36400 55123
tri 36400 54825 36698 55123 sw
tri 36698 54825 36996 55123 ne
rect 36996 54860 40911 55123
tri 40911 54860 41204 55154 sw
tri 41204 54860 41498 55154 ne
rect 41498 55152 43026 55154
tri 43026 55152 43186 55312 sw
tri 43318 55152 43478 55312 ne
rect 43478 55152 45298 55312
rect 41498 54860 43186 55152
tri 43186 54860 43478 55152 sw
tri 43478 54860 43770 55152 ne
rect 43770 55148 45298 55152
tri 45298 55148 45462 55312 sw
tri 45586 55148 45750 55312 ne
rect 45750 55185 49828 55312
tri 49828 55185 49955 55312 sw
tri 50154 55185 50280 55312 ne
rect 50280 55185 54396 55312
rect 45750 55148 49955 55185
rect 43770 54860 45462 55148
tri 45462 54860 45750 55148 sw
tri 45750 54860 46038 55148 ne
rect 46038 54860 49955 55148
tri 49955 54860 50280 55185 sw
tri 50280 54860 50606 55185 ne
rect 50606 55147 54396 55185
tri 54396 55147 54562 55312 sw
tri 54683 55147 54848 55312 ne
rect 54848 55147 56663 55312
rect 50606 54860 54562 55147
tri 54562 54860 54848 55147 sw
tri 54848 54860 55135 55147 ne
rect 55135 55144 56663 55147
tri 56663 55144 56831 55312 sw
tri 56947 55144 57115 55312 ne
rect 57115 55148 58927 55312
tri 58927 55148 59091 55312 sw
tri 59215 55148 59379 55312 ne
rect 59379 55148 61195 55312
rect 57115 55144 59091 55148
rect 55135 54860 56831 55144
tri 56831 54860 57115 55144 sw
tri 57115 54860 57399 55144 ne
rect 57399 54860 59091 55144
tri 59091 54860 59379 55148 sw
tri 59379 54860 59667 55148 ne
rect 59667 55114 61195 55148
tri 61195 55114 61393 55312 sw
tri 61481 55114 61679 55312 ne
rect 61679 55302 71000 55312
rect 61679 55114 70613 55302
rect 59667 54860 61393 55114
tri 61393 54860 61647 55114 sw
tri 61679 54860 61933 55114 ne
rect 61933 54860 70613 55114
rect 36996 54825 41204 54860
rect 33200 54688 36698 54825
tri 36698 54688 36835 54825 sw
tri 36996 54688 37133 54825 ne
rect 37133 54688 41204 54825
rect 33200 54390 36835 54688
tri 36835 54390 37133 54688 sw
tri 37133 54390 37431 54688 ne
rect 37431 54566 41204 54688
tri 41204 54566 41498 54860 sw
tri 41498 54566 41792 54860 ne
rect 41792 54772 43478 54860
tri 43478 54772 43566 54860 sw
tri 43770 54772 43858 54860 ne
rect 43858 54772 45750 54860
rect 41792 54566 43566 54772
rect 37431 54390 41498 54566
rect 33200 54092 37133 54390
tri 37133 54092 37431 54390 sw
tri 37431 54092 37730 54390 ne
rect 37730 54386 41498 54390
tri 41498 54386 41679 54566 sw
tri 41792 54386 41972 54566 ne
rect 41972 54480 43566 54566
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54768 45750 54772
tri 45750 54768 45842 54860 sw
tri 46038 54768 46130 54860 ne
rect 46130 54805 50280 54860
tri 50280 54805 50335 54860 sw
tri 50606 54805 50660 54860 ne
rect 50660 54847 54848 54860
tri 54848 54847 54862 54860 sw
tri 55135 54847 55148 54860 ne
rect 55148 54847 57115 54860
rect 50660 54805 54862 54847
rect 46130 54768 50335 54805
rect 44150 54480 45842 54768
tri 45842 54480 46130 54768 sw
tri 46130 54480 46418 54768 ne
rect 46418 54480 50335 54768
tri 50335 54480 50660 54805 sw
tri 50660 54480 50986 54805 ne
rect 50986 54560 54862 54805
tri 54862 54560 55148 54847 sw
tri 55148 54560 55435 54847 ne
rect 55435 54844 57115 54847
tri 57115 54844 57131 54860 sw
tri 57399 54844 57415 54860 ne
rect 57415 54848 59379 54860
tri 59379 54848 59391 54860 sw
tri 59667 54848 59679 54860 ne
rect 59679 54848 61647 54860
rect 57415 54844 59391 54848
rect 55435 54560 57131 54844
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54560 59391 54844
tri 59391 54560 59679 54848 sw
tri 59679 54560 59967 54848 ne
rect 59967 54846 61647 54848
tri 61647 54846 61661 54860 sw
tri 61933 54846 61947 54860 ne
rect 61947 54846 70613 54860
rect 59967 54560 61661 54846
tri 61661 54560 61947 54846 sw
tri 61947 54560 62233 54846 ne
rect 62233 54560 70613 54846
rect 50986 54480 55148 54560
tri 55148 54480 55228 54560 sw
tri 55435 54480 55515 54560 ne
rect 55515 54480 57415 54560
tri 57415 54480 57495 54560 sw
tri 57699 54480 57779 54560 ne
rect 57779 54480 59679 54560
tri 59679 54480 59759 54560 sw
tri 59967 54480 60047 54560 ne
rect 60047 54480 61947 54560
tri 61947 54480 62027 54560 sw
tri 62233 54480 62313 54560 ne
rect 62313 54480 70613 54560
rect 41972 54386 43858 54480
rect 37730 54092 41679 54386
tri 41679 54092 41972 54386 sw
tri 41972 54092 42266 54386 ne
rect 42266 54286 43858 54386
tri 43858 54286 44052 54480 sw
tri 44150 54286 44344 54480 ne
rect 44344 54286 46130 54480
tri 46130 54286 46324 54480 sw
tri 46418 54286 46612 54480 ne
rect 46612 54286 50660 54480
tri 50660 54286 50855 54480 sw
tri 50986 54286 51180 54480 ne
rect 51180 54286 55228 54480
tri 55228 54286 55423 54480 sw
tri 55515 54286 55709 54480 ne
rect 55709 54286 57495 54480
tri 57495 54286 57689 54480 sw
tri 57779 54286 57973 54480 ne
rect 57973 54286 59759 54480
tri 59759 54286 59953 54480 sw
tri 60047 54286 60241 54480 ne
rect 60241 54286 62027 54480
tri 62027 54286 62221 54480 sw
tri 62313 54286 62507 54480 ne
rect 62507 54286 70613 54480
rect 42266 54188 44052 54286
tri 44052 54188 44150 54286 sw
tri 44344 54188 44442 54286 ne
rect 44442 54188 46324 54286
rect 42266 54092 44150 54188
tri 44150 54092 44246 54188 sw
tri 44442 54092 44538 54188 ne
rect 44538 54092 46324 54188
tri 46324 54092 46518 54286 sw
tri 46612 54092 46806 54286 ne
rect 46806 54092 50855 54286
tri 50855 54092 51048 54286 sw
tri 51180 54092 51374 54286 ne
rect 51374 54273 55423 54286
tri 55423 54273 55435 54286 sw
tri 55709 54273 55722 54286 ne
rect 55722 54273 57689 54286
rect 51374 54092 55435 54273
tri 55435 54092 55616 54273 sw
tri 55722 54092 55903 54273 ne
rect 55903 54180 57689 54273
tri 57689 54180 57795 54286 sw
tri 57973 54180 58079 54286 ne
rect 58079 54180 59953 54286
tri 59953 54180 60059 54286 sw
tri 60241 54180 60347 54286 ne
rect 60347 54180 62221 54286
tri 62221 54180 62327 54286 sw
tri 62507 54180 62613 54286 ne
rect 62613 54180 70613 54286
rect 55903 54092 57795 54180
tri 57795 54092 57883 54180 sw
tri 58079 54092 58167 54180 ne
rect 58167 54092 60059 54180
tri 60059 54092 60147 54180 sw
tri 60347 54092 60435 54180 ne
rect 60435 54092 62327 54180
tri 62327 54092 62415 54180 sw
tri 62613 54092 62701 54180 ne
rect 62701 54102 70613 54180
rect 70669 54102 71000 55302
rect 62701 54092 71000 54102
rect 33200 54081 37431 54092
tri 33200 53991 33289 54081 ne
rect 33289 53991 37431 54081
tri 37431 53991 37532 54092 sw
tri 37730 53991 37830 54092 ne
rect 37830 53991 41972 54092
tri 41972 53991 42073 54092 sw
tri 42266 53991 42367 54092 ne
rect 42367 53991 44246 54092
tri 44246 53991 44347 54092 sw
tri 44538 53991 44639 54092 ne
rect 44639 53998 46518 54092
tri 46518 53998 46612 54092 sw
tri 46806 53998 46900 54092 ne
rect 46900 53998 51048 54092
rect 44639 53991 46612 53998
tri 46612 53991 46619 53998 sw
tri 46900 53991 46906 53998 ne
rect 46906 53991 51048 53998
tri 51048 53991 51149 54092 sw
tri 51374 53991 51474 54092 ne
rect 51474 53991 55616 54092
tri 55616 53991 55717 54092 sw
tri 55903 53991 56004 54092 ne
rect 56004 53991 57883 54092
tri 57883 53991 57984 54092 sw
tri 58167 53991 58268 54092 ne
rect 58268 53991 60147 54092
tri 60147 53991 60248 54092 sw
tri 60435 53991 60536 54092 ne
rect 60536 54000 62415 54092
tri 62415 54000 62507 54092 sw
tri 62701 54000 62793 54092 ne
rect 62793 54000 71000 54092
rect 60536 53991 62507 54000
tri 62507 53991 62516 54000 sw
tri 33000 53791 33200 53991 sw
tri 33289 53791 33489 53991 ne
rect 33489 53791 37532 53991
rect 30000 53732 33200 53791
tri 33200 53732 33259 53791 sw
tri 33489 53732 33549 53791 ne
rect 33549 53732 37532 53791
tri 37532 53732 37791 53991 sw
tri 37830 53732 38090 53991 ne
rect 38090 53732 42073 53991
tri 42073 53732 42332 53991 sw
tri 42367 53732 42626 53991 ne
rect 42626 53732 44347 53991
tri 44347 53732 44606 53991 sw
tri 44639 53732 44898 53991 ne
rect 44898 53732 46619 53991
tri 46619 53732 46878 53991 sw
tri 46906 53732 47166 53991 ne
rect 47166 53732 51149 53991
tri 51149 53732 51408 53991 sw
tri 51474 53732 51734 53991 ne
rect 51734 53732 55717 53991
tri 55717 53732 55976 53991 sw
tri 56004 53732 56263 53991 ne
rect 56263 53896 57984 53991
tri 57984 53896 58079 53991 sw
tri 58268 53896 58363 53991 ne
rect 58363 53896 60248 53991
rect 56263 53732 58079 53896
tri 58079 53732 58243 53896 sw
tri 58363 53732 58527 53896 ne
rect 58527 53800 60248 53896
tri 60248 53800 60439 53991 sw
tri 60536 53800 60727 53991 ne
rect 60727 53800 62516 53991
tri 62516 53800 62707 53991 sw
rect 58527 53732 60439 53800
tri 60439 53732 60507 53800 sw
tri 60727 53732 60795 53800 ne
rect 60795 53732 71000 53800
rect 30000 53443 33259 53732
tri 33259 53443 33549 53732 sw
tri 33549 53443 33838 53732 ne
rect 33838 53469 37791 53732
tri 37791 53469 38054 53732 sw
tri 38090 53469 38352 53732 ne
rect 38352 53469 42332 53732
rect 33838 53443 38054 53469
rect 30000 53232 33549 53443
tri 33549 53232 33760 53443 sw
tri 33838 53232 34049 53443 ne
rect 34049 53232 38054 53443
rect 30000 52943 33760 53232
tri 33760 52943 34049 53232 sw
tri 34049 52943 34338 53232 ne
rect 34338 53171 38054 53232
tri 38054 53171 38352 53469 sw
tri 38352 53171 38650 53469 ne
rect 38650 53465 42332 53469
tri 42332 53465 42600 53732 sw
tri 42626 53465 42893 53732 ne
rect 42893 53465 44606 53732
rect 38650 53171 42600 53465
tri 42600 53171 42893 53465 sw
tri 42893 53171 43187 53465 ne
rect 43187 53463 44606 53465
tri 44606 53463 44875 53732 sw
tri 44898 53463 45167 53732 ne
rect 45167 53463 46878 53732
rect 43187 53171 44875 53463
tri 44875 53171 45167 53463 sw
tri 45167 53171 45459 53463 ne
rect 45459 53459 46878 53463
tri 46878 53459 47151 53732 sw
tri 47166 53459 47439 53732 ne
rect 47439 53568 51408 53732
tri 51408 53568 51572 53732 sw
tri 51734 53568 51898 53732 ne
rect 51898 53568 55976 53732
rect 47439 53459 51572 53568
rect 45459 53171 47151 53459
tri 47151 53171 47439 53459 sw
tri 47439 53171 47726 53459 ne
rect 47726 53243 51572 53459
tri 51572 53243 51898 53568 sw
tri 51898 53243 52223 53568 ne
rect 52223 53529 55976 53568
tri 55976 53529 56179 53732 sw
tri 56263 53529 56466 53732 ne
rect 56466 53529 58243 53732
rect 52223 53243 56179 53529
tri 56179 53243 56466 53529 sw
tri 56466 53243 56752 53529 ne
rect 56752 53527 58243 53529
tri 58243 53527 58448 53732 sw
tri 58527 53527 58732 53732 ne
rect 58732 53527 60507 53732
rect 56752 53243 58448 53527
tri 58448 53243 58732 53527 sw
tri 58732 53243 59016 53527 ne
rect 59016 53512 60507 53527
tri 60507 53512 60727 53732 sw
tri 60795 53512 61015 53732 ne
rect 61015 53722 71000 53732
rect 61015 53512 70613 53722
rect 59016 53243 60727 53512
tri 60727 53243 60996 53512 sw
tri 61015 53243 61284 53512 ne
rect 61284 53243 70613 53512
rect 47726 53171 51898 53243
tri 51898 53171 51969 53243 sw
tri 52223 53171 52294 53243 ne
rect 52294 53171 56466 53243
tri 56466 53171 56537 53243 sw
tri 56752 53171 56824 53243 ne
rect 56824 53171 58732 53243
tri 58732 53171 58804 53243 sw
tri 59016 53171 59088 53243 ne
rect 59088 53171 60996 53243
tri 60996 53171 61068 53243 sw
tri 61284 53171 61356 53243 ne
rect 61356 53171 70613 53243
rect 34338 52952 38352 53171
tri 38352 52952 38572 53171 sw
tri 38650 52952 38870 53171 ne
rect 38870 52952 42893 53171
rect 34338 52943 38572 52952
rect 30000 52749 34049 52943
tri 30000 52653 30095 52749 ne
rect 30095 52653 34049 52749
tri 34049 52653 34338 52943 sw
tri 34338 52653 34627 52943 ne
rect 34627 52653 38572 52943
tri 38572 52653 38870 52952 sw
tri 38870 52653 39168 52952 ne
rect 39168 52880 42893 52952
tri 42893 52880 43184 53171 sw
tri 43187 52880 43478 53171 ne
rect 43478 52880 45167 53171
tri 45167 52880 45458 53171 sw
tri 45459 52880 45750 53171 ne
rect 45750 53168 47439 53171
tri 47439 53168 47442 53171 sw
tri 47726 53168 47730 53171 ne
rect 47730 53168 51969 53171
rect 45750 52880 47442 53168
tri 47442 52880 47730 53168 sw
tri 47730 52880 48018 53168 ne
rect 48018 52918 51969 53168
tri 51969 52918 52223 53171 sw
tri 52294 52918 52548 53171 ne
rect 52548 53167 56537 53171
tri 56537 53167 56542 53171 sw
tri 56824 53167 56828 53171 ne
rect 56828 53167 58804 53171
rect 52548 52918 56542 53167
rect 48018 52880 52223 52918
tri 52223 52880 52260 52918 sw
tri 52548 52880 52586 52918 ne
rect 52586 52880 56542 52918
tri 56542 52880 56828 53167 sw
tri 56828 52880 57115 53167 ne
rect 57115 53164 58804 53167
tri 58804 53164 58811 53171 sw
tri 59088 53164 59095 53171 ne
rect 59095 53168 61068 53171
tri 61068 53168 61071 53171 sw
tri 61356 53168 61359 53171 ne
rect 61359 53168 70613 53171
rect 59095 53164 61071 53168
rect 57115 52880 58811 53164
tri 58811 52880 59095 53164 sw
tri 59095 52880 59379 53164 ne
rect 59379 52880 61071 53164
tri 61071 52880 61359 53168 sw
tri 61359 52880 61647 53168 ne
rect 61647 52880 70613 53168
rect 39168 52653 43184 52880
tri 43184 52653 43411 52880 sw
tri 43478 52653 43705 52880 ne
rect 43705 52653 45458 52880
tri 45458 52653 45685 52880 sw
tri 45750 52653 45977 52880 ne
rect 45977 52653 47730 52880
tri 47730 52653 47957 52880 sw
tri 48018 52653 48244 52880 ne
rect 48244 52653 52260 52880
tri 52260 52653 52487 52880 sw
tri 52586 52653 52812 52880 ne
rect 52812 52653 56828 52880
tri 56828 52653 57055 52880 sw
tri 57115 52653 57342 52880 ne
rect 57342 52653 59095 52880
tri 59095 52653 59322 52880 sw
tri 59379 52653 59606 52880 ne
rect 59606 52653 61359 52880
tri 61359 52653 61586 52880 sw
tri 61647 52653 61874 52880 ne
rect 61874 52653 70613 52880
tri 29800 52512 29941 52653 sw
tri 30095 52512 30237 52653 ne
rect 30237 52512 34338 52653
tri 34338 52512 34479 52653 sw
tri 34627 52512 34769 52653 ne
rect 34769 52512 38870 52653
tri 38870 52512 39011 52653 sw
tri 39168 52512 39310 52653 ne
rect 39310 52586 43411 52653
tri 43411 52586 43478 52653 sw
tri 43705 52586 43772 52653 ne
rect 43772 52586 45685 52653
rect 39310 52512 43478 52586
tri 43478 52512 43552 52586 sw
tri 43772 52512 43846 52586 ne
rect 43846 52512 45685 52586
tri 45685 52512 45826 52653 sw
tri 45977 52512 46118 52653 ne
rect 46118 52512 47957 52653
tri 47957 52512 48098 52653 sw
tri 48244 52512 48386 52653 ne
rect 48386 52512 52487 52653
tri 52487 52512 52628 52653 sw
tri 52812 52512 52954 52653 ne
rect 52954 52580 57055 52653
tri 57055 52580 57128 52653 sw
tri 57342 52580 57415 52653 ne
rect 57415 52580 59322 52653
tri 59322 52580 59395 52653 sw
tri 59606 52580 59679 52653 ne
rect 59679 52580 61586 52653
tri 61586 52580 61659 52653 sw
tri 61874 52580 61947 52653 ne
rect 61947 52580 70613 52653
rect 52954 52512 57128 52580
tri 57128 52512 57196 52580 sw
tri 57415 52512 57483 52580 ne
rect 57483 52512 59395 52580
tri 59395 52512 59463 52580 sw
tri 59679 52512 59747 52580 ne
rect 59747 52512 61659 52580
tri 61659 52512 61727 52580 sw
tri 61947 52512 62015 52580 ne
rect 62015 52522 70613 52580
rect 70669 52522 71000 53722
rect 62015 52512 71000 52522
rect 26800 52453 29941 52512
tri 29941 52453 30000 52512 sw
tri 30237 52453 30295 52512 ne
rect 30295 52453 34479 52512
rect 26800 52158 30000 52453
tri 30000 52158 30295 52453 sw
tri 30295 52158 30590 52453 ne
rect 30590 52223 34479 52453
tri 34479 52223 34769 52512 sw
tri 34769 52223 35058 52512 ne
rect 35058 52427 39011 52512
tri 39011 52427 39097 52512 sw
tri 39310 52427 39395 52512 ne
rect 39395 52427 43552 52512
rect 35058 52223 39097 52427
rect 30590 52158 34769 52223
rect 26800 51910 30295 52158
tri 30295 51910 30543 52158 sw
tri 30590 51910 30838 52158 ne
rect 30838 51934 34769 52158
tri 34769 51934 35058 52223 sw
tri 35058 51934 35347 52223 ne
rect 35347 52128 39097 52223
tri 39097 52128 39395 52427 sw
tri 39395 52128 39693 52427 ne
rect 39693 52422 43552 52427
tri 43552 52422 43642 52512 sw
tri 43846 52422 43936 52512 ne
rect 43936 52500 45826 52512
tri 45826 52500 45838 52512 sw
tri 46118 52500 46130 52512 ne
rect 46130 52500 48098 52512
tri 48098 52500 48110 52512 sw
tri 48386 52500 48398 52512 ne
rect 48398 52500 52628 52512
tri 52628 52500 52640 52512 sw
tri 52954 52500 52966 52512 ne
rect 52966 52500 57196 52512
tri 57196 52500 57208 52512 sw
tri 57483 52500 57495 52512 ne
rect 57495 52500 59463 52512
tri 59463 52500 59475 52512 sw
tri 59747 52500 59759 52512 ne
rect 59759 52500 61727 52512
tri 61727 52500 61739 52512 sw
tri 62015 52500 62027 52512 ne
rect 62027 52500 71000 52512
rect 43936 52422 45838 52500
rect 39693 52128 43642 52422
tri 43642 52128 43936 52422 sw
tri 43936 52128 44230 52422 ne
rect 44230 52208 45838 52422
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52416 48110 52500
tri 48110 52416 48194 52500 sw
tri 48398 52416 48482 52500 ne
rect 48482 52454 52640 52500
tri 52640 52454 52687 52500 sw
tri 52966 52454 53012 52500 ne
rect 53012 52454 57208 52500
rect 48482 52416 52687 52454
rect 46422 52208 48194 52416
rect 44230 52128 46130 52208
tri 46130 52128 46210 52208 sw
tri 46422 52128 46502 52208 ne
rect 46502 52128 48194 52208
tri 48194 52128 48482 52416 sw
tri 48482 52128 48769 52416 ne
rect 48769 52128 52687 52416
tri 52687 52128 53012 52454 sw
tri 53012 52128 53337 52454 ne
rect 53337 52293 57208 52454
tri 57208 52293 57415 52500 sw
tri 57495 52293 57702 52500 ne
rect 57702 52484 59475 52500
tri 59475 52484 59491 52500 sw
tri 59759 52484 59775 52500 ne
rect 59775 52484 61739 52500
rect 57702 52293 59491 52484
rect 53337 52128 57415 52293
tri 57415 52128 57580 52293 sw
tri 57702 52128 57867 52293 ne
rect 57867 52200 59491 52293
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61739 52484
tri 61739 52400 61839 52500 sw
tri 62027 52400 62127 52500 ne
rect 62127 52400 71000 52500
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 57867 52128 59775 52200
tri 59775 52128 59847 52200 sw
tri 60059 52128 60131 52200 ne
rect 60131 52128 71000 52200
rect 35347 51934 39395 52128
rect 30838 51910 35058 51934
rect 26800 51615 30543 51910
tri 30543 51615 30838 51910 sw
tri 30838 51615 31133 51910 ne
rect 31133 51898 35058 51910
tri 35058 51898 35093 51934 sw
tri 35347 51898 35382 51934 ne
rect 35382 51898 39395 51934
rect 31133 51615 35093 51898
rect 26800 51411 30838 51615
tri 26800 51320 26891 51411 ne
rect 26891 51320 30838 51411
tri 30838 51320 31133 51615 sw
tri 31133 51320 31429 51615 ne
rect 31429 51609 35093 51615
tri 35093 51609 35382 51898 sw
tri 35382 51609 35671 51898 ne
rect 35671 51830 39395 51898
tri 39395 51830 39693 52128 sw
tri 39693 51830 39991 52128 ne
rect 39991 51835 43936 52128
tri 43936 51835 44230 52128 sw
tri 44230 51835 44523 52128 ne
rect 44523 51836 46210 52128
tri 46210 51836 46502 52128 sw
tri 46502 52018 46612 52128 ne
rect 46612 52018 48482 52128
tri 46612 51836 46794 52018 ne
rect 46794 51841 48482 52018
tri 48482 51841 48769 52128 sw
tri 48769 51841 49057 52128 ne
rect 49057 51841 53012 52128
rect 46794 51836 48769 51841
rect 44523 51835 46502 51836
rect 39991 51830 44230 51835
rect 35671 51618 39693 51830
tri 39693 51618 39905 51830 sw
tri 39991 51618 40203 51830 ne
rect 40203 51618 44230 51830
rect 35671 51609 39905 51618
rect 31429 51320 35382 51609
tri 35382 51320 35671 51609 sw
tri 35671 51320 35961 51609 ne
rect 35961 51320 39905 51609
tri 39905 51320 40203 51618 sw
tri 40203 51320 40502 51618 ne
rect 40502 51614 44230 51618
tri 44230 51614 44451 51835 sw
tri 44523 51614 44744 51835 ne
rect 44744 51726 46502 51835
tri 46502 51726 46612 51836 sw
tri 46794 51726 46904 51836 ne
rect 46904 51726 48769 51836
rect 44744 51614 46612 51726
rect 40502 51320 44451 51614
tri 44451 51320 44744 51614 sw
tri 44744 51320 45038 51614 ne
rect 45038 51612 46612 51614
tri 46612 51612 46726 51726 sw
tri 46904 51612 47018 51726 ne
rect 47018 51612 48769 51726
rect 45038 51320 46726 51612
tri 46726 51320 47018 51612 sw
tri 47018 51320 47310 51612 ne
rect 47310 51608 48769 51612
tri 48769 51608 49002 51841 sw
tri 49057 51608 49290 51841 ne
rect 49290 51803 53012 51841
tri 53012 51803 53337 52128 sw
tri 53337 51803 53662 52128 ne
rect 53662 51842 57580 52128
tri 57580 51842 57867 52128 sw
tri 57867 51842 58153 52128 ne
rect 58153 51916 59847 52128
tri 59847 51916 60059 52128 sw
tri 60131 51916 60343 52128 ne
rect 60343 51916 71000 52128
rect 58153 51842 60059 51916
rect 53662 51803 57867 51842
rect 49290 51645 53337 51803
tri 53337 51645 53495 51803 sw
tri 53662 51645 53820 51803 ne
rect 53820 51645 57867 51803
rect 49290 51608 53495 51645
rect 47310 51320 49002 51608
tri 49002 51320 49290 51608 sw
tri 49290 51320 49578 51608 ne
rect 49578 51320 53495 51608
tri 53495 51320 53820 51645 sw
tri 53820 51320 54146 51645 ne
rect 54146 51607 57867 51645
tri 57867 51607 58102 51842 sw
tri 58153 51607 58388 51842 ne
rect 58388 51632 60059 51842
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58388 51607 60343 51632
rect 54146 51320 58102 51607
tri 58102 51320 58388 51607 sw
tri 58388 51320 58675 51607 ne
rect 58675 51604 60343 51607
tri 60343 51604 60371 51632 sw
tri 60627 51604 60655 51632 ne
rect 60655 51604 71000 51632
rect 58675 51320 60371 51604
tri 60371 51320 60655 51604 sw
tri 60655 51320 60939 51604 ne
rect 60939 51320 71000 51604
tri 26600 51120 26800 51320 sw
tri 26891 51120 27091 51320 ne
rect 27091 51309 31133 51320
tri 31133 51309 31144 51320 sw
tri 31429 51309 31439 51320 ne
rect 31439 51309 35671 51320
rect 27091 51120 31144 51309
rect 25200 50942 26800 51120
tri 26800 50942 26978 51120 sw
tri 27091 50942 27269 51120 ne
rect 27269 51014 31144 51120
tri 31144 51014 31439 51309 sw
tri 31439 51014 31735 51309 ne
rect 31735 51081 35671 51309
tri 35671 51081 35911 51320 sw
tri 35961 51081 36200 51320 ne
rect 36200 51312 40203 51320
tri 40203 51312 40211 51320 sw
tri 40502 51312 40509 51320 ne
rect 40509 51312 44744 51320
rect 36200 51081 40211 51312
rect 31735 51014 35911 51081
tri 35911 51014 35977 51081 sw
tri 36200 51014 36267 51081 ne
rect 36267 51014 40211 51081
tri 40211 51014 40509 51312 sw
tri 40509 51014 40808 51312 ne
rect 40808 51308 44744 51312
tri 44744 51308 44757 51320 sw
tri 45038 51308 45050 51320 ne
rect 45050 51308 47018 51320
rect 40808 51014 44757 51308
tri 44757 51014 45050 51308 sw
tri 45050 51014 45344 51308 ne
rect 45344 51306 47018 51308
tri 47018 51306 47032 51320 sw
tri 47310 51306 47324 51320 ne
rect 47324 51306 49290 51320
rect 45344 51014 47032 51306
tri 47032 51014 47324 51306 sw
tri 47324 51014 47616 51306 ne
rect 47616 51302 49290 51306
tri 49290 51302 49308 51320 sw
tri 49578 51302 49596 51320 ne
rect 49596 51302 53820 51320
rect 47616 51014 49308 51302
tri 49308 51014 49596 51302 sw
tri 49596 51014 49884 51302 ne
rect 49884 51014 53820 51302
tri 53820 51014 54126 51320 sw
tri 54146 51014 54452 51320 ne
rect 54452 51301 58388 51320
tri 58388 51301 58408 51320 sw
tri 58675 51301 58694 51320 ne
rect 58694 51301 60655 51320
rect 54452 51014 58408 51301
tri 58408 51014 58694 51301 sw
tri 58694 51014 58981 51301 ne
rect 58981 51298 60655 51301
tri 60655 51298 60677 51320 sw
tri 60939 51298 60961 51320 ne
rect 60961 51298 71000 51320
rect 58981 51014 60677 51298
tri 60677 51014 60961 51298 sw
tri 60961 51014 61245 51298 ne
rect 61245 51014 71000 51298
rect 27269 50946 31439 51014
tri 31439 50946 31507 51014 sw
tri 31735 50946 31802 51014 ne
rect 31802 50946 35977 51014
rect 27269 50942 31507 50946
rect 25200 50740 26978 50942
tri 25200 50651 25289 50740 ne
rect 25289 50651 26978 50740
tri 26978 50651 27269 50942 sw
tri 27269 50651 27560 50942 ne
rect 27560 50651 31507 50942
tri 31507 50651 31802 50946 sw
tri 31802 50651 32098 50946 ne
rect 32098 50791 35977 50946
tri 35977 50791 36200 51014 sw
tri 36267 50791 36489 51014 ne
rect 36489 50949 40509 51014
tri 40509 50949 40574 51014 sw
tri 40808 50949 40872 51014 ne
rect 40872 50949 45050 51014
rect 36489 50791 40574 50949
rect 32098 50651 36200 50791
tri 36200 50651 36340 50791 sw
tri 36489 50651 36630 50791 ne
rect 36630 50651 40574 50791
tri 40574 50651 40872 50949 sw
tri 40872 50651 41171 50949 ne
rect 41171 50900 45050 50949
tri 45050 50900 45164 51014 sw
tri 45344 50900 45458 51014 ne
rect 45458 50900 47324 51014
tri 47324 50900 47438 51014 sw
tri 47616 50900 47730 51014 ne
rect 47730 50900 49596 51014
tri 49596 50900 49710 51014 sw
tri 49884 50900 49998 51014 ne
rect 49998 50900 54126 51014
tri 54126 50900 54240 51014 sw
tri 54452 50900 54566 51014 ne
rect 54566 50900 58694 51014
tri 58694 50900 58808 51014 sw
tri 58981 50900 59095 51014 ne
rect 59095 50900 60961 51014
tri 60961 50900 61075 51014 sw
tri 61245 50900 61359 51014 ne
rect 61359 50900 71000 51014
rect 41171 50651 45164 50900
tri 45164 50651 45413 50900 sw
tri 45458 50651 45707 50900 ne
rect 45707 50651 47438 50900
tri 47438 50651 47687 50900 sw
tri 47730 50651 47979 50900 ne
rect 47979 50651 49710 50900
tri 49710 50651 49959 50900 sw
tri 49998 50651 50247 50900 ne
rect 50247 50651 54240 50900
tri 54240 50651 54489 50900 sw
tri 54566 50651 54815 50900 ne
rect 54815 50651 58808 50900
tri 58808 50651 59057 50900 sw
tri 59095 50651 59344 50900 ne
rect 59344 50800 61075 50900
tri 61075 50800 61175 50900 sw
tri 61359 50800 61459 50900 ne
rect 61459 50800 71000 50900
rect 59344 50651 61175 50800
tri 61175 50651 61324 50800 sw
tri 25000 50451 25200 50651 sw
tri 25289 50451 25489 50651 ne
rect 25489 50451 27269 50651
rect 23600 50262 25200 50451
tri 25200 50262 25389 50451 sw
tri 25489 50262 25678 50451 ne
rect 25678 50360 27269 50451
tri 27269 50360 27560 50651 sw
tri 27560 50360 27851 50651 ne
rect 27851 50360 31802 50651
tri 31802 50360 32093 50651 sw
tri 32098 50360 32389 50651 ne
rect 32389 50649 36340 50651
tri 36340 50649 36342 50651 sw
tri 36630 50649 36631 50651 ne
rect 36631 50649 40872 50651
rect 32389 50360 36342 50649
tri 36342 50360 36631 50649 sw
tri 36631 50360 36921 50649 ne
rect 36921 50360 40872 50649
tri 40872 50360 41163 50651 sw
tri 41171 50360 41462 50651 ne
rect 41462 50606 45413 50651
tri 45413 50606 45458 50651 sw
tri 45707 50606 45752 50651 ne
rect 45752 50606 47687 50651
rect 41462 50360 45458 50606
tri 45458 50360 45704 50606 sw
tri 45752 50360 45998 50606 ne
rect 45998 50520 47687 50606
tri 47687 50520 47818 50651 sw
tri 47979 50520 48110 50651 ne
rect 48110 50520 49959 50651
tri 49959 50520 50090 50651 sw
tri 50247 50520 50378 50651 ne
rect 50378 50520 54489 50651
tri 54489 50520 54620 50651 sw
tri 54815 50520 54946 50651 ne
rect 54946 50600 59057 50651
tri 59057 50600 59108 50651 sw
tri 59344 50600 59395 50651 ne
rect 59395 50600 61324 50651
tri 61324 50600 61375 50651 sw
rect 54946 50520 59108 50600
tri 59108 50520 59188 50600 sw
tri 59395 50520 59475 50600 ne
rect 59475 50520 71000 50600
rect 45998 50360 47818 50520
tri 47818 50360 47978 50520 sw
tri 48110 50360 48270 50520 ne
rect 48270 50360 50090 50520
tri 50090 50360 50250 50520 sw
tri 50378 50360 50538 50520 ne
rect 50538 50360 54620 50520
tri 54620 50360 54780 50520 sw
tri 54946 50360 55106 50520 ne
rect 55106 50360 59188 50520
tri 59188 50360 59348 50520 sw
tri 59475 50360 59635 50520 ne
rect 59635 50360 71000 50520
rect 25678 50264 27560 50360
tri 27560 50264 27656 50360 sw
tri 27851 50264 27947 50360 ne
rect 27947 50269 32093 50360
tri 32093 50269 32185 50360 sw
tri 32389 50269 32480 50360 ne
rect 32480 50269 36631 50360
rect 27947 50264 32185 50269
rect 25678 50262 27656 50264
rect 23600 50071 25389 50262
tri 23600 49973 23698 50071 ne
rect 23698 49973 25389 50071
tri 25389 49973 25678 50262 sw
tri 25678 49973 25967 50262 ne
rect 25967 49973 27656 50262
tri 27656 49973 27947 50264 sw
tri 27947 49973 28237 50264 ne
rect 28237 49973 32185 50264
tri 32185 49973 32480 50269 sw
tri 32480 49973 32775 50269 ne
rect 32775 50263 36631 50269
tri 36631 50263 36729 50360 sw
tri 36921 50263 37018 50360 ne
rect 37018 50272 41163 50360
tri 41163 50272 41252 50360 sw
tri 41462 50272 41550 50360 ne
rect 41550 50272 45704 50360
rect 37018 50263 41252 50272
rect 32775 49973 36729 50263
tri 36729 49973 37018 50263 sw
tri 37018 49973 37307 50263 ne
rect 37307 49973 41252 50263
tri 41252 49973 41550 50272 sw
tri 41550 49973 41848 50272 ne
rect 41848 50267 45704 50272
tri 45704 50267 45797 50360 sw
tri 45998 50267 46091 50360 ne
rect 46091 50267 47978 50360
rect 41848 49973 45797 50267
tri 45797 49973 46091 50267 sw
tri 46091 49973 46385 50267 ne
rect 46385 50228 47978 50267
tri 47978 50228 48110 50360 sw
tri 48270 50228 48402 50360 ne
rect 48402 50330 50250 50360
tri 50250 50330 50280 50360 sw
tri 50538 50330 50567 50360 ne
rect 50567 50330 54780 50360
rect 48402 50228 50280 50330
rect 46385 50043 48110 50228
tri 48110 50043 48295 50228 sw
tri 48402 50043 48587 50228 ne
rect 48587 50043 50280 50228
tri 50280 50043 50567 50330 sw
tri 50567 50043 50855 50330 ne
rect 50855 50043 54780 50330
tri 54780 50043 55098 50360 sw
tri 55106 50043 55423 50360 ne
rect 55423 50313 59348 50360
tri 59348 50313 59395 50360 sw
tri 59635 50313 59682 50360 ne
rect 59682 50313 71000 50360
rect 55423 50043 59395 50313
tri 59395 50043 59666 50313 sw
tri 59682 50043 59952 50313 ne
rect 59952 50043 71000 50313
rect 46385 49973 48295 50043
tri 48295 49973 48365 50043 sw
tri 48587 49973 48657 50043 ne
rect 48657 49973 50567 50043
tri 50567 49973 50637 50043 sw
tri 50855 49973 50924 50043 ne
rect 50924 49973 55098 50043
tri 55098 49973 55167 50043 sw
tri 55423 49973 55492 50043 ne
rect 55492 49973 59666 50043
tri 59666 49973 59735 50043 sw
tri 59952 49973 60022 50043 ne
rect 60022 49973 71000 50043
tri 23400 49773 23600 49973 sw
tri 23698 49773 23898 49973 ne
rect 23898 49773 25678 49973
rect 20400 49476 23600 49773
tri 23600 49476 23898 49773 sw
tri 23898 49476 24195 49773 ne
rect 24195 49684 25678 49773
tri 25678 49684 25967 49973 sw
tri 25967 49684 26256 49973 ne
rect 26256 49684 27947 49973
rect 24195 49629 25967 49684
tri 25967 49629 26022 49684 sw
tri 26256 49629 26311 49684 ne
rect 26311 49683 27947 49684
tri 27947 49683 28237 49973 sw
tri 28237 49683 28528 49973 ne
rect 28528 49971 32480 49973
tri 32480 49971 32482 49973 sw
tri 32775 49971 32777 49973 ne
rect 32777 49971 37018 49973
tri 37018 49971 37020 49973 sw
tri 37307 49971 37309 49973 ne
rect 37309 49971 41550 49973
tri 41550 49971 41552 49973 sw
tri 41848 49971 41850 49973 ne
rect 41850 49971 46091 49973
tri 46091 49971 46093 49973 sw
tri 46385 49971 46387 49973 ne
rect 46387 49971 48365 49973
tri 48365 49971 48367 49973 sw
tri 48657 49971 48659 49973 ne
rect 48659 49971 50637 49973
tri 50637 49971 50639 49973 sw
tri 50924 49971 50926 49973 ne
rect 50926 49971 55167 49973
tri 55167 49971 55169 49973 sw
tri 55492 49971 55494 49973 ne
rect 55494 49971 59735 49973
tri 59735 49971 59737 49973 sw
tri 60022 49971 60024 49973 ne
rect 60024 49971 71000 49973
rect 28528 49749 32482 49971
tri 32482 49749 32705 49971 sw
tri 32777 49749 33000 49971 ne
rect 33000 49749 37020 49971
rect 28528 49683 32705 49749
rect 26311 49629 28237 49683
rect 24195 49476 26022 49629
rect 20400 49452 23898 49476
tri 23898 49452 23921 49476 sw
tri 24195 49452 24219 49476 ne
rect 24219 49452 26022 49476
rect 20400 49154 23921 49452
tri 23921 49154 24219 49452 sw
tri 24219 49154 24517 49452 ne
rect 24517 49340 26022 49452
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49438 28237 49629
tri 28237 49438 28482 49683 sw
tri 28528 49438 28773 49683 ne
rect 28773 49453 32705 49683
tri 32705 49453 33000 49749 sw
tri 33000 49453 33295 49749 ne
rect 33295 49682 37020 49749
tri 37020 49682 37309 49971 sw
tri 37309 49682 37599 49971 ne
rect 37599 49682 41552 49971
rect 33295 49507 37309 49682
tri 37309 49507 37485 49682 sw
tri 37599 49507 37774 49682 ne
rect 37774 49673 41552 49682
tri 41552 49673 41850 49971 sw
tri 41850 49673 42149 49971 ne
rect 42149 49678 46093 49971
tri 46093 49678 46387 49971 sw
tri 46387 49678 46680 49971 ne
rect 46680 49679 48367 49971
tri 48367 49679 48659 49971 sw
tri 48659 49679 48951 49971 ne
rect 48951 49755 50639 49971
tri 50639 49755 50855 49971 sw
tri 50926 49755 51142 49971 ne
rect 51142 49755 55169 49971
rect 48951 49679 50855 49755
rect 46680 49678 48659 49679
rect 42149 49673 46387 49678
rect 37774 49525 41850 49673
tri 41850 49525 41999 49673 sw
tri 42149 49525 42297 49673 ne
rect 42297 49525 46387 49673
rect 37774 49507 41999 49525
rect 33295 49453 37485 49507
rect 28773 49438 33000 49453
rect 26600 49340 28482 49438
rect 24517 49154 26311 49340
rect 20400 48857 24219 49154
tri 24219 48857 24517 49154 sw
tri 24517 48857 24814 49154 ne
rect 24814 49051 26311 49154
tri 26311 49051 26600 49340 sw
tri 26600 49140 26800 49340 ne
rect 26800 49147 28482 49340
tri 28482 49147 28773 49438 sw
tri 28773 49147 29063 49438 ne
rect 29063 49158 33000 49438
tri 33000 49158 33295 49453 sw
tri 33295 49158 33590 49453 ne
rect 33590 49218 37485 49453
tri 37485 49218 37774 49507 sw
tri 37774 49218 38063 49507 ne
rect 38063 49227 41999 49507
tri 41999 49227 42297 49525 sw
tri 42297 49227 42595 49525 ne
rect 42595 49516 46387 49525
tri 46387 49516 46549 49678 sw
tri 46680 49516 46842 49678 ne
rect 46842 49516 48659 49678
rect 42595 49227 46549 49516
rect 38063 49218 42297 49227
rect 33590 49158 37774 49218
rect 29063 49152 33295 49158
tri 33295 49152 33301 49158 sw
tri 33590 49152 33597 49158 ne
rect 33597 49152 37774 49158
rect 29063 49147 33301 49152
rect 26800 49140 28773 49147
tri 26800 49051 26889 49140 ne
rect 26889 49051 28773 49140
rect 24814 48857 26600 49051
tri 26600 48857 26794 49051 sw
tri 26889 48857 27083 49051 ne
rect 27083 48857 28773 49051
tri 28773 48857 29063 49147 sw
tri 29063 48857 29354 49147 ne
rect 29354 48857 33301 49147
tri 33301 48857 33597 49152 sw
tri 33597 48857 33892 49152 ne
rect 33892 48928 37774 49152
tri 37774 48928 38063 49218 sw
tri 38063 48928 38352 49218 ne
rect 38352 48928 42297 49218
tri 42297 48928 42595 49227 sw
tri 42595 48928 42893 49227 ne
rect 42893 49222 46549 49227
tri 46549 49222 46842 49516 sw
tri 46842 49222 47136 49516 ne
rect 47136 49512 48659 49516
tri 48659 49512 48826 49679 sw
tri 48951 49512 49118 49679 ne
rect 49118 49512 50855 49679
rect 47136 49222 48826 49512
rect 42893 48928 46842 49222
tri 46842 48928 47136 49222 sw
tri 47136 48928 47430 49222 ne
rect 47430 49220 48826 49222
tri 48826 49220 49118 49512 sw
tri 49118 49220 49410 49512 ne
rect 49410 49468 50855 49512
tri 50855 49468 51142 49755 sw
tri 51142 49468 51430 49755 ne
rect 51430 49646 55169 49755
tri 55169 49646 55494 49971 sw
tri 55494 49646 55820 49971 ne
rect 55820 49685 59737 49971
tri 59737 49685 60024 49971 sw
tri 60024 49685 60310 49971 ne
rect 60310 49685 71000 49971
rect 55820 49646 60024 49685
rect 51430 49468 55494 49646
rect 49410 49220 51142 49468
rect 47430 48928 49118 49220
tri 49118 48928 49410 49220 sw
tri 49410 48928 49702 49220 ne
rect 49702 49216 51142 49220
tri 51142 49216 51394 49468 sw
tri 51430 49216 51682 49468 ne
rect 51682 49325 55494 49468
tri 55494 49325 55815 49646 sw
tri 55820 49325 56140 49646 ne
rect 56140 49487 60024 49646
tri 60024 49487 60222 49685 sw
tri 60310 49487 60508 49685 ne
rect 60508 49487 71000 49685
rect 56140 49325 60222 49487
rect 51682 49216 55815 49325
rect 49702 48928 51394 49216
tri 51394 48928 51682 49216 sw
tri 51682 48928 51969 49216 ne
rect 51969 49000 55815 49216
tri 55815 49000 56140 49325 sw
tri 56140 49000 56466 49325 ne
rect 56466 49200 60222 49325
tri 60222 49200 60508 49487 sw
tri 60508 49200 60795 49487 ne
rect 60795 49200 71000 49487
rect 56466 49000 60508 49200
tri 60508 49000 60708 49200 sw
rect 51969 48928 56140 49000
tri 56140 48928 56212 49000 sw
tri 56466 48928 56537 49000 ne
rect 56537 48928 71000 49000
rect 33892 48857 38063 48928
tri 38063 48857 38135 48928 sw
tri 38352 48857 38424 48928 ne
rect 38424 48857 42595 48928
tri 42595 48857 42667 48928 sw
tri 42893 48857 42965 48928 ne
rect 42965 48920 47136 48928
tri 47136 48920 47144 48928 sw
tri 47430 48920 47438 48928 ne
rect 47438 48920 49410 48928
tri 49410 48920 49418 48928 sw
tri 49702 48920 49710 48928 ne
rect 49710 48920 51682 48928
tri 51682 48920 51690 48928 sw
tri 51969 48920 51978 48928 ne
rect 51978 48920 56212 48928
tri 56212 48920 56220 48928 sw
tri 56537 48920 56546 48928 ne
rect 56546 48920 71000 48928
rect 42965 48857 47144 48920
tri 47144 48857 47208 48920 sw
tri 47438 48857 47501 48920 ne
rect 47501 48857 49418 48920
tri 49418 48857 49481 48920 sw
tri 49710 48857 49773 48920 ne
rect 49773 48857 51690 48920
tri 51690 48857 51753 48920 sw
tri 51978 48857 52041 48920 ne
rect 52041 48857 56220 48920
tri 56220 48857 56284 48920 sw
tri 56546 48857 56609 48920 ne
rect 56609 48857 71000 48920
rect 20400 48731 24517 48857
tri 20400 48647 20483 48731 ne
rect 20483 48671 24517 48731
tri 24517 48671 24702 48857 sw
tri 24814 48760 24911 48857 ne
rect 24911 48851 26794 48857
tri 26794 48851 26800 48857 sw
tri 27083 48851 27089 48857 ne
rect 27089 48851 29063 48857
rect 24911 48760 26800 48851
tri 26800 48760 26891 48851 sw
tri 27089 48760 27180 48851 ne
rect 27180 48760 29063 48851
tri 29063 48760 29160 48857 sw
tri 29354 48760 29451 48857 ne
rect 29451 48760 33597 48857
tri 33597 48760 33693 48857 sw
tri 33892 48760 33989 48857 ne
rect 33989 48760 38135 48857
tri 38135 48760 38231 48857 sw
tri 38424 48760 38521 48857 ne
rect 38521 48760 42667 48857
tri 42667 48760 42763 48857 sw
tri 42965 48760 43062 48857 ne
rect 43062 48760 47208 48857
tri 47208 48760 47304 48857 sw
tri 47501 48760 47598 48857 ne
rect 47598 48760 49481 48857
tri 49481 48760 49578 48857 sw
tri 49773 48760 49870 48857 ne
rect 49870 48760 51753 48857
tri 51753 48760 51850 48857 sw
tri 52041 48760 52138 48857 ne
rect 52138 48760 56284 48857
tri 56284 48760 56380 48857 sw
tri 56609 48760 56706 48857 ne
rect 56706 48760 71000 48857
tri 24911 48671 25000 48760 ne
rect 25000 48671 26891 48760
rect 20483 48647 24702 48671
tri 24702 48647 24726 48671 sw
tri 25000 48647 25024 48671 ne
rect 25024 48647 26891 48671
tri 26891 48647 27004 48760 sw
tri 27180 48647 27293 48760 ne
rect 27293 48647 29160 48760
tri 29160 48647 29273 48760 sw
tri 29451 48647 29563 48760 ne
rect 29563 48647 33693 48760
tri 33693 48647 33806 48760 sw
tri 33989 48647 34101 48760 ne
rect 34101 48647 38231 48760
tri 38231 48647 38344 48760 sw
tri 38521 48647 38633 48760 ne
rect 38633 48647 42763 48760
tri 42763 48647 42876 48760 sw
tri 43062 48647 43174 48760 ne
rect 43174 48647 47304 48760
tri 47304 48647 47417 48760 sw
tri 47598 48647 47711 48760 ne
rect 47711 48647 49578 48760
tri 49578 48647 49691 48760 sw
tri 49870 48647 49983 48760 ne
rect 49983 48647 51850 48760
tri 51850 48647 51963 48760 sw
tri 52138 48647 52250 48760 ne
rect 52250 48675 56380 48760
tri 56380 48675 56466 48760 sw
tri 56706 48675 56791 48760 ne
rect 56791 48675 71000 48760
rect 52250 48647 56466 48675
tri 56466 48647 56493 48675 sw
tri 56791 48647 56818 48675 ne
rect 56818 48647 71000 48675
tri 20200 48447 20400 48647 sw
tri 20483 48447 20683 48647 ne
rect 20683 48447 24726 48647
rect 17200 48164 20400 48447
tri 20400 48164 20683 48447 sw
tri 20683 48164 20966 48447 ne
rect 20966 48373 24726 48447
tri 24726 48373 25000 48647 sw
tri 25024 48373 25298 48647 ne
rect 25298 48411 27004 48647
tri 27004 48411 27240 48647 sw
tri 27293 48411 27529 48647 ne
rect 27529 48411 29273 48647
tri 29273 48411 29509 48647 sw
tri 29563 48411 29800 48647 ne
rect 29800 48411 33806 48647
rect 25298 48380 27240 48411
tri 27240 48380 27271 48411 sw
tri 27529 48380 27560 48411 ne
rect 27560 48380 29509 48411
tri 29509 48380 29540 48411 sw
tri 29800 48380 29831 48411 ne
rect 29831 48380 33806 48411
tri 33806 48380 34073 48647 sw
tri 34101 48380 34369 48647 ne
rect 34369 48639 38344 48647
tri 38344 48639 38352 48647 sw
tri 38633 48639 38641 48647 ne
rect 38641 48639 42876 48647
rect 34369 48380 38352 48639
tri 38352 48380 38611 48639 sw
tri 38641 48380 38901 48639 ne
rect 38901 48380 42876 48639
tri 42876 48380 43143 48647 sw
tri 43174 48380 43442 48647 ne
rect 43442 48626 47417 48647
tri 47417 48626 47438 48647 sw
tri 47711 48626 47732 48647 ne
rect 47732 48626 49691 48647
rect 43442 48380 47438 48626
tri 47438 48380 47684 48626 sw
tri 47732 48380 47978 48626 ne
rect 47978 48540 49691 48626
tri 49691 48540 49798 48647 sw
tri 49983 48540 50090 48647 ne
rect 50090 48540 51963 48647
tri 51963 48540 52070 48647 sw
tri 52250 48540 52358 48647 ne
rect 52358 48540 56493 48647
tri 56493 48540 56600 48647 sw
tri 56818 48540 56926 48647 ne
rect 56926 48540 71000 48647
rect 47978 48380 49798 48540
tri 49798 48380 49958 48540 sw
tri 50090 48380 50250 48540 ne
rect 50250 48380 52070 48540
tri 52070 48380 52230 48540 sw
tri 52358 48380 52518 48540 ne
rect 52518 48380 56600 48540
tri 56600 48380 56760 48540 sw
tri 56926 48380 57086 48540 ne
rect 57086 48380 71000 48540
rect 25298 48373 27271 48380
rect 20966 48164 25000 48373
rect 17200 47881 20683 48164
tri 20683 47881 20966 48164 sw
tri 20966 47881 21250 48164 ne
rect 21250 48076 25000 48164
tri 25000 48076 25298 48373 sw
tri 25298 48076 25595 48373 ne
rect 25595 48091 27271 48373
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48120 29540 48380
tri 29540 48120 29800 48380 sw
tri 29831 48120 30091 48380 ne
rect 30091 48120 34073 48380
rect 27849 48091 29800 48120
rect 25595 48076 27560 48091
rect 21250 47907 25298 48076
tri 25298 47907 25467 48076 sw
tri 25595 47907 25764 48076 ne
rect 25764 47907 27560 48076
rect 21250 47881 25467 47907
rect 17200 47878 20966 47881
tri 20966 47878 20970 47881 sw
tri 21250 47878 21253 47881 ne
rect 21253 47878 25467 47881
rect 17200 47595 20970 47878
tri 20970 47595 21253 47878 sw
tri 21253 47595 21536 47878 ne
rect 21536 47609 25467 47878
tri 25467 47609 25764 47907 sw
tri 25764 47609 26062 47907 ne
rect 26062 47802 27560 47907
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 47829 29800 48091
tri 29800 47829 30091 48120 sw
tri 30091 47829 30381 48120 ne
rect 30381 48085 34073 48120
tri 34073 48085 34369 48380 sw
tri 34369 48085 34664 48380 ne
rect 34664 48091 38611 48380
tri 38611 48091 38901 48380 sw
tri 38901 48091 39190 48380 ne
rect 39190 48184 43143 48380
tri 43143 48184 43340 48380 sw
tri 43442 48184 43638 48380 ne
rect 43638 48184 47684 48380
rect 39190 48091 43340 48184
rect 34664 48085 38901 48091
rect 30381 47902 34369 48085
tri 34369 47902 34552 48085 sw
tri 34664 47902 34847 48085 ne
rect 34847 47902 38901 48085
rect 30381 47829 34552 47902
rect 28138 47802 30091 47829
rect 26062 47609 27849 47802
rect 21536 47595 25764 47609
rect 17200 47405 21253 47595
tri 17200 47311 17293 47405 ne
rect 17293 47311 21253 47405
tri 21253 47311 21536 47595 sw
tri 21536 47311 21819 47595 ne
rect 21819 47311 25764 47595
tri 25764 47311 26062 47609 sw
tri 26062 47311 26360 47609 ne
rect 26360 47600 27849 47609
tri 27849 47600 28051 47802 sw
tri 28138 47600 28340 47802 ne
rect 28340 47602 30091 47802
tri 30091 47602 30318 47829 sw
tri 30381 47602 30609 47829 ne
rect 30609 47607 34552 47829
tri 34552 47607 34847 47902 sw
tri 34847 47607 35142 47902 ne
rect 35142 47890 38901 47902
tri 38901 47890 39102 48091 sw
tri 39190 47890 39391 48091 ne
rect 39391 47890 43340 48091
rect 35142 47607 39102 47890
rect 30609 47602 34847 47607
rect 28340 47600 30318 47602
rect 26360 47311 28051 47600
tri 28051 47311 28340 47600 sw
tri 28340 47311 28629 47600 ne
rect 28629 47311 30318 47600
tri 30318 47311 30609 47602 sw
tri 30609 47311 30899 47602 ne
rect 30899 47311 34847 47602
tri 34847 47311 35142 47607 sw
tri 35142 47311 35437 47607 ne
rect 35437 47601 39102 47607
tri 39102 47601 39391 47890 sw
tri 39391 47601 39680 47890 ne
rect 39680 47886 43340 47890
tri 43340 47886 43638 48184 sw
tri 43638 47886 43936 48184 ne
rect 43936 48179 47684 48184
tri 47684 48179 47885 48380 sw
tri 47978 48179 48179 48380 ne
rect 48179 48248 49958 48380
tri 49958 48248 50090 48380 sw
tri 50250 48248 50382 48380 ne
rect 50382 48248 52230 48380
rect 48179 48179 50090 48248
rect 43936 47886 47885 48179
tri 47885 47886 48179 48179 sw
tri 48179 47886 48472 48179 ne
rect 48472 48178 50090 48179
tri 50090 48178 50160 48248 sw
tri 50382 48178 50452 48248 ne
rect 50452 48178 52230 48248
rect 48472 47886 50160 48178
tri 50160 47886 50452 48178 sw
tri 50452 47886 50744 48178 ne
rect 50744 48173 52230 48178
tri 52230 48173 52437 48380 sw
tri 52518 48173 52724 48380 ne
rect 52724 48211 56760 48380
tri 56760 48211 56930 48380 sw
tri 57086 48211 57255 48380 ne
rect 57255 48211 71000 48380
rect 52724 48173 56930 48211
rect 50744 47886 52437 48173
tri 52437 47886 52724 48173 sw
tri 52724 47886 53012 48173 ne
rect 53012 47886 56930 48173
tri 56930 47886 57255 48211 sw
tri 57255 47886 57580 48211 ne
rect 57580 47886 71000 48211
rect 39680 47601 43638 47886
rect 35437 47311 39391 47601
tri 39391 47311 39680 47601 sw
tri 39680 47311 39969 47601 ne
rect 39969 47587 43638 47601
tri 43638 47587 43936 47886 sw
tri 43936 47587 44234 47886 ne
rect 44234 47605 48179 47886
tri 48179 47605 48459 47886 sw
tri 48472 47605 48753 47886 ne
rect 48753 47605 50452 47886
rect 44234 47587 48459 47605
rect 39969 47311 43936 47587
tri 43936 47311 44212 47587 sw
tri 44234 47311 44510 47587 ne
rect 44510 47311 48459 47587
tri 48459 47311 48753 47605 sw
tri 48753 47311 49047 47605 ne
rect 49047 47603 50452 47605
tri 50452 47603 50735 47886 sw
tri 50744 47775 50855 47886 ne
rect 50855 47775 52724 47886
tri 50855 47603 51027 47775 ne
rect 51027 47603 52724 47775
rect 49047 47483 50735 47603
tri 50735 47483 50855 47603 sw
tri 51027 47483 51147 47603 ne
rect 51147 47599 52724 47603
tri 52724 47599 53011 47886 sw
tri 53012 47599 53299 47886 ne
rect 53299 47637 57255 47886
tri 57255 47637 57504 47886 sw
tri 57580 47637 57829 47886 ne
rect 57829 47637 71000 47886
rect 53299 47599 57504 47637
rect 51147 47483 53011 47599
rect 49047 47311 50855 47483
tri 50855 47311 51027 47483 sw
tri 51147 47311 51319 47483 ne
rect 51319 47311 53011 47483
tri 53011 47311 53299 47599 sw
tri 53299 47311 53586 47599 ne
rect 53586 47311 57504 47599
tri 57504 47311 57829 47637 sw
tri 57829 47311 58154 47637 ne
rect 58154 47311 71000 47637
tri 17000 47111 17200 47311 sw
tri 17293 47111 17493 47311 ne
rect 17493 47111 21536 47311
rect 14000 46993 17200 47111
tri 17200 46993 17319 47111 sw
tri 17493 46993 17612 47111 ne
rect 17612 47028 21536 47111
tri 21536 47028 21819 47311 sw
tri 21819 47028 22102 47311 ne
rect 22102 47078 26062 47311
tri 26062 47078 26296 47311 sw
tri 26360 47078 26593 47311 ne
rect 26593 47078 28340 47311
rect 22102 47028 26296 47078
rect 17612 46993 21819 47028
rect 14000 46700 17319 46993
tri 17319 46700 17612 46993 sw
tri 17612 46700 17905 46993 ne
rect 17905 46983 21819 46993
tri 21819 46983 21865 47028 sw
tri 22102 46983 22148 47028 ne
rect 22148 46983 26296 47028
rect 17905 46700 21865 46983
tri 21865 46700 22148 46983 sw
tri 22148 46700 22431 46983 ne
rect 22431 46780 26296 46983
tri 26296 46780 26593 47078 sw
tri 26593 46780 26891 47078 ne
rect 26891 47069 28340 47078
tri 28340 47069 28582 47311 sw
tri 28629 47069 28871 47311 ne
rect 28871 47071 30609 47311
tri 30609 47071 30849 47311 sw
tri 30899 47071 31140 47311 ne
rect 31140 47075 35142 47311
tri 35142 47075 35378 47311 sw
tri 35437 47075 35673 47311 ne
rect 35673 47075 39680 47311
rect 31140 47071 35378 47075
rect 28871 47069 30849 47071
rect 26891 46780 28582 47069
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46780 30849 47069
tri 30849 46780 31140 47071 sw
tri 31140 46780 31431 47071 ne
rect 31431 46780 35378 47071
tri 35378 46780 35673 47075 sw
tri 35673 46780 35969 47075 ne
rect 35969 47069 39680 47075
tri 39680 47069 39922 47311 sw
tri 39969 47069 40211 47311 ne
rect 40211 47078 44212 47311
tri 44212 47078 44445 47311 sw
tri 44510 47078 44743 47311 ne
rect 44743 47234 48753 47311
tri 48753 47234 48831 47311 sw
tri 49047 47234 49124 47311 ne
rect 49124 47234 51027 47311
rect 44743 47078 48831 47234
rect 40211 47069 44445 47078
rect 35969 46780 39922 47069
tri 39922 46780 40211 47069 sw
tri 40211 46780 40501 47069 ne
rect 40501 46780 44445 47069
tri 44445 46780 44743 47078 sw
tri 44743 46780 45042 47078 ne
rect 45042 46940 48831 47078
tri 48831 46940 49124 47234 sw
tri 49124 46940 49418 47234 ne
rect 49418 47232 51027 47234
tri 51027 47232 51106 47311 sw
tri 51319 47232 51398 47311 ne
rect 51398 47232 53299 47311
rect 49418 46940 51106 47232
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47228 53299 47232
tri 53299 47228 53382 47311 sw
tri 53586 47228 53670 47311 ne
rect 53670 47265 57829 47311
tri 57829 47265 57875 47311 sw
tri 58154 47265 58200 47311 ne
rect 58200 47265 71000 47311
rect 53670 47228 57875 47265
rect 51690 46940 53382 47228
tri 53382 46940 53670 47228 sw
tri 53670 46940 53958 47228 ne
rect 53958 46940 57875 47228
tri 57875 46940 58200 47265 sw
tri 58200 46940 58526 47265 ne
rect 58526 46940 71000 47265
rect 45042 46780 49124 46940
tri 49124 46780 49284 46940 sw
tri 49418 46780 49578 46940 ne
rect 49578 46780 51398 46940
tri 51398 46780 51558 46940 sw
tri 51690 46780 51850 46940 ne
rect 51850 46780 53670 46940
tri 53670 46780 53830 46940 sw
tri 53958 46780 54118 46940 ne
rect 54118 46780 58200 46940
tri 58200 46780 58360 46940 sw
tri 58526 46780 58686 46940 ne
rect 58686 46780 71000 46940
rect 22431 46700 26593 46780
tri 26593 46700 26674 46780 sw
tri 26891 46700 26971 46780 ne
rect 26971 46700 28871 46780
tri 28871 46700 28951 46780 sw
tri 29160 46700 29240 46780 ne
rect 29240 46771 31140 46780
tri 31140 46771 31149 46780 sw
tri 31431 46771 31439 46780 ne
rect 31439 46771 35673 46780
tri 35673 46771 35682 46780 sw
tri 35969 46771 35977 46780 ne
rect 35977 46771 40211 46780
tri 40211 46771 40220 46780 sw
tri 40501 46771 40509 46780 ne
rect 40509 46771 44743 46780
tri 44743 46771 44752 46780 sw
tri 45042 46771 45050 46780 ne
rect 45050 46771 49284 46780
tri 49284 46771 49293 46780 sw
tri 49578 46771 49587 46780 ne
rect 49587 46771 51558 46780
tri 51558 46771 51567 46780 sw
tri 51850 46771 51859 46780 ne
rect 51859 46771 53830 46780
tri 53830 46771 53839 46780 sw
tri 54118 46771 54126 46780 ne
rect 54126 46771 58360 46780
tri 58360 46771 58369 46780 sw
tri 58686 46771 58694 46780 ne
rect 58694 46771 71000 46780
rect 29240 46700 31149 46771
tri 31149 46700 31220 46771 sw
tri 31439 46700 31511 46771 ne
rect 31511 46700 35682 46771
tri 35682 46700 35754 46771 sw
tri 35977 46700 36049 46771 ne
rect 36049 46700 40220 46771
tri 40220 46700 40292 46771 sw
tri 40509 46700 40581 46771 ne
rect 40581 46700 44752 46771
tri 44752 46700 44824 46771 sw
tri 45050 46700 45122 46771 ne
rect 45122 46700 49293 46771
tri 49293 46700 49365 46771 sw
tri 49587 46700 49658 46771 ne
rect 49658 46700 51567 46771
tri 51567 46700 51638 46771 sw
tri 51859 46700 51930 46771 ne
rect 51930 46700 53839 46771
tri 53839 46700 53910 46771 sw
tri 54126 46700 54198 46771 ne
rect 54198 46700 58369 46771
tri 58369 46700 58441 46771 sw
tri 58694 46700 58766 46771 ne
rect 58766 46700 71000 46771
rect 14000 46406 17612 46700
tri 17612 46406 17905 46700 sw
tri 17905 46406 18198 46700 ne
rect 18198 46416 22148 46700
tri 22148 46416 22431 46700 sw
tri 22431 46416 22714 46700 ne
rect 22714 46482 26674 46700
tri 26674 46482 26891 46700 sw
tri 26971 46482 27189 46700 ne
rect 27189 46689 28951 46700
tri 28951 46689 28962 46700 sw
tri 29240 46689 29251 46700 ne
rect 29251 46689 31220 46700
rect 27189 46482 28962 46689
rect 22714 46416 26891 46482
rect 18198 46406 22431 46416
rect 14000 46335 17905 46406
tri 17905 46335 17976 46406 sw
tri 18198 46335 18269 46406 ne
rect 18269 46335 22431 46406
rect 14000 46069 17976 46335
tri 14000 44405 15664 46069 ne
rect 15664 46042 17976 46069
tri 17976 46042 18269 46335 sw
tri 18269 46042 18562 46335 ne
rect 18562 46315 22431 46335
tri 22431 46315 22532 46416 sw
tri 22714 46315 22815 46416 ne
rect 22815 46315 26891 46416
rect 18562 46042 22532 46315
rect 15664 45749 18269 46042
tri 18269 45749 18562 46042 sw
tri 18562 45749 18856 46042 ne
rect 18856 46032 22532 46042
tri 22532 46032 22815 46315 sw
tri 22815 46032 23098 46315 ne
rect 23098 46185 26891 46315
tri 26891 46185 27189 46482 sw
tri 27189 46185 27486 46482 ne
rect 27486 46400 28962 46482
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46481 31220 46689
tri 31220 46481 31439 46700 sw
tri 31511 46481 31730 46700 ne
rect 31730 46695 35754 46700
tri 35754 46695 35758 46700 sw
tri 36049 46695 36053 46700 ne
rect 36053 46695 40292 46700
rect 31730 46481 35758 46695
rect 29540 46400 31439 46481
tri 31439 46400 31520 46481 sw
tri 31730 46400 31811 46481 ne
rect 31811 46400 35758 46481
tri 35758 46400 36053 46695 sw
tri 36053 46400 36349 46695 ne
rect 36349 46689 40292 46695
tri 40292 46689 40302 46700 sw
tri 40581 46689 40591 46700 ne
rect 40591 46698 44824 46700
tri 44824 46698 44825 46700 sw
tri 45122 46698 45123 46700 ne
rect 45123 46698 49365 46700
rect 40591 46689 44825 46698
rect 36349 46400 40302 46689
tri 40302 46400 40591 46689 sw
tri 40591 46400 40881 46689 ne
rect 40881 46400 44825 46689
tri 44825 46400 45123 46698 sw
tri 45123 46400 45422 46698 ne
rect 45422 46646 49365 46698
tri 49365 46646 49418 46700 sw
tri 49658 46646 49712 46700 ne
rect 49712 46646 51638 46700
rect 45422 46400 49418 46646
tri 49418 46400 49664 46646 sw
tri 49712 46400 49958 46646 ne
rect 49958 46560 51638 46646
tri 51638 46560 51778 46700 sw
tri 51930 46560 52070 46700 ne
rect 52070 46560 53910 46700
tri 53910 46560 54050 46700 sw
tri 54198 46560 54338 46700 ne
rect 54338 46560 58441 46700
tri 58441 46560 58580 46700 sw
tri 58766 46560 58906 46700 ne
rect 58906 46560 71000 46700
rect 49958 46400 51778 46560
tri 51778 46400 51938 46560 sw
tri 52070 46400 52230 46560 ne
rect 52230 46400 54050 46560
tri 54050 46400 54210 46560 sw
tri 54338 46400 54498 46560 ne
rect 54498 46400 58580 46560
tri 58580 46400 58740 46560 sw
tri 58906 46400 59066 46560 ne
rect 59066 46400 71000 46560
rect 27486 46185 29251 46400
rect 23098 46047 27189 46185
tri 27189 46047 27327 46185 sw
tri 27486 46047 27624 46185 ne
rect 27624 46111 29251 46185
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46111 31520 46400
rect 27624 46047 29540 46111
rect 23098 46032 27327 46047
rect 18856 45749 22815 46032
tri 22815 45749 23098 46032 sw
tri 23098 45749 23382 46032 ne
rect 23382 45749 27327 46032
tri 27327 45749 27624 46047 sw
tri 27624 45749 27922 46047 ne
rect 27922 46038 29540 46047
tri 29540 46038 29613 46111 sw
tri 29829 46038 29902 46111 ne
rect 29902 46109 31520 46111
tri 31520 46109 31811 46400 sw
tri 31811 46109 32101 46400 ne
rect 32101 46109 36053 46400
rect 29902 46040 31811 46109
tri 31811 46040 31880 46109 sw
tri 32101 46040 32171 46109 ne
rect 32171 46105 36053 46109
tri 36053 46105 36349 46400 sw
tri 36349 46105 36644 46400 ne
rect 36644 46111 40591 46400
tri 40591 46111 40881 46400 sw
tri 40881 46111 41170 46400 ne
rect 41170 46111 45123 46400
rect 36644 46105 40881 46111
rect 32171 46044 36349 46105
tri 36349 46044 36409 46105 sw
tri 36644 46044 36704 46105 ne
rect 36704 46044 40881 46105
rect 32171 46040 36409 46044
rect 29902 46038 31880 46040
rect 27922 45749 29613 46038
tri 29613 45749 29902 46038 sw
tri 29902 45749 30191 46038 ne
rect 30191 45749 31880 46038
tri 31880 45749 32171 46040 sw
tri 32171 45749 32462 46040 ne
rect 32462 45749 36409 46040
tri 36409 45749 36704 46044 sw
tri 36704 45749 37000 46044 ne
rect 37000 46038 40881 46044
tri 40881 46038 40953 46111 sw
tri 41170 46038 41242 46111 ne
rect 41242 46102 45123 46111
tri 45123 46102 45422 46400 sw
tri 45422 46102 45720 46400 ne
rect 45720 46106 49664 46400
tri 49664 46106 49958 46400 sw
tri 49958 46106 50252 46400 ne
rect 50252 46268 51938 46400
tri 51938 46268 52070 46400 sw
tri 52230 46268 52362 46400 ne
rect 52362 46268 54210 46400
rect 50252 46106 52070 46268
rect 45720 46102 49958 46106
rect 41242 46047 45422 46102
tri 45422 46047 45476 46102 sw
tri 45720 46047 45774 46102 ne
rect 45774 46047 49958 46102
rect 41242 46038 45476 46047
rect 37000 45749 40953 46038
tri 40953 45749 41242 46038 sw
tri 41242 45749 41532 46038 ne
rect 41532 45749 45476 46038
tri 45476 45749 45774 46047 sw
tri 45774 45749 46073 46047 ne
rect 46073 46043 49958 46047
tri 49958 46043 50022 46106 sw
tri 50252 46043 50315 46106 ne
rect 50315 46043 52070 46106
rect 46073 45749 50022 46043
tri 50022 45749 50315 46043 sw
tri 50315 45749 50609 46043 ne
rect 50609 46041 52070 46043
tri 52070 46041 52297 46268 sw
tri 52362 46041 52589 46268 ne
rect 52589 46112 54210 46268
tri 54210 46112 54498 46400 sw
tri 54498 46112 54785 46400 ne
rect 54785 46325 58740 46400
tri 58740 46325 58815 46400 sw
tri 59066 46325 59140 46400 ne
rect 59140 46325 71000 46400
rect 54785 46112 58815 46325
rect 52589 46088 54498 46112
tri 54498 46088 54522 46112 sw
tri 54785 46088 54810 46112 ne
rect 54810 46088 58815 46112
rect 52589 46041 54522 46088
rect 50609 45800 52297 46041
tri 52297 45800 52538 46041 sw
tri 52589 45800 52830 46041 ne
rect 52830 45800 54522 46041
tri 54522 45800 54810 46088 sw
tri 54810 45800 55098 46088 ne
rect 55098 46000 58815 46088
tri 58815 46000 59140 46325 sw
tri 59140 46000 59466 46325 ne
rect 59466 46000 71000 46325
rect 55098 45800 59140 46000
tri 59140 45800 59340 46000 sw
rect 50609 45749 52538 45800
tri 52538 45749 52589 45800 sw
tri 52830 45749 52881 45800 ne
rect 52881 45749 54810 45800
tri 54810 45749 54861 45800 sw
tri 55098 45749 55149 45800 ne
rect 55149 45749 71000 45800
rect 15664 45657 18562 45749
tri 18562 45657 18655 45749 sw
tri 18856 45657 18948 45749 ne
rect 18948 45657 23098 45749
tri 23098 45657 23191 45749 sw
tri 23382 45657 23474 45749 ne
rect 23474 45657 27624 45749
tri 27624 45657 27717 45749 sw
tri 27922 45657 28014 45749 ne
rect 28014 45657 29902 45749
tri 29902 45657 29994 45749 sw
tri 30191 45657 30283 45749 ne
rect 30283 45657 32171 45749
tri 32171 45657 32263 45749 sw
tri 32462 45657 32554 45749 ne
rect 32554 45728 36704 45749
tri 36704 45728 36725 45749 sw
tri 37000 45728 37020 45749 ne
rect 37020 45728 41242 45749
tri 41242 45728 41263 45749 sw
tri 41532 45728 41552 45749 ne
rect 41552 45728 45774 45749
tri 45774 45728 45795 45749 sw
tri 46073 45728 46093 45749 ne
rect 46093 45728 50315 45749
tri 50315 45728 50336 45749 sw
tri 50609 45728 50630 45749 ne
rect 50630 45728 52589 45749
tri 52589 45728 52610 45749 sw
tri 52881 45728 52902 45749 ne
rect 52902 45728 54861 45749
tri 54861 45728 54882 45749 sw
tri 55149 45728 55169 45749 ne
rect 55169 45739 71000 45749
rect 55169 45728 70613 45739
rect 32554 45657 36725 45728
tri 36725 45657 36797 45728 sw
tri 37020 45657 37092 45728 ne
rect 37092 45657 41263 45728
tri 41263 45657 41335 45728 sw
tri 41552 45657 41624 45728 ne
rect 41624 45657 45795 45728
tri 45795 45657 45867 45728 sw
tri 46093 45657 46165 45728 ne
rect 46165 45657 50336 45728
tri 50336 45657 50408 45728 sw
tri 50630 45657 50701 45728 ne
rect 50701 45657 52610 45728
tri 52610 45657 52681 45728 sw
tri 52902 45657 52973 45728 ne
rect 52973 45657 54882 45728
tri 54882 45657 54953 45728 sw
tri 55169 45657 55241 45728 ne
rect 55241 45657 70613 45728
rect 15664 45364 18655 45657
tri 18655 45364 18948 45657 sw
tri 18948 45364 19241 45657 ne
rect 19241 45374 23191 45657
tri 23191 45374 23474 45657 sw
tri 23474 45374 23757 45657 ne
rect 23757 45374 27717 45657
rect 19241 45364 23474 45374
rect 15664 45070 18948 45364
tri 18948 45070 19241 45364 sw
tri 19241 45070 19534 45364 ne
rect 19534 45180 23474 45364
tri 23474 45180 23667 45374 sw
tri 23757 45180 23950 45374 ne
rect 23950 45359 27717 45374
tri 27717 45359 28014 45657 sw
tri 28014 45359 28312 45657 ne
rect 28312 45368 29994 45657
tri 29994 45368 30283 45657 sw
tri 30283 45368 30572 45657 ne
rect 30572 45368 32263 45657
rect 28312 45359 30283 45368
rect 23950 45180 28014 45359
rect 19534 45070 23667 45180
rect 15664 44991 19241 45070
tri 19241 44991 19320 45070 sw
tri 19534 44991 19614 45070 ne
rect 19614 44991 23667 45070
rect 15664 44698 19320 44991
tri 19320 44698 19614 44991 sw
tri 19614 44698 19907 44991 ne
rect 19907 44897 23667 44991
tri 23667 44897 23950 45180 sw
tri 23950 44897 24233 45180 ne
rect 24233 45098 28014 45180
tri 28014 45098 28276 45359 sw
tri 28312 45098 28573 45359 ne
rect 28573 45098 30283 45359
rect 24233 44897 28276 45098
rect 19907 44698 23950 44897
rect 15664 44405 19614 44698
tri 19614 44405 19907 44698 sw
tri 19907 44405 20200 44698 ne
rect 20200 44614 23950 44698
tri 23950 44614 24233 44897 sw
tri 24233 44614 24517 44897 ne
rect 24517 44800 28276 44897
tri 28276 44800 28573 45098 sw
tri 28573 44800 28871 45098 ne
rect 28871 45089 30283 45098
tri 30283 45089 30562 45368 sw
tri 30572 45089 30851 45368 ne
rect 30851 45366 32263 45368
tri 32263 45366 32554 45657 sw
tri 32554 45366 32844 45657 ne
rect 32844 45433 36797 45657
tri 36797 45433 37020 45657 sw
tri 37092 45433 37315 45657 ne
rect 37315 45433 41335 45657
rect 32844 45366 37020 45433
rect 30851 45091 32554 45366
tri 32554 45091 32829 45366 sw
tri 32844 45091 33120 45366 ne
rect 33120 45138 37020 45366
tri 37020 45138 37315 45433 sw
tri 37315 45138 37611 45433 ne
rect 37611 45368 41335 45433
tri 41335 45368 41624 45657 sw
tri 41624 45368 41913 45657 ne
rect 41913 45368 45867 45657
rect 37611 45138 41624 45368
rect 33120 45095 37315 45138
tri 37315 45095 37358 45138 sw
tri 37611 45095 37653 45138 ne
rect 37653 45095 41624 45138
rect 33120 45091 37358 45095
rect 30851 45089 32829 45091
rect 28871 44800 30562 45089
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 44800 32829 45089
tri 32829 44800 33120 45091 sw
tri 33120 44800 33411 45091 ne
rect 33411 44800 37358 45091
tri 37358 44800 37653 45095 sw
tri 37653 44800 37949 45095 ne
rect 37949 45089 41624 45095
tri 41624 45089 41902 45368 sw
tri 41913 45089 42191 45368 ne
rect 42191 45359 45867 45368
tri 45867 45359 46165 45657 sw
tri 46165 45359 46463 45657 ne
rect 46463 45363 50408 45657
tri 50408 45363 50701 45657 sw
tri 50701 45363 50995 45657 ne
rect 50995 45365 52681 45657
tri 52681 45365 52973 45657 sw
tri 52973 45365 53265 45657 ne
rect 53265 45512 54953 45657
tri 54953 45512 55098 45657 sw
tri 55241 45512 55385 45657 ne
rect 55385 45512 70613 45657
rect 53265 45365 55098 45512
rect 50995 45363 52973 45365
rect 46463 45359 50701 45363
rect 42191 45098 46165 45359
tri 46165 45098 46425 45359 sw
tri 46463 45098 46723 45359 ne
rect 46723 45254 50701 45359
tri 50701 45254 50811 45363 sw
tri 50995 45254 51104 45363 ne
rect 51104 45254 52973 45363
rect 46723 45098 50811 45254
rect 42191 45089 46425 45098
rect 37949 44800 41902 45089
tri 41902 44800 42191 45089 sw
tri 42191 44800 42481 45089 ne
rect 42481 44800 46425 45089
tri 46425 44800 46723 45098 sw
tri 46723 44800 47022 45098 ne
rect 47022 44960 50811 45098
tri 50811 44960 51104 45254 sw
tri 51104 44960 51398 45254 ne
rect 51398 45252 52973 45254
tri 52973 45252 53086 45365 sw
tri 53265 45252 53378 45365 ne
rect 53378 45252 55098 45365
rect 51398 44960 53086 45252
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45248 55098 45252
tri 55098 45248 55362 45512 sw
tri 55385 45248 55650 45512 ne
rect 55650 45248 70613 45512
rect 53670 44960 55362 45248
tri 55362 44960 55650 45248 sw
tri 55650 44960 55938 45248 ne
rect 55938 44960 70613 45248
rect 47022 44800 51104 44960
tri 51104 44800 51264 44960 sw
tri 51398 44800 51558 44960 ne
rect 51558 44800 53378 44960
tri 53378 44800 53538 44960 sw
tri 53670 44800 53830 44960 ne
rect 53830 44800 55650 44960
tri 55650 44800 55810 44960 sw
tri 55938 44800 56098 44960 ne
rect 56098 44800 70613 44960
rect 24517 44614 28573 44800
tri 28573 44614 28759 44800 sw
tri 28871 44614 29057 44800 ne
rect 29057 44614 30851 44800
tri 30851 44614 31037 44800 sw
tri 31140 44614 31326 44800 ne
rect 31326 44614 33120 44800
tri 33120 44614 33306 44800 sw
tri 33411 44614 33597 44800 ne
rect 33597 44614 37653 44800
tri 37653 44614 37839 44800 sw
tri 37949 44614 38135 44800 ne
rect 38135 44686 42191 44800
tri 42191 44686 42306 44800 sw
tri 42481 44686 42595 44800 ne
rect 42595 44686 46723 44800
tri 46723 44686 46838 44800 sw
tri 47022 44686 47136 44800 ne
rect 47136 44686 51264 44800
tri 51264 44686 51379 44800 sw
tri 51558 44686 51672 44800 ne
rect 51672 44686 53538 44800
tri 53538 44686 53652 44800 sw
tri 53830 44686 53944 44800 ne
rect 53944 44686 55810 44800
tri 55810 44686 55924 44800 sw
tri 56098 44686 56212 44800 ne
rect 56212 44686 70613 44800
rect 38135 44614 42306 44686
tri 42306 44614 42377 44686 sw
tri 42595 44614 42667 44686 ne
rect 42667 44614 46838 44686
tri 46838 44614 46909 44686 sw
tri 47136 44614 47208 44686 ne
rect 47208 44666 51379 44686
tri 51379 44666 51398 44686 sw
tri 51672 44666 51692 44686 ne
rect 51692 44666 53652 44686
rect 47208 44614 51398 44666
tri 51398 44614 51450 44666 sw
tri 51692 44614 51744 44666 ne
rect 51744 44614 53652 44666
tri 53652 44614 53724 44686 sw
tri 53944 44614 54016 44686 ne
rect 54016 44614 55924 44686
tri 55924 44614 55996 44686 sw
tri 56212 44614 56284 44686 ne
rect 56284 44614 70613 44686
rect 20200 44405 24233 44614
tri 15664 42457 17612 44405 ne
rect 17612 44111 19907 44405
tri 19907 44111 20200 44405 sw
tri 20200 44111 20493 44405 ne
rect 20493 44331 24233 44405
tri 24233 44331 24517 44614 sw
tri 24517 44331 24800 44614 ne
rect 24800 44502 28759 44614
tri 28759 44502 28871 44614 sw
tri 29057 44502 29169 44614 ne
rect 29169 44502 31037 44614
rect 24800 44331 28871 44502
rect 20493 44111 24517 44331
rect 17612 43818 20200 44111
tri 20200 43818 20493 44111 sw
tri 20493 43818 20786 44111 ne
rect 20786 44048 24517 44111
tri 24517 44048 24800 44331 sw
tri 24800 44048 25083 44331 ne
rect 25083 44205 28871 44331
tri 28871 44205 29169 44502 sw
tri 29169 44205 29466 44502 ne
rect 29466 44420 31037 44502
tri 31037 44420 31231 44614 sw
tri 31326 44501 31439 44614 ne
rect 31439 44501 33306 44614
tri 31439 44420 31520 44501 ne
rect 31520 44420 33306 44501
tri 33306 44420 33500 44614 sw
tri 33597 44420 33791 44614 ne
rect 33791 44420 37839 44614
tri 37839 44420 38033 44614 sw
tri 38135 44420 38329 44614 ne
rect 38329 44420 42377 44614
tri 42377 44420 42571 44614 sw
tri 42667 44420 42861 44614 ne
rect 42861 44420 46909 44614
tri 46909 44420 47103 44614 sw
tri 47208 44420 47402 44614 ne
rect 47402 44420 51450 44614
tri 51450 44420 51644 44614 sw
tri 51744 44420 51938 44614 ne
rect 51938 44580 53724 44614
tri 53724 44580 53758 44614 sw
tri 54016 44580 54050 44614 ne
rect 54050 44580 55996 44614
tri 55996 44580 56030 44614 sw
tri 56284 44580 56318 44614 ne
rect 56318 44580 70613 44614
rect 51938 44420 53758 44580
tri 53758 44420 53918 44580 sw
tri 54050 44420 54210 44580 ne
rect 54210 44420 56030 44580
tri 56030 44420 56190 44580 sw
tri 56318 44420 56478 44580 ne
rect 56478 44420 70613 44580
rect 29466 44212 31231 44420
tri 31231 44212 31439 44420 sw
tri 31520 44212 31728 44420 ne
rect 31728 44212 33500 44420
rect 29466 44205 31439 44212
rect 25083 44048 29169 44205
rect 20786 43818 24800 44048
rect 17612 43525 20493 43818
tri 20493 43525 20786 43818 sw
tri 20786 43525 21080 43818 ne
rect 21080 43764 24800 43818
tri 24800 43764 25083 44048 sw
tri 25083 43764 25366 44048 ne
rect 25366 43907 29169 44048
tri 29169 43907 29466 44205 sw
tri 29466 43907 29764 44205 ne
rect 29764 44131 31439 44205
tri 31439 44131 31520 44212 sw
tri 31728 44131 31809 44212 ne
rect 31809 44131 33500 44212
rect 29764 43907 31520 44131
rect 25366 43764 29466 43907
rect 21080 43715 25083 43764
tri 25083 43715 25133 43764 sw
tri 25366 43715 25416 43764 ne
rect 25416 43758 29466 43764
tri 29466 43758 29616 43907 sw
tri 29764 43758 29913 43907 ne
rect 29913 43842 31520 43907
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44129 33500 44131
tri 33500 44129 33791 44420 sw
tri 33791 44129 34081 44420 ne
rect 34081 44129 38033 44420
rect 32098 43842 33791 44129
rect 29913 43758 31809 43842
rect 25416 43715 29616 43758
rect 21080 43525 25133 43715
rect 17612 43451 20786 43525
tri 20786 43451 20860 43525 sw
tri 21080 43451 21153 43525 ne
rect 21153 43451 25133 43525
rect 17612 43158 20860 43451
tri 20860 43158 21153 43451 sw
tri 21153 43158 21446 43451 ne
rect 21446 43431 25133 43451
tri 25133 43431 25416 43715 sw
tri 25416 43431 25699 43715 ne
rect 25699 43460 29616 43715
tri 29616 43460 29913 43758 sw
tri 29913 43460 30211 43758 ne
rect 30211 43553 31809 43758
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43839 33791 43842
tri 33791 43839 34081 44129 sw
tri 34081 43839 34372 44129 ne
rect 34372 44125 38033 44129
tri 38033 44125 38329 44420 sw
tri 38329 44125 38624 44420 ne
rect 38624 44396 42571 44420
tri 42571 44396 42595 44420 sw
tri 42861 44396 42884 44420 ne
rect 42884 44396 47103 44420
rect 38624 44125 42595 44396
rect 34372 43839 38329 44125
rect 32387 43737 34081 43839
tri 34081 43737 34183 43839 sw
tri 34372 43737 34474 43839 ne
rect 34474 43830 38329 43839
tri 38329 43830 38624 44125 sw
tri 38624 43830 38919 44125 ne
rect 38919 44107 42595 44125
tri 42595 44107 42884 44396 sw
tri 42884 44107 43173 44396 ne
rect 43173 44122 47103 44396
tri 47103 44122 47402 44420 sw
tri 47402 44122 47700 44420 ne
rect 47700 44126 51644 44420
tri 51644 44126 51938 44420 sw
tri 51938 44126 52232 44420 ne
rect 52232 44288 53918 44420
tri 53918 44288 54050 44420 sw
tri 54210 44288 54342 44420 ne
rect 54342 44288 56190 44420
rect 52232 44126 54050 44288
rect 47700 44122 51938 44126
rect 43173 44107 47402 44122
rect 38919 43830 42884 44107
rect 34474 43751 38624 43830
tri 38624 43751 38703 43830 sw
tri 38919 43751 38998 43830 ne
rect 38998 43818 42884 43830
tri 42884 43818 43173 44107 sw
tri 43173 43818 43463 44107 ne
rect 43463 43941 47402 44107
tri 47402 43941 47582 44122 sw
tri 47700 43941 47881 44122 ne
rect 47881 43941 51938 44122
rect 43463 43818 47582 43941
rect 38998 43751 43173 43818
rect 34474 43737 38703 43751
rect 32387 43553 34183 43737
rect 30211 43460 32098 43553
rect 25699 43431 29913 43460
rect 21446 43158 25416 43431
rect 17612 42865 21153 43158
tri 21153 42865 21446 43158 sw
tri 21446 42865 21740 43158 ne
rect 21740 43148 25416 43158
tri 25416 43148 25699 43431 sw
tri 25699 43148 25982 43431 ne
rect 25982 43163 29913 43431
tri 29913 43163 30211 43460 sw
tri 30211 43163 30508 43460 ne
rect 30508 43443 32098 43460
tri 32098 43443 32208 43553 sw
tri 32387 43443 32497 43553 ne
rect 32497 43446 34183 43553
tri 34183 43446 34474 43737 sw
tri 34474 43446 34764 43737 ne
rect 34764 43455 38703 43737
tri 38703 43455 38998 43751 sw
tri 38998 43455 39293 43751 ne
rect 39293 43733 43173 43751
tri 43173 43733 43259 43818 sw
tri 43463 43733 43548 43818 ne
rect 43548 43733 47582 43818
rect 39293 43455 43259 43733
rect 34764 43446 38998 43455
rect 32497 43443 34474 43446
rect 30508 43163 32208 43443
rect 25982 43148 30211 43163
rect 21740 42865 25699 43148
tri 25699 42865 25982 43148 sw
tri 25982 42865 26266 43148 ne
rect 26266 42865 30211 43148
tri 30211 42865 30508 43163 sw
tri 30508 42865 30806 43163 ne
rect 30806 43154 32208 43163
tri 32208 43154 32497 43443 sw
tri 32497 43154 32786 43443 ne
rect 32786 43156 34474 43443
tri 34474 43156 34764 43446 sw
tri 34764 43156 35055 43446 ne
rect 35055 43160 38998 43446
tri 38998 43160 39293 43455 sw
tri 39293 43160 39588 43455 ne
rect 39588 43443 43259 43455
tri 43259 43443 43548 43733 sw
tri 43548 43443 43837 43733 ne
rect 43837 43643 47582 43733
tri 47582 43643 47881 43941 sw
tri 47881 43643 48179 43941 ne
rect 48179 43936 51938 43941
tri 51938 43936 52128 44126 sw
tri 52232 43936 52422 44126 ne
rect 52422 43996 54050 44126
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44132 56190 44288
tri 56190 44132 56478 44420 sw
tri 56478 44132 56765 44420 ne
rect 56765 44132 70613 44420
rect 54634 43996 56478 44132
rect 52422 43936 54342 43996
rect 48179 43643 52128 43936
tri 52128 43643 52422 43936 sw
tri 52422 43643 52715 43936 ne
rect 52715 43935 54342 43936
tri 54342 43935 54403 43996 sw
tri 54634 43935 54695 43996 ne
rect 54695 43935 56478 43996
rect 52715 43643 54403 43935
tri 54403 43643 54695 43935 sw
tri 54695 43643 54987 43935 ne
rect 54987 43930 56478 43935
tri 56478 43930 56680 44132 sw
tri 56765 43930 56967 44132 ne
rect 56967 43930 70613 44132
rect 54987 43643 56680 43930
tri 56680 43643 56967 43930 sw
tri 56967 43643 57255 43930 ne
rect 57255 43643 70613 43930
rect 43837 43443 47881 43643
rect 39588 43160 43548 43443
rect 35055 43156 39293 43160
rect 32786 43154 34764 43156
rect 30806 42865 32497 43154
tri 32497 42865 32786 43154 sw
tri 32786 42865 33075 43154 ne
rect 33075 42865 34764 43154
tri 34764 42865 35055 43156 sw
tri 35055 42865 35346 43156 ne
rect 35346 42865 39293 43156
tri 39293 42865 39588 43160 sw
tri 39588 42865 39884 43160 ne
rect 39884 43154 43548 43160
tri 43548 43154 43837 43443 sw
tri 43837 43154 44126 43443 ne
rect 44126 43345 47881 43443
tri 47881 43345 48179 43643 sw
tri 48179 43345 48477 43643 ne
rect 48477 43349 52422 43643
tri 52422 43349 52715 43643 sw
tri 52715 43349 53009 43643 ne
rect 53009 43351 54695 43643
tri 54695 43351 54987 43643 sw
tri 54987 43532 55098 43643 ne
rect 55098 43532 56967 43643
tri 55098 43351 55279 43532 ne
rect 55279 43355 56967 43532
tri 56967 43355 57255 43643 sw
tri 57255 43355 57542 43643 ne
rect 57542 43355 70613 43643
rect 55279 43351 57255 43355
rect 53009 43349 54987 43351
rect 48477 43345 52715 43349
rect 44126 43163 48179 43345
tri 48179 43163 48360 43345 sw
tri 48477 43163 48658 43345 ne
rect 48658 43274 52715 43345
tri 52715 43274 52791 43349 sw
tri 53009 43274 53084 43349 ne
rect 53084 43274 54987 43349
rect 48658 43163 52791 43274
rect 44126 43154 48360 43163
rect 39884 42865 43837 43154
tri 43837 42865 44126 43154 sw
tri 44126 42865 44416 43154 ne
rect 44416 42865 48360 43154
tri 48360 42865 48658 43163 sw
tri 48658 42865 48957 43163 ne
rect 48957 42980 52791 43163
tri 52791 42980 53084 43274 sw
tri 53084 42980 53378 43274 ne
rect 53378 43272 54987 43274
tri 54987 43272 55066 43351 sw
tri 55279 43272 55358 43351 ne
rect 55358 43272 57255 43351
rect 53378 43240 55066 43272
tri 55066 43240 55098 43272 sw
tri 55358 43240 55390 43272 ne
rect 55390 43268 57255 43272
tri 57255 43268 57342 43355 sw
tri 57542 43268 57630 43355 ne
rect 57630 43268 70613 43355
rect 55390 43240 57342 43268
rect 53378 42980 55098 43240
tri 55098 42980 55358 43240 sw
tri 55390 42980 55650 43240 ne
rect 55650 42980 57342 43240
tri 57342 42980 57630 43268 sw
tri 57630 42980 57918 43268 ne
rect 57918 42980 70613 43268
rect 48957 42865 53084 42980
tri 53084 42865 53199 42980 sw
tri 53378 42865 53493 42980 ne
rect 53493 42865 55358 42980
tri 55358 42865 55473 42980 sw
tri 55650 42865 55765 42980 ne
rect 55765 42865 57630 42980
tri 57630 42865 57745 42980 sw
tri 57918 42865 58033 42980 ne
rect 58033 42875 70613 42980
rect 70669 42875 71000 45739
rect 58033 42865 71000 42875
rect 17612 42800 21446 42865
tri 21446 42800 21511 42865 sw
tri 21740 42800 21804 42865 ne
rect 21804 42800 25982 42865
rect 17612 42507 21511 42800
tri 21511 42507 21804 42800 sw
tri 21804 42507 22098 42800 ne
rect 22098 42790 25982 42800
tri 25982 42790 26057 42865 sw
tri 26266 42790 26340 42865 ne
rect 26340 42820 30508 42865
tri 30508 42820 30553 42865 sw
tri 30806 42820 30851 42865 ne
rect 30851 42820 32786 42865
tri 32786 42820 32831 42865 sw
tri 33075 42820 33120 42865 ne
rect 33120 42820 35055 42865
tri 35055 42820 35100 42865 sw
tri 35346 42820 35391 42865 ne
rect 35391 42820 39588 42865
tri 39588 42820 39633 42865 sw
tri 39884 42820 39929 42865 ne
rect 39929 42820 44126 42865
tri 44126 42820 44171 42865 sw
tri 44416 42820 44461 42865 ne
rect 44461 42820 48658 42865
tri 48658 42820 48703 42865 sw
tri 48957 42820 49002 42865 ne
rect 49002 42820 53199 42865
tri 53199 42820 53244 42865 sw
tri 53493 42820 53538 42865 ne
rect 53538 42820 55473 42865
tri 55473 42820 55518 42865 sw
tri 55765 42820 55810 42865 ne
rect 55810 42820 57745 42865
tri 57745 42820 57790 42865 sw
tri 58033 42820 58078 42865 ne
rect 58078 42820 71000 42865
rect 26340 42790 30553 42820
rect 22098 42507 26057 42790
tri 26057 42507 26340 42790 sw
tri 26340 42507 26624 42790 ne
rect 26624 42522 30553 42790
tri 30553 42522 30851 42820 sw
tri 30851 42522 31149 42820 ne
rect 31149 42796 32831 42820
tri 32831 42796 32855 42820 sw
tri 33120 42796 33144 42820 ne
rect 33144 42819 35100 42820
tri 35100 42819 35101 42820 sw
tri 35391 42819 35392 42820 ne
rect 35392 42819 39633 42820
rect 33144 42796 35101 42819
rect 31149 42528 32855 42796
tri 32855 42528 33123 42796 sw
tri 33144 42528 33412 42796 ne
rect 33412 42528 35101 42796
tri 35101 42528 35392 42819 sw
tri 35392 42528 35682 42819 ne
rect 35682 42528 39633 42819
tri 39633 42528 39925 42820 sw
tri 39929 42528 40220 42820 ne
rect 40220 42818 44171 42820
tri 44171 42818 44174 42820 sw
tri 44461 42818 44463 42820 ne
rect 44463 42818 48703 42820
rect 40220 42528 44174 42818
tri 44174 42528 44463 42818 sw
tri 44463 42528 44752 42818 ne
rect 44752 42528 48703 42818
tri 48703 42528 48995 42820 sw
tri 49002 42528 49293 42820 ne
rect 49293 42686 53244 42820
tri 53244 42686 53378 42820 sw
tri 53538 42686 53672 42820 ne
rect 53672 42800 55518 42820
tri 55518 42800 55538 42820 sw
tri 55810 42800 55830 42820 ne
rect 55830 42800 57790 42820
tri 57790 42800 57810 42820 sw
tri 58078 42800 58098 42820 ne
rect 58098 42800 71000 42820
rect 53672 42686 55538 42800
rect 49293 42528 53378 42686
tri 53378 42528 53536 42686 sw
tri 53672 42528 53830 42686 ne
rect 53830 42600 55538 42686
tri 55538 42600 55738 42800 sw
tri 55830 42600 56030 42800 ne
rect 56030 42600 57810 42800
tri 57810 42600 58010 42800 sw
rect 53830 42528 55738 42600
tri 55738 42528 55810 42600 sw
tri 56030 42528 56102 42600 ne
rect 56102 42528 71000 42600
rect 31149 42522 33123 42528
rect 26624 42507 30851 42522
tri 30851 42507 30866 42522 sw
tri 31149 42507 31164 42522 ne
rect 31164 42507 33123 42522
tri 33123 42507 33144 42528 sw
tri 33412 42507 33433 42528 ne
rect 33433 42507 35392 42528
tri 35392 42507 35413 42528 sw
tri 35682 42507 35704 42528 ne
rect 35704 42507 39925 42528
tri 39925 42507 39946 42528 sw
tri 40220 42507 40242 42528 ne
rect 40242 42507 44463 42528
tri 44463 42507 44484 42528 sw
tri 44752 42507 44774 42528 ne
rect 44774 42507 48995 42528
tri 48995 42507 49016 42528 sw
tri 49293 42507 49315 42528 ne
rect 49315 42507 53536 42528
tri 53536 42507 53557 42528 sw
tri 53830 42507 53851 42528 ne
rect 53851 42507 55810 42528
tri 55810 42507 55831 42528 sw
tri 56102 42507 56123 42528 ne
rect 56123 42507 71000 42528
rect 17612 42457 21804 42507
tri 21804 42457 21855 42507 sw
tri 22098 42457 22148 42507 ne
rect 22148 42457 26340 42507
tri 26340 42457 26391 42507 sw
tri 26624 42457 26674 42507 ne
rect 26674 42457 30866 42507
tri 30866 42457 30917 42507 sw
tri 31164 42457 31214 42507 ne
rect 31214 42457 33144 42507
tri 33144 42457 33194 42507 sw
tri 33433 42457 33483 42507 ne
rect 33483 42457 35413 42507
tri 35413 42457 35463 42507 sw
tri 35704 42457 35754 42507 ne
rect 35754 42457 39946 42507
tri 39946 42457 39997 42507 sw
tri 40242 42457 40292 42507 ne
rect 40292 42457 44484 42507
tri 44484 42457 44535 42507 sw
tri 44774 42457 44824 42507 ne
rect 44824 42457 49016 42507
tri 49016 42457 49067 42507 sw
tri 49315 42457 49365 42507 ne
rect 49365 42457 53557 42507
tri 53557 42457 53608 42507 sw
tri 53851 42457 53901 42507 ne
rect 53901 42457 55831 42507
tri 55831 42457 55881 42507 sw
tri 56123 42457 56173 42507 ne
rect 56173 42497 71000 42507
rect 56173 42457 70613 42497
tri 17612 41414 18655 42457 ne
rect 18655 42164 21855 42457
tri 21855 42164 22148 42457 sw
tri 22148 42164 22441 42457 ne
rect 22441 42174 26391 42457
tri 26391 42174 26674 42457 sw
tri 26674 42174 26957 42457 ne
rect 26957 42174 30917 42457
rect 22441 42164 26674 42174
rect 18655 42000 22148 42164
tri 22148 42000 22311 42164 sw
tri 22441 42000 22604 42164 ne
rect 22604 42000 26674 42164
rect 18655 41707 22311 42000
tri 22311 41707 22604 42000 sw
tri 22604 41707 22897 42000 ne
rect 22897 41980 26674 42000
tri 26674 41980 26867 42174 sw
tri 26957 41980 27150 42174 ne
rect 27150 42159 30917 42174
tri 30917 42159 31214 42457 sw
tri 31214 42159 31512 42457 ne
rect 31512 42440 33194 42457
tri 33194 42440 33211 42457 sw
tri 33483 42440 33500 42457 ne
rect 33500 42440 35463 42457
tri 35463 42440 35480 42457 sw
tri 35754 42440 35771 42457 ne
rect 35771 42440 39997 42457
tri 39997 42440 40013 42457 sw
tri 40292 42440 40309 42457 ne
rect 40309 42440 44535 42457
tri 44535 42440 44551 42457 sw
tri 44824 42440 44841 42457 ne
rect 44841 42440 49067 42457
tri 49067 42440 49083 42457 sw
tri 49365 42440 49382 42457 ne
rect 49382 42440 53608 42457
tri 53608 42440 53624 42457 sw
tri 53901 42440 53918 42457 ne
rect 53918 42440 55881 42457
tri 55881 42440 55898 42457 sw
tri 56173 42440 56190 42457 ne
rect 56190 42440 70613 42457
rect 31512 42159 33211 42440
rect 27150 42009 31214 42159
tri 31214 42009 31364 42159 sw
tri 31512 42009 31662 42159 ne
rect 31662 42151 33211 42159
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42238 35480 42440
tri 35480 42238 35682 42440 sw
tri 35771 42238 35973 42440 ne
rect 35973 42238 40013 42440
rect 33789 42151 35682 42238
rect 31662 42009 33500 42151
rect 27150 41980 31364 42009
rect 22897 41707 26867 41980
rect 18655 41414 22604 41707
tri 22604 41414 22897 41707 sw
tri 22897 41414 23191 41707 ne
rect 23191 41697 26867 41707
tri 26867 41697 27150 41980 sw
tri 27150 41697 27433 41980 ne
rect 27433 41712 31364 41980
tri 31364 41712 31662 42009 sw
tri 31662 41712 31959 42009 ne
rect 31959 41862 33500 42009
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 41947 35682 42151
tri 35682 41947 35973 42238 sw
tri 35973 41947 36263 42238 ne
rect 36263 42145 40013 42238
tri 40013 42145 40309 42440 sw
tri 40309 42145 40604 42440 ne
rect 40604 42151 44551 42440
tri 44551 42151 44841 42440 sw
tri 44841 42151 45130 42440 ne
rect 45130 42151 49083 42440
rect 40604 42145 44841 42151
rect 36263 42076 40309 42145
tri 40309 42076 40377 42145 sw
tri 40604 42076 40673 42145 ne
rect 40673 42076 44841 42145
rect 36263 41947 40377 42076
rect 34078 41862 35973 41947
rect 31959 41712 33789 41862
rect 27433 41697 31662 41712
rect 23191 41414 27150 41697
tri 27150 41414 27433 41697 sw
tri 27433 41414 27717 41697 ne
rect 27717 41414 31662 41697
tri 31662 41414 31959 41712 sw
tri 31959 41414 32257 41712 ne
rect 32257 41703 33789 41712
tri 33789 41703 33948 41862 sw
tri 34078 41703 34237 41862 ne
rect 34237 41705 35973 41862
tri 35973 41705 36215 41947 sw
tri 36263 41705 36506 41947 ne
rect 36506 41781 40377 41947
tri 40377 41781 40673 42076 sw
tri 40673 41781 40968 42076 ne
rect 40968 42064 44841 42076
tri 44841 42064 44927 42151 sw
tri 45130 42064 45217 42151 ne
rect 45217 42142 49083 42151
tri 49083 42142 49382 42440 sw
tri 49382 42142 49680 42440 ne
rect 49680 42146 53624 42440
tri 53624 42146 53918 42440 sw
tri 53918 42146 54212 42440 ne
rect 54212 42308 55898 42440
tri 55898 42308 56030 42440 sw
tri 56190 42308 56322 42440 ne
rect 56322 42308 70613 42440
rect 54212 42146 56030 42308
rect 49680 42142 53918 42146
rect 45217 42082 49382 42142
tri 49382 42082 49441 42142 sw
tri 49680 42082 49740 42142 ne
rect 49740 42082 53918 42142
rect 45217 42064 49441 42082
rect 40968 41781 44927 42064
rect 36506 41705 40673 41781
rect 34237 41703 36215 41705
rect 32257 41414 33948 41703
tri 33948 41414 34237 41703 sw
tri 34237 41414 34526 41703 ne
rect 34526 41414 36215 41703
tri 36215 41414 36506 41705 sw
tri 36506 41414 36797 41705 ne
rect 36797 41486 40673 41705
tri 40673 41486 40968 41781 sw
tri 40968 41486 41263 41781 ne
rect 41263 41775 44927 41781
tri 44927 41775 45217 42064 sw
tri 45217 41775 45506 42064 ne
rect 45506 41784 49441 42064
tri 49441 41784 49740 42082 sw
tri 49740 41784 50038 42082 ne
rect 50038 42073 53918 42082
tri 53918 42073 53992 42146 sw
tri 54212 42073 54285 42146 ne
rect 54285 42073 56030 42146
rect 50038 41784 53992 42073
rect 45506 41775 49740 41784
rect 41263 41486 45217 41775
tri 45217 41486 45506 41775 sw
tri 45506 41486 45795 41775 ne
rect 45795 41486 49740 41775
tri 49740 41486 50038 41784 sw
tri 50038 41486 50336 41784 ne
rect 50336 41779 53992 41784
tri 53992 41779 54285 42073 sw
tri 54285 41779 54579 42073 ne
rect 54579 42016 56030 42073
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54579 41779 56322 42016
rect 50336 41486 54285 41779
tri 54285 41486 54579 41779 sw
tri 54579 41486 54872 41779 ne
rect 54872 41778 56322 41779
tri 56322 41778 56560 42016 sw
tri 56614 41778 56852 42016 ne
rect 56852 41778 70613 42016
rect 54872 41486 56560 41778
tri 56560 41486 56852 41778 sw
tri 56852 41486 57144 41778 ne
rect 57144 41486 70613 41778
rect 36797 41414 40968 41486
tri 40968 41414 41039 41486 sw
tri 41263 41414 41335 41486 ne
rect 41335 41414 45506 41486
tri 45506 41414 45577 41486 sw
tri 45795 41414 45867 41486 ne
rect 45867 41414 50038 41486
tri 50038 41414 50109 41486 sw
tri 50336 41414 50408 41486 ne
rect 50408 41414 54579 41486
tri 54579 41414 54650 41486 sw
tri 54872 41414 54944 41486 ne
rect 54944 41414 56852 41486
tri 56852 41414 56924 41486 sw
tri 57144 41414 57216 41486 ne
rect 57216 41414 70613 41486
tri 18655 38214 21855 41414 ne
rect 21855 41287 22897 41414
tri 22897 41287 23024 41414 sw
tri 23191 41287 23318 41414 ne
rect 23318 41287 27433 41414
tri 27433 41287 27560 41414 sw
tri 27717 41287 27844 41414 ne
rect 27844 41287 31959 41414
tri 31959 41287 32086 41414 sw
tri 32257 41287 32384 41414 ne
rect 32384 41287 34237 41414
tri 34237 41287 34364 41414 sw
tri 34526 41287 34653 41414 ne
rect 34653 41287 36506 41414
tri 36506 41287 36633 41414 sw
tri 36797 41287 36924 41414 ne
rect 36924 41287 41039 41414
tri 41039 41287 41166 41414 sw
tri 41335 41287 41462 41414 ne
rect 41462 41287 45577 41414
tri 45577 41287 45704 41414 sw
tri 45867 41287 45994 41414 ne
rect 45994 41287 50109 41414
tri 50109 41287 50236 41414 sw
tri 50408 41287 50535 41414 ne
rect 50535 41287 54650 41414
tri 54650 41287 54777 41414 sw
tri 54944 41287 55071 41414 ne
rect 55071 41287 56924 41414
tri 56924 41287 57051 41414 sw
tri 57216 41287 57343 41414 ne
rect 57343 41297 70613 41414
rect 70669 41297 71000 42497
rect 57343 41287 71000 41297
rect 21855 41121 23024 41287
tri 23024 41121 23191 41287 sw
tri 23318 41121 23484 41287 ne
rect 23484 41121 27560 41287
rect 21855 40828 23191 41121
tri 23191 40828 23484 41121 sw
tri 23484 40828 23777 41121 ne
rect 23777 41004 27560 41121
tri 27560 41004 27844 41287 sw
tri 27844 41004 28127 41287 ne
rect 28127 41138 32086 41287
tri 32086 41138 32236 41287 sw
tri 32384 41138 32533 41287 ne
rect 32533 41138 34364 41287
rect 28127 41004 32236 41138
rect 23777 40938 27844 41004
tri 27844 40938 27910 41004 sw
tri 28127 40938 28193 41004 ne
rect 28193 40938 32236 41004
rect 23777 40828 27910 40938
rect 21855 40534 23484 40828
tri 23484 40534 23777 40828 sw
tri 23777 40534 24070 40828 ne
rect 24070 40654 27910 40828
tri 27910 40654 28193 40938 sw
tri 28193 40654 28476 40938 ne
rect 28476 40840 32236 40938
tri 32236 40840 32533 41138 sw
tri 32533 40840 32831 41138 ne
rect 32831 41129 34364 41138
tri 34364 41129 34522 41287 sw
tri 34653 41129 34811 41287 ne
rect 34811 41131 36633 41287
tri 36633 41131 36789 41287 sw
tri 36924 41131 37080 41287 ne
rect 37080 41190 41166 41287
tri 41166 41190 41263 41287 sw
tri 41462 41190 41558 41287 ne
rect 41558 41190 45704 41287
rect 37080 41135 41263 41190
tri 41263 41135 41318 41190 sw
tri 41558 41135 41613 41190 ne
rect 41613 41135 45704 41190
rect 37080 41131 41318 41135
rect 34811 41129 36789 41131
rect 32831 40840 34522 41129
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 40840 36789 41129
tri 36789 40840 37080 41131 sw
tri 37080 40840 37371 41131 ne
rect 37371 40840 41318 41131
tri 41318 40840 41613 41135 sw
tri 41613 40840 41909 41135 ne
rect 41909 41129 45704 41135
tri 45704 41129 45862 41287 sw
tri 45994 41129 46151 41287 ne
rect 46151 41138 50236 41287
tri 50236 41138 50385 41287 sw
tri 50535 41138 50683 41287 ne
rect 50683 41138 54777 41287
rect 46151 41129 50385 41138
rect 41909 40840 45862 41129
tri 45862 40840 46151 41129 sw
tri 46151 40840 46441 41129 ne
rect 46441 40840 50385 41129
tri 50385 40840 50683 41138 sw
tri 50683 40840 50982 41138 ne
rect 50982 41000 54777 41138
tri 54777 41000 55064 41287 sw
tri 55071 41000 55358 41287 ne
rect 55358 41200 57051 41287
tri 57051 41200 57138 41287 sw
tri 57343 41200 57430 41287 ne
rect 57430 41200 71000 41287
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 50982 40840 55064 41000
tri 55064 40840 55224 41000 sw
tri 55358 40840 55518 41000 ne
rect 55518 40840 71000 41000
rect 28476 40654 32533 40840
rect 24070 40534 28193 40654
rect 21855 40241 23777 40534
tri 23777 40241 24070 40534 sw
tri 24070 40241 24363 40534 ne
rect 24363 40371 28193 40534
tri 28193 40371 28476 40654 sw
tri 28476 40371 28759 40654 ne
rect 28759 40542 32533 40654
tri 32533 40542 32831 40840 sw
tri 32831 40542 33129 40840 ne
rect 33129 40749 34811 40840
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40751 37080 40840
tri 37080 40751 37169 40840 sw
tri 37371 40751 37460 40840 ne
rect 37460 40755 41613 40840
tri 41613 40755 41698 40840 sw
tri 41909 40755 41993 40840 ne
rect 41993 40755 46151 40840
rect 37460 40751 41698 40755
rect 35191 40749 37169 40751
rect 33129 40542 34902 40749
rect 28759 40371 32831 40542
tri 32831 40371 33002 40542 sw
tri 33129 40371 33300 40542 ne
rect 33300 40460 34902 40542
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37169 40749
tri 37169 40460 37460 40751 sw
tri 37460 40460 37751 40751 ne
rect 37751 40460 41698 40751
tri 41698 40460 41993 40755 sw
tri 41993 40460 42289 40755 ne
rect 42289 40749 46151 40755
tri 46151 40749 46242 40840 sw
tri 46441 40749 46531 40840 ne
rect 46531 40758 50683 40840
tri 50683 40758 50765 40840 sw
tri 50982 40758 51063 40840 ne
rect 51063 40758 55224 40840
rect 46531 40749 50765 40758
rect 42289 40460 46242 40749
tri 46242 40460 46531 40749 sw
tri 46531 40460 46821 40749 ne
rect 46821 40460 50765 40749
tri 50765 40460 51063 40758 sw
tri 51063 40460 51362 40758 ne
rect 51362 40706 55224 40758
tri 55224 40706 55358 40840 sw
tri 55518 40706 55652 40840 ne
rect 55652 40706 71000 40840
rect 51362 40460 55358 40706
tri 55358 40460 55604 40706 sw
tri 55652 40460 55898 40706 ne
rect 55898 40460 71000 40706
rect 33300 40371 35191 40460
tri 35191 40371 35280 40460 sw
tri 35480 40371 35569 40460 ne
rect 35569 40371 37460 40460
tri 37460 40371 37549 40460 sw
tri 37751 40371 37839 40460 ne
rect 37839 40371 41993 40460
tri 41993 40371 42082 40460 sw
tri 42289 40371 42377 40460 ne
rect 42377 40443 46531 40460
tri 46531 40443 46549 40460 sw
tri 46821 40443 46838 40460 ne
rect 46838 40443 51063 40460
tri 51063 40443 51081 40460 sw
tri 51362 40443 51379 40460 ne
rect 51379 40443 55604 40460
tri 55604 40443 55622 40460 sw
tri 55898 40443 55915 40460 ne
rect 55915 40443 71000 40460
rect 42377 40371 46549 40443
tri 46549 40371 46620 40443 sw
tri 46838 40371 46909 40443 ne
rect 46909 40371 51081 40443
tri 51081 40371 51152 40443 sw
tri 51379 40371 51450 40443 ne
rect 51450 40371 55622 40443
tri 55622 40371 55693 40443 sw
tri 55915 40371 55987 40443 ne
rect 55987 40371 71000 40443
rect 24363 40241 28476 40371
rect 21855 40222 24070 40241
tri 24070 40222 24090 40241 sw
tri 24363 40222 24383 40241 ne
rect 24383 40222 28476 40241
rect 21855 39928 24090 40222
tri 24090 39928 24383 40222 sw
tri 24383 39928 24676 40222 ne
rect 24676 40088 28476 40222
tri 28476 40088 28759 40371 sw
tri 28759 40088 29043 40371 ne
rect 29043 40088 33002 40371
rect 24676 39928 28759 40088
rect 21855 39635 24383 39928
tri 24383 39635 24676 39928 sw
tri 24676 39635 24969 39928 ne
rect 24969 39805 28759 39928
tri 28759 39805 29043 40088 sw
tri 29043 39805 29326 40088 ne
rect 29326 40074 33002 40088
tri 33002 40074 33300 40371 sw
tri 33300 40074 33597 40371 ne
rect 33597 40171 35280 40371
tri 35280 40171 35480 40371 sw
tri 35569 40258 35682 40371 ne
rect 35682 40258 37549 40371
tri 35682 40171 35769 40258 ne
rect 35769 40171 37549 40258
rect 33597 40074 35480 40171
rect 29326 39937 33300 40074
tri 33300 39937 33436 40074 sw
tri 33597 39937 33734 40074 ne
rect 33734 39969 35480 40074
tri 35480 39969 35682 40171 sw
tri 35769 39969 35971 40171 ne
rect 35971 40081 37549 40171
tri 37549 40081 37839 40371 sw
tri 37839 40081 38130 40371 ne
rect 38130 40081 42082 40371
rect 35971 39969 37839 40081
rect 33734 39937 35682 39969
rect 29326 39805 33436 39937
rect 24969 39635 29043 39805
rect 21855 39342 24676 39635
tri 24676 39342 24969 39635 sw
tri 24969 39342 25263 39635 ne
rect 25263 39625 29043 39635
tri 29043 39625 29222 39805 sw
tri 29326 39625 29505 39805 ne
rect 29505 39640 33436 39805
tri 33436 39640 33734 39937 sw
tri 33734 39640 34031 39937 ne
rect 34031 39882 35682 39937
tri 35682 39882 35769 39969 sw
tri 35971 39882 36058 39969 ne
rect 36058 39923 37839 39969
tri 37839 39923 37997 40081 sw
tri 38130 39923 38287 40081 ne
rect 38287 40076 42082 40081
tri 42082 40076 42377 40371 sw
tri 42377 40076 42673 40371 ne
rect 42673 40154 46620 40371
tri 46620 40154 46838 40371 sw
tri 46909 40154 47127 40371 ne
rect 47127 40154 51152 40371
rect 42673 40076 46838 40154
rect 38287 39932 42377 40076
tri 42377 39932 42521 40076 sw
tri 42673 39932 42816 40076 ne
rect 42816 39932 46838 40076
rect 38287 39923 42521 39932
rect 36058 39882 37997 39923
rect 34031 39640 35769 39882
rect 29505 39625 33734 39640
rect 25263 39342 29222 39625
tri 29222 39342 29505 39625 sw
tri 29505 39342 29789 39625 ne
rect 29789 39342 33734 39625
tri 33734 39342 34031 39640 sw
tri 34031 39342 34329 39640 ne
rect 34329 39631 35769 39640
tri 35769 39631 36020 39882 sw
tri 36058 39631 36309 39882 ne
rect 36309 39633 37997 39882
tri 37997 39633 38287 39923 sw
tri 38287 39633 38578 39923 ne
rect 38578 39637 42521 39923
tri 42521 39637 42816 39932 sw
tri 42816 39637 43111 39932 ne
rect 43111 39864 46838 39932
tri 46838 39864 47127 40154 sw
tri 47127 39864 47416 40154 ne
rect 47416 40073 51152 40154
tri 51152 40073 51450 40371 sw
tri 51450 40073 51749 40371 ne
rect 51749 40078 55693 40371
tri 55693 40078 55987 40371 sw
tri 55987 40078 56280 40371 ne
rect 56280 40078 71000 40371
rect 51749 40073 55987 40078
rect 47416 39996 51450 40073
tri 51450 39996 51527 40073 sw
tri 51749 39996 51825 40073 ne
rect 51825 39996 55987 40073
rect 47416 39864 51527 39996
rect 43111 39637 47127 39864
rect 38578 39633 42816 39637
rect 36309 39631 38287 39633
rect 34329 39342 36020 39631
tri 36020 39342 36309 39631 sw
tri 36309 39342 36598 39631 ne
rect 36598 39342 38287 39631
tri 38287 39342 38578 39633 sw
tri 38578 39342 38869 39633 ne
rect 38869 39342 42816 39633
tri 42816 39342 43111 39637 sw
tri 43111 39342 43407 39637 ne
rect 43407 39631 47127 39637
tri 47127 39631 47360 39864 sw
tri 47416 39631 47649 39864 ne
rect 47649 39698 51527 39864
tri 51527 39698 51825 39996 sw
tri 51825 39698 52123 39996 ne
rect 52123 39894 55987 39996
tri 55987 39894 56171 40078 sw
tri 56280 39894 56464 40078 ne
rect 56464 39894 71000 40078
rect 52123 39698 56171 39894
rect 47649 39631 51825 39698
rect 43407 39342 47360 39631
tri 47360 39342 47649 39631 sw
tri 47649 39342 47939 39631 ne
rect 47939 39400 51825 39631
tri 51825 39400 52123 39698 sw
tri 52123 39400 52422 39698 ne
rect 52422 39600 56171 39698
tri 56171 39600 56464 39894 sw
tri 56464 39600 56758 39894 ne
rect 56758 39600 71000 39894
rect 52422 39400 56464 39600
tri 56464 39400 56664 39600 sw
rect 47939 39342 52123 39400
tri 52123 39342 52181 39400 sw
tri 52422 39342 52480 39400 ne
rect 52480 39342 71000 39400
rect 21855 39049 24969 39342
tri 24969 39049 25263 39342 sw
tri 25263 39049 25556 39342 ne
rect 25556 39059 29505 39342
tri 29505 39059 29789 39342 sw
tri 29789 39059 30072 39342 ne
rect 30072 39158 34031 39342
tri 34031 39158 34216 39342 sw
tri 34329 39158 34513 39342 ne
rect 34513 39158 36309 39342
rect 30072 39059 34216 39158
rect 25556 39049 29789 39059
rect 21855 38800 25263 39049
tri 25263 38800 25511 39049 sw
tri 25556 38800 25804 39049 ne
rect 25804 38800 29789 39049
rect 21855 38507 25511 38800
tri 25511 38507 25804 38800 sw
tri 25804 38507 26097 38800 ne
rect 26097 38780 29789 38800
tri 29789 38780 30067 39059 sw
tri 30072 38780 30350 39059 ne
rect 30350 38860 34216 39059
tri 34216 38860 34513 39158 sw
tri 34513 38860 34811 39158 ne
rect 34811 39149 36309 39158
tri 36309 39149 36502 39342 sw
tri 36598 39149 36791 39342 ne
rect 36791 39151 38578 39342
tri 38578 39151 38769 39342 sw
tri 38869 39151 39060 39342 ne
rect 39060 39155 43111 39342
tri 43111 39155 43298 39342 sw
tri 43407 39155 43593 39342 ne
rect 43593 39155 47649 39342
rect 39060 39151 43298 39155
rect 36791 39149 38769 39151
rect 34811 38860 36502 39149
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 38860 38769 39149
tri 38769 38860 39060 39151 sw
tri 39060 38860 39351 39151 ne
rect 39351 38860 43298 39151
tri 43298 38860 43593 39155 sw
tri 43593 38860 43889 39155 ne
rect 43889 39149 47649 39155
tri 47649 39149 47842 39342 sw
tri 47939 39149 48131 39342 ne
rect 48131 39149 52181 39342
rect 43889 38860 47842 39149
tri 47842 38860 48131 39149 sw
tri 48131 38860 48421 39149 ne
rect 48421 39102 52181 39149
tri 52181 39102 52422 39342 sw
tri 52480 39102 52720 39342 ne
rect 52720 39332 71000 39342
rect 52720 39102 70613 39332
rect 48421 38860 52422 39102
tri 52422 38860 52663 39102 sw
tri 52720 38860 52962 39102 ne
rect 52962 38860 70613 39102
rect 30350 38780 34513 38860
rect 26097 38507 30067 38780
rect 21855 38214 25804 38507
tri 25804 38214 26097 38507 sw
tri 26097 38214 26391 38507 ne
rect 26391 38497 30067 38507
tri 30067 38497 30350 38780 sw
tri 30350 38497 30633 38780 ne
rect 30633 38562 34513 38780
tri 34513 38562 34811 38860 sw
tri 34811 38562 35109 38860 ne
rect 35109 38769 36791 38860
tri 36791 38769 36882 38860 sw
tri 37080 38769 37171 38860 ne
rect 37171 38771 39060 38860
tri 39060 38771 39149 38860 sw
tri 39351 38771 39440 38860 ne
rect 39440 38775 43593 38860
tri 43593 38775 43678 38860 sw
tri 43889 38775 43973 38860 ne
rect 43973 38775 48131 38860
rect 39440 38771 43678 38775
rect 37171 38769 39149 38771
rect 35109 38562 36882 38769
rect 30633 38512 34811 38562
tri 34811 38512 34862 38562 sw
tri 35109 38512 35159 38562 ne
rect 35159 38512 36882 38562
rect 30633 38497 34862 38512
rect 26391 38214 30350 38497
tri 30350 38214 30633 38497 sw
tri 30633 38214 30917 38497 ne
rect 30917 38214 34862 38497
tri 34862 38214 35159 38512 sw
tri 35159 38214 35457 38512 ne
rect 35457 38480 36882 38512
tri 36882 38480 37171 38769 sw
tri 37171 38480 37460 38769 ne
rect 37460 38480 39149 38769
tri 39149 38480 39440 38771 sw
tri 39440 38480 39731 38771 ne
rect 39731 38480 43678 38771
tri 43678 38480 43973 38775 sw
tri 43973 38480 44269 38775 ne
rect 44269 38769 48131 38775
tri 48131 38769 48222 38860 sw
tri 48421 38769 48511 38860 ne
rect 48511 38778 52663 38860
tri 52663 38778 52745 38860 sw
tri 52962 38778 53043 38860 ne
rect 53043 38778 70613 38860
rect 48511 38769 52745 38778
rect 44269 38480 48222 38769
tri 48222 38480 48511 38769 sw
tri 48511 38480 48801 38769 ne
rect 48801 38480 52745 38769
tri 52745 38480 53043 38778 sw
tri 53043 38480 53342 38778 ne
rect 53342 38480 70613 38778
rect 35457 38286 37171 38480
tri 37171 38286 37365 38480 sw
tri 37460 38286 37654 38480 ne
rect 37654 38286 39440 38480
tri 39440 38286 39634 38480 sw
tri 39731 38286 39925 38480 ne
rect 39925 38286 43973 38480
tri 43973 38286 44168 38480 sw
tri 44269 38286 44463 38480 ne
rect 44463 38286 48511 38480
tri 48511 38286 48706 38480 sw
tri 48801 38286 48995 38480 ne
rect 48995 38286 53043 38480
tri 53043 38286 53238 38480 sw
tri 53342 38286 53536 38480 ne
rect 53536 38286 70613 38480
rect 35457 38214 37365 38286
tri 37365 38214 37437 38286 sw
tri 37654 38214 37726 38286 ne
rect 37726 38214 39634 38286
tri 39634 38214 39706 38286 sw
tri 39925 38214 39997 38286 ne
rect 39997 38214 44168 38286
tri 44168 38214 44239 38286 sw
tri 44463 38214 44535 38286 ne
rect 44535 38214 48706 38286
tri 48706 38214 48777 38286 sw
tri 48995 38214 49067 38286 ne
rect 49067 38214 53238 38286
tri 53238 38214 53309 38286 sw
tri 53536 38214 53608 38286 ne
rect 53608 38214 70613 38286
tri 21855 37171 22897 38214 ne
rect 22897 37921 26097 38214
tri 26097 37921 26391 38214 sw
tri 26391 37921 26684 38214 ne
rect 26684 37931 30633 38214
tri 30633 37931 30917 38214 sw
tri 30917 37931 31200 38214 ne
rect 31200 37931 35159 38214
rect 26684 37921 30917 37931
rect 22897 37758 26391 37921
tri 26391 37758 26554 37921 sw
tri 26684 37758 26847 37921 ne
rect 26847 37758 30917 37921
rect 22897 37464 26554 37758
tri 26554 37464 26847 37758 sw
tri 26847 37464 27140 37758 ne
rect 27140 37738 30917 37758
tri 30917 37738 31110 37931 sw
tri 31200 37738 31393 37931 ne
rect 31393 37916 35159 37931
tri 35159 37916 35457 38214 sw
tri 35457 37916 35755 38214 ne
rect 35755 38191 37437 38214
tri 37437 38191 37460 38214 sw
tri 37726 38191 37749 38214 ne
rect 37749 38191 39706 38214
rect 35755 37916 37460 38191
rect 31393 37766 35457 37916
tri 35457 37766 35607 37916 sw
tri 35755 37766 35905 37916 ne
rect 35905 37902 37460 37916
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 37995 39706 38191
tri 39706 37995 39925 38214 sw
tri 39997 37995 40216 38214 ne
rect 40216 37995 44239 38214
rect 38038 37902 39925 37995
rect 35905 37766 37749 37902
rect 31393 37738 35607 37766
rect 27140 37464 31110 37738
rect 22897 37171 26847 37464
tri 26847 37171 27140 37464 sw
tri 27140 37171 27433 37464 ne
rect 27433 37454 31110 37464
tri 31110 37454 31393 37738 sw
tri 31393 37454 31676 37738 ne
rect 31676 37469 35607 37738
tri 35607 37469 35905 37766 sw
tri 35905 37469 36202 37766 ne
rect 36202 37749 37749 37766
tri 37749 37749 37902 37902 sw
tri 38038 37749 38191 37902 ne
rect 38191 37749 39925 37902
rect 36202 37469 37902 37749
rect 31676 37454 35905 37469
rect 27433 37171 31393 37454
tri 31393 37171 31676 37454 sw
tri 31676 37171 31959 37454 ne
rect 31959 37171 35905 37454
tri 35905 37171 36202 37469 sw
tri 36202 37171 36500 37469 ne
rect 36500 37460 37902 37469
tri 37902 37460 38191 37749 sw
tri 38191 37460 38480 37749 ne
rect 38480 37704 39925 37749
tri 39925 37704 40216 37995 sw
tri 40216 37704 40506 37995 ne
rect 40506 37919 44239 37995
tri 44239 37919 44535 38214 sw
tri 44535 37919 44830 38214 ne
rect 44830 37925 48777 38214
tri 48777 37925 49067 38214 sw
tri 49067 37925 49356 38214 ne
rect 49356 37925 53309 38214
rect 44830 37919 49067 37925
rect 40506 37833 44535 37919
tri 44535 37833 44620 37919 sw
tri 44830 37833 44915 37919 ne
rect 44915 37833 49067 37919
rect 40506 37704 44620 37833
rect 38480 37462 40216 37704
tri 40216 37462 40458 37704 sw
tri 40506 37462 40749 37704 ne
rect 40749 37538 44620 37704
tri 44620 37538 44915 37833 sw
tri 44915 37538 45211 37833 ne
rect 45211 37821 49067 37833
tri 49067 37821 49170 37925 sw
tri 49356 37821 49459 37925 ne
rect 49459 37916 53309 37925
tri 53309 37916 53608 38214 sw
tri 53608 37916 53906 38214 ne
rect 53906 37916 70613 38214
rect 49459 37839 53608 37916
tri 53608 37839 53684 37916 sw
tri 53906 37839 53982 37916 ne
rect 53982 37839 70613 37916
rect 49459 37821 53684 37839
rect 45211 37538 49170 37821
rect 40749 37462 44915 37538
rect 38480 37460 40458 37462
rect 36500 37171 38191 37460
tri 38191 37171 38480 37460 sw
tri 38480 37171 38769 37460 ne
rect 38769 37171 40458 37460
tri 40458 37171 40749 37462 sw
tri 40749 37171 41039 37462 ne
rect 41039 37243 44915 37462
tri 44915 37243 45211 37538 sw
tri 45211 37243 45506 37538 ne
rect 45506 37532 49170 37538
tri 49170 37532 49459 37821 sw
tri 49459 37532 49749 37821 ne
rect 49749 37541 53684 37821
tri 53684 37541 53982 37839 sw
tri 53982 37541 54281 37839 ne
rect 54281 37541 70613 37839
rect 49749 37532 53982 37541
rect 45506 37243 49459 37532
tri 49459 37243 49749 37532 sw
tri 49749 37243 50038 37532 ne
rect 50038 37243 53982 37532
tri 53982 37243 54281 37541 sw
tri 54281 37243 54579 37541 ne
rect 54579 37243 70613 37541
rect 41039 37171 45211 37243
tri 45211 37171 45282 37243 sw
tri 45506 37171 45577 37243 ne
rect 45577 37171 49749 37243
tri 49749 37171 49820 37243 sw
tri 50038 37171 50109 37243 ne
rect 50109 37171 54281 37243
tri 54281 37171 54352 37243 sw
tri 54579 37171 54650 37243 ne
rect 54650 37171 70613 37243
tri 22897 33971 26097 37171 ne
rect 26097 36878 27140 37171
tri 27140 36878 27433 37171 sw
tri 27433 36878 27727 37171 ne
rect 27727 36888 31676 37171
tri 31676 36888 31959 37171 sw
tri 31959 36888 32243 37171 ne
rect 32243 36888 36202 37171
rect 27727 36878 31959 36888
rect 26097 36751 27433 36878
tri 27433 36751 27560 36878 sw
tri 27727 36751 27853 36878 ne
rect 27853 36751 31959 36878
rect 26097 36458 27560 36751
tri 27560 36458 27853 36751 sw
tri 27853 36458 28147 36751 ne
rect 28147 36741 31959 36751
tri 31959 36741 32106 36888 sw
tri 32243 36741 32389 36888 ne
rect 32389 36880 36202 36888
tri 36202 36880 36493 37171 sw
tri 36500 36880 36791 37171 ne
rect 36791 37169 38480 37171
tri 38480 37169 38482 37171 sw
tri 38769 37169 38771 37171 ne
rect 38771 37169 40749 37171
rect 36791 36880 38482 37169
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 36880 40749 37169
tri 40749 36880 41040 37171 sw
tri 41040 36880 41331 37171 ne
rect 41331 36948 45282 37171
tri 45282 36948 45506 37171 sw
tri 45577 36948 45801 37171 ne
rect 45801 37169 49820 37171
tri 49820 37169 49822 37171 sw
tri 50109 37169 50111 37171 ne
rect 50111 37169 54352 37171
rect 45801 36948 49822 37169
rect 41331 36880 45506 36948
tri 45506 36880 45573 36948 sw
tri 45801 36880 45869 36948 ne
rect 45869 36880 49822 36948
tri 49822 36880 50111 37169 sw
tri 50111 36880 50401 37169 ne
rect 50401 36880 54352 37169
tri 54352 36880 54643 37171 sw
tri 54650 36880 54942 37171 ne
rect 54942 36880 70613 37171
rect 32389 36741 36493 36880
rect 28147 36458 32106 36741
tri 32106 36458 32389 36741 sw
tri 32389 36458 32673 36741 ne
rect 32673 36582 36493 36741
tri 36493 36582 36791 36880 sw
tri 36791 36582 37089 36880 ne
rect 37089 36789 38771 36880
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36791 41040 36880
tri 41040 36791 41129 36880 sw
tri 41331 36791 41420 36880 ne
rect 41420 36795 45573 36880
tri 45573 36795 45658 36880 sw
tri 45869 36795 45953 36880 ne
rect 45953 36795 50111 36880
rect 41420 36791 45658 36795
rect 39151 36789 41129 36791
rect 37089 36582 38862 36789
rect 32673 36458 36791 36582
tri 36791 36458 36915 36582 sw
tri 37089 36458 37213 36582 ne
rect 37213 36500 38862 36582
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41129 36789
tri 41129 36500 41420 36791 sw
tri 41420 36500 41711 36791 ne
rect 41711 36500 45658 36791
tri 45658 36500 45953 36795 sw
tri 45953 36500 46249 36795 ne
rect 46249 36789 50111 36795
tri 50111 36789 50202 36880 sw
tri 50401 36789 50491 36880 ne
rect 50491 36798 54643 36880
tri 54643 36798 54725 36880 sw
tri 54942 36798 55023 36880 ne
rect 55023 36798 70613 36880
rect 50491 36789 54725 36798
rect 46249 36500 50202 36789
tri 50202 36500 50491 36789 sw
tri 50491 36500 50781 36789 ne
rect 50781 36500 54725 36789
tri 54725 36500 55023 36798 sw
tri 55023 36500 55322 36798 ne
rect 55322 36500 70613 36798
rect 37213 36458 39151 36500
tri 39151 36458 39193 36500 sw
tri 39440 36458 39482 36500 ne
rect 39482 36458 41420 36500
tri 41420 36458 41462 36500 sw
tri 41711 36458 41753 36500 ne
rect 41753 36458 45953 36500
tri 45953 36458 45995 36500 sw
tri 46249 36458 46291 36500 ne
rect 46291 36458 50491 36500
tri 50491 36458 50533 36500 sw
tri 50781 36458 50823 36500 ne
rect 50823 36458 55023 36500
tri 55023 36458 55065 36500 sw
tri 55322 36458 55364 36500 ne
rect 55364 36468 70613 36500
rect 70669 36468 71000 39332
rect 55364 36458 71000 36468
rect 26097 36435 27853 36458
tri 27853 36435 27876 36458 sw
tri 28147 36435 28169 36458 ne
rect 28169 36435 32389 36458
rect 26097 36142 27876 36435
tri 27876 36142 28169 36435 sw
tri 28169 36142 28463 36435 ne
rect 28463 36425 32389 36435
tri 32389 36425 32422 36458 sw
tri 32673 36425 32705 36458 ne
rect 32705 36440 36915 36458
tri 36915 36440 36934 36458 sw
tri 37213 36440 37231 36458 ne
rect 37231 36440 39193 36458
rect 32705 36425 36934 36440
rect 28463 36142 32422 36425
tri 32422 36142 32705 36425 sw
tri 32705 36142 32989 36425 ne
rect 32989 36142 36934 36425
tri 36934 36142 37231 36440 sw
tri 37231 36142 37529 36440 ne
rect 37529 36211 39193 36440
tri 39193 36211 39440 36458 sw
tri 39482 36211 39729 36458 ne
rect 39729 36433 41462 36458
tri 41462 36433 41487 36458 sw
tri 41753 36433 41778 36458 ne
rect 41778 36437 45995 36458
tri 45995 36437 46016 36458 sw
tri 46291 36437 46311 36458 ne
rect 46311 36437 50533 36458
rect 41778 36433 46016 36437
rect 39729 36211 41487 36433
rect 37529 36142 39440 36211
tri 39440 36142 39509 36211 sw
tri 39729 36142 39798 36211 ne
rect 39798 36142 41487 36211
tri 41487 36142 41778 36433 sw
tri 41778 36142 42069 36433 ne
rect 42069 36142 46016 36433
tri 46016 36142 46311 36437 sw
tri 46311 36142 46607 36437 ne
rect 46607 36200 50533 36437
tri 50533 36200 50791 36458 sw
tri 50823 36200 51081 36458 ne
rect 51081 36400 55065 36458
tri 55065 36400 55123 36458 sw
tri 55364 36400 55422 36458 ne
rect 55422 36400 71000 36458
rect 51081 36200 55123 36400
tri 55123 36200 55323 36400 sw
rect 46607 36142 50791 36200
tri 50791 36142 50849 36200 sw
tri 51081 36142 51139 36200 ne
rect 51139 36142 71000 36200
rect 26097 35849 28169 36142
tri 28169 35849 28463 36142 sw
tri 28463 35849 28756 36142 ne
rect 28756 36128 32705 36142
tri 32705 36128 32719 36142 sw
tri 32989 36128 33002 36142 ne
rect 33002 36128 37231 36142
tri 37231 36128 37245 36142 sw
tri 37529 36128 37543 36142 ne
rect 37543 36128 39509 36142
tri 39509 36128 39523 36142 sw
tri 39798 36128 39812 36142 ne
rect 39812 36128 41778 36142
tri 41778 36128 41792 36142 sw
tri 42069 36128 42082 36142 ne
rect 42082 36128 46311 36142
tri 46311 36128 46325 36142 sw
tri 46607 36128 46620 36142 ne
rect 46620 36128 50849 36142
tri 50849 36128 50863 36142 sw
tri 51139 36128 51152 36142 ne
rect 51152 36132 71000 36142
rect 51152 36128 70613 36132
rect 28756 35849 32719 36128
rect 26097 35556 28463 35849
tri 28463 35556 28756 35849 sw
tri 28756 35556 29049 35849 ne
rect 29049 35845 32719 35849
tri 32719 35845 33002 36128 sw
tri 33002 35845 33285 36128 ne
rect 33285 35845 37245 36128
rect 29049 35562 33002 35845
tri 33002 35562 33285 35845 sw
tri 33285 35562 33569 35845 ne
rect 33569 35831 37245 35845
tri 37245 35831 37543 36128 sw
tri 37543 35831 37840 36128 ne
rect 37840 35839 39523 36128
tri 39523 35839 39812 36128 sw
tri 39812 36015 39925 36128 ne
rect 39925 36015 41792 36128
tri 39925 35839 40101 36015 ne
rect 40101 35839 41792 36015
rect 37840 35831 39812 35839
rect 33569 35562 37543 35831
rect 29049 35556 33285 35562
rect 26097 35262 28756 35556
tri 28756 35262 29049 35556 sw
tri 29049 35262 29342 35556 ne
rect 29342 35279 33285 35556
tri 33285 35279 33569 35562 sw
tri 33569 35279 33852 35562 ne
rect 33852 35533 37543 35562
tri 37543 35533 37840 35831 sw
tri 37840 35533 38138 35831 ne
rect 38138 35726 39812 35831
tri 39812 35726 39925 35839 sw
tri 40101 35726 40214 35839 ne
rect 40214 35838 41792 35839
tri 41792 35838 42082 36128 sw
tri 42082 35838 42373 36128 ne
rect 42373 35838 46325 36128
rect 40214 35726 42082 35838
rect 38138 35550 39925 35726
tri 39925 35550 40101 35726 sw
tri 40214 35550 40390 35726 ne
rect 40390 35550 42082 35726
rect 38138 35533 40101 35550
rect 33852 35495 37840 35533
tri 37840 35495 37878 35533 sw
tri 38138 35495 38176 35533 ne
rect 38176 35495 40101 35533
rect 33852 35279 37878 35495
rect 29342 35262 33569 35279
rect 26097 35144 29049 35262
tri 29049 35144 29167 35262 sw
tri 29342 35144 29461 35262 ne
rect 29461 35144 33569 35262
rect 26097 34851 29167 35144
tri 29167 34851 29461 35144 sw
tri 29461 34851 29754 35144 ne
rect 29754 34996 33569 35144
tri 33569 34996 33852 35279 sw
tri 33852 34996 34135 35279 ne
rect 34135 35198 37878 35279
tri 37878 35198 38176 35495 sw
tri 38176 35198 38473 35495 ne
rect 38473 35478 40101 35495
tri 40101 35478 40173 35550 sw
tri 40390 35478 40462 35550 ne
rect 40462 35547 42082 35550
tri 42082 35547 42373 35838 sw
tri 42373 35547 42663 35838 ne
rect 42663 35833 46325 35838
tri 46325 35833 46620 36128 sw
tri 46620 35833 46915 36128 ne
rect 46915 35911 50863 36128
tri 50863 35911 51081 36128 sw
tri 51152 35911 51370 36128 ne
rect 51370 35911 70613 36128
rect 46915 35833 51081 35911
rect 42663 35547 46620 35833
rect 40462 35481 42373 35547
tri 42373 35481 42439 35547 sw
tri 42663 35481 42729 35547 ne
rect 42729 35538 46620 35547
tri 46620 35538 46915 35833 sw
tri 46915 35538 47211 35833 ne
rect 47211 35622 51081 35833
tri 51081 35622 51370 35911 sw
tri 51370 35622 51659 35911 ne
rect 51659 35622 70613 35911
rect 47211 35538 51370 35622
rect 42729 35490 46915 35538
tri 46915 35490 46963 35538 sw
tri 47211 35490 47258 35538 ne
rect 47258 35490 51370 35538
rect 42729 35481 46963 35490
rect 40462 35478 42439 35481
rect 38473 35198 40173 35478
rect 34135 34996 38176 35198
rect 29754 34851 33852 34996
rect 26097 34558 29461 34851
tri 29461 34558 29754 34851 sw
tri 29754 34558 30047 34851 ne
rect 30047 34821 33852 34851
tri 33852 34821 34027 34996 sw
tri 34135 34821 34310 34996 ne
rect 34310 34900 38176 34996
tri 38176 34900 38473 35198 sw
tri 38473 34900 38771 35198 ne
rect 38771 35189 40173 35198
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35191 42439 35478
tri 42439 35191 42729 35481 sw
tri 42729 35191 43020 35481 ne
rect 43020 35195 46963 35481
tri 46963 35195 47258 35490 sw
tri 47258 35195 47553 35490 ne
rect 47553 35478 51370 35490
tri 51370 35478 51513 35622 sw
tri 51659 35478 51802 35622 ne
rect 51802 35478 70613 35622
rect 47553 35195 51513 35478
rect 43020 35191 47258 35195
rect 40751 35189 42729 35191
rect 38771 34900 40462 35189
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34900 42729 35189
tri 42729 34900 43020 35191 sw
tri 43020 34900 43311 35191 ne
rect 43311 34900 47258 35191
tri 47258 34900 47553 35195 sw
tri 47553 34900 47849 35195 ne
rect 47849 35189 51513 35195
tri 51513 35189 51802 35478 sw
tri 51802 35189 52091 35478 ne
rect 52091 35189 70613 35478
rect 47849 34900 51802 35189
tri 51802 34900 52091 35189 sw
tri 52091 34900 52381 35189 ne
rect 52381 34900 70613 35189
rect 34310 34821 38473 34900
rect 30047 34558 34027 34821
rect 26097 34264 29754 34558
tri 29754 34264 30047 34558 sw
tri 30047 34264 30340 34558 ne
rect 30340 34538 34027 34558
tri 34027 34538 34310 34821 sw
tri 34310 34538 34593 34821 ne
rect 34593 34602 38473 34821
tri 38473 34602 38771 34900 sw
tri 38771 34602 39069 34900 ne
rect 39069 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34811 43020 34900
tri 43020 34811 43109 34900 sw
tri 43311 34811 43400 34900 ne
rect 43400 34815 47553 34900
tri 47553 34815 47638 34900 sw
tri 47849 34815 47933 34900 ne
rect 47933 34815 52091 34900
rect 43400 34811 47638 34815
rect 41131 34809 43109 34811
rect 39069 34602 40842 34809
rect 34593 34538 38771 34602
rect 30340 34264 34310 34538
rect 26097 33971 30047 34264
tri 30047 33971 30340 34264 sw
tri 30340 33971 30633 34264 ne
rect 30633 34254 34310 34264
tri 34310 34254 34593 34538 sw
tri 34593 34254 34876 34538 ne
rect 34876 34305 38771 34538
tri 38771 34305 39069 34602 sw
tri 39069 34305 39366 34602 ne
rect 39366 34520 40842 34602
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34520 43109 34809
tri 43109 34520 43400 34811 sw
tri 43400 34520 43691 34811 ne
rect 43691 34520 47638 34811
tri 47638 34520 47933 34815 sw
tri 47933 34520 48229 34815 ne
rect 48229 34809 52091 34815
tri 52091 34809 52182 34900 sw
tri 52381 34809 52471 34900 ne
rect 52471 34809 70613 34900
rect 48229 34520 52182 34809
tri 52182 34520 52471 34809 sw
tri 52471 34520 52761 34809 ne
rect 52761 34520 70613 34809
rect 39366 34305 41131 34520
rect 34876 34269 39069 34305
tri 39069 34269 39105 34305 sw
tri 39366 34269 39402 34305 ne
rect 39402 34269 41131 34305
rect 34876 34254 39105 34269
rect 30633 33971 34593 34254
tri 34593 33971 34876 34254 sw
tri 34876 33971 35159 34254 ne
rect 35159 33971 39105 34254
tri 39105 33971 39402 34269 sw
tri 39402 33971 39700 34269 ne
rect 39700 34231 41131 34269
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34333 43400 34520
tri 43400 34333 43587 34520 sw
tri 43691 34333 43877 34520 ne
rect 43877 34338 47933 34520
tri 47933 34338 48115 34520 sw
tri 48229 34338 48411 34520 ne
rect 48411 34338 52471 34520
rect 43877 34333 48115 34338
rect 41709 34231 43587 34333
rect 39700 34043 41420 34231
tri 41420 34043 41608 34231 sw
tri 41709 34043 41897 34231 ne
rect 41897 34043 43587 34231
tri 43587 34043 43877 34333 sw
tri 43877 34043 44168 34333 ne
rect 44168 34043 48115 34333
tri 48115 34043 48411 34338 sw
tri 48411 34043 48706 34338 ne
rect 48706 34332 52471 34338
tri 52471 34332 52659 34520 sw
tri 52761 34332 52949 34520 ne
rect 52949 34332 70613 34520
rect 48706 34043 52659 34332
tri 52659 34043 52949 34332 sw
tri 52949 34043 53238 34332 ne
rect 53238 34043 70613 34332
rect 39700 33971 41608 34043
tri 41608 33971 41680 34043 sw
tri 41897 33971 41969 34043 ne
rect 41969 33971 43877 34043
tri 43877 33971 43949 34043 sw
tri 44168 33971 44239 34043 ne
rect 44239 33971 48411 34043
tri 48411 33971 48482 34043 sw
tri 48706 33971 48777 34043 ne
rect 48777 33971 52949 34043
tri 52949 33971 53020 34043 sw
tri 53238 33971 53309 34043 ne
rect 53309 33971 70613 34043
tri 26097 32928 27140 33971 ne
rect 27140 33678 30340 33971
tri 30340 33678 30633 33971 sw
tri 30633 33678 30927 33971 ne
rect 30927 33688 34876 33971
tri 34876 33688 35159 33971 sw
tri 35159 33688 35443 33971 ne
rect 35443 33688 39402 33971
rect 30927 33678 35159 33688
rect 27140 33551 30633 33678
tri 30633 33551 30760 33678 sw
tri 30927 33551 31053 33678 ne
rect 31053 33551 35159 33678
rect 27140 33258 30760 33551
tri 30760 33258 31053 33551 sw
tri 31053 33258 31347 33551 ne
rect 31347 33541 35159 33551
tri 35159 33541 35306 33688 sw
tri 35443 33541 35589 33688 ne
rect 35589 33674 39402 33688
tri 39402 33674 39700 33971 sw
tri 39700 33674 39997 33971 ne
rect 39997 33682 41680 33971
tri 41680 33682 41969 33971 sw
tri 41969 33682 42258 33971 ne
rect 42258 33752 43949 33971
tri 43949 33752 44168 33971 sw
tri 44239 33752 44458 33971 ne
rect 44458 33752 48482 33971
rect 42258 33682 44168 33752
rect 39997 33674 41969 33682
rect 35589 33556 39700 33674
tri 39700 33556 39818 33674 sw
tri 39997 33556 40115 33674 ne
rect 40115 33556 41969 33674
rect 35589 33541 39818 33556
rect 31347 33258 35306 33541
tri 35306 33258 35589 33541 sw
tri 35589 33258 35873 33541 ne
rect 35873 33258 39818 33541
tri 39818 33258 40115 33556 sw
tri 40115 33258 40413 33556 ne
rect 40413 33547 41969 33556
tri 41969 33547 42104 33682 sw
tri 42258 33547 42393 33682 ne
rect 42393 33549 44168 33682
tri 44168 33549 44371 33752 sw
tri 44458 33549 44662 33752 ne
rect 44662 33676 48482 33752
tri 48482 33676 48777 33971 sw
tri 48777 33676 49073 33971 ne
rect 49073 33682 53020 33971
tri 53020 33682 53309 33971 sw
tri 53309 33682 53599 33971 ne
rect 53599 33682 70613 33971
rect 49073 33676 53309 33682
rect 44662 33553 48777 33676
tri 48777 33553 48900 33676 sw
tri 49073 33553 49195 33676 ne
rect 49195 33553 53309 33676
rect 44662 33549 48900 33553
rect 42393 33547 44371 33549
rect 40413 33258 42104 33547
tri 42104 33258 42393 33547 sw
tri 42393 33258 42682 33547 ne
rect 42682 33258 44371 33547
tri 44371 33258 44662 33549 sw
tri 44662 33258 44953 33549 ne
rect 44953 33258 48900 33549
tri 48900 33258 49195 33553 sw
tri 49195 33258 49491 33553 ne
rect 49491 33547 53309 33553
tri 53309 33547 53444 33682 sw
tri 53599 33547 53733 33682 ne
rect 53733 33547 70613 33682
rect 49491 33258 53444 33547
tri 53444 33258 53733 33547 sw
tri 53733 33258 54023 33547 ne
rect 54023 33268 70613 33547
rect 70669 33268 71000 36132
rect 54023 33258 71000 33268
rect 27140 33223 31053 33258
tri 31053 33223 31088 33258 sw
tri 31347 33223 31381 33258 ne
rect 31381 33223 35589 33258
rect 27140 32930 31088 33223
tri 31088 32930 31381 33223 sw
tri 31381 32930 31675 33223 ne
rect 31675 33213 35589 33223
tri 35589 33213 35634 33258 sw
tri 35873 33213 35917 33258 ne
rect 35917 33228 40115 33258
tri 40115 33228 40146 33258 sw
tri 40413 33228 40443 33258 ne
rect 40443 33228 42393 33258
rect 35917 33213 40146 33228
rect 31675 32930 35634 33213
tri 35634 32930 35917 33213 sw
tri 35917 32930 36201 33213 ne
rect 36201 32930 40146 33213
tri 40146 32930 40443 33228 sw
tri 40443 32930 40741 33228 ne
rect 40741 33219 42393 33228
tri 42393 33219 42432 33258 sw
tri 42682 33219 42721 33258 ne
rect 42721 33221 44662 33258
tri 44662 33221 44699 33258 sw
tri 44953 33221 44990 33258 ne
rect 44990 33221 49195 33258
rect 42721 33219 44699 33221
rect 40741 32930 42432 33219
tri 42432 32930 42721 33219 sw
tri 42721 32930 43010 33219 ne
rect 43010 32930 44699 33219
tri 44699 32930 44990 33221 sw
tri 44990 32930 45281 33221 ne
rect 45281 33000 49195 33221
tri 49195 33000 49453 33258 sw
tri 49491 33000 49749 33258 ne
rect 49749 33200 53733 33258
tri 53733 33200 53791 33258 sw
tri 54023 33200 54081 33258 ne
rect 54081 33200 71000 33258
rect 49749 33000 53791 33200
tri 53791 33000 53991 33200 sw
rect 45281 32930 49453 33000
tri 49453 32930 49523 33000 sw
tri 49749 32930 49819 33000 ne
rect 49819 32930 71000 33000
rect 27140 32928 31381 32930
tri 31381 32928 31383 32930 sw
tri 31675 32928 31676 32930 ne
rect 31676 32928 35917 32930
tri 35917 32928 35919 32930 sw
tri 36201 32928 36202 32930 ne
rect 36202 32928 40443 32930
tri 40443 32928 40445 32930 sw
tri 40741 32928 40743 32930 ne
rect 40743 32928 42721 32930
tri 42721 32928 42723 32930 sw
tri 43010 32928 43012 32930 ne
rect 43012 32928 44990 32930
tri 44990 32928 44992 32930 sw
tri 45281 32928 45282 32930 ne
rect 45282 32928 49523 32930
tri 49523 32928 49525 32930 sw
tri 49819 32928 49820 32930 ne
rect 49820 32928 71000 32930
tri 27140 29728 30340 32928 ne
rect 30340 32635 31383 32928
tri 31383 32635 31676 32928 sw
tri 31676 32635 31969 32928 ne
rect 31969 32645 35919 32928
tri 35919 32645 36202 32928 sw
tri 36202 32645 36485 32928 ne
rect 36485 32920 40445 32928
tri 40445 32920 40453 32928 sw
tri 40743 32920 40751 32928 ne
rect 40751 32920 42723 32928
tri 42723 32920 42731 32928 sw
tri 43012 32920 43020 32928 ne
rect 43020 32920 44992 32928
tri 44992 32920 45000 32928 sw
tri 45282 32920 45291 32928 ne
rect 45291 32920 49525 32928
tri 49525 32920 49533 32928 sw
tri 49820 32920 49829 32928 ne
rect 49829 32920 71000 32928
rect 36485 32645 40453 32920
rect 31969 32635 36202 32645
rect 30340 32342 31676 32635
tri 31676 32342 31969 32635 sw
tri 31969 32342 32263 32635 ne
rect 32263 32452 36202 32635
tri 36202 32452 36395 32645 sw
tri 36485 32452 36679 32645 ne
rect 36679 32622 40453 32645
tri 40453 32622 40751 32920 sw
tri 40751 32622 41049 32920 ne
rect 41049 32829 42731 32920
tri 42731 32829 42822 32920 sw
tri 43020 32829 43111 32920 ne
rect 43111 32831 45000 32920
tri 45000 32831 45089 32920 sw
tri 45291 32831 45380 32920 ne
rect 45380 32831 49533 32920
rect 43111 32829 45089 32831
rect 41049 32622 42822 32829
rect 36679 32452 40751 32622
rect 32263 32342 36395 32452
rect 30340 32049 31969 32342
tri 31969 32049 32263 32342 sw
tri 32263 32049 32556 32342 ne
rect 32556 32169 36395 32342
tri 36395 32169 36679 32452 sw
tri 36679 32169 36962 32452 ne
rect 36962 32325 40751 32452
tri 40751 32325 41049 32622 sw
tri 41049 32325 41346 32622 ne
rect 41346 32540 42822 32622
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45089 32829
tri 45089 32540 45380 32831 sw
tri 45380 32540 45671 32831 ne
rect 45671 32705 49533 32831
tri 49533 32705 49749 32920 sw
tri 49829 32705 50044 32920 ne
rect 50044 32705 70613 32920
rect 45671 32540 49749 32705
tri 49749 32540 49913 32705 sw
tri 50044 32540 50209 32705 ne
rect 50209 32540 70613 32705
rect 41346 32325 43111 32540
rect 36962 32183 41049 32325
tri 41049 32183 41190 32325 sw
tri 41346 32183 41488 32325 ne
rect 41488 32251 43111 32325
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32251 45380 32540
rect 41488 32183 43400 32251
rect 36962 32169 41190 32183
rect 32556 32049 36679 32169
rect 30340 31756 32263 32049
tri 32263 31756 32556 32049 sw
tri 32556 31756 32849 32049 ne
rect 32849 31886 36679 32049
tri 36679 31886 36962 32169 sw
tri 36962 31886 37245 32169 ne
rect 37245 31886 41190 32169
tri 41190 31886 41488 32183 sw
tri 41488 31886 41785 32183 ne
rect 41785 32175 43400 32183
tri 43400 32175 43476 32251 sw
tri 43689 32175 43765 32251 ne
rect 43765 32249 45380 32251
tri 45380 32249 45671 32540 sw
tri 45671 32249 45961 32540 ne
rect 45961 32249 49913 32540
rect 43765 32176 45671 32249
tri 45671 32176 45744 32249 sw
tri 45961 32176 46034 32249 ne
rect 46034 32245 49913 32249
tri 49913 32245 50209 32540 sw
tri 50209 32245 50504 32540 ne
rect 50504 32245 70613 32540
rect 46034 32181 50209 32245
tri 50209 32181 50273 32245 sw
tri 50504 32181 50568 32245 ne
rect 50568 32181 70613 32245
rect 46034 32176 50273 32181
rect 43765 32175 45744 32176
rect 41785 31886 43476 32175
tri 43476 31886 43765 32175 sw
tri 43765 31886 44054 32175 ne
rect 44054 31886 45744 32175
tri 45744 31886 46034 32176 sw
tri 46034 31886 46325 32176 ne
rect 46325 31886 50273 32176
tri 50273 31886 50568 32181 sw
tri 50568 31886 50863 32181 ne
rect 50863 31886 70613 32181
rect 32849 31756 36962 31886
rect 30340 31462 32556 31756
tri 32556 31462 32849 31756 sw
tri 32849 31462 33142 31756 ne
rect 33142 31602 36962 31756
tri 36962 31602 37245 31886 sw
tri 37245 31602 37528 31886 ne
rect 37528 31602 41488 31886
rect 33142 31462 37245 31602
rect 30340 31219 32849 31462
tri 32849 31219 33093 31462 sw
tri 33142 31219 33386 31462 ne
rect 33386 31319 37245 31462
tri 37245 31319 37528 31602 sw
tri 37528 31319 37811 31602 ne
rect 37811 31588 41488 31602
tri 41488 31588 41785 31886 sw
tri 41785 31588 42083 31886 ne
rect 42083 31597 43765 31886
tri 43765 31597 44054 31886 sw
tri 44054 31772 44168 31886 ne
rect 44168 31772 46034 31886
tri 44168 31597 44343 31772 ne
rect 44343 31597 46034 31772
rect 42083 31588 44054 31597
rect 37811 31535 41785 31588
tri 41785 31535 41838 31588 sw
tri 42083 31535 42136 31588 ne
rect 42136 31535 44054 31588
rect 37811 31319 41838 31535
rect 33386 31219 37528 31319
rect 30340 30926 33093 31219
tri 33093 30926 33386 31219 sw
tri 33386 30926 33679 31219 ne
rect 33679 31036 37528 31219
tri 37528 31036 37811 31319 sw
tri 37811 31036 38095 31319 ne
rect 38095 31238 41838 31319
tri 41838 31238 42136 31535 sw
tri 42136 31238 42433 31535 ne
rect 42433 31518 44054 31535
tri 44054 31518 44133 31597 sw
tri 44343 31518 44422 31597 ne
rect 44422 31595 46034 31597
tri 46034 31595 46325 31886 sw
tri 46325 31595 46616 31886 ne
rect 46616 31595 50568 31886
rect 44422 31521 46325 31595
tri 46325 31521 46399 31595 sw
tri 46616 31521 46689 31595 ne
rect 46689 31590 50568 31595
tri 50568 31590 50863 31886 sw
tri 50863 31590 51158 31886 ne
rect 51158 31590 70613 31886
rect 46689 31530 50863 31590
tri 50863 31530 50923 31590 sw
tri 51158 31530 51218 31590 ne
rect 51218 31530 70613 31590
rect 46689 31521 50923 31530
rect 44422 31518 46399 31521
rect 42433 31483 44133 31518
tri 44133 31483 44168 31518 sw
tri 44422 31483 44457 31518 ne
rect 44457 31483 46399 31518
rect 42433 31238 44168 31483
rect 38095 31036 42136 31238
rect 33679 30926 37811 31036
rect 30340 30632 33386 30926
tri 33386 30632 33679 30926 sw
tri 33679 30632 33972 30926 ne
rect 33972 30896 37811 30926
tri 37811 30896 37952 31036 sw
tri 38095 30896 38235 31036 ne
rect 38235 30940 42136 31036
tri 42136 30940 42433 31238 sw
tri 42433 30940 42731 31238 ne
rect 42731 31229 44168 31238
tri 44168 31229 44422 31483 sw
tri 44457 31229 44711 31483 ne
rect 44711 31231 46399 31483
tri 46399 31231 46689 31521 sw
tri 46689 31231 46980 31521 ne
rect 46980 31235 50923 31521
tri 50923 31235 51218 31530 sw
tri 51218 31235 51513 31530 ne
rect 51513 31235 70613 31530
rect 46980 31231 51218 31235
rect 44711 31229 46689 31231
rect 42731 30940 44422 31229
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 30940 46689 31229
tri 46689 30940 46980 31231 sw
tri 46980 30940 47271 31231 ne
rect 47271 30940 51218 31231
tri 51218 30940 51513 31235 sw
tri 51513 30940 51809 31235 ne
rect 51809 30940 70613 31235
rect 38235 30896 42433 30940
rect 33972 30632 37952 30896
rect 30340 30339 33679 30632
tri 33679 30339 33972 30632 sw
tri 33972 30339 34265 30632 ne
rect 34265 30612 37952 30632
tri 37952 30612 38235 30896 sw
tri 38235 30612 38518 30896 ne
rect 38518 30642 42433 30896
tri 42433 30642 42731 30940 sw
tri 42731 30642 43029 30940 ne
rect 43029 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30851 46980 30940
tri 46980 30851 47069 30940 sw
tri 47271 30851 47360 30940 ne
rect 47360 30855 51513 30940
tri 51513 30855 51598 30940 sw
tri 51809 30855 51893 30940 ne
rect 51893 30855 70613 30940
rect 47360 30851 51598 30855
rect 45091 30849 47069 30851
rect 43029 30642 44802 30849
rect 38518 30612 42731 30642
rect 34265 30339 38235 30612
rect 30340 30046 33972 30339
tri 33972 30046 34265 30339 sw
tri 34265 30046 34559 30339 ne
rect 34559 30329 38235 30339
tri 38235 30329 38518 30612 sw
tri 38518 30329 38801 30612 ne
rect 38801 30345 42731 30612
tri 42731 30345 43029 30642 sw
tri 43029 30345 43326 30642 ne
rect 43326 30560 44802 30642
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30560 47069 30849
tri 47069 30560 47360 30851 sw
tri 47360 30560 47651 30851 ne
rect 47651 30560 51598 30851
tri 51598 30560 51893 30855 sw
tri 51893 30560 52189 30855 ne
rect 52189 30560 70613 30855
rect 43326 30345 45091 30560
rect 38801 30344 43029 30345
tri 43029 30344 43030 30345 sw
tri 43326 30344 43327 30345 ne
rect 43327 30344 45091 30345
rect 38801 30329 43030 30344
rect 34559 30046 38518 30329
tri 38518 30046 38801 30329 sw
tri 38801 30046 39085 30329 ne
rect 39085 30046 43030 30329
tri 43030 30046 43327 30344 sw
tri 43327 30046 43625 30344 ne
rect 43625 30271 45091 30344
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30337 47360 30560
tri 47360 30337 47583 30560 sw
tri 47651 30337 47874 30560 ne
rect 47874 30341 51893 30560
tri 51893 30341 52112 30560 sw
tri 52189 30341 52407 30560 ne
rect 52407 30341 70613 30560
rect 47874 30337 52112 30341
rect 45669 30271 47583 30337
rect 43625 30046 45380 30271
tri 45380 30046 45605 30271 sw
tri 45669 30046 45894 30271 ne
rect 45894 30046 47583 30271
tri 47583 30046 47874 30337 sw
tri 47874 30046 48165 30337 ne
rect 48165 30046 52112 30337
tri 52112 30046 52407 30341 sw
tri 52407 30046 52703 30341 ne
rect 52703 30056 70613 30341
rect 70669 30056 71000 32920
rect 52703 30046 71000 30056
rect 30340 29762 34265 30046
tri 34265 29762 34549 30046 sw
tri 34559 29762 34843 30046 ne
rect 34843 30045 38801 30046
tri 38801 30045 38802 30046 sw
rect 39085 30045 43327 30046
rect 34843 29762 38802 30045
tri 38802 29762 39085 30045 sw
tri 39085 29762 39369 30045 ne
rect 39369 29762 43327 30045
tri 43327 29762 43611 30046 sw
tri 43625 29762 43909 30046 ne
rect 43909 29800 45605 30046
tri 45605 29800 45851 30046 sw
tri 45894 29800 46140 30046 ne
rect 46140 29800 47874 30046
tri 47874 29800 48120 30046 sw
tri 48165 29800 48411 30046 ne
rect 48411 30000 52407 30046
tri 52407 30000 52453 30046 sw
tri 52703 30000 52749 30046 ne
rect 52749 30000 71000 30046
rect 48411 29800 52453 30000
tri 52453 29800 52653 30000 sw
rect 43909 29762 45851 29800
tri 45851 29762 45889 29800 sw
tri 46140 29762 46178 29800 ne
rect 46178 29762 48120 29800
tri 48120 29762 48158 29800 sw
tri 48411 29762 48449 29800 ne
rect 48449 29762 71000 29800
rect 30340 29728 34549 29762
tri 34549 29728 34583 29762 sw
tri 34843 29728 34876 29762 ne
rect 34876 29728 39085 29762
tri 39085 29728 39119 29762 sw
tri 39369 29728 39402 29762 ne
rect 39402 29728 43611 29762
tri 43611 29728 43645 29762 sw
tri 43909 29728 43943 29762 ne
rect 43943 29728 45889 29762
tri 45889 29728 45923 29762 sw
tri 46178 29728 46212 29762 ne
rect 46212 29728 48158 29762
tri 48158 29728 48192 29762 sw
tri 48449 29728 48482 29762 ne
rect 48482 29752 71000 29762
rect 48482 29728 70613 29752
tri 30340 28686 31383 29728 ne
rect 31383 29435 34583 29728
tri 34583 29435 34876 29728 sw
tri 34876 29435 35169 29728 ne
rect 35169 29445 39119 29728
tri 39119 29445 39402 29728 sw
tri 39402 29445 39685 29728 ne
rect 39685 29445 43645 29728
rect 35169 29435 39402 29445
rect 31383 29272 34876 29435
tri 34876 29272 35039 29435 sw
tri 35169 29272 35333 29435 ne
rect 35333 29272 39402 29435
rect 31383 28979 35039 29272
tri 35039 28979 35333 29272 sw
tri 35333 28979 35626 29272 ne
rect 35626 29252 39402 29272
tri 39402 29252 39595 29445 sw
tri 39685 29252 39879 29445 ne
rect 39879 29431 43645 29445
tri 43645 29431 43943 29728 sw
tri 43943 29431 44240 29728 ne
rect 44240 29439 45923 29728
tri 45923 29439 46212 29728 sw
tri 46212 29439 46501 29728 ne
rect 46501 29509 48192 29728
tri 48192 29509 48411 29728 sw
tri 48482 29509 48701 29728 ne
rect 48701 29509 70613 29728
rect 46501 29439 48411 29509
rect 44240 29431 46212 29439
rect 39879 29258 43943 29431
tri 43943 29258 44116 29431 sw
tri 44240 29258 44413 29431 ne
rect 44413 29258 46212 29431
rect 39879 29252 44116 29258
rect 35626 28979 39595 29252
rect 31383 28686 35333 28979
tri 35333 28686 35626 28979 sw
tri 35626 28686 35919 28979 ne
rect 35919 28969 39595 28979
tri 39595 28969 39879 29252 sw
tri 39879 28969 40162 29252 ne
rect 40162 28969 44116 29252
rect 35919 28686 39879 28969
tri 39879 28686 40162 28969 sw
tri 40162 28686 40445 28969 ne
rect 40445 28960 44116 28969
tri 44116 28960 44413 29258 sw
tri 44413 28960 44711 29258 ne
rect 44711 29249 46212 29258
tri 46212 29249 46402 29439 sw
tri 46501 29249 46691 29439 ne
rect 46691 29251 48411 29439
tri 48411 29251 48669 29509 sw
tri 48701 29251 48960 29509 ne
rect 48960 29251 70613 29509
rect 46691 29249 48669 29251
rect 44711 28960 46402 29249
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 28960 48669 29249
tri 48669 28960 48960 29251 sw
tri 48960 28960 49251 29251 ne
rect 49251 28960 70613 29251
rect 40445 28686 44413 28960
tri 44413 28686 44688 28960 sw
tri 44711 28686 44985 28960 ne
rect 44985 28686 46691 28960
tri 46691 28686 46965 28960 sw
tri 46980 28686 47254 28960 ne
rect 47254 28686 48960 28960
tri 48960 28686 49234 28960 sw
tri 49251 28686 49525 28960 ne
rect 49525 28686 70613 28960
tri 31383 25486 34583 28686 ne
rect 34583 28392 35626 28686
tri 35626 28392 35919 28686 sw
tri 35919 28392 36212 28686 ne
rect 36212 28402 40162 28686
tri 40162 28402 40445 28686 sw
tri 40445 28402 40728 28686 ne
rect 40728 28662 44688 28686
tri 44688 28662 44711 28686 sw
tri 44985 28662 45009 28686 ne
rect 45009 28662 46965 28686
rect 40728 28402 44711 28662
rect 36212 28392 40445 28402
rect 34583 28099 35919 28392
tri 35919 28099 36212 28392 sw
tri 36212 28099 36505 28392 ne
rect 36505 28209 40445 28392
tri 40445 28209 40638 28402 sw
tri 40728 28209 40921 28402 ne
rect 40921 28365 44711 28402
tri 44711 28365 45009 28662 sw
tri 45009 28365 45306 28662 ne
rect 45306 28580 46965 28662
tri 46965 28580 47071 28686 sw
tri 47254 28580 47360 28686 ne
rect 47360 28580 49234 28686
tri 49234 28580 49340 28686 sw
tri 49525 28580 49631 28686 ne
rect 49631 28580 70613 28686
rect 45306 28365 47071 28580
rect 40921 28238 45009 28365
tri 45009 28238 45135 28365 sw
tri 45306 28238 45433 28365 ne
rect 45433 28291 47071 28365
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28291 49340 28580
rect 45433 28238 47360 28291
rect 40921 28209 45135 28238
rect 36505 28099 40638 28209
rect 34583 27806 36212 28099
tri 36212 27806 36505 28099 sw
tri 36505 27806 36799 28099 ne
rect 36799 27926 40638 28099
tri 40638 27926 40921 28209 sw
tri 40921 27926 41205 28209 ne
rect 41205 27940 45135 28209
tri 45135 27940 45433 28238 sw
tri 45433 27940 45731 28238 ne
rect 45731 28002 47360 28238
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28289 49340 28291
tri 49340 28289 49631 28580 sw
tri 49631 28289 49921 28580 ne
rect 49921 28289 70613 28580
rect 47938 28224 49631 28289
tri 49631 28224 49696 28289 sw
tri 49921 28224 49987 28289 ne
rect 49987 28224 70613 28289
rect 47938 28002 49696 28224
rect 45731 27940 47649 28002
rect 41205 27926 45433 27940
rect 36799 27806 40921 27926
rect 34583 27758 36505 27806
tri 36505 27758 36554 27806 sw
tri 36799 27758 36847 27806 ne
rect 36847 27758 40921 27806
rect 34583 27464 36554 27758
tri 36554 27464 36847 27758 sw
tri 36847 27464 37140 27758 ne
rect 37140 27643 40921 27758
tri 40921 27643 41205 27926 sw
tri 41205 27643 41488 27926 ne
rect 41488 27643 45433 27926
tri 45433 27643 45731 27940 sw
tri 45731 27643 46028 27940 ne
rect 46028 27932 47649 27940
tri 47649 27932 47719 28002 sw
tri 47938 27932 48008 28002 ne
rect 48008 27933 49696 28002
tri 49696 27933 49987 28224 sw
tri 49987 27933 50277 28224 ne
rect 50277 27933 70613 28224
rect 48008 27932 49987 27933
rect 46028 27643 47719 27932
tri 47719 27643 48008 27932 sw
tri 48008 27643 48297 27932 ne
rect 48297 27643 49987 27932
tri 49987 27643 50277 27933 sw
tri 50277 27643 50568 27933 ne
rect 50568 27643 70613 27933
rect 37140 27464 41205 27643
rect 34583 27171 36847 27464
tri 36847 27171 37140 27464 sw
tri 37140 27171 37433 27464 ne
rect 37433 27360 41205 27464
tri 41205 27360 41488 27643 sw
tri 41488 27360 41771 27643 ne
rect 41771 27360 45731 27643
rect 37433 27171 41488 27360
rect 34583 26878 37140 27171
tri 37140 26878 37433 27171 sw
tri 37433 26878 37727 27171 ne
rect 37727 27161 41488 27171
tri 41488 27161 41686 27360 sw
tri 41771 27161 41969 27360 ne
rect 41969 27345 45731 27360
tri 45731 27345 46028 27643 sw
tri 46028 27345 46326 27643 ne
rect 46326 27354 48008 27643
tri 48008 27354 48297 27643 sw
tri 48297 27529 48411 27643 ne
rect 48411 27529 50277 27643
tri 48411 27354 48586 27529 ne
rect 48586 27354 50277 27529
rect 46326 27345 48297 27354
rect 41969 27278 46028 27345
tri 46028 27278 46096 27345 sw
tri 46326 27278 46393 27345 ne
rect 46393 27278 48297 27345
rect 41969 27161 46096 27278
rect 37727 26878 41686 27161
tri 41686 26878 41969 27161 sw
tri 41969 26878 42253 27161 ne
rect 42253 26980 46096 27161
tri 46096 26980 46393 27278 sw
tri 46393 26980 46691 27278 ne
rect 46691 27269 48297 27278
tri 48297 27269 48382 27354 sw
tri 48586 27269 48671 27354 ne
rect 48671 27352 50277 27354
tri 50277 27352 50568 27643 sw
tri 50568 27352 50858 27643 ne
rect 50858 27352 70613 27643
rect 48671 27271 50568 27352
tri 50568 27271 50649 27352 sw
tri 50858 27271 50940 27352 ne
rect 50940 27271 70613 27352
rect 48671 27269 50649 27271
rect 46691 27240 48382 27269
tri 48382 27240 48411 27269 sw
tri 48671 27240 48700 27269 ne
rect 48700 27240 50649 27269
rect 46691 26980 48411 27240
tri 48411 26980 48671 27240 sw
tri 48700 26980 48960 27240 ne
rect 48960 26980 50649 27240
tri 50649 26980 50940 27271 sw
tri 50940 26980 51231 27271 ne
rect 51231 26980 70613 27271
rect 42253 26878 46393 26980
tri 46393 26878 46495 26980 sw
tri 46691 26878 46793 26980 ne
rect 46793 26878 48671 26980
tri 48671 26878 48773 26980 sw
tri 48960 26878 49062 26980 ne
rect 49062 26878 50940 26980
tri 50940 26878 51042 26980 sw
tri 51231 26878 51333 26980 ne
rect 51333 26888 70613 26980
rect 70669 26888 71000 29752
rect 51333 26878 71000 26888
rect 34583 26585 37433 26878
tri 37433 26585 37727 26878 sw
tri 37727 26585 38020 26878 ne
rect 38020 26595 41969 26878
tri 41969 26595 42253 26878 sw
tri 42253 26595 42536 26878 ne
rect 42536 26682 46495 26878
tri 46495 26682 46691 26878 sw
tri 46793 26682 46989 26878 ne
rect 46989 26800 48773 26878
tri 48773 26800 48851 26878 sw
tri 49062 26800 49140 26878 ne
rect 49140 26800 51042 26878
tri 51042 26800 51120 26878 sw
tri 51333 26800 51411 26878 ne
rect 51411 26800 71000 26878
rect 46989 26682 48851 26800
rect 42536 26595 46691 26682
rect 38020 26585 42253 26595
rect 34583 26292 37727 26585
tri 37727 26292 38020 26585 sw
tri 38020 26292 38313 26585 ne
rect 38313 26312 42253 26585
tri 42253 26312 42536 26595 sw
tri 42536 26312 42819 26595 ne
rect 42819 26385 46691 26595
tri 46691 26385 46989 26682 sw
tri 46989 26385 47286 26682 ne
rect 47286 26600 48851 26682
tri 48851 26600 49051 26800 sw
tri 49140 26600 49340 26800 ne
rect 49340 26600 51120 26800
tri 51120 26600 51320 26800 sw
rect 47286 26385 49051 26600
rect 42819 26312 46989 26385
rect 38313 26292 42536 26312
rect 34583 26072 38020 26292
tri 38020 26072 38239 26292 sw
tri 38313 26072 38533 26292 ne
rect 38533 26072 42536 26292
rect 34583 25779 38239 26072
tri 38239 25779 38533 26072 sw
tri 38533 25779 38826 26072 ne
rect 38826 26052 42536 26072
tri 42536 26052 42795 26312 sw
tri 42819 26052 43079 26312 ne
rect 43079 26087 46989 26312
tri 46989 26087 47286 26385 sw
tri 47286 26087 47584 26385 ne
rect 47584 26311 49051 26385
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47584 26087 49340 26311
rect 43079 26081 47286 26087
tri 47286 26081 47293 26087 sw
tri 47584 26081 47590 26087 ne
rect 47590 26081 49340 26087
rect 43079 26052 47293 26081
rect 38826 25779 42795 26052
rect 34583 25486 38533 25779
tri 38533 25486 38826 25779 sw
tri 38826 25486 39119 25779 ne
rect 39119 25769 42795 25779
tri 42795 25769 43079 26052 sw
tri 43079 25769 43362 26052 ne
rect 43362 25783 47293 26052
tri 47293 25783 47590 26081 sw
tri 47590 25783 47888 26081 ne
rect 47888 26022 49340 26081
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47888 25783 49629 26022
rect 43362 25769 47590 25783
rect 39119 25486 43079 25769
tri 43079 25486 43362 25769 sw
tri 43362 25486 43645 25769 ne
rect 43645 25486 47590 25769
tri 47590 25486 47888 25783 sw
tri 47888 25486 48185 25783 ne
rect 48185 25775 49629 25783
tri 49629 25775 49876 26022 sw
tri 49918 25775 50165 26022 ne
rect 50165 25775 71000 26022
rect 48185 25486 49876 25775
tri 49876 25486 50165 25775 sw
tri 50165 25486 50454 25775 ne
rect 50454 25486 71000 25775
tri 34583 24443 35626 25486 ne
rect 35626 25209 38826 25486
tri 38826 25209 39102 25486 sw
tri 39119 25209 39395 25486 ne
rect 39395 25209 43362 25486
rect 35626 24916 39102 25209
tri 39102 24916 39395 25209 sw
tri 39395 24916 39689 25209 ne
rect 39689 25202 43362 25209
tri 43362 25202 43645 25486 sw
tri 43645 25202 43928 25486 ne
rect 43928 25298 47888 25486
tri 47888 25298 48076 25486 sw
tri 48185 25298 48373 25486 ne
rect 48373 25298 50165 25486
rect 43928 25202 48076 25298
rect 39689 25199 43645 25202
tri 43645 25199 43648 25202 sw
tri 43928 25199 43931 25202 ne
rect 43931 25199 48076 25202
rect 39689 24916 43648 25199
tri 43648 24916 43931 25199 sw
tri 43931 24916 44215 25199 ne
rect 44215 25000 48076 25199
tri 48076 25000 48373 25298 sw
tri 48373 25000 48671 25298 ne
rect 48671 25200 50165 25298
tri 50165 25200 50451 25486 sw
tri 50454 25200 50740 25486 ne
rect 50740 25200 71000 25486
rect 48671 25000 50451 25200
tri 50451 25000 50651 25200 sw
rect 44215 24916 48373 25000
tri 48373 24916 48457 25000 sw
tri 48671 24916 48755 25000 ne
rect 48755 24916 71000 25000
rect 35626 24736 39395 24916
tri 39395 24736 39575 24916 sw
tri 39689 24736 39869 24916 ne
rect 39869 24736 43931 24916
rect 35626 24443 39575 24736
tri 39575 24443 39869 24736 sw
tri 39869 24443 40162 24736 ne
rect 40162 24726 43931 24736
tri 43931 24726 44121 24916 sw
tri 44215 24726 44405 24916 ne
rect 44405 24726 48457 24916
rect 40162 24443 44121 24726
tri 44121 24443 44405 24726 sw
tri 44405 24443 44688 24726 ne
rect 44688 24702 48457 24726
tri 48457 24702 48671 24916 sw
tri 48755 24702 48969 24916 ne
rect 48969 24906 71000 24916
rect 48969 24702 70613 24906
rect 44688 24443 48671 24702
tri 48671 24443 48931 24702 sw
tri 48969 24443 49228 24702 ne
rect 49228 24443 70613 24702
tri 35626 21243 38826 24443 ne
rect 38826 24150 39869 24443
tri 39869 24150 40162 24443 sw
tri 40162 24150 40455 24443 ne
rect 40455 24160 44405 24443
tri 44405 24160 44688 24443 sw
tri 44688 24160 44971 24443 ne
rect 44971 24160 48931 24443
rect 40455 24150 44688 24160
rect 38826 23989 40162 24150
tri 40162 23989 40322 24150 sw
tri 40455 23989 40615 24150 ne
rect 40615 23989 44688 24150
rect 38826 23696 40322 23989
tri 40322 23696 40615 23989 sw
tri 40615 23696 40909 23989 ne
rect 40909 23979 44688 23989
tri 44688 23979 44868 24160 sw
tri 44971 23979 45151 24160 ne
rect 45151 24145 48931 24160
tri 48931 24145 49228 24443 sw
tri 49228 24145 49526 24443 ne
rect 49526 24145 70613 24443
rect 45151 23994 49228 24145
tri 49228 23994 49380 24145 sw
tri 49526 23994 49677 24145 ne
rect 49677 23994 70613 24145
rect 45151 23979 49380 23994
rect 40909 23696 44868 23979
tri 44868 23696 45151 23979 sw
tri 45151 23696 45435 23979 ne
rect 45435 23696 49380 23979
tri 49380 23696 49677 23994 sw
tri 49677 23696 49975 23994 ne
rect 49975 23706 70613 23994
rect 70669 23706 71000 24906
rect 49975 23696 71000 23706
rect 38826 23403 40615 23696
tri 40615 23403 40909 23696 sw
tri 40909 23403 41202 23696 ne
rect 41202 23683 45151 23696
tri 45151 23683 45164 23696 sw
tri 45435 23683 45447 23696 ne
rect 45447 23683 49677 23696
rect 41202 23403 45164 23683
rect 38826 23110 40909 23403
tri 40909 23110 41202 23403 sw
tri 41202 23400 41205 23403 ne
rect 41205 23400 45164 23403
tri 45164 23400 45447 23683 sw
tri 45447 23400 45731 23683 ne
rect 45731 23600 49677 23683
tri 49677 23600 49773 23696 sw
tri 49975 23600 50071 23696 ne
rect 50071 23600 71000 23696
rect 45731 23400 49773 23600
tri 49773 23400 49973 23600 sw
tri 41205 23110 41495 23400 ne
rect 41495 23117 45447 23400
tri 45447 23117 45731 23400 sw
tri 45731 23117 46014 23400 ne
rect 46014 23117 71000 23400
rect 41495 23110 45731 23117
rect 38826 22816 41202 23110
tri 41202 22816 41495 23110 sw
tri 41495 22816 41788 23110 ne
rect 41788 22834 45731 23110
tri 45731 22834 46014 23117 sw
tri 46014 22834 46297 23117 ne
rect 46297 22834 71000 23117
rect 41788 22816 46014 22834
rect 38826 22523 41495 22816
tri 41495 22523 41788 22816 sw
tri 41788 22523 42081 22816 ne
rect 42081 22550 46014 22816
tri 46014 22550 46297 22834 sw
tri 46297 22550 46580 22834 ne
rect 46580 22550 71000 22834
rect 42081 22523 46297 22550
rect 38826 22416 41788 22523
tri 41788 22416 41896 22523 sw
tri 42081 22416 42189 22523 ne
rect 42189 22416 46297 22523
rect 38826 22122 41896 22416
tri 41896 22122 42189 22416 sw
tri 42189 22122 42482 22416 ne
rect 42482 22267 46297 22416
tri 46297 22267 46580 22550 sw
tri 46580 22267 46863 22550 ne
rect 46863 22267 71000 22550
rect 42482 22122 46580 22267
rect 38826 21829 42189 22122
tri 42189 21829 42482 22122 sw
tri 42482 21829 42775 22122 ne
rect 42775 22092 46580 22122
tri 46580 22092 46755 22267 sw
tri 46863 22092 47038 22267 ne
rect 47038 22092 71000 22267
rect 42775 21829 46755 22092
rect 38826 21536 42482 21829
tri 42482 21536 42775 21829 sw
tri 42775 21536 43069 21829 ne
rect 43069 21809 46755 21829
tri 46755 21809 47038 22092 sw
tri 47038 21809 47321 22092 ne
rect 47321 21809 71000 22092
rect 43069 21536 47038 21809
rect 38826 21243 42775 21536
tri 42775 21243 43069 21536 sw
tri 43069 21243 43362 21536 ne
rect 43362 21526 47038 21536
tri 47038 21526 47321 21809 sw
tri 47321 21526 47605 21809 ne
rect 47605 21526 71000 21809
rect 43362 21243 47321 21526
tri 47321 21243 47605 21526 sw
tri 47605 21243 47888 21526 ne
rect 47888 21243 71000 21526
tri 38826 20200 39869 21243 ne
rect 39869 20950 43069 21243
tri 43069 20950 43362 21243 sw
tri 43362 20950 43655 21243 ne
rect 43655 20960 47605 21243
tri 47605 20960 47888 21243 sw
tri 47888 20960 48171 21243 ne
rect 48171 20960 71000 21243
rect 43655 20950 47888 20960
rect 39869 20786 43362 20950
tri 43362 20786 43525 20950 sw
tri 43655 20786 43818 20950 ne
rect 43818 20786 47888 20950
rect 39869 20493 43525 20786
tri 43525 20493 43818 20786 sw
tri 43818 20493 44111 20786 ne
rect 44111 20683 47888 20786
tri 47888 20683 48164 20960 sw
tri 48171 20683 48447 20960 ne
rect 48447 20683 71000 20960
rect 44111 20493 48164 20683
rect 39869 20200 43818 20493
tri 43818 20200 44111 20493 sw
tri 44111 20200 44405 20493 ne
rect 44405 20400 48164 20493
tri 48164 20400 48447 20683 sw
tri 48447 20400 48731 20683 ne
rect 48731 20400 71000 20683
rect 44405 20200 48447 20400
tri 48447 20200 48647 20400 sw
tri 39869 17000 43069 20200 ne
rect 43069 19907 44111 20200
tri 44111 19907 44405 20200 sw
tri 44405 19907 44698 20200 ne
rect 44698 19907 71000 20200
rect 43069 19614 44405 19907
tri 44405 19614 44698 19907 sw
tri 44698 19614 44991 19907 ne
rect 44991 19614 71000 19907
rect 43069 19320 44698 19614
tri 44698 19320 44991 19614 sw
tri 44991 19320 45284 19614 ne
rect 45284 19320 71000 19614
rect 43069 19027 44991 19320
tri 44991 19027 45284 19320 sw
tri 45284 19027 45577 19320 ne
rect 45577 19027 71000 19320
rect 43069 18734 45284 19027
tri 45284 18734 45577 19027 sw
tri 45577 18734 45871 19027 ne
rect 45871 18734 71000 19027
rect 43069 18666 45577 18734
tri 45577 18666 45645 18734 sw
tri 45871 18666 45939 18734 ne
rect 45939 18666 71000 18734
rect 43069 18373 45645 18666
tri 45645 18373 45939 18666 sw
tri 45939 18373 46232 18666 ne
rect 46232 18373 71000 18666
rect 43069 18080 45939 18373
tri 45939 18080 46232 18373 sw
tri 46232 18080 46525 18373 ne
rect 46525 18080 71000 18373
rect 43069 17786 46232 18080
tri 46232 17786 46525 18080 sw
tri 46525 17786 46818 18080 ne
rect 46818 17786 71000 18080
rect 43069 17493 46525 17786
tri 46525 17493 46818 17786 sw
tri 46818 17493 47111 17786 ne
rect 47111 17493 71000 17786
rect 43069 17200 46818 17493
tri 46818 17200 47111 17493 sw
tri 47111 17200 47405 17493 ne
rect 47405 17200 71000 17493
rect 43069 17000 47111 17200
tri 47111 17000 47311 17200 sw
tri 43069 14000 46069 17000 ne
rect 46069 14000 71000 17000
use M1_PSUB_CDNS_406619561340  M1_PSUB_CDNS_406619561340_0
timestamp 1669390400
transform -1 0 58007 0 -1 13194
box 0 0 1 1
use M1_PSUB_CDNS_406619561341  M1_PSUB_CDNS_406619561341_0
timestamp 1669390400
transform 0 -1 69871 1 0 70385
box 0 0 1 1
use M1_PSUB_CDNS_406619561342  M1_PSUB_CDNS_406619561342_0
timestamp 1669390400
transform 1 0 70235 0 1 69871
box 0 0 1 1
use M1_PSUB_CDNS_406619561343  M1_PSUB_CDNS_406619561343_0
timestamp 1669390400
transform 0 -1 70899 1 0 41649
box 0 0 1 1
use M1_PSUB_CDNS_406619561343  M1_PSUB_CDNS_406619561343_1
timestamp 1669390400
transform 1 0 41636 0 1 70900
box 0 0 1 1
use M1_PSUB_CDNS_406619561344  M1_PSUB_CDNS_406619561344_0
timestamp 1669390400
transform 0 -1 13194 1 0 58004
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_0
timestamp 1669390400
transform 1 0 44693 0 1 13385
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_1
timestamp 1669390400
transform 1 0 44561 0 1 13517
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_2
timestamp 1669390400
transform 1 0 44429 0 1 13649
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_3
timestamp 1669390400
transform 1 0 44297 0 1 13781
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_4
timestamp 1669390400
transform 1 0 44165 0 1 13913
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_5
timestamp 1669390400
transform 1 0 44033 0 1 14045
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_6
timestamp 1669390400
transform 1 0 43901 0 1 14177
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_7
timestamp 1669390400
transform 1 0 43769 0 1 14309
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_8
timestamp 1669390400
transform 1 0 43637 0 1 14441
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_9
timestamp 1669390400
transform 1 0 43505 0 1 14573
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_10
timestamp 1669390400
transform 1 0 43373 0 1 14705
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_11
timestamp 1669390400
transform 1 0 43241 0 1 14837
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_12
timestamp 1669390400
transform 1 0 43109 0 1 14969
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_13
timestamp 1669390400
transform 1 0 42845 0 1 15233
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_14
timestamp 1669390400
transform 1 0 42713 0 1 15365
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_15
timestamp 1669390400
transform 1 0 42581 0 1 15497
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_16
timestamp 1669390400
transform 1 0 42449 0 1 15629
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_17
timestamp 1669390400
transform 1 0 42317 0 1 15761
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_18
timestamp 1669390400
transform 1 0 42185 0 1 15893
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_19
timestamp 1669390400
transform 1 0 42977 0 1 15101
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_20
timestamp 1669390400
transform 1 0 44873 0 1 13233
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_21
timestamp 1669390400
transform 1 0 38885 0 1 19193
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_22
timestamp 1669390400
transform 1 0 38753 0 1 19325
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_23
timestamp 1669390400
transform 1 0 38621 0 1 19457
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_24
timestamp 1669390400
transform 1 0 38489 0 1 19589
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_25
timestamp 1669390400
transform 1 0 38357 0 1 19721
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_26
timestamp 1669390400
transform 1 0 33869 0 1 24209
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_27
timestamp 1669390400
transform 1 0 34001 0 1 24077
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_28
timestamp 1669390400
transform 1 0 34133 0 1 23945
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_29
timestamp 1669390400
transform 1 0 34265 0 1 23813
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_30
timestamp 1669390400
transform 1 0 34397 0 1 23681
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_31
timestamp 1669390400
transform 1 0 34529 0 1 23549
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_32
timestamp 1669390400
transform 1 0 34661 0 1 23417
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_33
timestamp 1669390400
transform 1 0 34793 0 1 23285
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_34
timestamp 1669390400
transform 1 0 33209 0 1 24869
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_35
timestamp 1669390400
transform 1 0 41261 0 1 16817
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_36
timestamp 1669390400
transform 1 0 36245 0 1 21833
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_37
timestamp 1669390400
transform 1 0 37301 0 1 20777
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_38
timestamp 1669390400
transform 1 0 37169 0 1 20909
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_39
timestamp 1669390400
transform 1 0 37037 0 1 21041
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_40
timestamp 1669390400
transform 1 0 36905 0 1 21173
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_41
timestamp 1669390400
transform 1 0 36773 0 1 21305
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_42
timestamp 1669390400
transform 1 0 36641 0 1 21437
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_43
timestamp 1669390400
transform 1 0 36509 0 1 21569
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_44
timestamp 1669390400
transform 1 0 36377 0 1 21701
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_45
timestamp 1669390400
transform 1 0 32945 0 1 25133
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_46
timestamp 1669390400
transform 1 0 32813 0 1 25265
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_47
timestamp 1669390400
transform 1 0 32681 0 1 25397
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_48
timestamp 1669390400
transform 1 0 32549 0 1 25529
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_49
timestamp 1669390400
transform 1 0 32417 0 1 25661
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_50
timestamp 1669390400
transform 1 0 32285 0 1 25793
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_51
timestamp 1669390400
transform 1 0 32153 0 1 25925
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_52
timestamp 1669390400
transform 1 0 32021 0 1 26057
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_53
timestamp 1669390400
transform 1 0 31889 0 1 26189
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_54
timestamp 1669390400
transform 1 0 31757 0 1 26321
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_55
timestamp 1669390400
transform 1 0 31625 0 1 26453
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_56
timestamp 1669390400
transform 1 0 31493 0 1 26585
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_57
timestamp 1669390400
transform 1 0 31361 0 1 26717
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_58
timestamp 1669390400
transform 1 0 31229 0 1 26849
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_59
timestamp 1669390400
transform 1 0 33077 0 1 25001
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_60
timestamp 1669390400
transform 1 0 30965 0 1 27113
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_61
timestamp 1669390400
transform 1 0 30833 0 1 27245
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_62
timestamp 1669390400
transform 1 0 30701 0 1 27377
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_63
timestamp 1669390400
transform 1 0 39017 0 1 19061
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_64
timestamp 1669390400
transform 1 0 31097 0 1 26981
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_65
timestamp 1669390400
transform 1 0 36113 0 1 21965
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_66
timestamp 1669390400
transform 1 0 35981 0 1 22097
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_67
timestamp 1669390400
transform 1 0 35849 0 1 22229
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_68
timestamp 1669390400
transform 1 0 35717 0 1 22361
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_69
timestamp 1669390400
transform 1 0 35585 0 1 22493
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_70
timestamp 1669390400
transform 1 0 35453 0 1 22625
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_71
timestamp 1669390400
transform 1 0 35321 0 1 22757
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_72
timestamp 1669390400
transform 1 0 35189 0 1 22889
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_73
timestamp 1669390400
transform 1 0 34925 0 1 23153
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_74
timestamp 1669390400
transform 1 0 41921 0 1 16157
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_75
timestamp 1669390400
transform 1 0 41789 0 1 16289
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_76
timestamp 1669390400
transform 1 0 41657 0 1 16421
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_77
timestamp 1669390400
transform 1 0 41525 0 1 16553
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_78
timestamp 1669390400
transform 1 0 41393 0 1 16685
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_79
timestamp 1669390400
transform 1 0 39281 0 1 18797
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_80
timestamp 1669390400
transform 1 0 41129 0 1 16949
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_81
timestamp 1669390400
transform 1 0 40997 0 1 17081
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_82
timestamp 1669390400
transform 1 0 40865 0 1 17213
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_83
timestamp 1669390400
transform 1 0 40733 0 1 17345
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_84
timestamp 1669390400
transform 1 0 40601 0 1 17477
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_85
timestamp 1669390400
transform 1 0 40469 0 1 17609
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_86
timestamp 1669390400
transform 1 0 40337 0 1 17741
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_87
timestamp 1669390400
transform 1 0 40205 0 1 17873
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_88
timestamp 1669390400
transform 1 0 40073 0 1 18005
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_89
timestamp 1669390400
transform 1 0 39941 0 1 18137
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_90
timestamp 1669390400
transform 1 0 39809 0 1 18269
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_91
timestamp 1669390400
transform 1 0 39677 0 1 18401
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_92
timestamp 1669390400
transform 1 0 39545 0 1 18533
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_93
timestamp 1669390400
transform 1 0 38225 0 1 19853
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_94
timestamp 1669390400
transform 1 0 38093 0 1 19985
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_95
timestamp 1669390400
transform 1 0 37961 0 1 20117
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_96
timestamp 1669390400
transform 1 0 37829 0 1 20249
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_97
timestamp 1669390400
transform 1 0 37697 0 1 20381
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_98
timestamp 1669390400
transform 1 0 37565 0 1 20513
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_99
timestamp 1669390400
transform 1 0 37433 0 1 20645
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_100
timestamp 1669390400
transform 1 0 39413 0 1 18665
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_101
timestamp 1669390400
transform 1 0 35057 0 1 23021
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_102
timestamp 1669390400
transform 1 0 39149 0 1 18929
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_103
timestamp 1669390400
transform 1 0 33341 0 1 24737
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_104
timestamp 1669390400
transform 1 0 33473 0 1 24605
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_105
timestamp 1669390400
transform 1 0 33605 0 1 24473
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_106
timestamp 1669390400
transform 1 0 33737 0 1 24341
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_107
timestamp 1669390400
transform 1 0 23045 0 1 35033
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_108
timestamp 1669390400
transform 1 0 23309 0 1 34769
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_109
timestamp 1669390400
transform 1 0 23441 0 1 34637
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_110
timestamp 1669390400
transform 1 0 23573 0 1 34505
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_111
timestamp 1669390400
transform 1 0 23705 0 1 34373
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_112
timestamp 1669390400
transform 1 0 23837 0 1 34241
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_113
timestamp 1669390400
transform 1 0 23969 0 1 34109
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_114
timestamp 1669390400
transform 1 0 24101 0 1 33977
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_115
timestamp 1669390400
transform 1 0 24233 0 1 33845
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_116
timestamp 1669390400
transform 1 0 24365 0 1 33713
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_117
timestamp 1669390400
transform 1 0 24497 0 1 33581
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_118
timestamp 1669390400
transform 1 0 24629 0 1 33449
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_119
timestamp 1669390400
transform 1 0 24761 0 1 33317
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_120
timestamp 1669390400
transform 1 0 25025 0 1 33053
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_121
timestamp 1669390400
transform 1 0 23177 0 1 34901
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_122
timestamp 1669390400
transform 1 0 22913 0 1 35165
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_123
timestamp 1669390400
transform 1 0 22781 0 1 35297
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_124
timestamp 1669390400
transform 1 0 22649 0 1 35429
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_125
timestamp 1669390400
transform 1 0 22517 0 1 35561
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_126
timestamp 1669390400
transform 1 0 22385 0 1 35693
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_127
timestamp 1669390400
transform 1 0 22253 0 1 35825
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_128
timestamp 1669390400
transform 1 0 22121 0 1 35957
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_129
timestamp 1669390400
transform 1 0 21989 0 1 36089
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_130
timestamp 1669390400
transform 1 0 21857 0 1 36221
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_131
timestamp 1669390400
transform 1 0 21725 0 1 36353
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_132
timestamp 1669390400
transform 1 0 21593 0 1 36485
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_133
timestamp 1669390400
transform 1 0 21461 0 1 36617
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_134
timestamp 1669390400
transform 1 0 21329 0 1 36749
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_135
timestamp 1669390400
transform 1 0 21065 0 1 37013
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_136
timestamp 1669390400
transform 1 0 24893 0 1 33185
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_137
timestamp 1669390400
transform 1 0 18557 0 1 39521
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_138
timestamp 1669390400
transform 1 0 18425 0 1 39653
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_139
timestamp 1669390400
transform 1 0 18293 0 1 39785
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_140
timestamp 1669390400
transform 1 0 18161 0 1 39917
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_141
timestamp 1669390400
transform 1 0 16973 0 1 41105
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_142
timestamp 1669390400
transform 1 0 18029 0 1 40049
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_143
timestamp 1669390400
transform 1 0 17897 0 1 40181
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_144
timestamp 1669390400
transform 1 0 17765 0 1 40313
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_145
timestamp 1669390400
transform 1 0 17633 0 1 40445
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_146
timestamp 1669390400
transform 1 0 17501 0 1 40577
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_147
timestamp 1669390400
transform 1 0 17369 0 1 40709
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_148
timestamp 1669390400
transform 1 0 27401 0 1 30677
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_149
timestamp 1669390400
transform 1 0 27269 0 1 30809
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_150
timestamp 1669390400
transform 1 0 27137 0 1 30941
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_151
timestamp 1669390400
transform 1 0 21197 0 1 36881
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_152
timestamp 1669390400
transform 1 0 26873 0 1 31205
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_153
timestamp 1669390400
transform 1 0 26741 0 1 31337
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_154
timestamp 1669390400
transform 1 0 26609 0 1 31469
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_155
timestamp 1669390400
transform 1 0 26477 0 1 31601
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_156
timestamp 1669390400
transform 1 0 26345 0 1 31733
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_157
timestamp 1669390400
transform 1 0 26213 0 1 31865
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_158
timestamp 1669390400
transform 1 0 26081 0 1 31997
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_159
timestamp 1669390400
transform 1 0 25949 0 1 32129
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_160
timestamp 1669390400
transform 1 0 25817 0 1 32261
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_161
timestamp 1669390400
transform 1 0 25685 0 1 32393
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_162
timestamp 1669390400
transform 1 0 25553 0 1 32525
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_163
timestamp 1669390400
transform 1 0 25421 0 1 32657
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_164
timestamp 1669390400
transform 1 0 25289 0 1 32789
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_165
timestamp 1669390400
transform 1 0 25157 0 1 32921
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_166
timestamp 1669390400
transform 1 0 27005 0 1 31073
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_167
timestamp 1669390400
transform 1 0 17105 0 1 40973
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_168
timestamp 1669390400
transform 1 0 16841 0 1 41237
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_169
timestamp 1669390400
transform 1 0 16709 0 1 41369
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_170
timestamp 1669390400
transform 1 0 16577 0 1 41501
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_171
timestamp 1669390400
transform 1 0 16445 0 1 41633
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_172
timestamp 1669390400
transform 1 0 16313 0 1 41765
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_173
timestamp 1669390400
transform 1 0 16181 0 1 41897
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_174
timestamp 1669390400
transform 1 0 19085 0 1 38993
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_175
timestamp 1669390400
transform 1 0 20933 0 1 37145
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_176
timestamp 1669390400
transform 1 0 20801 0 1 37277
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_177
timestamp 1669390400
transform 1 0 20669 0 1 37409
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_178
timestamp 1669390400
transform 1 0 20537 0 1 37541
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_179
timestamp 1669390400
transform 1 0 20405 0 1 37673
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_180
timestamp 1669390400
transform 1 0 20273 0 1 37805
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_181
timestamp 1669390400
transform 1 0 20141 0 1 37937
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_182
timestamp 1669390400
transform 1 0 20009 0 1 38069
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_183
timestamp 1669390400
transform 1 0 19877 0 1 38201
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_184
timestamp 1669390400
transform 1 0 19745 0 1 38333
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_185
timestamp 1669390400
transform 1 0 19613 0 1 38465
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_186
timestamp 1669390400
transform 1 0 19481 0 1 38597
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_187
timestamp 1669390400
transform 1 0 19349 0 1 38729
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_188
timestamp 1669390400
transform 1 0 19217 0 1 38861
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_189
timestamp 1669390400
transform 1 0 17237 0 1 40841
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_190
timestamp 1669390400
transform 1 0 18953 0 1 39125
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_191
timestamp 1669390400
transform 1 0 18821 0 1 39257
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_192
timestamp 1669390400
transform 1 0 18689 0 1 39389
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_193
timestamp 1669390400
transform 1 0 29117 0 1 28961
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_194
timestamp 1669390400
transform 1 0 28853 0 1 29225
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_195
timestamp 1669390400
transform 1 0 28589 0 1 29489
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_196
timestamp 1669390400
transform 1 0 28457 0 1 29621
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_197
timestamp 1669390400
transform 1 0 28325 0 1 29753
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_198
timestamp 1669390400
transform 1 0 28193 0 1 29885
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_199
timestamp 1669390400
transform 1 0 28061 0 1 30017
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_200
timestamp 1669390400
transform 1 0 27929 0 1 30149
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_201
timestamp 1669390400
transform 1 0 27797 0 1 30281
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_202
timestamp 1669390400
transform 1 0 27665 0 1 30413
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_203
timestamp 1669390400
transform 1 0 28721 0 1 29357
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_204
timestamp 1669390400
transform 1 0 28985 0 1 29093
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_205
timestamp 1669390400
transform 1 0 29249 0 1 28829
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_206
timestamp 1669390400
transform 1 0 30437 0 1 27641
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_207
timestamp 1669390400
transform 1 0 30305 0 1 27773
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_208
timestamp 1669390400
transform 1 0 30173 0 1 27905
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_209
timestamp 1669390400
transform 1 0 30041 0 1 28037
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_210
timestamp 1669390400
transform 1 0 29909 0 1 28169
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_211
timestamp 1669390400
transform 1 0 29777 0 1 28301
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_212
timestamp 1669390400
transform 1 0 29645 0 1 28433
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_213
timestamp 1669390400
transform 1 0 29513 0 1 28565
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_214
timestamp 1669390400
transform 1 0 29381 0 1 28697
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_215
timestamp 1669390400
transform 1 0 27533 0 1 30545
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_216
timestamp 1669390400
transform 1 0 30569 0 1 27509
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_217
timestamp 1669390400
transform 1 0 13673 0 1 44405
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_218
timestamp 1669390400
transform 1 0 13541 0 1 44537
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_219
timestamp 1669390400
transform 1 0 13409 0 1 44669
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_220
timestamp 1669390400
transform 1 0 13277 0 1 44801
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_221
timestamp 1669390400
transform 1 0 15125 0 1 42953
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_222
timestamp 1669390400
transform 1 0 15917 0 1 42161
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_223
timestamp 1669390400
transform 1 0 15785 0 1 42293
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_224
timestamp 1669390400
transform 1 0 15653 0 1 42425
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_225
timestamp 1669390400
transform 1 0 15521 0 1 42557
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_226
timestamp 1669390400
transform 1 0 15389 0 1 42689
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_227
timestamp 1669390400
transform 1 0 15257 0 1 42821
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_228
timestamp 1669390400
transform 1 0 14993 0 1 43085
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_229
timestamp 1669390400
transform 1 0 14861 0 1 43217
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_230
timestamp 1669390400
transform 1 0 14729 0 1 43349
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_231
timestamp 1669390400
transform 1 0 14597 0 1 43481
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_232
timestamp 1669390400
transform 1 0 14465 0 1 43613
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_233
timestamp 1669390400
transform 1 0 14333 0 1 43745
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_234
timestamp 1669390400
transform 1 0 14201 0 1 43877
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_235
timestamp 1669390400
transform 1 0 14069 0 1 44009
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_236
timestamp 1669390400
transform 1 0 13937 0 1 44141
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_237
timestamp 1669390400
transform 1 0 13805 0 1 44273
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_238
timestamp 1669390400
transform 1 0 16049 0 1 42029
box 0 0 1 1
use M1_PSUB_CDNS_406619561345  M1_PSUB_CDNS_406619561345_239
timestamp 1669390400
transform 1 0 42053 0 1 16025
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_0
timestamp 1669390400
transform 1 0 70641 0 1 24306
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_1
timestamp 1669390400
transform 1 0 70641 0 1 56310
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_2
timestamp 1669390400
transform 1 0 70641 0 1 54702
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_3
timestamp 1669390400
transform 1 0 70641 0 1 53122
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_4
timestamp 1669390400
transform 1 0 70641 0 1 67516
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_5
timestamp 1669390400
transform 1 0 70641 0 1 59520
box 0 0 1 1
use M3_M2_CDNS_406619561346  M3_M2_CDNS_406619561346_6
timestamp 1669390400
transform 1 0 70641 0 1 41897
box 0 0 1 1
use M3_M2_CDNS_406619561347  M3_M2_CDNS_406619561347_0
timestamp 1669390400
transform 1 0 70641 0 1 37900
box 0 0 1 1
use M3_M2_CDNS_406619561347  M3_M2_CDNS_406619561347_1
timestamp 1669390400
transform 1 0 70641 0 1 28320
box 0 0 1 1
use M3_M2_CDNS_406619561347  M3_M2_CDNS_406619561347_2
timestamp 1669390400
transform 1 0 70641 0 1 31488
box 0 0 1 1
use M3_M2_CDNS_406619561347  M3_M2_CDNS_406619561347_3
timestamp 1669390400
transform 1 0 70641 0 1 34700
box 0 0 1 1
use M3_M2_CDNS_406619561347  M3_M2_CDNS_406619561347_4
timestamp 1669390400
transform 1 0 70641 0 1 44307
box 0 0 1 1
use polygon00001  polygon00001_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 13108 13108 46414 45051
use polygon00002  polygon00002_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 0 0 1 1
use polygon00003  polygon00003_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 0 0 1 1
use polygon00004  polygon00004_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 14000 14000 71000 71000
use polygon00005  polygon00005_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 17200 17200 71000 71000
use polygon00006  polygon00006_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 20400 20400 71000 71000
use polygon00007  polygon00007_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 26800 26800 71000 71000
use polygon00008  polygon00008_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 30000 30000 71000 71000
use polygon00009  polygon00009_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 33200 33200 71000 71000
use polygon00010  polygon00010_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 36400 36400 71000 71000
use polygon00011  polygon00011_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 42800 42800 71000 71000
use polygon00012  polygon00012_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 46000 46000 71000 71000
use polygon00013  polygon00013_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 68400 68400 71000 71000
use polygon00014  polygon00014_0
timestamp 1669648928
transform 1 0 0 0 1 0
box 68400 68400 71000 71000
<< labels >>
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 6504834
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 6486408
string path 1687.500 1775.000 1687.500 1710.075 1710.075 1687.500 1775.000 1687.500 
<< end >>
