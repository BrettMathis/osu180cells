magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 240 120
<< mvndiff >>
rect -88 83 0 120
rect -88 37 -75 83
rect -29 37 0 83
rect -88 0 0 37
rect 240 83 328 120
rect 240 37 269 83
rect 315 37 328 83
rect 240 0 328 37
<< mvndiffc >>
rect -75 37 -29 83
rect 269 37 315 83
<< polysilicon >>
rect 0 120 240 164
rect 0 -44 240 0
<< metal1 >>
rect -75 83 -29 120
rect -75 0 -29 37
rect 269 83 315 120
rect 269 0 315 37
<< labels >>
flabel metal1 s -52 60 -52 60 0 FreeSans 200 0 0 0 S
flabel metal1 s 292 60 292 60 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 853342
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 852318
<< end >>
