magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< obsv1 >>
rect 0 0 86372 53776
<< obsv2 >>
rect 0 0 86372 53776
<< metal3 >>
rect 1401 52976 2401 53776
rect 2626 53168 3626 53776
rect 4137 52976 5137 53776
rect 5362 53168 6362 53776
rect 6801 52976 7801 53776
rect 8026 53168 9026 53776
rect 9537 52976 10537 53776
rect 10762 53168 11762 53776
rect 12201 52976 13201 53776
rect 13426 53168 14426 53776
rect 14937 52976 15937 53776
rect 16162 53168 17162 53776
rect 17601 52976 18601 53776
rect 18826 53168 19826 53776
rect 20653 52976 21653 53776
rect 22258 53168 23258 53776
rect 23483 52976 24483 53776
rect 25158 53168 26158 53776
rect 26572 52976 27572 53776
rect 27877 53168 28877 53776
rect 29273 53168 30273 53776
rect 30710 52976 31710 53776
rect 32381 53168 33381 53776
rect 34024 53168 35024 53776
rect 35415 52976 36415 53776
rect 36948 53168 37948 53776
rect 38585 52976 39585 53776
rect 39882 53168 40882 53776
rect 41230 52976 42230 53776
rect 42430 53168 43430 53776
rect 43713 53168 44713 53776
rect 45069 52976 46069 53776
rect 46313 52976 47313 53776
rect 47538 53168 48538 53776
rect 48901 52976 49901 53776
rect 50465 53168 51465 53776
rect 52569 52976 53569 53776
rect 54262 52976 55262 53776
rect 55990 53168 56990 53776
rect 57547 52976 58547 53776
rect 58791 53168 59791 53776
rect 60977 52976 61977 53776
rect 62202 53168 63202 53776
rect 63713 52976 64713 53776
rect 64938 53168 65938 53776
rect 66377 52976 67377 53776
rect 67602 53168 68602 53776
rect 69113 52976 70113 53776
rect 70338 53168 71338 53776
rect 71777 52976 72777 53776
rect 73002 53168 74002 53776
rect 74513 52976 75513 53776
rect 75738 53168 76738 53776
rect 77177 52976 78177 53776
rect 78402 53168 79402 53776
rect 80229 52976 81229 53776
rect 81834 53168 82834 53776
rect 83059 52976 84059 53776
rect 84666 52976 85666 53776
rect 0 51976 86372 52976
rect 0 51626 1014 51776
rect 0 51528 27779 51626
rect 58791 51576 59517 51591
rect 85358 51576 86372 51776
rect 58791 51528 86372 51576
rect 0 51327 86372 51528
rect 0 51226 27779 51327
rect 30402 51326 54622 51327
rect 58791 51276 86372 51327
rect 0 51076 1014 51226
rect 58791 51258 59517 51276
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49726 27272 49776
rect 30403 49726 54622 49728
rect 59421 49726 86372 49776
rect 0 49526 86372 49726
rect 0 49476 27272 49526
rect 59421 49476 86372 49526
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47926 27272 47976
rect 30403 47926 54622 47928
rect 59421 47926 86372 47976
rect 0 47726 86372 47926
rect 0 47676 27272 47726
rect 59421 47676 86372 47726
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46126 27272 46176
rect 30403 46126 54622 46128
rect 59421 46126 86372 46176
rect 0 45926 86372 46126
rect 0 45876 27272 45926
rect 59421 45876 86372 45926
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44326 27272 44376
rect 30403 44326 54622 44328
rect 59421 44326 86372 44376
rect 0 44126 86372 44326
rect 0 44076 27272 44126
rect 59421 44076 86372 44126
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42526 27272 42576
rect 30403 42526 54622 42528
rect 59421 42526 86372 42576
rect 0 42326 86372 42526
rect 0 42276 27272 42326
rect 59421 42276 86372 42326
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40726 27272 40776
rect 30403 40726 54622 40728
rect 59421 40726 86372 40776
rect 0 40526 86372 40726
rect 0 40476 27272 40526
rect 59421 40476 86372 40526
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38926 27272 38976
rect 30403 38926 54622 38928
rect 59421 38926 86372 38976
rect 0 38726 86372 38926
rect 0 38676 27272 38726
rect 59421 38676 86372 38726
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37126 27272 37176
rect 30403 37126 54622 37128
rect 59421 37126 86372 37176
rect 0 36926 86372 37126
rect 0 36876 27272 36926
rect 59421 36876 86372 36926
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 84666 35776 86372 36476
rect 0 34536 27828 35326
rect 57369 34536 86372 35326
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 32318 27214 34124
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 32315 86372 34124
rect 57908 32199 58351 32315
rect 26772 31486 58351 32199
rect 26772 29714 58351 30105
rect 84666 29714 86372 32315
rect 0 29430 86372 29714
rect 0 26890 26070 28416
rect 26772 27382 58351 29430
rect 0 26435 27828 26890
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 58785 26890 86372 28416
rect 57295 26435 86372 26890
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 0 23380 1706 23938
rect 26770 23380 58348 24278
rect 84666 23380 86372 23938
rect 0 23370 86372 23380
rect 0 22938 27214 23370
rect 27387 22291 57677 23199
rect 57908 22938 86372 23370
rect 57908 22937 83763 22938
rect 27387 22282 27826 22291
rect 0 21827 27826 22282
rect 56078 22282 57677 22291
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 21827 86372 22282
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 19969 86372 20739
rect 0 18016 24250 19969
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 61807 16784 86372 17730
rect 24111 16597 27828 16598
rect 0 15015 27828 16597
rect 46982 15015 86372 16784
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14936 51760 14966
rect 0 14491 47683 14936
rect 0 14329 45977 14491
rect 0 14328 24250 14329
rect 24047 14178 27214 14179
rect 0 13461 27214 14178
rect 0 12846 1706 13461
rect 24047 12934 27214 13461
rect 27387 13760 45977 14329
rect 57295 14328 86372 14968
rect 57295 14327 83763 14328
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13245 49775 13760
rect 29478 13243 49775 13245
rect 41493 13078 49775 13243
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12574 34761 12846
rect 50228 13461 86372 13866
rect 50228 12846 58421 13461
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12574 86372 12846
rect 0 12046 86372 12574
rect 0 12036 24250 12046
rect 26772 12036 86372 12046
rect 26772 12035 84999 12036
rect 26772 11844 58351 12035
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 10176 27828 11491
rect 29478 11697 58351 11844
rect 29478 10756 41516 11697
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 34741 9972 41516 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 10740 86372 11491
rect 24047 9515 28729 9516
rect 0 8154 28729 9515
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 6982 27828 7595
rect 28178 7652 28729 8154
rect 41857 9502 51430 10420
rect 57295 10176 86372 10740
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 41857 9165 55482 9502
rect 29513 7900 41397 8582
rect 28178 7084 34622 7652
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8888 55482 9165
rect 50922 7596 57736 8888
rect 57909 9514 62278 9516
rect 83361 9514 86372 9515
rect 57909 8154 86372 9514
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7392 86372 7595
rect 34860 6984 86372 7392
rect 34860 6592 55482 6984
rect 57295 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 0 5766 34622 6177
rect 23687 5629 27214 5630
rect 0 5175 27214 5629
rect 29458 5665 34622 5766
rect 50922 6199 55482 6592
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 50922 5766 86372 6198
rect 50922 5605 55482 5766
rect 0 5174 24250 5175
rect 0 5173 3011 5174
rect 0 4515 1712 5173
rect 57909 5629 62429 5630
rect 57909 5175 86372 5629
rect 61802 5174 86372 5175
rect 83361 5173 86372 5174
rect 57909 4619 62429 4621
rect 23909 4515 62429 4619
rect 84660 4515 86372 5173
rect 0 4166 86372 4515
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3772 61215 3875
rect 0 3524 86372 3772
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 0 2854 1000 3420
rect 60886 3420 86372 3524
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
<< obsm3 >>
rect 0 53032 1345 53776
rect 2457 53112 2570 53776
rect 3682 53112 4081 53776
rect 2457 53032 4081 53112
rect 5193 53112 5306 53776
rect 6418 53112 6745 53776
rect 5193 53032 6745 53112
rect 7857 53112 7970 53776
rect 9082 53112 9481 53776
rect 7857 53032 9481 53112
rect 10593 53112 10706 53776
rect 11818 53112 12145 53776
rect 10593 53032 12145 53112
rect 13257 53112 13370 53776
rect 14482 53112 14881 53776
rect 13257 53032 14881 53112
rect 15993 53112 16106 53776
rect 17218 53112 17545 53776
rect 15993 53032 17545 53112
rect 18657 53112 18770 53776
rect 19882 53112 20597 53776
rect 18657 53032 20597 53112
rect 21709 53112 22202 53776
rect 23314 53112 23427 53776
rect 21709 53032 23427 53112
rect 24539 53112 25102 53776
rect 26214 53112 26516 53776
rect 24539 53032 26516 53112
rect 27628 53112 27821 53776
rect 28933 53112 29217 53776
rect 30329 53112 30654 53776
rect 27628 53032 30654 53112
rect 31766 53112 32325 53776
rect 33437 53112 33968 53776
rect 35080 53112 35359 53776
rect 31766 53032 35359 53112
rect 36471 53112 36892 53776
rect 38004 53112 38529 53776
rect 36471 53032 38529 53112
rect 39641 53112 39826 53776
rect 40938 53112 41174 53776
rect 39641 53032 41174 53112
rect 42286 53112 42374 53776
rect 43486 53112 43657 53776
rect 44769 53112 45013 53776
rect 42286 53032 45013 53112
rect 46125 53032 46257 53776
rect 47369 53112 47482 53776
rect 48594 53112 48845 53776
rect 47369 53032 48845 53112
rect 49957 53112 50409 53776
rect 51521 53112 52513 53776
rect 49957 53032 52513 53112
rect 53625 53032 54206 53776
rect 55318 53112 55934 53776
rect 57046 53112 57491 53776
rect 55318 53032 57491 53112
rect 58603 53112 58735 53776
rect 59847 53112 60921 53776
rect 58603 53032 60921 53112
rect 62033 53112 62146 53776
rect 63258 53112 63657 53776
rect 62033 53032 63657 53112
rect 64769 53112 64882 53776
rect 65994 53112 66321 53776
rect 64769 53032 66321 53112
rect 67433 53112 67546 53776
rect 68658 53112 69057 53776
rect 67433 53032 69057 53112
rect 70169 53112 70282 53776
rect 71394 53112 71721 53776
rect 70169 53032 71721 53112
rect 72833 53112 72946 53776
rect 74058 53112 74457 53776
rect 72833 53032 74457 53112
rect 75569 53112 75682 53776
rect 76794 53112 77121 53776
rect 75569 53032 77121 53112
rect 78233 53112 78346 53776
rect 79458 53112 80173 53776
rect 78233 53032 80173 53112
rect 81285 53112 81778 53776
rect 82890 53112 83003 53776
rect 81285 53032 83003 53112
rect 84115 53032 84610 53776
rect 85722 53032 86372 53776
rect 0 51832 86372 51920
rect 1070 51682 85302 51832
rect 27835 51647 85302 51682
rect 27835 51584 58735 51647
rect 59573 51632 85302 51647
rect 27835 51270 30346 51271
rect 54678 51270 58735 51271
rect 27835 51202 58735 51270
rect 59573 51202 85302 51220
rect 27835 51170 85302 51202
rect 1070 51020 85302 51170
rect 0 50932 86372 51020
rect 1762 50120 84610 50932
rect 0 50032 86372 50120
rect 1070 49832 85302 50032
rect 27328 49784 59365 49832
rect 27328 49782 30347 49784
rect 54678 49782 59365 49784
rect 27328 49420 59365 49470
rect 1070 49220 85302 49420
rect 0 49132 86372 49220
rect 1762 48320 84610 49132
rect 0 48232 86372 48320
rect 1070 48032 85302 48232
rect 27328 47984 59365 48032
rect 27328 47982 30347 47984
rect 54678 47982 59365 47984
rect 27328 47620 59365 47670
rect 1070 47420 85302 47620
rect 0 47332 86372 47420
rect 1762 46520 84610 47332
rect 0 46432 86372 46520
rect 1070 46232 85302 46432
rect 27328 46184 59365 46232
rect 27328 46182 30347 46184
rect 54678 46182 59365 46184
rect 27328 45820 59365 45870
rect 1070 45620 85302 45820
rect 0 45532 86372 45620
rect 1762 44720 84610 45532
rect 0 44632 86372 44720
rect 1070 44432 85302 44632
rect 27328 44384 59365 44432
rect 27328 44382 30347 44384
rect 54678 44382 59365 44384
rect 27328 44020 59365 44070
rect 1070 43820 85302 44020
rect 0 43732 86372 43820
rect 1762 42920 84610 43732
rect 0 42832 86372 42920
rect 1070 42632 85302 42832
rect 27328 42584 59365 42632
rect 27328 42582 30347 42584
rect 54678 42582 59365 42584
rect 27328 42220 59365 42270
rect 1070 42020 85302 42220
rect 0 41932 86372 42020
rect 1762 41120 84610 41932
rect 0 41032 86372 41120
rect 1070 40832 85302 41032
rect 27328 40784 59365 40832
rect 27328 40782 30347 40784
rect 54678 40782 59365 40784
rect 27328 40420 59365 40470
rect 1070 40220 85302 40420
rect 0 40132 86372 40220
rect 1762 39320 84610 40132
rect 0 39232 86372 39320
rect 1070 39032 85302 39232
rect 27328 38984 59365 39032
rect 27328 38982 30347 38984
rect 54678 38982 59365 38984
rect 27328 38620 59365 38670
rect 1070 38420 85302 38620
rect 0 38332 86372 38420
rect 1762 37520 84610 38332
rect 0 37432 86372 37520
rect 1070 37232 85302 37432
rect 27328 37184 59365 37232
rect 27328 37182 30347 37184
rect 54678 37182 59365 37184
rect 27328 36820 59365 36870
rect 1070 36620 85302 36820
rect 0 36532 86372 36620
rect 1762 35720 84610 36532
rect 0 35382 86372 35720
rect 27884 34480 57313 35382
rect 0 34182 86372 34480
rect 0 34181 2039 34182
rect 2244 34181 86372 34182
rect 25141 34180 61797 34181
rect 72439 34180 72597 34181
rect 27270 32262 57852 34180
rect 25141 32260 57852 32262
rect 3067 32259 57852 32260
rect 1762 32255 57852 32259
rect 1762 31430 26716 32255
rect 58407 31430 84610 32259
rect 1762 30161 84610 31430
rect 1762 29770 26716 30161
rect 58407 29770 84610 30161
rect 0 28472 26716 29374
rect 26126 27326 26716 28472
rect 58407 28472 86372 29374
rect 58407 27326 58729 28472
rect 26126 26946 58729 27326
rect 27884 26379 57239 26946
rect 0 26378 6865 26379
rect 8219 26378 17665 26379
rect 19019 26378 66441 26379
rect 67795 26378 77241 26379
rect 78595 26378 86372 26379
rect 0 24334 86372 26378
rect 0 23994 26714 24334
rect 1762 23436 26714 23994
rect 58404 23994 86372 24334
rect 58404 23436 84610 23994
rect 27270 23255 57852 23314
rect 27270 22882 27331 23255
rect 0 22338 27331 22882
rect 57733 22881 57852 23255
rect 83819 22881 86372 22882
rect 57733 22338 86372 22881
rect 1070 21770 23980 21771
rect 27882 21770 56022 22235
rect 83819 21770 85302 21771
rect 1070 21764 85302 21770
rect 1070 21763 44376 21764
rect 1070 21681 29465 21763
rect 1070 21226 29457 21681
rect 0 20795 29457 21226
rect 55701 21226 85302 21764
rect 55701 20795 86372 21226
rect 24306 17960 61751 19913
rect 0 17959 61769 17960
rect 83819 17959 86372 17960
rect 0 17786 86372 17959
rect 23734 16840 61751 17786
rect 23734 16654 46926 16840
rect 23734 16653 24055 16654
rect 27884 15071 46926 16654
rect 55701 14910 57239 14912
rect 51816 14880 57239 14910
rect 47739 14435 57239 14880
rect 24306 14272 27331 14273
rect 0 14235 27331 14272
rect 0 14234 23991 14235
rect 1762 12903 23991 13405
rect 27270 13189 27331 14235
rect 46033 14271 57239 14435
rect 83819 14271 86372 14272
rect 46033 14235 86372 14271
rect 46033 14234 83113 14235
rect 84277 14234 86372 14235
rect 46033 14233 61751 14234
rect 72485 14233 72551 14234
rect 46033 14073 61717 14233
rect 46033 13922 59770 14073
rect 46033 13816 50172 13922
rect 60082 13922 61717 14073
rect 27270 13187 29422 13189
rect 27270 13022 41437 13187
rect 49831 13022 50172 13816
rect 27270 12990 50172 13022
rect 1762 12902 23765 12903
rect 34817 12630 50172 12990
rect 58477 12902 59770 13405
rect 60082 12903 84610 13405
rect 60082 12902 83113 12903
rect 84277 12902 84610 12903
rect 24306 11980 26716 11990
rect 0 11788 26716 11980
rect 85055 11979 86372 11980
rect 0 11549 29422 11788
rect 3067 11547 23991 11549
rect 27884 10700 29422 11549
rect 58407 11641 86372 11979
rect 27884 10120 34685 10700
rect 0 10119 2173 10120
rect 0 10118 2193 10119
rect 24306 10118 34685 10120
rect 0 9916 34685 10118
rect 41572 11583 86372 11641
rect 41572 10684 42205 11583
rect 57792 11549 86372 11583
rect 57792 11547 61769 11549
rect 41572 10476 57239 10684
rect 41572 9916 41801 10476
rect 0 9572 41801 9916
rect 0 9571 23991 9572
rect 24306 8097 28122 8098
rect 3067 8096 28122 8097
rect 0 7652 28122 8096
rect 3067 7651 23569 7652
rect 27884 7028 28122 7652
rect 28785 9109 41801 9572
rect 51486 10120 57239 10476
rect 51486 10119 61749 10120
rect 51486 10117 61769 10119
rect 84538 10117 86372 10120
rect 51486 9572 86372 10117
rect 51486 9558 57853 9572
rect 62334 9571 86372 9572
rect 62334 9570 83305 9571
rect 28785 8638 50866 9109
rect 28785 7844 29457 8638
rect 28785 7708 34804 7844
rect 27884 6926 29481 7028
rect 1070 6925 2170 6926
rect 1070 6924 2193 6925
rect 24306 6924 29481 6926
rect 1070 6688 29481 6924
rect 34678 6688 34804 7708
rect 1070 6629 34804 6688
rect 41453 7448 50866 8638
rect 55538 8944 57853 9558
rect 57792 8098 57853 8944
rect 57792 8097 61746 8098
rect 57792 8096 61769 8097
rect 57792 7652 86372 8096
rect 62803 7651 83305 7652
rect 1070 6255 29402 6629
rect 3067 6254 23631 6255
rect 41453 6121 50866 6536
rect 0 5686 29402 5710
rect 0 5685 23631 5686
rect 27270 5609 29402 5686
rect 34678 5609 50866 6121
rect 27270 5549 50866 5609
rect 55538 6926 57239 6928
rect 55538 6925 61746 6926
rect 55538 6924 61769 6925
rect 84843 6924 85302 6926
rect 55538 6255 85302 6924
rect 62485 6254 83305 6255
rect 55538 5686 86372 5710
rect 55538 5549 57853 5686
rect 62485 5685 86372 5686
rect 27270 5119 57853 5549
rect 24306 5118 61746 5119
rect 3067 5117 83305 5118
rect 1768 4677 84604 5117
rect 1768 4675 57853 4677
rect 1768 4571 23853 4675
rect 62485 4571 84604 4677
rect 59379 4108 61732 4110
rect 24397 4004 61732 4108
rect 0 3932 86372 4004
rect 0 3931 27382 3932
rect 27834 3931 28708 3932
rect 28950 3931 41718 3932
rect 41960 3931 42243 3932
rect 42485 3931 46817 3932
rect 47059 3931 47265 3932
rect 47507 3931 47713 3932
rect 47955 3931 48161 3932
rect 48403 3931 57289 3932
rect 0 3828 23853 3931
rect 61271 3828 86372 3932
rect 24397 3365 60830 3468
rect 3067 3364 60830 3365
rect 1056 2910 85302 3364
rect 0 2288 86372 2446
rect 0 0 650 1176
rect 1762 0 1983 1176
rect 3095 0 3386 1176
rect 4498 988 5786 1176
rect 4498 0 4586 988
rect 5698 0 5786 988
rect 6898 0 6986 1176
rect 8098 0 8186 1176
rect 9298 988 10586 1176
rect 9298 0 9386 988
rect 10498 0 10586 988
rect 11698 0 12387 1176
rect 13499 0 14186 1176
rect 15298 988 16586 1176
rect 15298 0 15386 988
rect 16498 0 16586 988
rect 17698 0 17786 1176
rect 18898 0 18986 1176
rect 20098 988 21854 1176
rect 20098 0 20186 988
rect 21298 0 21854 988
rect 22966 0 23054 1176
rect 24166 0 24354 1176
rect 25466 0 25654 1176
rect 26766 0 26954 1176
rect 28066 0 28254 1176
rect 29366 0 29554 1176
rect 30666 988 35975 1176
rect 30666 0 31268 988
rect 32380 0 32966 988
rect 34078 0 34775 988
rect 35887 0 35975 988
rect 37087 988 39172 1176
rect 37087 0 37972 988
rect 39084 0 39172 988
rect 40284 988 42377 1176
rect 40284 0 41177 988
rect 42289 0 42377 988
rect 43489 988 44777 1176
rect 43489 0 43577 988
rect 44689 0 44777 988
rect 45889 988 47177 1176
rect 45889 0 45977 988
rect 47089 0 47177 988
rect 48289 0 48510 1176
rect 49622 0 49820 1176
rect 50932 988 54402 1176
rect 50932 0 51177 988
rect 52289 0 52422 988
rect 53534 0 54402 988
rect 55514 0 55702 1176
rect 56814 0 57002 1176
rect 58114 0 58302 1176
rect 59414 0 59602 1176
rect 60714 0 60902 1176
rect 62014 0 62239 1176
rect 63351 988 65362 1176
rect 63351 0 64162 988
rect 65274 0 65362 988
rect 66474 0 66562 1176
rect 67674 0 67762 1176
rect 68874 988 70162 1176
rect 68874 0 68962 988
rect 70074 0 70162 988
rect 71274 0 71961 1176
rect 73073 0 73762 1176
rect 74874 988 76162 1176
rect 74874 0 74962 988
rect 76074 0 76162 988
rect 77274 0 77362 1176
rect 78474 0 78562 1176
rect 79674 988 80962 1176
rect 79674 0 79762 988
rect 80874 0 80962 988
rect 82074 0 82363 1176
rect 83475 0 84610 1176
rect 85722 0 86372 1176
<< labels >>
rlabel metal2 s 34243 0 34467 200 6 A[0]
port 7 nsew signal input
rlabel metal2 s 32552 0 32776 200 6 A[1]
port 6 nsew signal input
rlabel metal2 s 30859 0 31083 200 6 A[2]
port 5 nsew signal input
rlabel metal2 s 56265 0 56489 200 6 A[3]
port 4 nsew signal input
rlabel metal2 s 55164 0 55388 200 6 A[4]
port 3 nsew signal input
rlabel metal2 s 54417 0 54641 200 6 A[5]
port 2 nsew signal input
rlabel metal2 s 53772 0 53996 200 6 A[6]
port 1 nsew signal input
rlabel metal2 s 50342 0 50566 200 6 CEN
port 8 nsew signal input
rlabel metal2 s 27936 0 28160 200 6 CLK
port 9 nsew signal input
rlabel metal2 s 1864 0 2088 200 6 D[0]
port 17 nsew signal input
rlabel metal2 s 12206 0 12430 200 6 D[1]
port 16 nsew signal input
rlabel metal2 s 13454 0 13678 200 6 D[2]
port 15 nsew signal input
rlabel metal2 s 23795 0 24019 200 6 D[3]
port 14 nsew signal input
rlabel metal2 s 61447 0 61671 200 6 D[4]
port 13 nsew signal input
rlabel metal2 s 71782 0 72006 200 6 D[5]
port 12 nsew signal input
rlabel metal2 s 73030 0 73254 200 6 D[6]
port 11 nsew signal input
rlabel metal2 s 83372 0 83596 200 6 D[7]
port 10 nsew signal input
rlabel metal2 s 40588 0 40812 200 6 GWEN
port 18 nsew signal input
rlabel metal2 s 3380 0 3604 200 6 Q[0]
port 26 nsew signal output
rlabel metal2 s 11533 0 11757 200 6 Q[1]
port 25 nsew signal output
rlabel metal2 s 14127 0 14351 200 6 Q[2]
port 24 nsew signal output
rlabel metal2 s 22279 0 22503 200 6 Q[3]
port 23 nsew signal output
rlabel metal2 s 62958 0 63182 200 6 Q[4]
port 22 nsew signal output
rlabel metal2 s 71109 0 71333 200 6 Q[5]
port 21 nsew signal output
rlabel metal2 s 73703 0 73927 200 6 Q[6]
port 20 nsew signal output
rlabel metal2 s 81855 0 82079 200 6 Q[7]
port 19 nsew signal output
rlabel metal2 s 2539 0 2763 200 6 WEN[0]
port 36 nsew signal input
rlabel metal2 s 12604 0 12828 200 6 WEN[1]
port 35 nsew signal input
rlabel metal2 s 13054 0 13278 200 6 WEN[2]
port 34 nsew signal input
rlabel metal2 s 23404 0 23628 200 6 WEN[3]
port 33 nsew signal input
rlabel metal2 s 62115 0 62339 200 6 WEN[4]
port 32 nsew signal input
rlabel metal2 s 72180 0 72404 200 6 WEN[5]
port 31 nsew signal input
rlabel metal2 s 72630 0 72854 200 6 WEN[6]
port 30 nsew signal input
rlabel metal2 s 82695 0 82919 200 6 WEN[7]
port 29 nsew signal input
rlabel metal3 s 0 50176 1706 50876 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 48376 1706 49076 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 46576 1706 47276 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 44776 1706 45476 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 42976 1706 43676 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 41176 1706 41876 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 39376 1706 40076 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 37576 1706 38276 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 35776 1706 36476 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 8152 3011 9515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 8153 24250 9515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 28178 7084 28729 9516 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24047 8154 28729 9516 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29537 6744 34622 7652 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 28178 7084 34622 7652 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 1401 51976 2401 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 4137 51976 5137 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 6801 51976 7801 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 9537 51976 10537 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 12201 51976 13201 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 14937 51976 15937 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 17601 51976 18601 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 20653 51976 21653 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23483 51976 24483 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26572 51976 27572 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 30710 51976 31710 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 35415 51976 36415 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 38585 51976 39585 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 41230 51976 42230 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 45069 51976 46069 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 46313 51976 47313 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 48901 51976 49901 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 52569 51976 53569 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 54262 51976 55262 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57547 51976 58547 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 60977 51976 61977 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 63713 51976 64713 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 66377 51976 67377 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 69113 51976 70113 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 71777 51976 72777 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 74513 51976 75513 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 77177 51976 78177 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 80229 51976 81229 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83059 51976 84059 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 51976 85666 53776 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 51976 86372 52976 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 50176 86372 50876 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 48376 86372 49076 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 46576 86372 47276 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 44776 86372 45476 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 42976 86372 43676 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 41176 86372 41876 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 39376 86372 40076 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 37576 86372 38276 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 35776 86372 36476 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 29430 1706 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 2095 32315 2188 34126 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 32315 3011 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 32316 25085 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 32318 27214 34124 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26772 31486 58351 32199 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26772 27382 58351 30105 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57908 31486 58351 34124 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61853 32315 72383 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57908 32315 86372 34124 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 29430 86372 29714 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 29430 86372 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 72653 32315 86372 34125 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 22938 1706 23938 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 22938 27214 23380 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26770 23370 58348 24278 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57908 22937 83763 23380 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57908 22938 86372 23380 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 22938 86372 23938 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 18016 24250 20739 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29513 19969 55645 21625 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29521 19969 55645 21707 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 44432 19969 55645 21708 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61825 18015 83763 20739 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61807 18016 86372 20739 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 19969 86372 20739 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 12036 1706 14178 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23821 12046 34761 12847 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 13461 27214 14178 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 12036 24250 12846 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24047 12046 27214 14179 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24047 12046 34761 12934 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 34741 9972 41516 12574 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29478 10756 41516 12574 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29478 11697 58351 12574 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26772 11844 58351 12574 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 50228 12035 58421 13866 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 59826 12035 60026 14017 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 50228 13461 86372 13866 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61807 13461 72429 14178 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61773 13461 86372 14177 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83169 12035 84221 12847 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83169 13461 84221 14179 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 50228 12036 86372 12846 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 26772 12035 84999 12574 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 12036 86372 14178 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 72607 13461 86372 14178 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61802 8153 86372 9514 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 8154 62278 9516 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61825 8152 86372 9514 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83361 8152 86372 9515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 4060 1712 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 5173 3011 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 5174 24250 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 4060 24341 4515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 6 VDD
port 27 nsew power bidirectional
rlabel metal3 s 2626 53168 3626 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 4642 0 5642 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 5362 53168 6362 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 8026 53168 9026 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 9442 0 10442 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 10762 53168 11762 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 13426 53168 14426 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 15442 0 16442 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 16162 53168 17162 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 18826 53168 19826 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 20242 0 21242 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 22258 53168 23258 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 25158 53168 26158 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 34536 27828 35326 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 6921 26434 8163 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 17721 26434 18963 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 26435 26070 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 26435 27828 26890 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 10176 3011 11493 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2249 10174 24250 11491 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2229 10175 24250 11491 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24047 10176 27828 11493 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27877 53168 28877 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29273 53168 30273 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 31324 0 32324 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 32381 53168 33381 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 33022 0 34022 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34024 53168 35024 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34831 0 35831 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 36948 53168 37948 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 38028 0 39028 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 39882 53168 40882 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41233 0 42233 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42430 53168 43430 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 43633 0 44633 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 43713 53168 44713 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46033 0 47033 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47538 53168 48538 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50465 53168 51465 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 51233 0 52233 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 52478 0 53478 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 55990 53168 56990 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58791 53168 59791 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 62202 53168 63202 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 64218 0 65218 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 64938 53168 65938 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 67602 53168 68602 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 69018 0 70018 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 70338 53168 71338 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 73002 53168 74002 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 75018 0 76018 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 75738 53168 76738 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 78402 53168 79402 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 79818 0 80818 932 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 81834 53168 82834 53776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 51076 1014 51776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 51226 27779 51626 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30402 51326 54622 51528 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 51327 86372 51528 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58791 51258 59517 51591 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58791 51276 86372 51576 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 51076 86372 51776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 49276 1014 49976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 49476 27272 49776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 49526 86372 49726 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 49476 86372 49776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 49276 86372 49976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 47476 1014 48176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 47676 27272 47976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 47726 86372 47926 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 47676 86372 47976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 47476 86372 48176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 45676 1014 46376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 45876 27272 46176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 45926 86372 46126 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 45876 86372 46176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 45676 86372 46376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 44076 27272 44376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 44126 86372 44326 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42326 86372 42526 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40526 86372 40726 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38726 86372 38926 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36926 86372 37126 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57369 34536 86372 35326 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8888 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 6982 86372 7595 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 6 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 6 VSS
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 53776
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2348210
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2298636
<< end >>
