magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 111 64 123
rect 11 70 16 111
rect 28 76 33 104
rect 28 70 41 76
rect 46 70 51 111
rect 13 44 23 50
rect 11 12 16 36
rect 28 19 33 70
rect 45 12 50 36
rect 0 0 64 12
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 9 112 19 118
rect 33 112 43 118
rect 10 111 18 112
rect 34 111 42 112
rect 32 76 40 77
rect 31 70 41 76
rect 32 69 40 70
rect 13 43 23 51
rect 10 11 18 12
rect 34 11 42 12
rect 9 5 19 11
rect 33 5 43 11
rect 10 4 18 5
rect 34 4 42 5
<< labels >>
rlabel metal2 s 13 43 23 51 6 A
port 1 nsew signal input
rlabel metal1 s 13 44 23 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 46 70 51 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 64 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 0 50 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 64 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 32 69 40 77 6 Y
port 2 nsew signal output
rlabel metal2 s 31 70 41 76 6 Y
port 2 nsew signal output
rlabel metal1 s 28 19 33 104 6 Y
port 2 nsew signal output
rlabel metal1 s 28 70 41 76 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 64 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 179234
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 174146
<< end >>
