magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 578 69 698 333
rect 772 69 892 333
<< mvpmos >>
rect 144 573 244 939
rect 348 573 448 939
rect 588 647 688 939
rect 792 647 892 939
<< mvndiff >>
rect 36 320 124 333
rect 36 180 49 320
rect 95 180 124 320
rect 36 69 124 180
rect 244 285 348 333
rect 244 239 273 285
rect 319 239 348 285
rect 244 69 348 239
rect 468 320 578 333
rect 468 180 497 320
rect 543 180 578 320
rect 468 69 578 180
rect 698 69 772 333
rect 892 320 980 333
rect 892 180 921 320
rect 967 180 980 320
rect 892 69 980 180
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 348 939
rect 448 861 588 939
rect 448 721 477 861
rect 523 721 588 861
rect 448 647 588 721
rect 688 861 792 939
rect 688 721 717 861
rect 763 721 792 861
rect 688 647 792 721
rect 892 861 980 939
rect 892 721 921 861
rect 967 721 980 861
rect 892 647 980 721
rect 448 573 528 647
<< mvndiffc >>
rect 49 180 95 320
rect 273 239 319 285
rect 497 180 543 320
rect 921 180 967 320
<< mvpdiffc >>
rect 69 721 115 861
rect 477 721 523 861
rect 717 721 763 861
rect 921 721 967 861
<< polysilicon >>
rect 144 939 244 983
rect 348 939 448 983
rect 588 939 688 983
rect 792 939 892 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 377 244 454
rect 124 333 244 377
rect 348 500 448 573
rect 348 454 377 500
rect 423 454 448 500
rect 348 377 448 454
rect 588 500 688 647
rect 588 454 601 500
rect 647 454 688 500
rect 588 377 688 454
rect 792 500 892 647
rect 792 454 809 500
rect 855 454 892 500
rect 792 377 892 454
rect 348 333 468 377
rect 578 333 698 377
rect 772 333 892 377
rect 124 25 244 69
rect 348 25 468 69
rect 578 25 698 69
rect 772 25 892 69
<< polycontact >>
rect 157 454 203 500
rect 377 454 423 500
rect 601 454 647 500
rect 809 454 855 500
<< metal1 >>
rect 0 918 1120 1098
rect 69 861 115 918
rect 69 710 115 721
rect 477 861 523 872
rect 477 664 523 721
rect 717 861 763 918
rect 717 710 763 721
rect 921 861 967 872
rect 921 664 967 721
rect 254 618 967 664
rect 142 500 203 542
rect 142 454 157 500
rect 142 443 203 454
rect 49 320 95 331
rect 254 285 319 618
rect 366 500 434 542
rect 366 454 377 500
rect 423 454 434 500
rect 590 500 658 542
rect 590 454 601 500
rect 647 454 658 500
rect 798 500 866 542
rect 798 454 809 500
rect 855 454 866 500
rect 254 239 273 285
rect 254 228 319 239
rect 497 320 543 331
rect 95 180 497 182
rect 49 136 543 180
rect 921 320 967 331
rect 921 90 967 180
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 366 454 434 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 142 443 203 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 590 454 658 542 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 798 454 866 542 0 FreeSans 200 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 921 90 967 331 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 921 664 967 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
rlabel metal1 s 477 664 523 872 1 ZN
port 5 nsew default output
rlabel metal1 s 254 618 967 664 1 ZN
port 5 nsew default output
rlabel metal1 s 254 228 319 618 1 ZN
port 5 nsew default output
rlabel metal1 s 717 710 763 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 202482
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 198866
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
