magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 568 822
<< polysilicon >>
rect -31 681 88 754
rect 193 681 312 754
rect -31 -74 89 -1
rect 193 -74 313 -1
use pmos_5p04310590548731_128x8m81  pmos_5p04310590548731_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 802
<< properties >>
string GDS_END 316344
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 315902
<< end >>
