magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -71 66 71 71
rect -71 -66 -66 66
rect 66 -66 71 66
rect -71 -71 71 -66
<< via2 >>
rect -66 -66 66 66
<< metal3 >>
rect -71 66 71 71
rect -71 -66 -66 66
rect 66 -66 71 66
rect -71 -71 71 -66
<< properties >>
string GDS_END 524536
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 523828
<< end >>
