magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 2016 844
rect 48 563 116 724
rect 497 540 543 676
rect 934 563 1002 724
rect 1393 540 1439 676
rect 1820 563 1888 724
rect 234 517 774 540
rect 1130 517 1439 540
rect 26 470 1439 517
rect 26 219 86 470
rect 330 360 1683 424
rect 1812 312 1884 451
rect 159 265 1884 312
rect 1608 244 1884 265
rect 26 173 1546 219
rect 36 60 108 127
rect 273 106 319 173
rect 486 60 554 127
rect 721 106 767 173
rect 934 60 1002 127
rect 1169 106 1215 173
rect 1500 152 1546 173
rect 1382 60 1450 127
rect 1500 106 1682 152
rect 1828 60 1900 127
rect 0 -60 2016 60
<< labels >>
rlabel metal1 s 330 360 1683 424 6 A1
port 1 nsew default input
rlabel metal1 s 1812 312 1884 451 6 A2
port 2 nsew default input
rlabel metal1 s 159 265 1884 312 6 A2
port 2 nsew default input
rlabel metal1 s 1608 244 1884 265 6 A2
port 2 nsew default input
rlabel metal1 s 1393 540 1439 676 6 ZN
port 3 nsew default output
rlabel metal1 s 497 540 543 676 6 ZN
port 3 nsew default output
rlabel metal1 s 1130 517 1439 540 6 ZN
port 3 nsew default output
rlabel metal1 s 234 517 774 540 6 ZN
port 3 nsew default output
rlabel metal1 s 26 470 1439 517 6 ZN
port 3 nsew default output
rlabel metal1 s 26 219 86 470 6 ZN
port 3 nsew default output
rlabel metal1 s 26 173 1546 219 6 ZN
port 3 nsew default output
rlabel metal1 s 1500 152 1546 173 6 ZN
port 3 nsew default output
rlabel metal1 s 1169 152 1215 173 6 ZN
port 3 nsew default output
rlabel metal1 s 721 152 767 173 6 ZN
port 3 nsew default output
rlabel metal1 s 273 152 319 173 6 ZN
port 3 nsew default output
rlabel metal1 s 1500 106 1682 152 6 ZN
port 3 nsew default output
rlabel metal1 s 1169 106 1215 152 6 ZN
port 3 nsew default output
rlabel metal1 s 721 106 767 152 6 ZN
port 3 nsew default output
rlabel metal1 s 273 106 319 152 6 ZN
port 3 nsew default output
rlabel metal1 s 0 724 2016 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1820 563 1888 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 934 563 1002 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 48 563 116 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1828 60 1900 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 36 60 108 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2016 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 733360
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 729006
<< end >>
