magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 147 64 159
rect 11 106 16 147
rect 28 93 33 140
rect 46 106 51 147
rect 28 91 37 93
rect 28 85 40 91
rect 28 82 37 85
rect 13 67 23 73
rect 11 9 16 33
rect 28 16 33 82
rect 45 9 50 33
rect 0 -3 64 9
<< metal2 >>
rect 10 154 18 155
rect 9 148 19 154
rect 10 147 18 148
rect 30 84 40 92
rect 13 66 23 74
rect 10 8 18 9
rect 9 2 19 8
rect 10 1 18 2
<< labels >>
rlabel metal2 s 13 66 23 74 6 A
port 1 nsew signal input
rlabel metal1 s 13 67 23 73 6 A
port 1 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 46 106 51 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 147 64 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 -3 50 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 -3 64 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 30 84 40 92 6 Y
port 2 nsew signal output
rlabel metal1 s 28 16 33 140 6 Y
port 2 nsew signal output
rlabel metal1 s 28 82 37 93 6 Y
port 2 nsew signal output
rlabel metal1 s 28 85 40 91 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 64 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 174128
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 169808
<< end >>
