magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect -17 147 95 159
rect 11 106 16 147
rect 28 100 33 140
rect 45 106 50 147
rect 62 100 67 140
rect 79 106 84 147
rect 28 94 70 100
rect 4 80 14 86
rect 28 43 33 94
rect 62 43 67 94
rect 28 38 67 43
rect 11 9 16 33
rect 28 16 33 38
rect 45 9 50 33
rect 62 16 67 38
rect 79 9 84 33
rect -17 -3 95 9
<< obsm1 >>
rect -6 61 -1 140
rect -6 55 23 61
rect -6 16 -1 55
<< metal2 >>
rect -7 154 1 155
rect 17 154 25 155
rect 41 154 49 155
rect 65 154 73 155
rect -8 148 2 154
rect 16 148 26 154
rect 40 148 50 154
rect 64 148 74 154
rect -7 147 1 148
rect 17 147 25 148
rect 41 147 49 148
rect 65 147 73 148
rect 60 100 70 101
rect 59 94 70 100
rect 60 93 70 94
rect 5 86 13 87
rect 4 80 14 86
rect 5 79 13 80
rect -7 8 1 9
rect 17 8 25 9
rect 41 8 49 9
rect 65 8 73 9
rect -8 2 2 8
rect 16 2 26 8
rect 40 2 50 8
rect 64 2 74 8
rect -7 1 1 2
rect 17 1 25 2
rect 41 1 49 2
rect 65 1 73 2
<< labels >>
rlabel metal2 s 5 79 13 87 6 A
port 1 nsew signal input
rlabel metal2 s 4 80 14 86 6 A
port 1 nsew signal input
rlabel metal1 s 4 80 14 86 6 A
port 1 nsew signal input
rlabel metal2 s -7 147 1 155 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s -8 148 2 154 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 17 147 25 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 16 148 26 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 41 147 49 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 40 148 50 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 65 147 73 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 64 148 74 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 45 106 50 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 79 106 84 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s -17 147 95 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s -7 1 1 9 4 VSS
port 6 nsew ground bidirectional
rlabel metal2 s -8 2 2 8 4 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 17 1 25 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 16 2 26 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 41 1 49 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 40 2 50 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 65 1 73 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 64 2 74 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 -3 50 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 79 -3 84 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s -17 -3 95 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 59 94 70 100 6 Y
port 2 nsew signal output
rlabel metal2 s 60 93 70 101 6 Y
port 2 nsew signal output
rlabel metal1 s 28 16 33 140 6 Y
port 2 nsew signal output
rlabel metal1 s 28 38 67 43 6 Y
port 2 nsew signal output
rlabel metal1 s 62 16 67 140 6 Y
port 2 nsew signal output
rlabel metal1 s 28 94 70 100 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX -17 -3 95 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 130302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 121374
<< end >>
