magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 4342 870
<< pwell >>
rect -86 -86 4342 352
<< mvnmos >>
rect 124 156 244 232
rect 348 156 468 232
rect 660 156 780 232
rect 884 156 1004 232
rect 1108 156 1228 232
rect 1332 156 1452 232
rect 1556 156 1676 232
rect 1780 156 1900 232
rect 2232 156 2352 229
rect 2475 156 2595 229
rect 2872 156 2992 229
rect 3096 156 3216 229
rect 3320 156 3440 229
rect 3544 156 3664 229
rect 3768 156 3888 229
rect 3992 156 4112 229
<< mvpmos >>
rect 124 472 224 628
rect 424 472 524 628
rect 628 472 728 628
rect 884 472 984 628
rect 1148 472 1248 628
rect 1352 472 1452 628
rect 1556 472 1656 628
rect 1760 472 1860 628
rect 2220 509 2320 628
rect 2496 509 2596 628
rect 2892 509 2992 628
rect 3116 509 3216 628
rect 3320 509 3420 628
rect 3524 509 3624 628
rect 3768 509 3868 628
rect 3992 509 4092 628
<< mvndiff >>
rect 36 215 124 232
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 232
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 215 660 232
rect 468 169 525 215
rect 571 169 660 215
rect 468 156 660 169
rect 780 215 884 232
rect 780 169 809 215
rect 855 169 884 215
rect 780 156 884 169
rect 1004 215 1108 232
rect 1004 169 1033 215
rect 1079 169 1108 215
rect 1004 156 1108 169
rect 1228 215 1332 232
rect 1228 169 1257 215
rect 1303 169 1332 215
rect 1228 156 1332 169
rect 1452 215 1556 232
rect 1452 169 1481 215
rect 1527 169 1556 215
rect 1452 156 1556 169
rect 1676 215 1780 232
rect 1676 169 1705 215
rect 1751 169 1780 215
rect 1676 156 1780 169
rect 1900 215 1988 232
rect 1900 169 1929 215
rect 1975 169 1988 215
rect 1900 156 1988 169
rect 2082 215 2232 229
rect 2082 169 2095 215
rect 2141 169 2232 215
rect 2082 156 2232 169
rect 2352 215 2475 229
rect 2352 169 2381 215
rect 2427 169 2475 215
rect 2352 156 2475 169
rect 2595 215 2684 229
rect 2595 169 2625 215
rect 2671 169 2684 215
rect 2595 156 2684 169
rect 2784 216 2872 229
rect 2784 170 2797 216
rect 2843 170 2872 216
rect 2784 156 2872 170
rect 2992 216 3096 229
rect 2992 170 3021 216
rect 3067 170 3096 216
rect 2992 156 3096 170
rect 3216 216 3320 229
rect 3216 170 3245 216
rect 3291 170 3320 216
rect 3216 156 3320 170
rect 3440 216 3544 229
rect 3440 170 3469 216
rect 3515 170 3544 216
rect 3440 156 3544 170
rect 3664 216 3768 229
rect 3664 170 3693 216
rect 3739 170 3768 216
rect 3664 156 3768 170
rect 3888 216 3992 229
rect 3888 170 3917 216
rect 3963 170 3992 216
rect 3888 156 3992 170
rect 4112 216 4200 229
rect 4112 170 4141 216
rect 4187 170 4200 216
rect 4112 156 4200 170
<< mvpdiff >>
rect 36 579 124 628
rect 36 533 49 579
rect 95 533 124 579
rect 36 472 124 533
rect 224 579 424 628
rect 224 533 253 579
rect 299 533 424 579
rect 224 472 424 533
rect 524 605 628 628
rect 524 559 553 605
rect 599 559 628 605
rect 524 472 628 559
rect 728 574 884 628
rect 728 528 797 574
rect 843 528 884 574
rect 728 472 884 528
rect 984 615 1148 628
rect 984 569 1035 615
rect 1081 569 1148 615
rect 984 472 1148 569
rect 1248 574 1352 628
rect 1248 528 1277 574
rect 1323 528 1352 574
rect 1248 472 1352 528
rect 1452 615 1556 628
rect 1452 569 1481 615
rect 1527 569 1556 615
rect 1452 472 1556 569
rect 1656 574 1760 628
rect 1656 528 1685 574
rect 1731 528 1760 574
rect 1656 472 1760 528
rect 1860 615 1976 628
rect 1860 569 1917 615
rect 1963 569 1976 615
rect 1860 472 1976 569
rect 2085 590 2220 628
rect 2085 544 2098 590
rect 2144 544 2220 590
rect 2085 509 2220 544
rect 2320 590 2496 628
rect 2320 544 2367 590
rect 2413 544 2496 590
rect 2320 509 2496 544
rect 2596 590 2684 628
rect 2596 544 2625 590
rect 2671 544 2684 590
rect 2596 509 2684 544
rect 2804 574 2892 628
rect 2804 528 2817 574
rect 2863 528 2892 574
rect 2804 509 2892 528
rect 2992 615 3116 628
rect 2992 569 3041 615
rect 3087 569 3116 615
rect 2992 509 3116 569
rect 3216 574 3320 628
rect 3216 528 3245 574
rect 3291 528 3320 574
rect 3216 509 3320 528
rect 3420 574 3524 628
rect 3420 528 3449 574
rect 3495 528 3524 574
rect 3420 509 3524 528
rect 3624 609 3768 628
rect 3624 563 3676 609
rect 3722 563 3768 609
rect 3624 509 3768 563
rect 3868 609 3992 628
rect 3868 563 3897 609
rect 3943 563 3992 609
rect 3868 509 3992 563
rect 4092 609 4180 628
rect 4092 563 4121 609
rect 4167 563 4180 609
rect 4092 509 4180 563
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 525 169 571 215
rect 809 169 855 215
rect 1033 169 1079 215
rect 1257 169 1303 215
rect 1481 169 1527 215
rect 1705 169 1751 215
rect 1929 169 1975 215
rect 2095 169 2141 215
rect 2381 169 2427 215
rect 2625 169 2671 215
rect 2797 170 2843 216
rect 3021 170 3067 216
rect 3245 170 3291 216
rect 3469 170 3515 216
rect 3693 170 3739 216
rect 3917 170 3963 216
rect 4141 170 4187 216
<< mvpdiffc >>
rect 49 533 95 579
rect 253 533 299 579
rect 553 559 599 605
rect 797 528 843 574
rect 1035 569 1081 615
rect 1277 528 1323 574
rect 1481 569 1527 615
rect 1685 528 1731 574
rect 1917 569 1963 615
rect 2098 544 2144 590
rect 2367 544 2413 590
rect 2625 544 2671 590
rect 2817 528 2863 574
rect 3041 569 3087 615
rect 3245 528 3291 574
rect 3449 528 3495 574
rect 3676 563 3722 609
rect 3897 563 3943 609
rect 4121 563 4167 609
<< polysilicon >>
rect 628 720 3420 760
rect 124 628 224 672
rect 424 628 524 672
rect 628 628 728 720
rect 884 628 984 672
rect 1148 628 1248 672
rect 1352 628 1452 672
rect 1556 628 1656 672
rect 1760 628 1860 672
rect 2220 628 2320 672
rect 2496 628 2596 672
rect 2892 628 2992 672
rect 3116 628 3216 672
rect 3320 628 3420 720
rect 3524 720 4092 760
rect 3524 628 3624 720
rect 3768 628 3868 672
rect 3992 628 4092 720
rect 124 394 224 472
rect 124 348 141 394
rect 187 380 224 394
rect 424 439 524 472
rect 424 393 451 439
rect 497 393 524 439
rect 628 412 728 472
rect 424 380 524 393
rect 187 348 244 380
rect 124 232 244 348
rect 572 372 728 412
rect 884 408 984 472
rect 884 394 1004 408
rect 572 332 612 372
rect 348 292 612 332
rect 884 348 928 394
rect 974 348 1004 394
rect 1148 364 1248 472
rect 1352 364 1452 472
rect 1556 364 1656 472
rect 1760 364 1860 472
rect 2220 409 2320 509
rect 2496 468 2596 509
rect 2496 422 2509 468
rect 2555 449 2596 468
rect 2892 449 2992 509
rect 2555 422 2992 449
rect 3116 426 3216 509
rect 2496 409 2992 422
rect 2220 369 2448 409
rect 660 311 780 324
rect 348 232 468 292
rect 660 265 679 311
rect 725 265 780 311
rect 660 232 780 265
rect 884 232 1004 348
rect 1108 351 2172 364
rect 1108 305 2113 351
rect 2159 305 2172 351
rect 2400 361 2448 369
rect 2400 348 2777 361
rect 2400 321 2718 348
rect 1108 304 2172 305
rect 1108 232 1228 304
rect 1332 232 1452 304
rect 1556 232 1676 304
rect 1780 292 2172 304
rect 2232 308 2352 321
rect 1780 232 1900 292
rect 2232 262 2293 308
rect 2339 262 2352 308
rect 2232 229 2352 262
rect 2475 302 2718 321
rect 2764 302 2777 348
rect 2475 289 2777 302
rect 2475 229 2595 289
rect 2872 229 2992 409
rect 3096 414 3216 426
rect 3096 368 3130 414
rect 3176 368 3216 414
rect 3096 229 3216 368
rect 3320 405 3420 509
rect 3524 465 3624 509
rect 3768 431 3868 509
rect 3768 412 3888 431
rect 3320 392 3712 405
rect 3320 352 3653 392
rect 3544 346 3653 352
rect 3699 346 3712 392
rect 3544 333 3712 346
rect 3768 366 3801 412
rect 3847 366 3888 412
rect 3320 229 3440 273
rect 3544 229 3664 333
rect 3768 229 3888 366
rect 3992 355 4092 509
rect 3992 229 4112 355
rect 124 112 244 156
rect 348 112 468 156
rect 660 64 780 156
rect 884 112 1004 156
rect 1108 112 1228 156
rect 1332 112 1452 156
rect 1556 112 1676 156
rect 1780 112 1900 156
rect 2232 112 2352 156
rect 2475 112 2595 156
rect 2872 112 2992 156
rect 3096 112 3216 156
rect 3320 64 3440 156
rect 3544 112 3664 156
rect 3768 112 3888 156
rect 3992 64 4112 156
rect 660 24 4112 64
<< polycontact >>
rect 141 348 187 394
rect 451 393 497 439
rect 928 348 974 394
rect 2509 422 2555 468
rect 679 265 725 311
rect 2113 305 2159 351
rect 2293 262 2339 308
rect 2718 302 2764 348
rect 3130 368 3176 414
rect 3653 346 3699 392
rect 3801 366 3847 412
<< metal1 >>
rect 0 724 4256 844
rect 49 579 95 724
rect 542 620 947 666
rect 542 605 610 620
rect 542 594 553 605
rect 252 579 299 590
rect 49 515 95 533
rect 141 394 202 567
rect 187 348 202 394
rect 49 215 95 226
rect 141 205 202 348
rect 252 533 253 579
rect 252 215 299 533
rect 345 559 553 594
rect 599 559 610 605
rect 345 548 610 559
rect 345 314 391 548
rect 786 528 797 574
rect 843 528 855 574
rect 451 439 740 450
rect 497 393 740 439
rect 451 360 740 393
rect 345 268 458 314
rect 408 215 458 268
rect 660 311 740 360
rect 660 265 679 311
rect 725 265 740 311
rect 660 248 740 265
rect 786 215 855 528
rect 901 523 947 620
rect 1024 615 1092 724
rect 1024 569 1035 615
rect 1081 569 1092 615
rect 1151 632 1424 678
rect 1151 523 1197 632
rect 901 476 1197 523
rect 1246 574 1323 585
rect 1246 528 1277 574
rect 1246 430 1323 528
rect 1378 523 1424 632
rect 1470 615 1538 724
rect 1470 569 1481 615
rect 1527 569 1538 615
rect 1584 631 1860 678
rect 1584 523 1630 631
rect 1378 476 1630 523
rect 1685 574 1768 585
rect 1731 528 1768 574
rect 1685 430 1768 528
rect 1814 523 1860 631
rect 1906 615 1974 724
rect 1906 569 1917 615
rect 1963 569 1974 615
rect 2098 590 2144 601
rect 2098 523 2144 544
rect 1814 476 2144 523
rect 2190 544 2367 590
rect 2413 544 2424 590
rect 252 169 273 215
rect 319 169 330 215
rect 408 169 525 215
rect 571 169 582 215
rect 786 169 809 215
rect 49 60 95 169
rect 786 156 855 169
rect 901 394 1151 430
rect 901 348 928 394
rect 974 360 1151 394
rect 1246 360 1768 430
rect 974 348 987 360
rect 901 110 987 348
rect 1033 215 1079 232
rect 1033 60 1079 169
rect 1246 215 1320 360
rect 1246 169 1257 215
rect 1303 169 1320 215
rect 1246 120 1320 169
rect 1481 215 1527 232
rect 1481 60 1527 169
rect 1685 215 1768 360
rect 1685 169 1705 215
rect 1751 169 1768 215
rect 1685 120 1768 169
rect 1929 215 1975 232
rect 1929 60 1975 169
rect 2021 226 2067 476
rect 2190 364 2236 544
rect 2481 468 2555 664
rect 2481 430 2509 468
rect 2113 351 2236 364
rect 2159 305 2236 351
rect 2113 292 2236 305
rect 2021 215 2144 226
rect 2021 169 2095 215
rect 2141 169 2144 215
rect 2190 215 2236 292
rect 2282 422 2509 430
rect 2282 354 2555 422
rect 2625 632 2966 678
rect 2625 590 2671 632
rect 2282 308 2355 354
rect 2282 262 2293 308
rect 2339 262 2355 308
rect 2282 261 2355 262
rect 2625 215 2671 544
rect 2190 169 2381 215
rect 2427 169 2438 215
rect 2021 158 2144 169
rect 2625 156 2671 169
rect 2717 574 2863 585
rect 2717 528 2817 574
rect 2717 515 2863 528
rect 2920 523 2966 632
rect 3029 615 3098 724
rect 3029 569 3041 615
rect 3087 569 3098 615
rect 3148 632 3515 678
rect 3148 523 3194 632
rect 2717 348 2767 515
rect 2920 476 3194 523
rect 3245 574 3291 585
rect 2815 414 3195 426
rect 2815 368 3130 414
rect 3176 368 3195 414
rect 2815 356 3195 368
rect 2717 302 2718 348
rect 2764 302 2767 348
rect 2717 229 2767 302
rect 2717 216 2863 229
rect 2717 170 2797 216
rect 2843 170 2863 216
rect 2717 159 2863 170
rect 3021 216 3067 229
rect 3021 60 3067 170
rect 3245 216 3291 528
rect 3245 156 3291 170
rect 3449 574 3515 632
rect 3886 609 3954 724
rect 3495 528 3515 574
rect 3449 216 3515 528
rect 3449 170 3469 216
rect 3561 563 3676 609
rect 3722 563 3733 609
rect 3886 563 3897 609
rect 3943 563 3954 609
rect 4120 609 4187 628
rect 4120 563 4121 609
rect 4167 563 4187 609
rect 3561 216 3607 563
rect 4120 517 4187 563
rect 3653 471 4187 517
rect 3653 392 3699 471
rect 3745 412 4083 424
rect 3745 366 3801 412
rect 3847 366 4083 412
rect 3745 356 4083 366
rect 3653 335 3699 346
rect 3917 216 3963 229
rect 3561 170 3693 216
rect 3739 170 3750 216
rect 3449 156 3515 170
rect 3917 60 3963 170
rect 4141 216 4187 471
rect 4141 156 4187 170
rect 0 -60 4256 60
<< labels >>
flabel metal1 s 3745 356 4083 424 0 FreeSans 400 0 0 0 I0
port 1 nsew default input
flabel metal1 s 1929 229 1975 232 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 0 724 4256 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 141 205 202 567 0 FreeSans 400 0 0 0 I2
port 3 nsew default input
flabel metal1 s 2815 356 3195 426 0 FreeSans 400 0 0 0 I1
port 2 nsew default input
flabel metal1 s 451 360 740 450 0 FreeSans 400 0 0 0 S0
port 5 nsew default input
flabel metal1 s 901 360 1151 430 0 FreeSans 400 0 0 0 I3
port 4 nsew default input
flabel metal1 s 2481 430 2555 664 0 FreeSans 400 0 0 0 S1
port 6 nsew default input
flabel metal1 s 1685 430 1768 585 0 FreeSans 400 0 0 0 Z
port 7 nsew default output
rlabel metal1 s 901 110 987 360 1 I3
port 4 nsew default input
rlabel metal1 s 660 248 740 360 1 S0
port 5 nsew default input
rlabel metal1 s 2282 354 2555 430 1 S1
port 6 nsew default input
rlabel metal1 s 2282 261 2355 354 1 S1
port 6 nsew default input
rlabel metal1 s 1246 430 1323 585 1 Z
port 7 nsew default output
rlabel metal1 s 1246 360 1768 430 1 Z
port 7 nsew default output
rlabel metal1 s 1685 120 1768 360 1 Z
port 7 nsew default output
rlabel metal1 s 1246 120 1320 360 1 Z
port 7 nsew default output
rlabel metal1 s 3886 569 3954 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3029 569 3098 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1906 569 1974 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1470 569 1538 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1024 569 1092 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 569 95 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3886 563 3954 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 563 95 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 515 95 563 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1481 229 1527 232 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1033 229 1079 232 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3917 226 3963 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3021 226 3067 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1929 226 1975 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1481 226 1527 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1033 226 1079 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3917 60 3963 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3021 60 3067 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1929 60 1975 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1481 60 1527 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1033 60 1079 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string GDS_END 685642
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 677120
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
