magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< obsm1 >>
rect -32 13108 15032 69957
<< metal2 >>
rect 272 69800 2172 70000
rect 2752 69800 4802 70000
rect 5122 69800 7172 70000
rect 7828 69800 9878 70000
rect 10198 69800 12248 70000
rect 12828 69800 14728 70000
<< obsm2 >>
rect 0 69740 212 69800
rect 2232 69740 2692 69800
rect 4862 69740 5062 69800
rect 7232 69740 7768 69800
rect 9938 69740 10138 69800
rect 12308 69740 12768 69800
rect 14788 69740 15000 69800
rect 0 0 15000 69740
<< metal3 >>
rect 0 68400 200 69678
rect 0 66800 2502 68200
rect 0 65200 200 66600
rect 14800 68400 15000 69678
rect 12498 66800 15000 68200
rect 0 63600 200 65000
rect 14800 65200 15000 66600
rect 14800 63600 15000 65000
rect 0 62000 2313 63400
rect 2369 62000 15000 63400
rect 0 60400 200 61800
rect 0 58800 2502 60200
rect 0 57200 200 58600
rect 14800 60400 15000 61800
rect 12498 58800 15000 60200
rect 0 55600 2502 57000
rect 0 54000 2502 55400
rect 0 52400 2502 53800
rect 14800 57200 15000 58600
rect 12498 55600 15000 57000
rect 12498 54000 15000 55400
rect 12498 52400 15000 53800
rect 0 50800 2313 52200
rect 2369 50800 15000 52200
rect 0 49200 200 50600
rect 0 46000 200 49000
rect 14800 49200 15000 50600
rect 0 42800 2502 45800
rect 0 41200 2502 42600
rect 0 39600 200 41000
rect 14800 46000 15000 49000
rect 12498 42800 15000 45800
rect 12498 41200 15000 42600
rect 0 36400 2502 39400
rect 0 33200 2502 36200
rect 0 30000 2502 33000
rect 0 26800 2502 29800
rect 0 25200 200 26600
rect 14800 39600 15000 41000
rect 12498 36400 15000 39400
rect 12498 33200 15000 36200
rect 12498 30000 15000 33000
rect 12498 26800 15000 29800
rect 0 23600 2502 25000
rect 0 20400 200 23400
rect 14800 25200 15000 26600
rect 12498 23600 15000 25000
rect 0 17200 200 20200
rect 0 14000 200 17000
rect 14800 20400 15000 23400
rect 14800 17200 15000 20200
rect 14800 14000 15000 17000
<< obsm3 >>
rect 560 68560 14440 69678
rect 2862 66440 12138 68560
rect 560 63760 14440 66440
rect 560 60560 14440 61640
rect 2862 58440 12138 60560
rect 560 57360 14440 58440
rect 2862 52560 12138 57360
rect 560 46160 14440 50440
rect 2862 40840 12138 46160
rect 560 39760 14440 40840
rect 2862 26440 12138 39760
rect 560 25360 14440 26440
rect 2862 23240 12138 25360
rect 560 13640 14440 23240
rect 200 0 14800 13640
<< labels >>
rlabel metal3 s 12498 23600 15000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 36400 15000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 33200 15000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 30000 15000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 26800 15000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 42800 15000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 41200 15000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 55600 15000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 54000 15000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 52400 15000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 58800 15000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 12498 66800 15000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 66800 2502 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 2502 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 2502 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 2502 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 2502 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 2502 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 2502 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 2502 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 2502 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 2502 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 2502 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 2502 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 20400 15000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 17200 15000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 14000 15000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 25200 15000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 39600 15000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 46000 15000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 49200 15000 50600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 57200 15000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 60400 15000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 63600 15000 65000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 65200 15000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 68400 15000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 272 69800 2172 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 2752 69800 4802 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 5122 69800 7172 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 7828 69800 9878 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 10198 69800 12248 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 12828 69800 14728 70000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 2369 50800 15000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 2369 62000 15000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 62000 2313 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 2313 52200 6 VDD
port 3 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD POWER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4240138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4238430
<< end >>
