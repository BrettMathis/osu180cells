magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 672 844
rect 49 528 95 724
rect 244 536 334 678
rect 503 586 549 724
rect 244 472 536 536
rect 126 341 430 424
rect 476 295 536 472
rect 279 244 536 295
rect 49 60 95 190
rect 279 106 325 244
rect 503 60 549 190
rect 0 -60 672 60
<< labels >>
rlabel metal1 s 126 341 430 424 6 I
port 1 nsew default input
rlabel metal1 s 244 536 334 678 6 ZN
port 2 nsew default output
rlabel metal1 s 244 472 536 536 6 ZN
port 2 nsew default output
rlabel metal1 s 476 295 536 472 6 ZN
port 2 nsew default output
rlabel metal1 s 279 244 536 295 6 ZN
port 2 nsew default output
rlabel metal1 s 279 106 325 244 6 ZN
port 2 nsew default output
rlabel metal1 s 0 724 672 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 503 586 549 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 586 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 528 95 586 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 503 60 549 190 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 190 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 672 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 469870
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 467434
<< end >>
