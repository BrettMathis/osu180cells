magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect 22205 9106 22518 9125
rect 22205 8971 22453 9106
rect 22434 8966 22453 8971
rect 22499 8966 22518 9106
rect 22434 8947 22518 8966
rect 22205 7482 22573 7583
rect 22205 7436 22454 7482
rect 22500 7436 22573 7482
rect 22205 7429 22573 7436
rect 22381 7325 22573 7429
rect 22205 7318 22573 7325
rect 22205 7272 22454 7318
rect 22500 7272 22573 7318
rect 22205 7171 22573 7272
rect 22205 5682 22573 5783
rect 22205 5636 22454 5682
rect 22500 5636 22573 5682
rect 22205 5629 22573 5636
rect 22381 5525 22573 5629
rect 22205 5518 22573 5525
rect 22205 5472 22454 5518
rect 22500 5472 22573 5518
rect 22205 5371 22573 5472
rect 22205 3882 22573 3983
rect 22205 3836 22454 3882
rect 22500 3836 22573 3882
rect 22205 3829 22573 3836
rect 22381 3725 22573 3829
rect 22205 3718 22573 3725
rect 22205 3672 22454 3718
rect 22500 3672 22573 3718
rect 22205 3571 22573 3672
rect 22205 2082 22573 2183
rect 22205 2036 22454 2082
rect 22500 2036 22573 2082
rect 22205 2029 22573 2036
rect 22381 1925 22573 2029
rect 22205 1918 22573 1925
rect 22205 1872 22454 1918
rect 22500 1872 22573 1918
rect 22205 1771 22573 1872
rect 22381 522 22573 568
rect 22381 476 22454 522
rect 22500 476 22573 522
rect 22381 383 22573 476
rect 22205 358 22573 383
rect 22205 312 22454 358
rect 22500 312 22573 358
rect 22205 229 22573 312
<< polycontact >>
rect 22453 8966 22499 9106
rect 22454 7436 22500 7482
rect 22454 7272 22500 7318
rect 22454 5636 22500 5682
rect 22454 5472 22500 5518
rect 22454 3836 22500 3882
rect 22454 3672 22500 3718
rect 22454 2036 22500 2082
rect 22454 1872 22500 1918
rect 22454 476 22500 522
rect 22454 312 22500 358
<< metal1 >>
rect 22438 9106 22514 9117
rect 22438 9105 22453 9106
rect 22499 9105 22514 9106
rect 22438 8845 22450 9105
rect 22502 8845 22514 9105
rect 22438 8833 22514 8845
rect 22413 7514 22537 7554
rect 22413 7462 22449 7514
rect 22501 7462 22537 7514
rect 22413 7436 22454 7462
rect 22500 7436 22537 7462
rect 22413 7318 22537 7436
rect 22413 7296 22454 7318
rect 22500 7296 22537 7318
rect 22413 7244 22449 7296
rect 22501 7244 22537 7296
rect 22413 7204 22537 7244
rect 22413 5710 22537 5750
rect 22413 5658 22449 5710
rect 22501 5658 22537 5710
rect 22413 5636 22454 5658
rect 22500 5636 22537 5658
rect 22413 5518 22537 5636
rect 22413 5492 22454 5518
rect 22500 5492 22537 5518
rect 22413 5440 22449 5492
rect 22501 5440 22537 5492
rect 22413 5400 22537 5440
rect 22413 3914 22537 3954
rect 22413 3862 22449 3914
rect 22501 3862 22537 3914
rect 22413 3836 22454 3862
rect 22500 3836 22537 3862
rect 22413 3718 22537 3836
rect 22413 3696 22454 3718
rect 22500 3696 22537 3718
rect 22413 3644 22449 3696
rect 22501 3644 22537 3696
rect 22413 3604 22537 3644
rect 22413 2110 22537 2150
rect 22413 2058 22449 2110
rect 22501 2058 22537 2110
rect 22413 2036 22454 2058
rect 22500 2036 22537 2058
rect 22413 1918 22537 2036
rect 22413 1892 22454 1918
rect 22500 1892 22537 1918
rect 22413 1840 22449 1892
rect 22501 1840 22537 1892
rect 22413 1800 22537 1840
rect 22421 522 22533 559
rect 22421 476 22454 522
rect 22500 476 22533 522
rect 22421 457 22533 476
rect 22421 301 22449 457
rect 22501 301 22533 457
rect 22421 276 22533 301
<< via1 >>
rect 22450 8966 22453 9105
rect 22453 8966 22499 9105
rect 22499 8966 22502 9105
rect 22450 8845 22502 8966
rect 22449 7482 22501 7514
rect 22449 7462 22454 7482
rect 22454 7462 22500 7482
rect 22500 7462 22501 7482
rect 22449 7272 22454 7296
rect 22454 7272 22500 7296
rect 22500 7272 22501 7296
rect 22449 7244 22501 7272
rect 22449 5682 22501 5710
rect 22449 5658 22454 5682
rect 22454 5658 22500 5682
rect 22500 5658 22501 5682
rect 22449 5472 22454 5492
rect 22454 5472 22500 5492
rect 22500 5472 22501 5492
rect 22449 5440 22501 5472
rect 22449 3882 22501 3914
rect 22449 3862 22454 3882
rect 22454 3862 22500 3882
rect 22500 3862 22501 3882
rect 22449 3672 22454 3696
rect 22454 3672 22500 3696
rect 22500 3672 22501 3696
rect 22449 3644 22501 3672
rect 22449 2082 22501 2110
rect 22449 2058 22454 2082
rect 22454 2058 22500 2082
rect 22500 2058 22501 2082
rect 22449 1872 22454 1892
rect 22454 1872 22500 1892
rect 22500 1872 22501 1892
rect 22449 1840 22501 1872
rect 22449 358 22501 457
rect 22449 312 22454 358
rect 22454 312 22500 358
rect 22500 312 22501 358
rect 22449 301 22501 312
<< metal2 >>
rect 22412 9258 22537 9277
rect 22412 9098 22448 9258
rect 22504 9098 22537 9258
rect 22412 8845 22450 9098
rect 22502 8845 22537 9098
rect 22412 7514 22537 8845
rect 22412 7462 22449 7514
rect 22501 7462 22537 7514
rect 22412 7296 22537 7462
rect 22412 7244 22449 7296
rect 22501 7244 22537 7296
rect 22412 5710 22537 7244
rect 22412 5658 22449 5710
rect 22501 5658 22537 5710
rect 22412 5492 22537 5658
rect 22412 5440 22449 5492
rect 22501 5440 22537 5492
rect 22412 3914 22537 5440
rect 22412 3862 22449 3914
rect 22501 3862 22537 3914
rect 22412 3696 22537 3862
rect 22412 3644 22449 3696
rect 22501 3644 22537 3696
rect 22412 2110 22537 3644
rect 22412 2058 22449 2110
rect 22501 2058 22537 2110
rect 22412 1892 22537 2058
rect 22412 1840 22449 1892
rect 22501 1840 22537 1892
rect 22412 457 22537 1840
rect 22412 301 22449 457
rect 22501 301 22537 457
rect 22412 261 22537 301
rect 22412 101 22447 261
rect 22503 101 22537 261
rect 22412 76 22537 101
<< via2 >>
rect 22448 9105 22504 9258
rect 22448 9098 22450 9105
rect 22450 9098 22502 9105
rect 22502 9098 22504 9105
rect 22447 101 22503 261
<< metal3 >>
rect -636 9258 22538 9277
rect -636 9098 22448 9258
rect 22504 9098 22538 9258
rect -636 9077 22538 9098
rect -636 261 22540 277
rect -636 101 22447 261
rect 22503 101 22540 261
rect -636 77 22540 101
use 018SRAM_cell1_64x8m81  018SRAM_cell1_64x8m81_0
timestamp 1669390400
transform -1 0 22262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_64x8m81  018SRAM_cell1_64x8m81_1
timestamp 1669390400
transform -1 0 22262 0 -1 9177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_0
timestamp 1669390400
transform -1 0 22262 0 1 1977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_1
timestamp 1669390400
transform -1 0 22262 0 1 3777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_2
timestamp 1669390400
transform -1 0 22262 0 1 5577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_3
timestamp 1669390400
transform -1 0 22262 0 1 7377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_4
timestamp 1669390400
transform -1 0 22262 0 -1 7377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_5
timestamp 1669390400
transform -1 0 22262 0 -1 5577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_6
timestamp 1669390400
transform -1 0 22262 0 -1 1977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_64x8m81  018SRAM_cell1_cutPC_64x8m81_7
timestamp 1669390400
transform -1 0 22262 0 -1 3777
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_0
timestamp 1669390400
transform -1 0 16862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_1
timestamp 1669390400
transform -1 0 17462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_2
timestamp 1669390400
transform -1 0 18662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_3
timestamp 1669390400
transform -1 0 18062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_4
timestamp 1669390400
transform -1 0 19262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_5
timestamp 1669390400
transform -1 0 19862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_6
timestamp 1669390400
transform -1 0 20462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_7
timestamp 1669390400
transform -1 0 21062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_8
timestamp 1669390400
transform -1 0 15662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_9
timestamp 1669390400
transform -1 0 15062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_10
timestamp 1669390400
transform -1 0 14462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_11
timestamp 1669390400
transform -1 0 13862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_12
timestamp 1669390400
transform -1 0 12662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_13
timestamp 1669390400
transform -1 0 13262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_14
timestamp 1669390400
transform -1 0 12062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_15
timestamp 1669390400
transform -1 0 11462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_16
timestamp 1669390400
transform -1 0 6662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_17
timestamp 1669390400
transform -1 0 7862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_18
timestamp 1669390400
transform -1 0 7262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_19
timestamp 1669390400
transform -1 0 8462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_20
timestamp 1669390400
transform -1 0 9062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_21
timestamp 1669390400
transform -1 0 9662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_22
timestamp 1669390400
transform -1 0 10262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_23
timestamp 1669390400
transform -1 0 4862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_24
timestamp 1669390400
transform -1 0 4262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_25
timestamp 1669390400
transform -1 0 3662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_26
timestamp 1669390400
transform -1 0 3062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_27
timestamp 1669390400
transform -1 0 1862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_28
timestamp 1669390400
transform -1 0 2462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_29
timestamp 1669390400
transform -1 0 1262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_30
timestamp 1669390400
transform -1 0 662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_64x8m81  018SRAM_cell1_dummy_64x8m81_31
timestamp 1669390400
transform -1 0 6062 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_0
timestamp 1669390400
transform -1 0 16262 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_1
timestamp 1669390400
transform -1 0 10862 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_2
timestamp 1669390400
transform -1 0 5462 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_3
timestamp 1669390400
transform -1 0 62 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_4
timestamp 1669390400
transform -1 0 62 0 -1 9177
box -68 -68 668 968
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_5
timestamp 1669390400
transform 1 0 21062 0 1 177
box -68 -68 668 968
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_0
timestamp 1669390400
transform 1 0 22477 0 -1 417
box 0 0 1 1
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_1
timestamp 1669390400
transform 1 0 22477 0 -1 7377
box 0 0 1 1
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_2
timestamp 1669390400
transform 1 0 22477 0 -1 5577
box 0 0 1 1
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_3
timestamp 1669390400
transform 1 0 22477 0 -1 1977
box 0 0 1 1
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_4
timestamp 1669390400
transform 1 0 22477 0 -1 3777
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1669390400
transform 1 0 22476 0 1 9036
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1669390400
transform 1 0 22475 0 -1 3779
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1669390400
transform 1 0 22475 0 -1 1975
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_2
timestamp 1669390400
transform 1 0 22475 0 -1 5575
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_3
timestamp 1669390400
transform 1 0 22475 0 -1 7379
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_0
timestamp 1669390400
transform 1 0 22475 0 1 379
box 0 0 1 1
use M2_M14310589983233_64x8m81  M2_M14310589983233_64x8m81_0
timestamp 1669390400
transform 1 0 22476 0 1 8975
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_0
timestamp 1669390400
transform 1 0 22475 0 1 181
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_1
timestamp 1669390400
transform 1 0 22476 0 1 9178
box 0 0 1 1
use new_dummyrow_unit_01_64x8m81  new_dummyrow_unit_01_64x8m81_0
timestamp 1669390400
transform 1 0 0 0 -1 9354
box -6 109 10930 1145
use new_dummyrow_unit_64x8m81  new_dummyrow_unit_64x8m81_0
timestamp 1669390400
transform 1 0 10800 0 -1 9354
box -6 109 10930 1145
<< labels >>
rlabel metal3 s 22196 1995 22196 1995 4 VSS
rlabel metal3 s 22196 1070 22196 1070 4 VDD
<< properties >>
string GDS_END 1246418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1241284
<< end >>
