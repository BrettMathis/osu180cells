* NGSPICE file created from gf180mcu_fd_ip_sram__sram512x8m8wm1.ext - technology: gf180mcuC

.subckt x018SRAM_cell1_dummy_512x8m81 a_n36_52# m2_90_n50# a_246_342# m2_390_n50#
+ a_246_712# m3_n36_330# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_cutPC_512x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt array16_512_dummy_01_512x8m81 018SRAM_cell1_cutPC_512x8m81_43/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_10/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_49/a_246_342# 018SRAM_cell1_cutPC_512x8m81_2/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_55/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_44/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_59/a_246_342# 018SRAM_cell1_cutPC_512x8m81_3/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_28/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_56/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_4/a_246_712# 018SRAM_cell1_cutPC_512x8m81_48/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_4/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_57/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_37/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_24/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_57/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_58/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_1/a_246_342# 018SRAM_cell1_cutPC_512x8m81_1/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_5/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_20/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_53/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_59/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_6/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_40/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_41/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_10/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_8/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_7/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_38/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_53/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_45/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_42/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_20/a_246_342# 018SRAM_cell1_cutPC_512x8m81_36/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_34/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_8/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_42/a_246_712# 018SRAM_cell1_cutPC_512x8m81_9/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_2/a_246_342# 018SRAM_cell1_cutPC_512x8m81_9/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_43/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_30/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_2/a_246_712# 018SRAM_cell1_cutPC_512x8m81_32/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_30/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_5/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_63/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_40/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_19/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_44/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_40/a_246_712# 018SRAM_cell1_cutPC_512x8m81_11/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_50/a_246_342# 018SRAM_cell1_cutPC_512x8m81_45/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_1/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_48/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_15/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_7/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_47/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_52/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_60/a_246_342# 018SRAM_cell1_cutPC_512x8m81_21/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_46/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_35/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_44/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_11/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_41/a_246_712# 018SRAM_cell1_cutPC_512x8m81_31/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_3/a_246_342# 018SRAM_cell1_cutPC_512x8m81_47/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_61/a_246_712# 018SRAM_cell1_cutPC_512x8m81_3/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_9/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_48/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_29/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_40/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_41/a_246_342# 018SRAM_cell1_cutPC_512x8m81_49/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_12/a_246_342# 018SRAM_cell1_cutPC_512x8m81_51/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_25/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_58/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_30/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_51/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_31/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_61/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_22/a_246_342# 018SRAM_cell1_cutPC_512x8m81_21/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_34/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_54/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_32/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_4/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_32/a_246_342# 018SRAM_cell1_cutPC_512x8m81_50/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_39/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_33/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_42/a_246_342# 018SRAM_cell1_cutPC_512x8m81_35/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_34/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_52/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_13/a_246_342# 018SRAM_cell1_cutPC_512x8m81_43/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_50/a_246_712# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_62/a_246_342# 018SRAM_cell1_cutPC_512x8m81_35/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_23/a_246_342# 018SRAM_cell1_cutPC_512x8m81_33/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_62/a_246_712# 018SRAM_cell1_cutPC_512x8m81_6/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_31/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_39/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_5/a_246_342# 018SRAM_cell1_cutPC_512x8m81_33/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_36/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_5/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_0/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_16/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_49/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_60/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_2/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_43/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_37/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_53/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_14/a_246_342# 018SRAM_cell1_cutPC_512x8m81_38/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_45/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_12/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_4/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_49/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_39/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_63/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_24/a_246_342# 018SRAM_cell1_cutPC_512x8m81_20/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_38/a_246_712# 018SRAM_cell1_cutPC_512x8m81_41/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_21/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_6/a_246_342# 018SRAM_cell1_cutPC_512x8m81_34/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_6/a_246_712# 018SRAM_cell1_cutPC_512x8m81_26/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_59/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_44/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_22/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_44/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_23/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_22/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_54/a_246_342# 018SRAM_cell1_cutPC_512x8m81_15/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_55/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_53/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_48/a_246_712# 018SRAM_cell1_cutPC_512x8m81_24/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_25/a_246_342# 018SRAM_cell1_cutPC_512x8m81_51/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_37/a_246_712# 018SRAM_cell1_cutPC_512x8m81_7/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_25/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_35/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_2/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_32/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_7/a_246_712# 018SRAM_cell1_cutPC_512x8m81_36/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_26/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_45/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_32/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_7/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_27/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_55/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_16/a_246_342# 018SRAM_cell1_cutPC_512x8m81_8/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_45/a_246_712# 018SRAM_cell1_cutPC_512x8m81_60/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_28/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_26/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_41/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_17/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_61/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_3/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_36/a_246_712# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_29/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_8/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_36/a_246_342# 018SRAM_cell1_cutPC_512x8m81_10/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_61/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_61/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_3/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_46/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_13/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_46/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_62/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_11/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_12/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_56/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_17/a_246_342# 018SRAM_cell1_cutPC_512x8m81_42/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_63/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_51/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_47/a_246_712# 018SRAM_cell1_cutPC_512x8m81_13/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_27/a_246_342# 018SRAM_cell1_cutPC_512x8m81_40/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_35/a_246_712# 018SRAM_cell1_cutPC_512x8m81_27/a_n36_52#
+ VSS 018SRAM_cell1_cutPC_512x8m81_14/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_37/a_246_342# 018SRAM_cell1_cutPC_512x8m81_9/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_23/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_56/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_15/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_47/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_42/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_52/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_16/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_52/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_57/a_246_342# 018SRAM_cell1_cutPC_512x8m81_18/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_50/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_62/w_n68_622#
+ 018SRAM_cell1_cutPC_512x8m81_17/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_28/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_39/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_34/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_37/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_18/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_50/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_38/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_5/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_33/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_8/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_19/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_51/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_48/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_58/a_246_342# 018SRAM_cell1_cutPC_512x8m81_18/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_4/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_62/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_52/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_19/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_49/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_43/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_29/a_246_342# 018SRAM_cell1_cutPC_512x8m81_53/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_38/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_0/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_47/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_cutPC_512x8m81_14/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_33/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_0/a_246_342# 018SRAM_cell1_cutPC_512x8m81_39/a_246_342#
+ 018SRAM_cell1_cutPC_512x8m81_1/m3_n36_330# VSUBS 018SRAM_cell1_cutPC_512x8m81_54/m3_n36_330#
+ 018SRAM_cell1_cutPC_512x8m81_6/w_n68_622# 018SRAM_cell1_cutPC_512x8m81_0/a_246_712#
X018SRAM_cell1_cutPC_512x8m81_3 018SRAM_cell1_cutPC_512x8m81_3/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_3/a_246_342# 018SRAM_cell1_cutPC_512x8m81_3/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_3/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_3/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_4 018SRAM_cell1_cutPC_512x8m81_4/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_4/a_246_342# 018SRAM_cell1_cutPC_512x8m81_4/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_4/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_4/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_5 018SRAM_cell1_cutPC_512x8m81_5/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_5/a_246_342# 018SRAM_cell1_cutPC_512x8m81_5/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_5/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_5/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_6 018SRAM_cell1_cutPC_512x8m81_6/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_6/a_246_342# 018SRAM_cell1_cutPC_512x8m81_6/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_6/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_6/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_7 018SRAM_cell1_cutPC_512x8m81_7/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_7/a_246_342# 018SRAM_cell1_cutPC_512x8m81_7/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_7/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_7/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_9 018SRAM_cell1_cutPC_512x8m81_9/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_9/a_246_342# 018SRAM_cell1_cutPC_512x8m81_9/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_9/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_9/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_8 018SRAM_cell1_cutPC_512x8m81_8/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_8/a_246_342# 018SRAM_cell1_cutPC_512x8m81_8/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_8/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_8/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_60 018SRAM_cell1_cutPC_512x8m81_60/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_60/a_246_342# 018SRAM_cell1_cutPC_512x8m81_3/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_60/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_3/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_50 018SRAM_cell1_cutPC_512x8m81_50/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_50/a_246_342# 018SRAM_cell1_cutPC_512x8m81_50/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_50/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_50/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_61 018SRAM_cell1_cutPC_512x8m81_61/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_61/a_246_342# 018SRAM_cell1_cutPC_512x8m81_61/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_61/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_61/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_40 018SRAM_cell1_cutPC_512x8m81_40/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_40/a_246_342# 018SRAM_cell1_cutPC_512x8m81_40/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_40/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_40/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_51 018SRAM_cell1_cutPC_512x8m81_51/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_51/a_246_342# 018SRAM_cell1_cutPC_512x8m81_51/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_51/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_51/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_62 018SRAM_cell1_cutPC_512x8m81_62/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_62/a_246_342# 018SRAM_cell1_cutPC_512x8m81_62/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_62/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_62/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_30 018SRAM_cell1_cutPC_512x8m81_30/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_30/a_246_342# 018SRAM_cell1_cutPC_512x8m81_32/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_30/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_32/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_41 018SRAM_cell1_cutPC_512x8m81_41/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_41/a_246_342# 018SRAM_cell1_cutPC_512x8m81_41/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_41/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_41/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_52 018SRAM_cell1_cutPC_512x8m81_52/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_52/a_246_342# 018SRAM_cell1_cutPC_512x8m81_52/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_52/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_52/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_63 018SRAM_cell1_cutPC_512x8m81_63/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_63/a_246_342# 018SRAM_cell1_cutPC_512x8m81_2/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_63/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_2/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_42 018SRAM_cell1_cutPC_512x8m81_42/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_42/a_246_342# 018SRAM_cell1_cutPC_512x8m81_42/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_42/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_42/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_20 018SRAM_cell1_cutPC_512x8m81_20/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_20/a_246_342# 018SRAM_cell1_cutPC_512x8m81_42/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_20/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_42/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_53 018SRAM_cell1_cutPC_512x8m81_53/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_53/a_246_342# 018SRAM_cell1_cutPC_512x8m81_53/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_53/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_53/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_31 018SRAM_cell1_cutPC_512x8m81_31/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_31/a_246_342# 018SRAM_cell1_cutPC_512x8m81_61/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_31/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_61/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_32 018SRAM_cell1_cutPC_512x8m81_32/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_32/a_246_342# 018SRAM_cell1_cutPC_512x8m81_32/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_32/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_32/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_21 018SRAM_cell1_cutPC_512x8m81_21/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_21/a_246_342# 018SRAM_cell1_cutPC_512x8m81_41/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_21/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_41/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_43 018SRAM_cell1_cutPC_512x8m81_43/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_43/a_246_342# 018SRAM_cell1_cutPC_512x8m81_43/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_43/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_43/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_10 018SRAM_cell1_cutPC_512x8m81_10/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_10/a_246_342# 018SRAM_cell1_cutPC_512x8m81_53/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_10/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_53/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_54 018SRAM_cell1_cutPC_512x8m81_54/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_54/a_246_342# 018SRAM_cell1_cutPC_512x8m81_9/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_54/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_9/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_33 018SRAM_cell1_cutPC_512x8m81_33/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_33/a_246_342# 018SRAM_cell1_cutPC_512x8m81_33/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_33/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_33/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_22 018SRAM_cell1_cutPC_512x8m81_22/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_22/a_246_342# 018SRAM_cell1_cutPC_512x8m81_40/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_22/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_40/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_44 018SRAM_cell1_cutPC_512x8m81_44/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_44/a_246_342# 018SRAM_cell1_cutPC_512x8m81_44/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_44/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_44/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_11 018SRAM_cell1_cutPC_512x8m81_11/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_11/a_246_342# 018SRAM_cell1_cutPC_512x8m81_52/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_11/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_52/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_55 018SRAM_cell1_cutPC_512x8m81_55/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_55/a_246_342# 018SRAM_cell1_cutPC_512x8m81_8/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_55/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_8/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_34 018SRAM_cell1_cutPC_512x8m81_34/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_34/a_246_342# 018SRAM_cell1_cutPC_512x8m81_34/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_34/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_34/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_23 018SRAM_cell1_cutPC_512x8m81_23/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_23/a_246_342# 018SRAM_cell1_cutPC_512x8m81_39/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_23/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_39/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_45 018SRAM_cell1_cutPC_512x8m81_45/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_45/a_246_342# 018SRAM_cell1_cutPC_512x8m81_45/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_45/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_45/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_12 018SRAM_cell1_cutPC_512x8m81_12/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_12/a_246_342# 018SRAM_cell1_cutPC_512x8m81_51/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_12/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_51/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_56 018SRAM_cell1_cutPC_512x8m81_56/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_56/a_246_342# 018SRAM_cell1_cutPC_512x8m81_7/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_56/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_7/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_35 018SRAM_cell1_cutPC_512x8m81_35/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_35/a_246_342# 018SRAM_cell1_cutPC_512x8m81_35/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_35/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_35/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_36 018SRAM_cell1_cutPC_512x8m81_36/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_36/a_246_342# 018SRAM_cell1_cutPC_512x8m81_36/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_36/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_36/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_25 018SRAM_cell1_cutPC_512x8m81_25/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_25/a_246_342# 018SRAM_cell1_cutPC_512x8m81_37/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_25/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_37/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_24 018SRAM_cell1_cutPC_512x8m81_24/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_24/a_246_342# 018SRAM_cell1_cutPC_512x8m81_38/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_24/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_38/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_47 018SRAM_cell1_cutPC_512x8m81_47/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_47/a_246_342# 018SRAM_cell1_cutPC_512x8m81_47/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_47/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_47/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_46 018SRAM_cell1_cutPC_512x8m81_46/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_46/a_246_342# 018SRAM_cell1_cutPC_512x8m81_0/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_46/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_14 018SRAM_cell1_cutPC_512x8m81_14/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_14/a_246_342# 018SRAM_cell1_cutPC_512x8m81_49/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_14/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_49/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_13 018SRAM_cell1_cutPC_512x8m81_13/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_13/a_246_342# 018SRAM_cell1_cutPC_512x8m81_50/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_13/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_50/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_57 018SRAM_cell1_cutPC_512x8m81_57/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_57/a_246_342# 018SRAM_cell1_cutPC_512x8m81_6/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_57/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_6/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_58 018SRAM_cell1_cutPC_512x8m81_58/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_58/a_246_342# 018SRAM_cell1_cutPC_512x8m81_5/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_58/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_5/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_26 018SRAM_cell1_cutPC_512x8m81_26/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_26/a_246_342# 018SRAM_cell1_cutPC_512x8m81_36/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_26/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_36/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_37 018SRAM_cell1_cutPC_512x8m81_37/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_37/a_246_342# 018SRAM_cell1_cutPC_512x8m81_37/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_37/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_37/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_48 018SRAM_cell1_cutPC_512x8m81_48/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_48/a_246_342# 018SRAM_cell1_cutPC_512x8m81_48/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_48/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_48/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_15 018SRAM_cell1_cutPC_512x8m81_15/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_15/a_246_342# 018SRAM_cell1_cutPC_512x8m81_48/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_15/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_48/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_59 018SRAM_cell1_cutPC_512x8m81_59/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_59/a_246_342# 018SRAM_cell1_cutPC_512x8m81_4/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_59/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_4/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_27 018SRAM_cell1_cutPC_512x8m81_27/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_27/a_246_342# 018SRAM_cell1_cutPC_512x8m81_35/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_27/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_35/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_38 018SRAM_cell1_cutPC_512x8m81_38/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_38/a_246_342# 018SRAM_cell1_cutPC_512x8m81_38/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_38/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_38/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_16 018SRAM_cell1_cutPC_512x8m81_16/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_16/a_246_342# 018SRAM_cell1_cutPC_512x8m81_45/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_16/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_45/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_49 018SRAM_cell1_cutPC_512x8m81_49/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_49/a_246_342# 018SRAM_cell1_cutPC_512x8m81_49/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_49/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_49/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_28 018SRAM_cell1_cutPC_512x8m81_28/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_28/a_246_342# 018SRAM_cell1_cutPC_512x8m81_34/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_28/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_34/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_39 018SRAM_cell1_cutPC_512x8m81_39/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_39/a_246_342# 018SRAM_cell1_cutPC_512x8m81_39/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_39/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_39/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_17 018SRAM_cell1_cutPC_512x8m81_17/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_17/a_246_342# 018SRAM_cell1_cutPC_512x8m81_47/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_17/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_47/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_29 018SRAM_cell1_cutPC_512x8m81_29/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_29/a_246_342# 018SRAM_cell1_cutPC_512x8m81_33/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_29/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_33/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_18 018SRAM_cell1_cutPC_512x8m81_18/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_18/a_246_342# 018SRAM_cell1_cutPC_512x8m81_44/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_18/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_44/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_19 018SRAM_cell1_cutPC_512x8m81_19/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_19/a_246_342# 018SRAM_cell1_cutPC_512x8m81_43/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_19/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_43/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_0 018SRAM_cell1_cutPC_512x8m81_0/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_0/a_246_342# 018SRAM_cell1_cutPC_512x8m81_0/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_0/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_1 018SRAM_cell1_cutPC_512x8m81_1/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_1/a_246_342# 018SRAM_cell1_cutPC_512x8m81_1/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_1/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
X018SRAM_cell1_cutPC_512x8m81_2 018SRAM_cell1_cutPC_512x8m81_2/a_n36_52# 018SRAM_cell1_cutPC_512x8m81_9/a_444_n42#
+ 018SRAM_cell1_cutPC_512x8m81_2/a_246_342# 018SRAM_cell1_cutPC_512x8m81_2/a_246_712#
+ 018SRAM_cell1_cutPC_512x8m81_2/m3_n36_330# 018SRAM_cell1_cutPC_512x8m81_9/a_36_n42#
+ 018SRAM_cell1_cutPC_512x8m81_2/w_n68_622# VSUBS x018SRAM_cell1_cutPC_512x8m81
.ends

.subckt new_dummyrowunit01_512x8m81 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50# VSUBS
X018SRAM_cell1_dummy_512x8m81_13 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_14 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_15 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_0 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_1 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_2 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_3 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_4 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_5 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_6 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_7 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_8 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_9 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_10 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_11 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_12 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
.ends

.subckt new_dummyrow_unit_512x8m81 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ 018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ VSUBS
X018SRAM_cell1_dummy_512x8m81_13 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_14 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_15 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_0 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_1 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_2 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_3 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_4 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_5 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_6 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_7 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_8 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_9 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_10 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_11 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_12 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
.ends

.subckt x018SRAM_cell1_512x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt ldummy_512x4_512x8m81 array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_20/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_1/m3_n36_330#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_17/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/a_246_342# 018SRAM_cell1_dummy_512x8m81_21/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_16/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_18/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_59/a_246_342# 018SRAM_cell1_dummy_512x8m81_22/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/a_246_712# 018SRAM_cell1_dummy_512x8m81_26/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_19/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/w_n68_622# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_23/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/w_n68_622#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/m3_n36_330#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_24/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/VSS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/m3_n36_330#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_25/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_17/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_26/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_54/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/a_246_712# 018SRAM_cell1_dummy_512x8m81_27/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_1/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_20/a_246_342# 018SRAM_cell1_dummy_512x8m81_27/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_55/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/m3_n36_330#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_30/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_28/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_56/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/a_246_342# 018SRAM_cell1_dummy_512x8m81_29/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_57/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_18/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_11/a_246_342# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_58/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/a_246_712# 018SRAM_cell1_dummy_512x8m81_28/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_60/a_246_342# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_21/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_59/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/w_n68_622#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_31/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/a_246_712# 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_19/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/a_246_342# 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_12/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_29/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_16/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_22/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/a_246_712#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_17/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/m3_n36_330#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_18/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_46/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_19/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_13/a_246_342# 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/a_246_712#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_62/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_23/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/a_246_712# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_30/m3_n36_330#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_31/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_14/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/a_246_712# 018SRAM_cell1_dummy_512x8m81_20/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_63/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_24/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/a_246_712# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/a_246_712# 018SRAM_cell1_dummy_512x8m81_30/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_54/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_15/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/a_246_712# 018SRAM_cell1_dummy_512x8m81_21/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_25/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/a_246_712#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_31/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/w_n68_622#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_20/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_16/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_55/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_21/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/a_246_712#
+ 018SRAM_cell1_dummy_512x8m81_22/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_22/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_26/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/a_246_712#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/a_246_712#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_23/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/w_n68_622#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_24/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_46/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_56/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_25/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_17/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_23/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/a_246_712#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_26/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_27/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/w_n68_622# 018SRAM_cell1_dummy_512x8m81_30/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/w_n68_622# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/a_246_712# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_27/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_31/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_28/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/a_246_342#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_60/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_29/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_18/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_57/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_10/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/w_n68_622#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/w_n68_622# 018SRAM_cell1_dummy_512x8m81_24/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_11/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_28/a_246_342# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_62/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/w_n68_622# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_12/m3_n36_330# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_390_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_63/m3_n36_330# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_13/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/a_246_342#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_58/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_14/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_19/a_246_342# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_25/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/a_246_712#
+ 018SRAM_cell1_512x8m81_1/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_15/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_29/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/w_n68_622# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/m3_n36_330#
+ VSUBS new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_90_n50# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_16/m3_n36_330#
X018SRAM_cell1_dummy_512x8m81_13 VSUBS 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_24 VSUBS 018SRAM_cell1_dummy_512x8m81_24/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_24/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_14 VSUBS 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_25 VSUBS 018SRAM_cell1_dummy_512x8m81_25/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_25/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_15 VSUBS 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_26 VSUBS 018SRAM_cell1_dummy_512x8m81_26/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_26/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_16 VSUBS 018SRAM_cell1_dummy_512x8m81_16/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_16/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_27 VSUBS 018SRAM_cell1_dummy_512x8m81_27/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_27/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
Xarray16_512_dummy_01_512x8m81_0 VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_55/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_59/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/m3_n36_330# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_56/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_57/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/w_n68_622#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_58/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_1/a_246_342# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/m3_n36_330# VSUBS
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_59/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_10/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/m3_n36_330#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_20/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/w_n68_622#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/a_246_712# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_30/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/a_246_712#
+ VSUBS VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/a_246_342#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_11/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/m3_n36_330#
+ VSUBS VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_60/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_21/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_46/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/w_n68_622#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_31/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/m3_n36_330# VSUBS
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_12/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/a_246_342# VSUBS
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_30/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_31/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_22/a_246_342#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/w_n68_622#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/a_246_342#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/a_246_342# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_13/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/a_246_712# 018SRAM_cell1_512x8m81_1/a_444_n42#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_62/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_23/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/w_n68_622#
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/w_n68_622# VSUBS
+ VSUBS VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_14/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/m3_n36_330#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_4/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_63/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_24/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_20/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/a_246_712#
+ VSUBS 018SRAM_cell1_512x8m81_1/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_21/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/a_246_712# VSUBS
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_22/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_44/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_23/m3_n36_330# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_54/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_15/a_246_342#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_24/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_25/a_246_342# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_25/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_2/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_32/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_7/a_246_712# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_26/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/a_246_342#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_27/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_55/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_16/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_45/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_60/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_28/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_26/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_41/w_n68_622#
+ VSUBS VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/a_246_712#
+ 018SRAM_cell1_512x8m81_1/a_36_n42# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_29/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_8/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_36/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_10/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_61/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_3/w_n68_622#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_46/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_62/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_11/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_12/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_56/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_17/a_246_342# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_63/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_13/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_27/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_40/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_35/a_246_712# VSUBS
+ array16_512_dummy_01_512x8m81_0/VSS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_14/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_37/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_9/a_246_712# VSUBS
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_15/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_47/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_42/w_n68_622#
+ VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_16/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_57/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_18/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/w_n68_622#
+ 018SRAM_cell1_512x8m81_0/w_n68_622# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_17/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_28/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_34/a_246_712# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_18/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_50/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_5/w_n68_622#
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_19/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_51/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_48/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_58/a_246_342# VSUBS
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_52/m3_n36_330#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_19/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_49/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_43/a_246_712# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_29/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_53/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_38/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/m3_n36_330# VSUBS
+ VSUBS VSUBS array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_33/a_246_712#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/a_246_342# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_39/a_246_342#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_1/m3_n36_330# VSUBS
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_54/m3_n36_330# array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_6/w_n68_622#
+ array16_512_dummy_01_512x8m81_0/018SRAM_cell1_cutPC_512x8m81_0/a_246_712# array16_512_dummy_01_512x8m81
X018SRAM_cell1_dummy_512x8m81_17 VSUBS 018SRAM_cell1_dummy_512x8m81_17/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_17/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_28 VSUBS 018SRAM_cell1_dummy_512x8m81_28/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_28/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_18 VSUBS 018SRAM_cell1_dummy_512x8m81_18/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_18/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_29 VSUBS 018SRAM_cell1_dummy_512x8m81_29/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_29/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_19 VSUBS 018SRAM_cell1_dummy_512x8m81_19/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_19/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
Xnew_dummyrowunit01_512x8m81_0 new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_390_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_90_n50#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_90_n50# VSUBS 018SRAM_cell1_512x8m81_1/w_n68_622#
+ new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_90_n50# new_dummyrowunit01_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ VSUBS new_dummyrowunit01_512x8m81
X018SRAM_cell1_dummy_512x8m81_0 VSUBS 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_1 VSUBS 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_2 VSUBS 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
Xnew_dummyrow_unit_512x8m81_0 new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_4/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_5/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_6/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_390_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_10/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_11/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_12/m2_90_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_2/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ VSUBS new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_15/m2_90_n50# new_dummyrow_unit_512x8m81_0/018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ VSUBS new_dummyrow_unit_512x8m81
X018SRAM_cell1_dummy_512x8m81_3 VSUBS 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_4 VSUBS 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_5 VSUBS 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_6 VSUBS 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_30 VSUBS 018SRAM_cell1_dummy_512x8m81_30/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_30/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_7 VSUBS 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_31 VSUBS 018SRAM_cell1_dummy_512x8m81_31/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_31/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_20 VSUBS 018SRAM_cell1_dummy_512x8m81_20/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_20/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_8 VSUBS 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_10 VSUBS 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_21 VSUBS 018SRAM_cell1_dummy_512x8m81_21/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_21/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_9 VSUBS 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_11 VSUBS 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_22 VSUBS 018SRAM_cell1_dummy_512x8m81_22/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_22/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_512x8m81_0 VSUBS 018SRAM_cell1_512x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS
+ x018SRAM_cell1_512x8m81
X018SRAM_cell1_dummy_512x8m81_12 VSUBS 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_23 VSUBS 018SRAM_cell1_dummy_512x8m81_23/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_512x8m81_23/m2_390_n50# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_512x8m81_1 VSUBS 018SRAM_cell1_512x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_512x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_512x8m81
.ends

.subckt dcap_103_novia_512x8m81 w_n203_44# a_n67_185# a_73_103#
X0 a_n67_185# a_73_103# a_n67_185# w_n203_44# pmos_3p3 w=2.275u l=2.365u
.ends

.subckt pmos_5p04310591302020_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46897196_512x8m81 pmos_5p04310591302020_512x8m81_0/D a_193_n74#
+ w_n286_n142# pmos_5p04310591302020_512x8m81_0/S a_n31_n74#
Xpmos_5p04310591302020_512x8m81_0 w_n286_n142# pmos_5p04310591302020_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302020_512x8m81_0/S a_193_n74# pmos_5p04310591302020_512x8m81
.ends

.subckt nmos_5p04310591302015_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46553132_512x8m81 nmos_5p04310591302015_512x8m81_0/D nmos_5p04310591302015_512x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310591302015_512x8m81_0 nmos_5p04310591302015_512x8m81_0/D a_n31_n74# nmos_5p04310591302015_512x8m81_0/S
+ VSUBS nmos_5p04310591302015_512x8m81
.ends

.subckt nmos_5p04310591302017_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_1p2$$46550060_512x8m81 a_1537_n74# a_1313_n74# nmos_5p04310591302017_512x8m81_0/S
+ a_193_n74# a_1089_n74# nmos_5p04310591302017_512x8m81_0/D a_865_n74# a_n31_n74#
+ a_641_n74# a_417_n74# VSUBS
Xnmos_5p04310591302017_512x8m81_0 nmos_5p04310591302017_512x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310591302017_512x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310591302017_512x8m81
.ends

.subckt pmos_5p04310591302014_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46285868_512x8m81 pmos_5p04310591302014_512x8m81_0/S w_n286_n142#
+ a_n31_n73# pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n286_n142# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt pmos_5p04310591302013_512x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46286892_512x8m81 pmos_5p04310591302013_512x8m81_0/D a_193_n73#
+ a_n31_n73# a_417_n73# w_n286_n142# pmos_5p04310591302013_512x8m81_0/S
Xpmos_5p04310591302013_512x8m81_0 w_n286_n142# pmos_5p04310591302013_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302013_512x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310591302013_512x8m81
.ends

.subckt nmos_5p04310591302010_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$46551084_512x8m81 nmos_5p04310591302010_512x8m81_0/D a_n31_n73#
+ nmos_5p04310591302010_512x8m81_0/S VSUBS
Xnmos_5p04310591302010_512x8m81_0 nmos_5p04310591302010_512x8m81_0/D a_n31_n73# nmos_5p04310591302010_512x8m81_0/S
+ VSUBS nmos_5p04310591302010_512x8m81
.ends

.subckt pmos_5p04310591302019_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46898220_512x8m81 pmos_5p04310591302019_512x8m81_0/S w_n286_n142#
+ a_n31_n74# pmos_5p04310591302019_512x8m81_0/D
Xpmos_5p04310591302019_512x8m81_0 w_n286_n142# pmos_5p04310591302019_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302019_512x8m81_0/S pmos_5p04310591302019_512x8m81
.ends

.subckt pmos_5p04310591302021_512x8m81 w_n208_n120# D a_0_n44# a_672_n44# S a_448_n44#
+ a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46896172_512x8m81 a_668_n74# a_193_n74# pmos_5p04310591302021_512x8m81_0/S
+ w_n286_n142# a_n31_n74# pmos_5p04310591302021_512x8m81_0/D a_417_n74#
Xpmos_5p04310591302021_512x8m81_0 w_n286_n142# pmos_5p04310591302021_512x8m81_0/D
+ a_n31_n74# a_668_n74# pmos_5p04310591302021_512x8m81_0/S a_417_n74# a_193_n74# pmos_5p04310591302021_512x8m81
.ends

.subckt nmos_5p04310591302012_512x8m81 D a_0_n44# a_672_n44# S a_448_n44# a_224_n44#
+ VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45107244_512x8m81 a_193_n73# nmos_5p04310591302012_512x8m81_0/S
+ a_n31_n73# a_641_n73# a_417_n73# nmos_5p04310591302012_512x8m81_0/D VSUBS
Xnmos_5p04310591302012_512x8m81_0 nmos_5p04310591302012_512x8m81_0/D a_n31_n73# a_641_n73#
+ nmos_5p04310591302012_512x8m81_0/S a_417_n73# a_193_n73# VSUBS nmos_5p04310591302012_512x8m81
.ends

.subckt pmos_5p04310591302018_512x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46549036_512x8m81 pmos_5p04310591302018_512x8m81_0/D a_193_n74#
+ w_n286_n142# pmos_5p04310591302018_512x8m81_0/S a_1089_n74# a_865_n74# a_n31_n74#
+ a_641_n74# a_417_n74#
Xpmos_5p04310591302018_512x8m81_0 w_n286_n142# pmos_5p04310591302018_512x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310591302018_512x8m81_0/S a_417_n74# a_193_n74#
+ a_1089_n74# pmos_5p04310591302018_512x8m81
.ends

.subckt nmos_5p04310591302016_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46552108_512x8m81 a_1089_n74# a_865_n74# a_641_n74# a_n31_n74# a_417_n74#
+ a_193_n74# a_1537_n74# nmos_5p04310591302016_512x8m81_0/S a_1313_n74# nmos_5p04310591302016_512x8m81_0/D
+ VSUBS
Xnmos_5p04310591302016_512x8m81_0 nmos_5p04310591302016_512x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310591302016_512x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310591302016_512x8m81
.ends

.subckt sa_512x8m81 qp wep se pcb vss d
Xpmos_1p2$$46897196_512x8m81_1 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ se d d se pmos_1p2$$46897196_512x8m81
Xpmos_1p2$$46897196_512x8m81_2 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ se d d se pmos_1p2$$46897196_512x8m81
Xpmos_1p2$$46897196_512x8m81_3 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ se d d se pmos_1p2$$46897196_512x8m81
Xnmos_1p2$$46553132_512x8m81_0 vss pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ vss vss nmos_1p2$$46553132_512x8m81
Xnmos_1p2$$46550060_512x8m81_0 se se vss se se nmos_1p2$$46552108_512x8m81_0/nmos_5p04310591302016_512x8m81_0/D
+ se se se se vss nmos_1p2$$46550060_512x8m81
Xnmos_1p2$$46553132_512x8m81_1 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_512x8m81
Xpmos_1p2$$46285868_512x8m81_0 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ d pcb pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46285868_512x8m81
Xpmos_1p2$$46286892_512x8m81_0 d pcb pcb pcb d d pmos_1p2$$46286892_512x8m81
Xnmos_1p2$$46551084_512x8m81_0 vss pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ qp vss nmos_1p2$$46551084_512x8m81
Xpmos_1p2$$46898220_512x8m81_0 d d d pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81
Xpmos_1p2$$46898220_512x8m81_1 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ d d d pmos_1p2$$46898220_512x8m81
Xpmos_1p2$$46896172_512x8m81_0 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ d pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S d pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46896172_512x8m81
Xnmos_1p2$$45107244_512x8m81_0 qp qp pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ qp qp vss vss nmos_1p2$$45107244_512x8m81
Xpmos_1p2$$46549036_512x8m81_0 qp pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ d d pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S qp qp pmos_1p2$$46549036_512x8m81
Xpmos_1p2$$46897196_512x8m81_0 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ se d d se pmos_1p2$$46897196_512x8m81
Xnmos_1p2$$46552108_512x8m81_0 pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S pmos_1p2$$46898220_512x8m81_1/pmos_5p04310591302019_512x8m81_0/S
+ nmos_1p2$$46552108_512x8m81_0/nmos_5p04310591302016_512x8m81_0/D vss nmos_1p2$$46552108_512x8m81
.ends

.subckt nmos_5p0431059130205_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_1p2$$46883884_512x8m81 nmos_5p0431059130205_512x8m81_0/S a_n31_n73# nmos_5p0431059130205_512x8m81_0/D
+ VSUBS
Xnmos_5p0431059130205_512x8m81_0 nmos_5p0431059130205_512x8m81_0/D a_n31_n73# nmos_5p0431059130205_512x8m81_0/S
+ VSUBS nmos_5p0431059130205_512x8m81
.ends

.subckt pmos_5p0431059130206_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_1p2$$46885932_512x8m81 pmos_5p0431059130206_512x8m81_0/D a_193_n73# a_n31_n74#
+ w_n286_n141# pmos_5p0431059130206_512x8m81_0/S
Xpmos_5p0431059130206_512x8m81_0 w_n286_n141# pmos_5p0431059130206_512x8m81_0/D a_n31_n74#
+ pmos_5p0431059130206_512x8m81_0/S a_193_n73# pmos_5p0431059130206_512x8m81
.ends

.subckt pmos_5p0431059130209_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_5p0431059130208_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$46563372_512x8m81 nmos_5p0431059130208_512x8m81_0/D a_n31_n74# nmos_5p0431059130208_512x8m81_0/S
+ VSUBS
Xnmos_5p0431059130208_512x8m81_0 nmos_5p0431059130208_512x8m81_0/D a_n31_n74# nmos_5p0431059130208_512x8m81_0/S
+ VSUBS nmos_5p0431059130208_512x8m81
.ends

.subckt pmos_5p0431059130203_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_1p2$$46273580_512x8m81 pmos_5p0431059130203_512x8m81_0/S a_193_n74# a_n31_n74#
+ pmos_5p0431059130203_512x8m81_0/D w_n286_n142#
Xpmos_5p0431059130203_512x8m81_0 w_n286_n142# pmos_5p0431059130203_512x8m81_0/D a_n31_n74#
+ pmos_5p0431059130203_512x8m81_0/S a_193_n74# pmos_5p0431059130203_512x8m81
.ends

.subckt nmos_5p04310591302011_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_5p0431059130204_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.61u l=0.6u
.ends

.subckt pmos_1p2$$46887980_512x8m81 pmos_5p0431059130204_512x8m81_0/S a_n31_n74# pmos_5p0431059130204_512x8m81_0/D
+ w_n286_n142#
Xpmos_5p0431059130204_512x8m81_0 w_n286_n142# pmos_5p0431059130204_512x8m81_0/D a_n31_n74#
+ pmos_5p0431059130204_512x8m81_0/S pmos_5p0431059130204_512x8m81
.ends

.subckt nmos_5p0431059130207_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=13.61u l=0.6u
.ends

.subckt nmos_1p2$$46884908_512x8m81 nmos_5p0431059130207_512x8m81_0/S nmos_5p0431059130207_512x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p0431059130207_512x8m81_0 nmos_5p0431059130207_512x8m81_0/D a_n31_n74# nmos_5p0431059130207_512x8m81_0/S
+ VSUBS nmos_5p0431059130207_512x8m81
.ends

.subckt pmos_5p0431059130201_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.81u l=0.6u
.ends

.subckt pmos_1p2$$46889004_512x8m81 pmos_5p0431059130201_512x8m81_0/D w_n286_n142#
+ a_n31_n74# pmos_5p0431059130201_512x8m81_0/S
Xpmos_5p0431059130201_512x8m81_0 w_n286_n142# pmos_5p0431059130201_512x8m81_0/D a_n31_n74#
+ pmos_5p0431059130201_512x8m81_0/S pmos_5p0431059130201_512x8m81
.ends

.subckt din_512x8m81 d db datain wep men m1_164_8068# pmos_5p0431059130201_512x8m81_0/D
+ vdd vss
Xnmos_1p2$$46883884_512x8m81_0 db wep pmos_5p0431059130209_512x8m81_0/S vss nmos_1p2$$46883884_512x8m81
Xnmos_1p2$$46883884_512x8m81_1 pmos_5p0431059130209_512x8m81_0/S pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ vss vss nmos_1p2$$46883884_512x8m81
Xnmos_1p2$$46883884_512x8m81_2 d wep pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ vss nmos_1p2$$46883884_512x8m81
Xpmos_1p2$$46885932_512x8m81_0 nmos_5p04310591302011_512x8m81_1/D pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ men vdd pmos_5p0431059130206_512x8m81_0/S pmos_1p2$$46885932_512x8m81
Xpmos_5p0431059130209_512x8m81_0 vdd vdd pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ pmos_5p0431059130209_512x8m81_0/S pmos_5p0431059130209_512x8m81
Xnmos_1p2$$46563372_512x8m81_0 pmos_5p0431059130206_512x8m81_0/S pmos_5p0431059130201_512x8m81_0/S
+ vss vss nmos_1p2$$46563372_512x8m81
Xnmos_1p2$$46563372_512x8m81_1 pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ men vss vss nmos_1p2$$46563372_512x8m81
Xpmos_1p2$$46273580_512x8m81_0 vdd men men pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ vdd pmos_1p2$$46273580_512x8m81
Xpmos_1p2$$46273580_512x8m81_1 vdd pmos_5p0431059130201_512x8m81_0/S pmos_5p0431059130201_512x8m81_0/S
+ pmos_5p0431059130206_512x8m81_0/S vdd pmos_1p2$$46273580_512x8m81
Xpmos_5p0431059130206_512x8m81_0 vdd vdd datain pmos_5p0431059130206_512x8m81_0/S
+ pmos_5p0431059130206_512x8m81_0/S pmos_5p0431059130206_512x8m81
Xnmos_5p04310591302011_512x8m81_0 vss datain pmos_5p0431059130206_512x8m81_0/S pmos_5p0431059130206_512x8m81_0/S
+ vss nmos_5p04310591302011_512x8m81
Xnmos_5p04310591302011_512x8m81_1 nmos_5p04310591302011_512x8m81_1/D pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ pmos_5p0431059130206_512x8m81_0/S men vss nmos_5p04310591302011_512x8m81
Xpmos_1p2$$46887980_512x8m81_0 vdd pmos_5p0431059130201_512x8m81_0/S pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ vdd pmos_1p2$$46887980_512x8m81
Xnmos_5p04310591302010_512x8m81_0 vss nmos_5p04310591302011_512x8m81_1/D pmos_5p0431059130201_512x8m81_0/S
+ vss nmos_5p04310591302010_512x8m81
Xnmos_1p2$$46884908_512x8m81_0 vss pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ pmos_5p0431059130201_512x8m81_0/S vss nmos_1p2$$46884908_512x8m81
Xpmos_1p2$$46889004_512x8m81_0 pmos_1p2$$46889004_512x8m81_0/pmos_5p0431059130201_512x8m81_0/D
+ vdd a_500_6666# d pmos_1p2$$46889004_512x8m81
Xpmos_1p2$$46889004_512x8m81_1 pmos_5p0431059130209_512x8m81_0/S vdd a_500_6666# db
+ pmos_1p2$$46889004_512x8m81
Xpmos_5p0431059130201_512x8m81_0 vdd pmos_5p0431059130201_512x8m81_0/D nmos_5p04310591302011_512x8m81_1/D
+ pmos_5p0431059130201_512x8m81_0/S pmos_5p0431059130201_512x8m81
X0 vdd wep a_500_6666# vdd pmos_3p3 w=1.485u l=0.6u
X1 a_500_6666# wep vss vss nmos_3p3 w=1.14u l=0.6u
X2 a_500_6666# wep vdd vdd pmos_3p3 w=1.485u l=0.6u
.ends

.subckt nmos_5p04310591302034_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.44u l=0.6u
.ends

.subckt pmos_5p04310591302024_512x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46282796_512x8m81 a_193_n74# pmos_5p04310591302024_512x8m81_0/D
+ a_865_n74# a_n31_n74# a_641_n74# a_417_n74# w_n286_n142# pmos_5p04310591302024_512x8m81_0/S
Xpmos_5p04310591302024_512x8m81_0 w_n286_n142# pmos_5p04310591302024_512x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310591302024_512x8m81_0/S a_417_n74# a_193_n74#
+ pmos_5p04310591302024_512x8m81
.ends

.subckt nmos_5p04310591302033_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310591302023_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.6u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310591302036_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_1p2$$45101100_512x8m81 nmos_5p04310591302036_512x8m81_0/S a_193_n74#
+ a_865_n74# a_n31_n74# a_641_n74# a_417_n74# nmos_5p04310591302036_512x8m81_0/D VSUBS
Xnmos_5p04310591302036_512x8m81_0 nmos_5p04310591302036_512x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310591302036_512x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310591302036_512x8m81
.ends

.subckt nmos_5p04310591302032_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_5p04310591302026_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45102124_512x8m81 a_1313_n74# nmos_5p04310591302026_512x8m81_0/D
+ a_193_n74# a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# nmos_5p04310591302026_512x8m81_0/S
+ a_417_n74# VSUBS
Xnmos_5p04310591302026_512x8m81_0 nmos_5p04310591302026_512x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310591302026_512x8m81_0/S a_417_n74# a_193_n74# a_1313_n74#
+ a_1089_n74# VSUBS nmos_5p04310591302026_512x8m81
.ends

.subckt nmos_5p04310591302037_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
.ends

.subckt nmos_1p2$$45103148_512x8m81 nmos_5p04310591302037_512x8m81_0/S a_865_n73#
+ nmos_5p04310591302037_512x8m81_0/D a_193_n74# a_1089_n74# a_n31_n74# a_641_n74#
+ a_417_n74# VSUBS
Xnmos_5p04310591302037_512x8m81_0 nmos_5p04310591302037_512x8m81_0/D a_n31_n74# a_865_n73#
+ a_641_n74# nmos_5p04310591302037_512x8m81_0/S a_417_n74# a_193_n74# a_1089_n74#
+ VSUBS nmos_5p04310591302037_512x8m81
.ends

.subckt pmos_5p04310591302022_512x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
.ends

.subckt pmos_1p2$$46283820_512x8m81 a_641_n74# a_1985_n74# a_1761_n74# a_417_n74#
+ a_1537_n74# a_1313_n74# pmos_5p04310591302022_512x8m81_0/S w_n286_n142# a_193_n74#
+ pmos_5p04310591302022_512x8m81_0/D a_1089_n74# a_865_n74# a_n31_n74#
Xpmos_5p04310591302022_512x8m81_0 w_n286_n142# pmos_5p04310591302022_512x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310591302022_512x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310591302022_512x8m81
.ends

.subckt nmos_5p04310591302029_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.61u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.61u l=0.6u
.ends

.subckt nmos_1p2$$45100076_512x8m81 nmos_5p04310591302029_512x8m81_0/S a_193_n74#
+ nmos_5p04310591302029_512x8m81_0/D a_n31_n74# VSUBS
Xnmos_5p04310591302029_512x8m81_0 nmos_5p04310591302029_512x8m81_0/D a_n31_n74# nmos_5p04310591302029_512x8m81_0/S
+ a_193_n74# VSUBS nmos_5p04310591302029_512x8m81
.ends

.subckt nmos_5p04310591302028_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310591302038_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310591302031_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.41u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.41u l=0.6u
.ends

.subckt pmos_1p2$$46287916_512x8m81 pmos_5p04310591302031_512x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310591302031_512x8m81_0/S
Xpmos_5p04310591302031_512x8m81_0 w_n286_n142# pmos_5p04310591302031_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302031_512x8m81_0/S a_193_n74# pmos_5p04310591302031_512x8m81
.ends

.subckt pmos_5p04310591302027_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310591302035_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$46284844_512x8m81 pmos_5p04310591302035_512x8m81_0/S a_n31_n74#
+ pmos_5p04310591302035_512x8m81_0/D w_n286_n142# a_193_n74#
Xpmos_5p04310591302035_512x8m81_0 w_n286_n142# pmos_5p04310591302035_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302035_512x8m81_0/S a_193_n74# pmos_5p04310591302035_512x8m81
.ends

.subckt pmos_5p04310591302025_512x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$46281772_512x8m81 pmos_5p04310591302025_512x8m81_0/D a_n31_n73#
+ w_n286_n142# pmos_5p04310591302025_512x8m81_0/S a_193_n73# a_417_n73#
Xpmos_5p04310591302025_512x8m81_0 w_n286_n142# pmos_5p04310591302025_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302025_512x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310591302025_512x8m81
.ends

.subckt pmos_5p04310591302030_512x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
.ends

.subckt pmos_1p2$$45095980_512x8m81 pmos_5p04310591302030_512x8m81_0/S a_193_n74#
+ pmos_5p04310591302030_512x8m81_0/D a_1089_n74# a_865_n74# a_n31_n74# a_641_n74#
+ a_1985_n74# a_1761_n74# a_417_n74# w_n286_n142# a_1537_n74# a_1313_n74#
Xpmos_5p04310591302030_512x8m81_0 w_n286_n142# pmos_5p04310591302030_512x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310591302030_512x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310591302030_512x8m81
.ends

.subckt sacntl_2_512x8m81 men pcb a_4718_983# nmos_5p04310591302023_512x8m81_1/D pmos_5p04310591302027_512x8m81_2/S
+ a_4560_1922# a_2796_670# se pmos_5p04310591302027_512x8m81_1/S pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ vdd vss
Xnmos_5p04310591302034_512x8m81_0 nmos_5p04310591302034_512x8m81_0/D pmos_5p04310591302027_512x8m81_1/S
+ vss vss nmos_5p04310591302034_512x8m81
Xpmos_1p2$$46285868_512x8m81_0 nmos_5p04310591302028_512x8m81_1/S vdd pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ vdd pmos_1p2$$46285868_512x8m81
Xpmos_1p2$$46282796_512x8m81_0 men pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ men men men men vdd vdd pmos_1p2$$46282796_512x8m81
Xnmos_5p04310591302033_512x8m81_0 vss pmos_5p04310591302027_512x8m81_0/S pmos_5p04310591302038_512x8m81_0/S
+ vss nmos_5p04310591302033_512x8m81
Xnmos_5p04310591302023_512x8m81_0 vss a_2796_670# pmos_5p04310591302027_512x8m81_0/S
+ pmos_5p04310591302027_512x8m81_0/S vss nmos_5p04310591302023_512x8m81
Xnmos_5p04310591302023_512x8m81_1 nmos_5p04310591302023_512x8m81_1/D pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ pmos_5p04310591302027_512x8m81_1/S vss vss nmos_5p04310591302023_512x8m81
Xnmos_5p04310591302023_512x8m81_2 vss pmos_5p04310591302027_512x8m81_1/S pmos_5p04310591302027_512x8m81_2/S
+ pmos_5p04310591302027_512x8m81_2/S vss nmos_5p04310591302023_512x8m81
Xnmos_1p2$$45101100_512x8m81_0 vss men men men men men pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ vss nmos_1p2$$45101100_512x8m81
Xnmos_5p04310591302032_512x8m81_0 nmos_5p04310591302032_512x8m81_0/D nmos_5p04310591302034_512x8m81_0/D
+ vss nmos_5p04310591302034_512x8m81_0/D vss nmos_5p04310591302032_512x8m81
Xpmos_1p2$$46286892_512x8m81_0 nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302032_512x8m81_0/D
+ nmos_5p04310591302032_512x8m81_0/D nmos_5p04310591302032_512x8m81_0/D vdd vdd pmos_1p2$$46286892_512x8m81
Xnmos_5p04310591302012_512x8m81_0 se nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S
+ vss nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S vss nmos_5p04310591302012_512x8m81
Xnmos_1p2$$45102124_512x8m81_0 pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pcb pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S vss pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ vss nmos_1p2$$45102124_512x8m81
Xnmos_1p2$$45103148_512x8m81_0 vss nmos_5p04310591302034_512x8m81_0/D pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S
+ nmos_5p04310591302034_512x8m81_0/D pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D nmos_5p04310591302028_512x8m81_1/S
+ nmos_5p04310591302028_512x8m81_1/S vss nmos_1p2$$45103148_512x8m81
Xpmos_1p2$$46283820_512x8m81_0 pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S vdd vdd pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pcb pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46283820_512x8m81
Xnmos_1p2$$45100076_512x8m81_0 vss pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S
+ vss nmos_1p2$$45100076_512x8m81
Xnmos_5p04310591302028_512x8m81_0 nmos_5p04310591302028_512x8m81_1/D nmos_5p04310591302032_512x8m81_0/D
+ nmos_5p04310591302032_512x8m81_0/D nmos_5p04310591302032_512x8m81_0/D vss nmos_5p04310591302032_512x8m81_0/D
+ nmos_5p04310591302032_512x8m81_0/D vss nmos_5p04310591302028_512x8m81
Xnmos_5p04310591302028_512x8m81_1 nmos_5p04310591302028_512x8m81_1/D pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ nmos_5p04310591302028_512x8m81_1/S pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D vss nmos_5p04310591302028_512x8m81
Xpmos_5p04310591302038_512x8m81_0 vdd vdd pmos_5p04310591302027_512x8m81_0/S pmos_5p04310591302038_512x8m81_0/S
+ pmos_5p04310591302038_512x8m81
Xpmos_1p2$$46287916_512x8m81_0 nmos_5p04310591302032_512x8m81_0/D nmos_5p04310591302034_512x8m81_0/D
+ vdd nmos_5p04310591302034_512x8m81_0/D vdd pmos_1p2$$46287916_512x8m81
Xpmos_5p04310591302027_512x8m81_0 vdd vdd a_2796_670# pmos_5p04310591302027_512x8m81_0/S
+ pmos_5p04310591302027_512x8m81_0/S pmos_5p04310591302027_512x8m81
Xpmos_1p2$$46284844_512x8m81_0 vdd pmos_5p04310591302027_512x8m81_1/S nmos_5p04310591302034_512x8m81_0/D
+ vdd pmos_5p04310591302027_512x8m81_1/S pmos_1p2$$46284844_512x8m81
Xpmos_1p2$$46281772_512x8m81_0 vdd pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S
+ vdd pmos_1p2$$46281772_512x8m81_0/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S
+ pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S pmos_1p2$$46281772_512x8m81
Xpmos_5p04310591302027_512x8m81_1 vdd vdd pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ pmos_5p04310591302027_512x8m81_1/S vss pmos_5p04310591302027_512x8m81
Xpmos_5p04310591302027_512x8m81_2 vdd vdd pmos_5p04310591302027_512x8m81_1/S pmos_5p04310591302027_512x8m81_2/S
+ pmos_5p04310591302027_512x8m81_2/S pmos_5p04310591302027_512x8m81
Xpmos_1p2$$46281772_512x8m81_1 vdd pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ vdd pmos_1p2$$46281772_512x8m81_1/pmos_5p04310591302025_512x8m81_0/S nmos_5p04310591302034_512x8m81_0/D
+ nmos_5p04310591302028_512x8m81_1/S pmos_1p2$$46281772_512x8m81
Xpmos_1p2$$45095980_512x8m81_0 vdd nmos_5p04310591302028_512x8m81_1/S se nmos_5p04310591302028_512x8m81_1/S
+ nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S
+ nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S
+ vdd nmos_5p04310591302028_512x8m81_1/S nmos_5p04310591302028_512x8m81_1/S pmos_1p2$$45095980_512x8m81
.ends

.subckt pmos_1p2$$202586156_512x8m81 pmos_5p04310591302014_512x8m81_0/S w_n286_n141#
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n286_n141# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt pmos_1p2$$202583084_512x8m81 pmos_5p04310591302035_512x8m81_0/S pmos_5p04310591302035_512x8m81_0/D
+ a_193_n74# w_n286_n142# a_n31_n74#
Xpmos_5p04310591302035_512x8m81_0 w_n286_n142# pmos_5p04310591302035_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302035_512x8m81_0/S a_193_n74# pmos_5p04310591302035_512x8m81
.ends

.subckt nmos_5p04310591302042_512x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.8u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
.ends

.subckt pmos_5p04310591302043_512x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_1p2$$202587180_512x8m81 pmos_5p04310591302014_512x8m81_0/S w_n286_n141#
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n286_n141# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt nmos_5p04310591302040_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.37u l=0.6u
.ends

.subckt pmos_5p04310591302041_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$202594348_512x8m81 a_n31_n73# nmos_5p04310591302040_512x8m81_0/D
+ nmos_5p04310591302040_512x8m81_0/S VSUBS
Xnmos_5p04310591302040_512x8m81_0 nmos_5p04310591302040_512x8m81_0/D a_n31_n73# nmos_5p04310591302040_512x8m81_0/S
+ VSUBS nmos_5p04310591302040_512x8m81
.ends

.subckt nmos_1p2$$202598444_512x8m81 nmos_5p04310591302010_512x8m81_0/D nmos_5p04310591302010_512x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310591302010_512x8m81_0 nmos_5p04310591302010_512x8m81_0/D a_n31_n74# nmos_5p04310591302010_512x8m81_0/S
+ VSUBS nmos_5p04310591302010_512x8m81
.ends

.subckt nmos_1p2$$202595372_512x8m81 nmos_5p0431059130208_512x8m81_0/D a_n31_n73#
+ nmos_5p0431059130208_512x8m81_0/S VSUBS
Xnmos_5p0431059130208_512x8m81_0 nmos_5p0431059130208_512x8m81_0/D a_n31_n73# nmos_5p0431059130208_512x8m81_0/S
+ VSUBS nmos_5p0431059130208_512x8m81
.ends

.subckt nmos_5p04310591302039_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$202596396_512x8m81 nmos_5p0431059130208_512x8m81_0/D a_n31_n73#
+ nmos_5p0431059130208_512x8m81_0/S VSUBS
Xnmos_5p0431059130208_512x8m81_0 nmos_5p0431059130208_512x8m81_0/D a_n31_n73# nmos_5p0431059130208_512x8m81_0/S
+ VSUBS nmos_5p0431059130208_512x8m81
.ends

.subckt pmos_1p2$$202584108_512x8m81 a_n31_n74# pmos_5p04310591302014_512x8m81_0/S
+ w_n286_n141# pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n286_n141# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt pmos_1p2$$202585132_512x8m81 w_n256_n141# pmos_5p04310591302014_512x8m81_0/S
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n256_n141# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt wen_wm1_512x8m81 GWEN wep wen men vss vdd
Xpmos_5p04310591302035_512x8m81_0 vdd pmos_5p04310591302035_512x8m81_0/D pmos_5p04310591302020_512x8m81_0/S
+ vdd pmos_5p04310591302020_512x8m81_0/S pmos_5p04310591302035_512x8m81
Xpmos_1p2$$202586156_512x8m81_0 pmos_5p04310591302041_512x8m81_0/D vdd nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S
+ vdd pmos_1p2$$202586156_512x8m81
Xpmos_1p2$$202583084_512x8m81_0 vdd pmos_1p2$$202583084_512x8m81_0/pmos_5p04310591302035_512x8m81_0/D
+ nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D vdd nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ pmos_1p2$$202583084_512x8m81
Xpmos_5p04310591302014_512x8m81_0 vdd pmos_5p04310591302014_512x8m81_2/S wen vdd pmos_5p04310591302014_512x8m81
Xnmos_5p04310591302042_512x8m81_0 wep pmos_5p04310591302035_512x8m81_0/D vss pmos_5p04310591302035_512x8m81_0/D
+ pmos_5p04310591302035_512x8m81_0/D vss nmos_5p04310591302042_512x8m81
Xpmos_5p04310591302043_512x8m81_0 vdd wep pmos_5p04310591302035_512x8m81_0/D vdd pmos_5p04310591302035_512x8m81_0/D
+ pmos_5p04310591302035_512x8m81_0/D pmos_5p04310591302043_512x8m81
Xpmos_5p04310591302014_512x8m81_1 vdd nmos_5p0431059130208_512x8m81_1/D nmos_5p0431059130208_512x8m81_2/D
+ vdd pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302014_512x8m81_2 vdd nmos_5p0431059130208_512x8m81_2/D GWEN pmos_5p04310591302014_512x8m81_2/S
+ pmos_5p04310591302014_512x8m81
Xpmos_1p2$$202587180_512x8m81_0 nmos_5p0431059130208_512x8m81_1/D vdd nmos_5p0431059130208_512x8m81_3/D
+ pmos_5p04310591302041_512x8m81_0/S pmos_1p2$$202587180_512x8m81
Xpmos_5p04310591302014_512x8m81_3 vdd pmos_5p04310591302014_512x8m81_5/S men vdd pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302014_512x8m81_4 vdd nmos_5p0431059130208_512x8m81_3/D pmos_5p04310591302014_512x8m81_5/D
+ vdd pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302014_512x8m81_5 vdd pmos_5p04310591302014_512x8m81_5/D vss pmos_5p04310591302014_512x8m81_5/S
+ pmos_5p04310591302014_512x8m81
Xnmos_5p04310591302040_512x8m81_0 pmos_5p04310591302035_512x8m81_0/D pmos_5p04310591302020_512x8m81_0/S
+ vss vss nmos_5p04310591302040_512x8m81
Xpmos_5p04310591302041_512x8m81_0 vdd pmos_5p04310591302041_512x8m81_0/D pmos_5p04310591302014_512x8m81_5/D
+ pmos_5p04310591302041_512x8m81_0/S pmos_5p04310591302041_512x8m81
Xnmos_5p04310591302040_512x8m81_1 pmos_5p04310591302014_512x8m81_5/D men vss vss nmos_5p04310591302040_512x8m81
Xnmos_5p0431059130208_512x8m81_0 vss GWEN nmos_5p0431059130208_512x8m81_2/D vss nmos_5p0431059130208_512x8m81
Xnmos_1p2$$202594348_512x8m81_0 nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ vss pmos_1p2$$202583084_512x8m81_0/pmos_5p04310591302035_512x8m81_0/D vss nmos_1p2$$202594348_512x8m81
Xnmos_5p04310591302040_512x8m81_2 vss vss pmos_5p04310591302014_512x8m81_5/D vss nmos_5p04310591302040_512x8m81
Xnmos_5p04310591302010_512x8m81_0 vss nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ pmos_5p04310591302020_512x8m81_0/S vss nmos_5p04310591302010_512x8m81
Xnmos_5p0431059130208_512x8m81_1 nmos_5p0431059130208_512x8m81_1/D nmos_5p0431059130208_512x8m81_2/D
+ vss vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_2 nmos_5p0431059130208_512x8m81_2/D wen vss vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_3 nmos_5p0431059130208_512x8m81_3/D pmos_5p04310591302014_512x8m81_5/D
+ vss vss nmos_5p0431059130208_512x8m81
Xnmos_1p2$$202598444_512x8m81_0 pmos_5p04310591302041_512x8m81_0/S nmos_5p0431059130208_512x8m81_1/D
+ pmos_5p04310591302014_512x8m81_5/D vss nmos_1p2$$202598444_512x8m81
Xpmos_5p04310591302020_512x8m81_0 vdd men nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ pmos_5p04310591302020_512x8m81_0/S nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ pmos_5p04310591302020_512x8m81
Xnmos_1p2$$202595372_512x8m81_0 pmos_5p04310591302041_512x8m81_0/D nmos_5p0431059130208_512x8m81_3/D
+ pmos_5p04310591302041_512x8m81_0/S vss nmos_1p2$$202595372_512x8m81
Xnmos_1p2$$202595372_512x8m81_1 vss pmos_5p04310591302041_512x8m81_0/S nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S
+ vss nmos_1p2$$202595372_512x8m81
Xnmos_5p04310591302039_512x8m81_0 men pmos_1p2$$202583084_512x8m81_0/pmos_5p04310591302035_512x8m81_0/D
+ pmos_5p04310591302020_512x8m81_0/S pmos_1p2$$202583084_512x8m81_0/pmos_5p04310591302035_512x8m81_0/D
+ vss nmos_5p04310591302039_512x8m81
Xnmos_1p2$$202596396_512x8m81_0 nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S vss vss nmos_1p2$$202596396_512x8m81
Xnmos_1p2$$202596396_512x8m81_1 vss nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S
+ pmos_5p04310591302041_512x8m81_0/D vss nmos_1p2$$202596396_512x8m81
Xpmos_1p2$$202584108_512x8m81_0 pmos_5p04310591302041_512x8m81_0/S nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S
+ vdd vdd pmos_1p2$$202584108_512x8m81
Xpmos_1p2$$202585132_512x8m81_0 vdd vdd nmos_1p2$$202595372_512x8m81_1/nmos_5p0431059130208_512x8m81_0/S
+ nmos_1p2$$202596396_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D pmos_1p2$$202585132_512x8m81
.ends

.subckt nmos_5p0431059130202_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.57u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.57u l=0.6u
.ends

.subckt nmos_5p0431059130200_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.81u l=0.6u
.ends

.subckt nmos_1p2$$47119404_512x8m81 nmos_5p0431059130200_512x8m81_0/S a_n31_n74# VSUBS
+ nmos_5p0431059130200_512x8m81_0/D
Xnmos_5p0431059130200_512x8m81_0 nmos_5p0431059130200_512x8m81_0/D a_n31_n74# nmos_5p0431059130200_512x8m81_0/S
+ VSUBS nmos_5p0431059130200_512x8m81
.ends

.subckt ypass_gate_a_512x8m81 vss b bb db ypass d pcb a_222_11191# a_n4_11191# m3_n1_4331#
+ a_447_11191# vdd a_222_10416# m3_n1_1708# a_n4_10416# m3_n1_1160# m3_n1_2030# pmos_5p0431059130201_512x8m81_1/D
+ m3_n1_3366# a_447_10416# m3_n1_2352# m3_n1_3688# m3_n1_4009# m3_n1_2674#
Xnmos_5p0431059130202_512x8m81_0 nmos_5p0431059130202_512x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059130202_512x8m81
Xnmos_1p2$$47119404_512x8m81_0 b ypass vss d nmos_1p2$$47119404_512x8m81
Xnmos_1p2$$47119404_512x8m81_1 bb ypass vss pmos_5p0431059130201_512x8m81_1/D nmos_1p2$$47119404_512x8m81
Xpmos_1p2$$46889004_512x8m81_0 d vdd nmos_5p0431059130202_512x8m81_0/D b pmos_1p2$$46889004_512x8m81
Xpmos_5p0431059130201_512x8m81_0 vdd b pcb bb pmos_5p0431059130201_512x8m81
Xpmos_5p0431059130201_512x8m81_1 vdd pmos_5p0431059130201_512x8m81_1/D nmos_5p0431059130202_512x8m81_0/D
+ bb pmos_5p0431059130201_512x8m81
X0 nmos_5p0431059130202_512x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd ypass nmos_5p0431059130202_512x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X2 a_447_11191# pcb a_222_11191# vdd pmos_3p3 w=3.41u l=0.6u
X3 a_222_11191# pcb a_n4_11191# vdd pmos_3p3 w=3.41u l=0.6u
X4 a_447_10416# pcb a_222_10416# vdd pmos_3p3 w=3.41u l=0.6u
X5 a_222_10416# pcb a_n4_10416# vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt ypass_gate_512x8m81 vss b bb db ypass d pcb m3_n1_4331# vdd m3_n1_1708# m3_n1_1160#
+ m3_n1_2030# m3_n1_3366# m3_n1_2352# m3_n1_3688# m3_n1_4009# m3_n1_2674#
Xnmos_5p0431059130202_512x8m81_0 nmos_5p0431059130202_512x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059130202_512x8m81
Xnmos_1p2$$47119404_512x8m81_0 b ypass vss d nmos_1p2$$47119404_512x8m81
Xnmos_1p2$$47119404_512x8m81_1 bb ypass vss db nmos_1p2$$47119404_512x8m81
Xpmos_1p2$$46889004_512x8m81_0 d vdd nmos_5p0431059130202_512x8m81_0/D b pmos_1p2$$46889004_512x8m81
Xpmos_5p0431059130201_512x8m81_0 vdd b pcb bb pmos_5p0431059130201_512x8m81
Xpmos_5p0431059130201_512x8m81_1 vdd db nmos_5p0431059130202_512x8m81_0/D bb pmos_5p0431059130201_512x8m81
X0 nmos_5p0431059130202_512x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd ypass nmos_5p0431059130202_512x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt mux821_512x8m81 ypass_gate_512x8m81_1/d ypass_gate_512x8m81_0/ypass a_656_7735#
+ ypass_gate_512x8m81_1/ypass ypass_gate_a_512x8m81_0/db ypass_gate_512x8m81_2/ypass
+ ypass_gate_a_512x8m81_0/a_222_11191# ypass_gate_512x8m81_3/d ypass_gate_512x8m81_4/b
+ ypass_gate_512x8m81_3/ypass ypass_gate_512x8m81_4/ypass ypass_gate_512x8m81_5/d
+ ypass_gate_512x8m81_5/ypass ypass_gate_512x8m81_6/ypass ypass_gate_512x8m81_6/m3_n1_2030#
+ ypass_gate_512x8m81_5/db ypass_gate_a_512x8m81_0/ypass ypass_gate_a_512x8m81_0/a_447_11191#
+ ypass_gate_512x8m81_6/m3_n1_3366# ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688#
+ ypass_gate_512x8m81_0/d ypass_gate_512x8m81_6/m3_n1_4009# ypass_gate_512x8m81_6/m3_n1_2674#
+ ypass_gate_512x8m81_2/d ypass_gate_a_512x8m81_0/a_222_10416# ypass_gate_512x8m81_4/d
+ ypass_gate_512x8m81_6/d a_4992_424# ypass_gate_a_512x8m81_0/a_447_10416# ypass_gate_512x8m81_6/m3_n1_4331#
+ ypass_gate_512x8m81_6/pcb ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/db ypass_gate_a_512x8m81_0/d
+ ypass_gate_512x8m81_4/db ypass_gate_512x8m81_6/vss ypass_gate_a_512x8m81_0/b ypass_gate_512x8m81_6/m3_n1_1708#
Xypass_gate_a_512x8m81_0 ypass_gate_512x8m81_6/vss ypass_gate_a_512x8m81_0/b ypass_gate_a_512x8m81_0/bb
+ ypass_gate_a_512x8m81_0/db ypass_gate_a_512x8m81_0/ypass ypass_gate_a_512x8m81_0/d
+ ypass_gate_512x8m81_6/pcb ypass_gate_a_512x8m81_0/a_222_11191# ypass_gate_512x8m81_6/vdd
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_a_512x8m81_0/a_447_11191# ypass_gate_512x8m81_6/vdd
+ ypass_gate_a_512x8m81_0/a_222_10416# ypass_gate_512x8m81_6/m3_n1_1708# ypass_gate_512x8m81_6/vdd
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_1/db
+ ypass_gate_512x8m81_6/m3_n1_3366# ypass_gate_a_512x8m81_0/a_447_10416# ypass_gate_512x8m81_6/m3_n1_2352#
+ ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009# ypass_gate_512x8m81_6/m3_n1_2674#
+ ypass_gate_a_512x8m81
Xypass_gate_512x8m81_0 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_0/b ypass_gate_512x8m81_0/bb
+ ypass_gate_512x8m81_4/db ypass_gate_512x8m81_0/ypass ypass_gate_512x8m81_0/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_1 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_1/b ypass_gate_512x8m81_1/bb
+ ypass_gate_512x8m81_1/db ypass_gate_512x8m81_1/ypass ypass_gate_512x8m81_1/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_2 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_2/b ypass_gate_512x8m81_2/bb
+ ypass_gate_512x8m81_5/db ypass_gate_512x8m81_2/ypass ypass_gate_512x8m81_2/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_3 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_3/b ypass_gate_512x8m81_3/bb
+ ypass_gate_512x8m81_6/db ypass_gate_512x8m81_3/ypass ypass_gate_512x8m81_3/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_4 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_4/b ypass_gate_512x8m81_4/bb
+ ypass_gate_512x8m81_4/db ypass_gate_512x8m81_4/ypass ypass_gate_512x8m81_4/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_5 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_5/b ypass_gate_512x8m81_5/bb
+ ypass_gate_512x8m81_5/db ypass_gate_512x8m81_5/ypass ypass_gate_512x8m81_5/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
Xypass_gate_512x8m81_6 ypass_gate_512x8m81_6/vss ypass_gate_512x8m81_6/b ypass_gate_512x8m81_6/bb
+ ypass_gate_512x8m81_6/db ypass_gate_512x8m81_6/ypass ypass_gate_512x8m81_6/d ypass_gate_512x8m81_6/pcb
+ ypass_gate_512x8m81_6/m3_n1_4331# ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_1708#
+ ypass_gate_512x8m81_6/vdd ypass_gate_512x8m81_6/m3_n1_2030# ypass_gate_512x8m81_6/m3_n1_3366#
+ ypass_gate_512x8m81_6/m3_n1_2352# ypass_gate_512x8m81_6/m3_n1_3688# ypass_gate_512x8m81_6/m3_n1_4009#
+ ypass_gate_512x8m81_6/m3_n1_2674# ypass_gate_512x8m81
.ends

.subckt nmos_5p04310591302045_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310591302044_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310591302052_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.6u l=0.6u
.ends

.subckt nmos_5p04310591302050_512x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310591302051_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.67u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$171625516_512x8m81 pmos_5p0431059130203_512x8m81_0/S a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p0431059130203_512x8m81_0/D pmos_5p0431059130203_512x8m81_0/w_n208_n120#
Xpmos_5p0431059130203_512x8m81_0 pmos_5p0431059130203_512x8m81_0/w_n208_n120# pmos_5p0431059130203_512x8m81_0/D
+ a_n31_n74# pmos_5p0431059130203_512x8m81_0/S a_193_n74# pmos_5p0431059130203_512x8m81
.ends

.subckt pmos_5p04310591302049_512x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
.ends

.subckt pmos_5p04310591302048_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.5u l=0.6u
.ends

.subckt nmos_5p04310591302046_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
.ends

.subckt pmos_5p04310591302047_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4u l=0.6u
.ends

.subckt outbuf_oe_512x8m81 qp qn se q GWE a_4913_n316# vss vdd
Xnmos_5p04310591302045_512x8m81_1 pmos_5p04310591302051_512x8m81_0/D qn nmos_5p04310591302045_512x8m81_1/S
+ qn vss nmos_5p04310591302045_512x8m81
Xnmos_5p04310591302044_512x8m81_0 vss pmos_5p04310591302047_512x8m81_0/S pmos_5p04310591302048_512x8m81_0/S
+ vss nmos_5p04310591302044_512x8m81
Xnmos_5p04310591302033_512x8m81_0 pmos_5p04310591302038_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ vss vss nmos_5p04310591302033_512x8m81
Xnmos_5p04310591302052_512x8m81_0 vss GWE pmos_5p04310591302047_512x8m81_0/S vss nmos_5p04310591302052_512x8m81
Xpmos_5p04310591302014_512x8m81_0 vdd nmos_5p0431059130208_512x8m81_0/D se vdd pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302013_512x8m81_0 vdd nmos_5p0431059130208_512x8m81_1/S se pmos_5p04310591302051_512x8m81_0/D
+ se se pmos_5p04310591302013_512x8m81
Xnmos_5p04310591302050_512x8m81_0 nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_0/D
+ pmos_5p04310591302051_512x8m81_0/D nmos_5p0431059130208_512x8m81_0/D nmos_5p0431059130208_512x8m81_0/D
+ vss nmos_5p04310591302050_512x8m81
Xpmos_5p04310591302051_512x8m81_0 vdd pmos_5p04310591302051_512x8m81_0/D qp pmos_5p04310591302051_512x8m81_1/S
+ qp pmos_5p04310591302051_512x8m81
Xpmos_5p04310591302051_512x8m81_1 vdd vdd pmos_5p04310591302048_512x8m81_0/S pmos_5p04310591302051_512x8m81_1/S
+ pmos_5p04310591302048_512x8m81_0/S pmos_5p04310591302051_512x8m81
Xnmos_5p0431059130208_512x8m81_0 nmos_5p0431059130208_512x8m81_0/D se vss vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_1 vss pmos_5p04310591302038_512x8m81_0/D nmos_5p0431059130208_512x8m81_1/S
+ vss nmos_5p0431059130208_512x8m81
Xpmos_1p2$$171625516_512x8m81_0 vdd pmos_5p04310591302038_512x8m81_0/D vdd pmos_5p04310591302038_512x8m81_0/D
+ nmos_5p0431059130208_512x8m81_1/S vdd pmos_1p2$$171625516_512x8m81
Xpmos_5p04310591302049_512x8m81_0 vdd vdd pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ pmos_5p04310591302051_512x8m81_0/D q pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302049_512x8m81
Xpmos_5p04310591302048_512x8m81_0 vdd vdd pmos_5p04310591302047_512x8m81_0/S pmos_5p04310591302048_512x8m81_0/S
+ pmos_5p04310591302048_512x8m81
Xpmos_5p04310591302038_512x8m81_0 vdd pmos_5p04310591302038_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ vdd pmos_5p04310591302038_512x8m81
Xnmos_5p04310591302046_512x8m81_0 vss pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ pmos_5p04310591302051_512x8m81_0/D q pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ pmos_5p04310591302051_512x8m81_0/D vss nmos_5p04310591302046_512x8m81
Xpmos_5p04310591302047_512x8m81_0 vdd vdd GWE pmos_5p04310591302047_512x8m81_0/S pmos_5p04310591302047_512x8m81
Xnmos_5p04310591302045_512x8m81_0 vss pmos_5p04310591302047_512x8m81_0/S nmos_5p04310591302045_512x8m81_1/S
+ pmos_5p04310591302047_512x8m81_0/S vss nmos_5p04310591302045_512x8m81
.ends

.subckt saout_m2_512x8m81 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWEN GWE bb[6] b[0] datain q pcb WEN a_5189_27176# a_5414_27176# a_5189_27951#
+ a_5414_27951# bb[5] b[4] bb[7] bb[2] sacntl_2_512x8m81_0/a_4718_983# mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass
+ b[7] mux821_512x8m81_0/a_4992_424# b[5] men b[6] mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass
+ wen_wm1_512x8m81_0/GWEN b[1] bb[4] b[2] wen_wm1_512x8m81_0/vdd mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b
+ bb[3] mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass b[3] vdd mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass
+ bb[1] sa_512x8m81_0/wep mux821_512x8m81_0/a_656_7735# mux821_512x8m81_0/ypass_gate_512x8m81_6/vdd
+ mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass sacntl_2_512x8m81_0/a_4560_1922# vss
+ sa_512x8m81_0/pcb mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass outbuf_oe_512x8m81_0/a_4913_n316#
+ sacntl_2_512x8m81_0/vdd bb[0] mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass
Xsa_512x8m81_0 sa_512x8m81_0/qp sa_512x8m81_0/wep sa_512x8m81_0/se sa_512x8m81_0/pcb
+ vss vdd sa_512x8m81
Xdin_512x8m81_0 vdd vdd datain sa_512x8m81_0/wep men sa_512x8m81_0/pcb vdd vdd vss
+ din_512x8m81
Xsacntl_2_512x8m81_0 men sa_512x8m81_0/pcb sacntl_2_512x8m81_0/a_4718_983# vss sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_2/S
+ sacntl_2_512x8m81_0/a_4560_1922# sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_2/S
+ sa_512x8m81_0/se sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_1/S sacntl_2_512x8m81_0/pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ sacntl_2_512x8m81_0/vdd vss sacntl_2_512x8m81
Xwen_wm1_512x8m81_0 wen_wm1_512x8m81_0/GWEN sa_512x8m81_0/wep wen_wm1_512x8m81_0/wen
+ men vss wen_wm1_512x8m81_0/vdd wen_wm1_512x8m81
Xmux821_512x8m81_0 vdd mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass mux821_512x8m81_0/a_656_7735#
+ mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass vdd mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass
+ a_5189_27951# vdd mux821_512x8m81_0/ypass_gate_512x8m81_4/b mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass vdd mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass
+ vdd mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass a_5414_27951# mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass
+ vdd mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass
+ vdd a_5189_27176# vdd vdd mux821_512x8m81_0/a_4992_424# a_5414_27176# mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass
+ sa_512x8m81_0/pcb mux821_512x8m81_0/ypass_gate_512x8m81_6/vdd vdd vdd vdd vss mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b
+ mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass mux821_512x8m81
Xoutbuf_oe_512x8m81_0 sa_512x8m81_0/qp sa_512x8m81_0/qp sa_512x8m81_0/se q GWE outbuf_oe_512x8m81_0/a_4913_n316#
+ vss vdd outbuf_oe_512x8m81
.ends

.subckt x018SRAM_cell1_2x_512x8m81 018SRAM_cell1_512x8m81_1/a_246_342# 018SRAM_cell1_512x8m81_1/a_246_712#
+ 018SRAM_cell1_512x8m81_0/m3_n36_330# 018SRAM_cell1_512x8m81_1/m3_n36_330# 018SRAM_cell1_512x8m81_0/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_0/a_n36_52# 018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_512x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_512x8m81_0/a_246_342# 018SRAM_cell1_512x8m81_0/a_246_712#
+ 018SRAM_cell1_512x8m81_1/a_444_n42#
X018SRAM_cell1_512x8m81_1 018SRAM_cell1_512x8m81_1/a_n36_52# 018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_512x8m81_1/a_246_342# 018SRAM_cell1_512x8m81_1/a_246_712# 018SRAM_cell1_512x8m81_1/m3_n36_330#
+ 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_512x8m81
X018SRAM_cell1_512x8m81_0 018SRAM_cell1_512x8m81_0/a_n36_52# 018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_512x8m81_0/a_246_342# 018SRAM_cell1_512x8m81_0/a_246_712# 018SRAM_cell1_512x8m81_0/m3_n36_330#
+ 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_512x8m81
.ends

.subckt Cell_array8x8_512x8m81 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42# VSUBS 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
X018SRAM_cell1_2x_512x8m81_0[0|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[0|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[1|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[2|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[3|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[4|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[5|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[6|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[7|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[8|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[9|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[10|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[11|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[12|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[13|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[14|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[15|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[16|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[17|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[18|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[19|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[20|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[21|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[22|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[23|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[24|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[25|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[26|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[27|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[28|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[29|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[30|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0[31|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_0[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[0|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[1|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[2|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[3|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[4|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[5|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[6|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[7|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[8|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[9|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[10|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[11|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[12|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[13|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[14|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[15|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[16|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[17|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[18|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[19|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[20|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[21|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[22|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[23|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[24|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[25|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[26|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[27|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[28|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[29|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[30|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1[31|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_1[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[0|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[1|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[2|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[3|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[4|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[5|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[6|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[7|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[8|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[9|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[10|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[11|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[12|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[13|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[14|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[15|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[16|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[17|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[18|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[19|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[20|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[21|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[22|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[23|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[24|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[25|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[26|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[27|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[28|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[29|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[30|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3[31|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_3[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|0] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|0]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|1] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|1]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|2] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|2]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|3] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|3]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|4] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|4]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|5] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|5]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|6] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|6]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[0|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[0]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[1|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[1]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[2|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[2]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[3|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[3]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[4|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[4]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[5|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[5]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[6|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[6]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[7|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[7]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[8|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[8]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[9|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[10|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[10]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[11|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[11]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[12|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[12]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[13|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[13]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[14|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[14]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[15|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[15]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[16|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[16]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[17|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[17]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[18|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[18]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[19|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[19]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[20|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[20]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[21|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[21]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[22|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[22]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[23|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[23]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[24|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[24]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[25|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[25]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[26|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[26]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[27|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[27]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[28|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[28]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[29|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[29]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[30|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[30]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2[31|7] VSUBS 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52#
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_0/a_n36_52# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_36_n42#
+ 018SRAM_strap1_2x_512x8m81_3[31]/018SRAM_strap1_512x8m81_1/a_n36_52# VSUBS VSUBS
+ 018SRAM_strap1_2x_512x8m81_3[9]/018SRAM_strap1_512x8m81_1/w_n68_622# 018SRAM_cell1_2x_512x8m81_2[9|7]/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
.ends

.subckt saout_R_m2_512x8m81 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6]
+ ypass[7] ypass[0] GWE GWEN datain b[0] q bb[1] pcb WEN wen_wm1_512x8m81_0/wen mux821_512x8m81_0/ypass_gate_512x8m81_4/b
+ bb[2] b[3] mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass bb[0] bb[5] sacntl_2_512x8m81_0/a_4718_983#
+ men b[7] a_5189_27169# a_5414_27169# a_5189_27944# a_5414_27944# b[2] b[1] wen_wm1_512x8m81_0/GWEN
+ b[6] bb[3] b[5] mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass wen_wm1_512x8m81_0/vdd
+ bb[4] b[4] mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass vdd mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass
+ bb[6] sa_512x8m81_0/wep mux821_512x8m81_0/a_656_7735# mux821_512x8m81_0/ypass_gate_512x8m81_6/vdd
+ mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass
+ sacntl_2_512x8m81_0/a_4560_1922# mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass vss
+ sa_512x8m81_0/pcb mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass outbuf_oe_512x8m81_0/a_4913_n316#
+ sacntl_2_512x8m81_0/vdd bb[7]
Xsa_512x8m81_0 sa_512x8m81_0/qp sa_512x8m81_0/wep sa_512x8m81_0/se sa_512x8m81_0/pcb
+ vss vdd sa_512x8m81
Xdin_512x8m81_0 vdd vdd datain sa_512x8m81_0/wep men sa_512x8m81_0/pcb vdd vdd vss
+ din_512x8m81
Xsacntl_2_512x8m81_0 men sa_512x8m81_0/pcb sacntl_2_512x8m81_0/a_4718_983# vss sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_2/S
+ sacntl_2_512x8m81_0/a_4560_1922# sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_2/S
+ sa_512x8m81_0/se sacntl_2_512x8m81_0/pmos_5p04310591302027_512x8m81_1/S sacntl_2_512x8m81_0/pmos_1p2$$46282796_512x8m81_0/pmos_5p04310591302024_512x8m81_0/D
+ sacntl_2_512x8m81_0/vdd vss sacntl_2_512x8m81
Xwen_wm1_512x8m81_0 wen_wm1_512x8m81_0/GWEN sa_512x8m81_0/wep wen_wm1_512x8m81_0/wen
+ men vss wen_wm1_512x8m81_0/vdd wen_wm1_512x8m81
Xmux821_512x8m81_0 vdd mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass mux821_512x8m81_0/a_656_7735#
+ mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass vdd mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass
+ a_5189_27944# vdd mux821_512x8m81_0/ypass_gate_512x8m81_4/b mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass vdd mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass mux821_512x8m81_0/ypass_gate_512x8m81_6/ypass
+ vdd mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass a_5414_27944# mux821_512x8m81_0/ypass_gate_512x8m81_0/ypass
+ mux821_512x8m81_0/ypass_gate_512x8m81_2/ypass mux821_512x8m81_0/ypass_gate_512x8m81_4/ypass
+ vdd mux821_512x8m81_0/ypass_gate_512x8m81_1/ypass mux821_512x8m81_0/ypass_gate_512x8m81_5/ypass
+ vdd a_5189_27169# vdd vdd mux821_512x8m81_0/a_4992_424# a_5414_27169# mux821_512x8m81_0/ypass_gate_a_512x8m81_0/ypass
+ sa_512x8m81_0/pcb mux821_512x8m81_0/ypass_gate_512x8m81_6/vdd vdd vdd vdd vss mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b
+ mux821_512x8m81_0/ypass_gate_512x8m81_3/ypass mux821_512x8m81
Xoutbuf_oe_512x8m81_0 sa_512x8m81_0/qp sa_512x8m81_0/qp sa_512x8m81_0/se q GWE outbuf_oe_512x8m81_0/a_4913_n316#
+ vss vdd outbuf_oe_512x8m81
.ends

.subckt col_512a_512x8m81 WL[3] ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] GWE WL[2]
+ WL[1] WL[32] WL[31] WL[30] WL[29] WL[24] WL[23] WL[22] WL[21] WL[57] WL[56] WL[20]
+ WL[19] WL[58] WL[59] WL[49] WL[48] WL[12] WL[11] WL[50] WL[51] WL[41] WL[40] WL[10]
+ WL[9] WL[42] WL[43] WL[35] WL[34] WL[8] WL[39] WL[37] WL[7] WL[33] WL[6] WL[38]
+ WL[36] WL[5] WL[47] WL[45] WL[4] WL[46] WL[44] WL[18] WL[55] WL[53] WL[17] WL[54]
+ WL[52] WL[16] WL[63] WL[61] WL[15] WL[14] WL[62] WL[60] WL[13] WL[28] WL[27] WL[26]
+ WL[0] ypass[2] WL[25] b[10] b[13] b[16] b[22] b[31] din[1] din[3] din[2] din[0]
+ q[0] q[1] q[2] q[3] b[17] bb[10] bb[11] bb[12] bb[14] bb[15] bb[16] bb[22] bb[23]
+ bb[25] bb[31] b[27] b[0] b[18] pcb[0] pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1]
+ WEN[0] a_15501_29383# m3_n1102_31970# saout_R_m2_512x8m81_0/wen_wm1_512x8m81_0/wen
+ a_15261_28608# saout_m2_512x8m81_1/GWEN a_4701_29383# b[8] b[2] a_4461_28608# bb[3]
+ a_15501_28608# saout_R_m2_512x8m81_0/mux821_512x8m81_0/ypass_gate_512x8m81_4/b b[4]
+ ypass[6] ypass[7] bb[5] bb[26] a_15261_29383# b[11] bb[0] bb[19] b[1] saout_m2_512x8m81_1/sa_512x8m81_0/pcb
+ bb[24] bb[9] bb[21] b[24] bb[2] b[6] a_4701_28608# b[3] saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ bb[18] b[30] b[20] bb[8] bb[4] b[19] bb[29] saout_m2_512x8m81_0/WEN b[23] b[14]
+ b[5] bb[20] b[29] b[28] b[25] saout_m2_512x8m81_0/pcb bb[13] men saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb
+ saout_R_m2_512x8m81_1/sa_512x8m81_0/pcb bb[28] bb[7] bb[17] bb[6] bb[1] b[21] b[26]
+ bb[27] b[12] b[9] a_4461_29383# b[15] bb[30] VDD b[7] VSS
Xsaout_m2_512x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] saout_m2_512x8m81_1/GWEN GWE bb[14] b[8] saout_m2_512x8m81_1/datain saout_m2_512x8m81_1/q
+ saout_m2_512x8m81_1/pcb saout_m2_512x8m81_1/WEN a_15036_28608# a_15261_28608# a_15036_29383#
+ a_15261_29383# bb[13] b[12] bb[15] bb[10] saout_m2_512x8m81_1/sacntl_2_512x8m81_0/a_4718_983#
+ ypass[7] b[15] VSS b[13] men b[14] ypass[0] saout_m2_512x8m81_1/GWEN b[9] bb[12]
+ b[10] VDD saout_m2_512x8m81_1/mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b bb[11]
+ ypass[1] b[11] VDD ypass[4] bb[9] saout_m2_512x8m81_1/sa_512x8m81_0/wep saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ VDD ypass[2] VSS VSS saout_m2_512x8m81_1/sa_512x8m81_0/pcb ypass[3] VSS VDD bb[8]
+ ypass[5] ypass[6] saout_m2_512x8m81
XCell_array8x8_512x8m81_0 bb[26] bb[12] WL[6] bb[16] WL[2] b[17] WL[8] b[4] b[18]
+ bb[18] b[25] b[31] bb[15] b[11] WL[1] WL[12] b[19] b[14] WL[3] b[5] bb[20] WL[14]
+ bb[13] bb[6] b[21] b[12] bb[5] bb[19] bb[24] b[7] bb[30] WL[7] bb[22] bb[10] bb[31]
+ bb[11] WL[18] b[23] b[30] WL[9] b[10] WL[4] bb[29] WL[28] WL[47] bb[9] WL[5] WL[10]
+ WL[58] WL[42] b[6] b[28] WL[11] b[0] WL[16] WL[30] WL[61] WL[49] b[20] b[8] WL[13]
+ b[2] b[29] WL[35] b[9] b[15] bb[27] bb[0] WL[23] WL[37] WL[15] WL[21] WL[60] b[22]
+ b[26] b[16] WL[34] WL[53] WL[46] b[1] WL[32] WL[25] WL[17] WL[33] bb[25] WL[44]
+ WL[36] WL[55] bb[2] b[27] WL[48] WL[27] WL[39] bb[7] bb[1] bb[21] WL[19] WL[20]
+ b[24] bb[3] bb[28] WL[38] WL[51] bb[8] WL[56] WL[62] b[3] bb[14] WL[29] WL[50] WL[24]
+ WL[43] WL[57] WL[63] b[13] WL[22] WL[59] bb[4] WL[41] WL[40] WL[54] bb[23] WL[31]
+ bb[17] VSS WL[26] WL[45] WL[52] WL[0] VDD Cell_array8x8_512x8m81
Xsaout_R_m2_512x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWE saout_m2_512x8m81_1/GWEN saout_R_m2_512x8m81_0/datain b[0] saout_R_m2_512x8m81_0/q
+ bb[1] saout_R_m2_512x8m81_0/pcb saout_R_m2_512x8m81_0/WEN saout_R_m2_512x8m81_0/wen_wm1_512x8m81_0/wen
+ saout_R_m2_512x8m81_0/mux821_512x8m81_0/ypass_gate_512x8m81_4/b bb[2] b[3] ypass[7]
+ bb[0] bb[5] VSS men b[7] a_15727_28608# a_15501_28608# a_15727_29383# a_15501_29383#
+ b[2] b[1] saout_m2_512x8m81_1/GWEN b[6] bb[3] b[5] ypass[0] VDD bb[4] b[4] ypass[1]
+ VDD ypass[4] bb[6] saout_R_m2_512x8m81_0/sa_512x8m81_0/wep saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ VDD ypass[2] ypass[5] VSS ypass[6] VSS saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb ypass[3]
+ VSS VDD bb[7] saout_R_m2_512x8m81
Xsaout_R_m2_512x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWE saout_m2_512x8m81_1/GWEN saout_R_m2_512x8m81_1/datain b[16] saout_R_m2_512x8m81_1/q
+ bb[17] saout_R_m2_512x8m81_1/pcb saout_R_m2_512x8m81_1/WEN saout_R_m2_512x8m81_1/wen_wm1_512x8m81_0/wen
+ saout_R_m2_512x8m81_1/mux821_512x8m81_0/ypass_gate_512x8m81_4/b bb[18] b[19] ypass[7]
+ bb[16] bb[21] VSS men b[23] a_4927_28608# a_4701_28608# a_4927_29383# a_4701_29383#
+ b[18] b[17] saout_m2_512x8m81_1/GWEN b[22] bb[19] b[21] ypass[0] VDD bb[20] b[20]
+ ypass[1] VDD ypass[4] bb[22] saout_R_m2_512x8m81_1/sa_512x8m81_0/wep saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ VDD ypass[2] ypass[5] VSS ypass[6] VSS saout_R_m2_512x8m81_1/sa_512x8m81_0/pcb ypass[3]
+ VSS VDD bb[23] saout_R_m2_512x8m81
Xsaout_m2_512x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] saout_m2_512x8m81_1/GWEN GWE bb[30] b[24] saout_m2_512x8m81_0/datain saout_m2_512x8m81_0/q
+ saout_m2_512x8m81_0/pcb saout_m2_512x8m81_0/WEN a_4236_28608# a_4461_28608# a_4236_29383#
+ a_4461_29383# bb[29] b[28] bb[31] bb[26] saout_m2_512x8m81_0/sacntl_2_512x8m81_0/a_4718_983#
+ ypass[7] b[31] saout_m2_512x8m81_0/mux821_512x8m81_0/a_4992_424# b[29] men b[30]
+ ypass[0] saout_m2_512x8m81_1/GWEN b[25] bb[28] b[26] VDD saout_m2_512x8m81_0/mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b
+ bb[27] ypass[1] b[27] VDD ypass[4] bb[25] saout_m2_512x8m81_0/sa_512x8m81_0/wep
+ saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# VDD ypass[2] VSS VSS saout_m2_512x8m81_0/pcb
+ ypass[3] VSS VDD bb[24] ypass[5] ypass[6] saout_m2_512x8m81
.ends

.subckt lcol4_512_512x8m81 WL[32] WL[33] WL[34] WL[38] WL[39] WL[35] WL[36] WL[37]
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51]
+ WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63]
+ WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+ WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+ WL[0] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] men ypass[0] ypass[1] ypass[2] ypass[3]
+ ypass[4] ypass[5] ypass[6] ypass[7] VSS GWEN GWE din[0] din[1] din[3] din[2] q[0]
+ q[1] q[2] q[3] pcb[2] pcb[3] pcb[0] pcb[1] vdd WEN[3] WEN[2] WEN[1] WEN[0] col_512a_512x8m81_0/WL[62]
+ col_512a_512x8m81_0/WL[29] col_512a_512x8m81_0/WL[46] col_512a_512x8m81_0/WL[63]
+ col_512a_512x8m81_0/a_15261_28608# col_512a_512x8m81_0/WL[47] col_512a_512x8m81_0/WL[48]
+ col_512a_512x8m81_0/saout_R_m2_512x8m81_0/wen_wm1_512x8m81_0/wen col_512a_512x8m81_0/WL[49]
+ col_512a_512x8m81_0/WL[10] col_512a_512x8m81_0/WL[11] col_512a_512x8m81_0/WL[12]
+ col_512a_512x8m81_0/WL[13] col_512a_512x8m81_0/WL[30] col_512a_512x8m81_0/WL[14]
+ col_512a_512x8m81_0/WL[31] col_512a_512x8m81_0/a_4701_29383# col_512a_512x8m81_0/WL[15]
+ col_512a_512x8m81_0/WL[32] col_512a_512x8m81_0/WL[0] col_512a_512x8m81_0/WL[16]
+ col_512a_512x8m81_0/WL[33] col_512a_512x8m81_0/WL[1] col_512a_512x8m81_0/WL[50]
+ col_512a_512x8m81_0/a_15501_28608# col_512a_512x8m81_0/WL[17] col_512a_512x8m81_0/WL[34]
+ col_512a_512x8m81_0/WL[2] col_512a_512x8m81_0/WL[51] col_512a_512x8m81_0/WL[18]
+ col_512a_512x8m81_0/WL[35] col_512a_512x8m81_0/a_4461_28608# col_512a_512x8m81_0/WL[3]
+ col_512a_512x8m81_0/WL[52] col_512a_512x8m81_0/WL[19] col_512a_512x8m81_0/WL[36]
+ col_512a_512x8m81_0/WL[53] col_512a_512x8m81_0/WL[4] col_512a_512x8m81_0/WL[37]
+ col_512a_512x8m81_0/WL[54] col_512a_512x8m81_0/WL[5] col_512a_512x8m81_0/WL[38]
+ col_512a_512x8m81_0/WL[6] col_512a_512x8m81_0/WL[55] col_512a_512x8m81_0/WL[39]
+ col_512a_512x8m81_0/WL[7] col_512a_512x8m81_0/WL[56] col_512a_512x8m81_0/a_15261_29383#
+ col_512a_512x8m81_0/WL[8] col_512a_512x8m81_0/WL[57] col_512a_512x8m81_0/WL[58]
+ col_512a_512x8m81_0/WL[9] col_512a_512x8m81_0/WL[59] col_512a_512x8m81_0/saout_m2_512x8m81_0/WEN
+ col_512a_512x8m81_0/men col_512a_512x8m81_0/saout_m2_512x8m81_1/sa_512x8m81_0/pcb
+ col_512a_512x8m81_0/WL[20] col_512a_512x8m81_0/WL[21] col_512a_512x8m81_0/ypass[0]
+ col_512a_512x8m81_0/GWE col_512a_512x8m81_0/a_4701_28608# col_512a_512x8m81_0/WL[22]
+ col_512a_512x8m81_0/ypass[1] col_512a_512x8m81_0/WL[23] col_512a_512x8m81_0/WL[40]
+ col_512a_512x8m81_0/ypass[2] col_512a_512x8m81_0/saout_m2_512x8m81_1/GWEN col_512a_512x8m81_0/WL[24]
+ col_512a_512x8m81_0/WL[41] col_512a_512x8m81_0/ypass[3] col_512a_512x8m81_0/WL[25]
+ ldummy_512x4_512x8m81_0/array16_512_dummy_01_512x8m81_0/VSS col_512a_512x8m81_0/saout_m2_512x8m81_0/pcb
+ col_512a_512x8m81_0/WL[42] col_512a_512x8m81_0/ypass[4] col_512a_512x8m81_0/WL[26]
+ col_512a_512x8m81_0/ypass[5] col_512a_512x8m81_0/WL[43] col_512a_512x8m81_0/WL[60]
+ col_512a_512x8m81_0/saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# col_512a_512x8m81_0/a_15501_29383#
+ col_512a_512x8m81_0/saout_R_m2_512x8m81_1/sa_512x8m81_0/pcb col_512a_512x8m81_0/saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb
+ col_512a_512x8m81_0/WL[27] col_512a_512x8m81_0/ypass[6] col_512a_512x8m81_0/WL[44]
+ col_512a_512x8m81_0/WL[61] col_512a_512x8m81_0/WL[28] VDD col_512a_512x8m81_0/ypass[7]
+ col_512a_512x8m81_0/WL[45] col_512a_512x8m81_0/a_4461_29383# VSUBS
Xldummy_512x4_512x8m81_0 VSUBS col_512a_512x8m81_0/b[19] col_512a_512x8m81_0/WL[63]
+ col_512a_512x8m81_0/b[2] col_512a_512x8m81_0/WL[33] VSUBS col_512a_512x8m81_0/bb[18]
+ VDD col_512a_512x8m81_0/WL[1] col_512a_512x8m81_0/bb[23] col_512a_512x8m81_0/WL[37]
+ VSUBS col_512a_512x8m81_0/b[17] col_512a_512x8m81_0/bb[7] col_512a_512x8m81_0/WL[26]
+ VDD col_512a_512x8m81_0/WL[5] VDD col_512a_512x8m81_0/b[26] VSUBS col_512a_512x8m81_0/WL[39]
+ VDD col_512a_512x8m81_0/bb[22] col_512a_512x8m81_0/bb[16] col_512a_512x8m81_0/WL[24]
+ VDD VDD col_512a_512x8m81_0/b[16] col_512a_512x8m81_0/WL[7] col_512a_512x8m81_0/bb[13]
+ col_512a_512x8m81_0/bb[20] col_512a_512x8m81_0/bb[24] col_512a_512x8m81_0/WL[22]
+ ldummy_512x4_512x8m81_0/array16_512_dummy_01_512x8m81_0/VSS col_512a_512x8m81_0/WL[9]
+ col_512a_512x8m81_0/bb[1] col_512a_512x8m81_0/b[25] col_512a_512x8m81_0/b[21] col_512a_512x8m81_0/WL[20]
+ col_512a_512x8m81_0/WL[11] col_512a_512x8m81_0/b[22] col_512a_512x8m81_0/b[19] VSUBS
+ col_512a_512x8m81_0/bb[26] col_512a_512x8m81_0/WL[18] col_512a_512x8m81_0/b[6] VDD
+ VDD col_512a_512x8m81_0/WL[13] VDD col_512a_512x8m81_0/bb[27] col_512a_512x8m81_0/b[11]
+ VSUBS VSUBS col_512a_512x8m81_0/b[27] col_512a_512x8m81_0/bb[18] col_512a_512x8m81_0/WL[16]
+ VDD col_512a_512x8m81_0/WL[15] col_512a_512x8m81_0/b[24] VDD col_512a_512x8m81_0/b[13]
+ col_512a_512x8m81_0/b[12] col_512a_512x8m81_0/b[17] VSUBS col_512a_512x8m81_0/b[29]
+ col_512a_512x8m81_0/WL[14] col_512a_512x8m81_0/WL[17] VDD col_512a_512x8m81_0/bb[12]
+ col_512a_512x8m81_0/b[0] VSUBS col_512a_512x8m81_0/bb[28] col_512a_512x8m81_0/bb[16]
+ col_512a_512x8m81_0/b[1] col_512a_512x8m81_0/WL[12] VDD col_512a_512x8m81_0/b[20]
+ col_512a_512x8m81_0/bb[14] col_512a_512x8m81_0/bb[24] VSUBS VSUBS col_512a_512x8m81_0/b[4]
+ col_512a_512x8m81_0/WL[10] col_512a_512x8m81_0/bb[0] VDD VDD VDD col_512a_512x8m81_0/bb[29]
+ col_512a_512x8m81_0/b[7] VSUBS VSUBS col_512a_512x8m81_0/b[25] VSUBS col_512a_512x8m81_0/WL[8]
+ col_512a_512x8m81_0/bb[8] col_512a_512x8m81_0/WL[46] VDD VDD col_512a_512x8m81_0/bb[25]
+ VDD col_512a_512x8m81_0/bb[6] col_512a_512x8m81_0/b[14] col_512a_512x8m81_0/bb[26]
+ VSUBS col_512a_512x8m81_0/b[9] col_512a_512x8m81_0/WL[44] VDD col_512a_512x8m81_0/bb[4]
+ col_512a_512x8m81_0/b[8] VSUBS col_512a_512x8m81_0/bb[10] col_512a_512x8m81_0/WL[42]
+ col_512a_512x8m81_0/bb[21] col_512a_512x8m81_0/b[5] VSUBS col_512a_512x8m81_0/b[31]
+ VSUBS col_512a_512x8m81_0/WL[40] col_512a_512x8m81_0/bb[5] VDD col_512a_512x8m81_0/b[3]
+ col_512a_512x8m81_0/b[28] VSUBS VSUBS col_512a_512x8m81_0/b[23] VDD VSUBS col_512a_512x8m81_0/WL[38]
+ VDD VDD col_512a_512x8m81_0/b[26] col_512a_512x8m81_0/bb[2] col_512a_512x8m81_0/bb[15]
+ col_512a_512x8m81_0/bb[22] VSUBS col_512a_512x8m81_0/WL[36] col_512a_512x8m81_0/bb[9]
+ VSUBS col_512a_512x8m81_0/bb[20] col_512a_512x8m81_0/WL[32] col_512a_512x8m81_0/b[21]
+ col_512a_512x8m81_0/bb[27] VSUBS col_512a_512x8m81_0/WL[34] VSUBS col_512a_512x8m81_0/bb[3]
+ VDD VDD col_512a_512x8m81_0/b[11] VSUBS VSUBS VSUBS col_512a_512x8m81_0/WL[30] VDD
+ VDD col_512a_512x8m81_0/b[13] col_512a_512x8m81_0/bb[7] col_512a_512x8m81_0/WL[28]
+ VSUBS col_512a_512x8m81_0/WL[61] col_512a_512x8m81_0/b[10] col_512a_512x8m81_0/bb[12]
+ VSUBS col_512a_512x8m81_0/WL[3] col_512a_512x8m81_0/bb[1] col_512a_512x8m81_0/bb[14]
+ col_512a_512x8m81_0/bb[29] VSUBS VSUBS col_512a_512x8m81_0/WL[62] col_512a_512x8m81_0/b[2]
+ VDD VDD col_512a_512x8m81_0/bb[19] col_512a_512x8m81_0/b[15] VSUBS VSUBS VDD VSUBS
+ col_512a_512x8m81_0/WL[60] VDD col_512a_512x8m81_0/b[22] VDD col_512a_512x8m81_0/b[30]
+ col_512a_512x8m81_0/b[7] VSUBS col_512a_512x8m81_0/WL[58] VSUBS col_512a_512x8m81_0/WL[56]
+ VDD col_512a_512x8m81_0/b[0] col_512a_512x8m81_0/b[28] VSUBS col_512a_512x8m81_0/WL[54]
+ VSUBS VDD VDD col_512a_512x8m81_0/b[18] VSUBS VSUBS col_512a_512x8m81_0/WL[52] VDD
+ col_512a_512x8m81_0/b[20] VDD col_512a_512x8m81_0/bb[15] col_512a_512x8m81_0/WL[50]
+ VSUBS VDD col_512a_512x8m81_0/b[6] col_512a_512x8m81_0/bb[6] VSUBS col_512a_512x8m81_0/WL[41]
+ col_512a_512x8m81_0/WL[48] col_512a_512x8m81_0/b[8] col_512a_512x8m81_0/bb[4] col_512a_512x8m81_0/b[30]
+ VSUBS VSUBS col_512a_512x8m81_0/WL[43] col_512a_512x8m81_0/bb[11] VDD VDD col_512a_512x8m81_0/bb[17]
+ col_512a_512x8m81_0/b[5] VSUBS col_512a_512x8m81_0/WL[45] VDD VSUBS VDD VDD col_512a_512x8m81_0/bb[21]
+ VDD col_512a_512x8m81_0/b[3] VSUBS col_512a_512x8m81_0/WL[47] VDD col_512a_512x8m81_0/b[4]
+ col_512a_512x8m81_0/bb[2] col_512a_512x8m81_0/WL[49] VSUBS col_512a_512x8m81_0/bb[9]
+ col_512a_512x8m81_0/b[1] col_512a_512x8m81_0/bb[31] VSUBS col_512a_512x8m81_0/WL[51]
+ VSUBS col_512a_512x8m81_0/bb[13] VDD col_512a_512x8m81_0/b[16] VDD col_512a_512x8m81_0/bb[0]
+ VSUBS col_512a_512x8m81_0/WL[53] VSUBS VDD col_512a_512x8m81_0/bb[30] VDD col_512a_512x8m81_0/bb[19]
+ VDD col_512a_512x8m81_0/bb[8] col_512a_512x8m81_0/WL[55] VSUBS col_512a_512x8m81_0/b[15]
+ col_512a_512x8m81_0/b[27] col_512a_512x8m81_0/bb[5] col_512a_512x8m81_0/b[9] col_512a_512x8m81_0/WL[57]
+ VSUBS col_512a_512x8m81_0/b[29] VDD col_512a_512x8m81_0/WL[6] col_512a_512x8m81_0/b[10]
+ col_512a_512x8m81_0/bb[10] col_512a_512x8m81_0/bb[23] col_512a_512x8m81_0/WL[59]
+ VSUBS VSUBS col_512a_512x8m81_0/WL[19] col_512a_512x8m81_0/b[12] VDD col_512a_512x8m81_0/bb[28]
+ col_512a_512x8m81_0/WL[4] VDD col_512a_512x8m81_0/b[24] VSUBS col_512a_512x8m81_0/WL[21]
+ VSUBS col_512a_512x8m81_0/bb[30] VDD col_512a_512x8m81_0/WL[0] VDD col_512a_512x8m81_0/b[18]
+ VDD VSUBS col_512a_512x8m81_0/WL[23] col_512a_512x8m81_0/b[31] col_512a_512x8m81_0/WL[2]
+ col_512a_512x8m81_0/bb[3] col_512a_512x8m81_0/WL[25] VSUBS col_512a_512x8m81_0/b[23]
+ col_512a_512x8m81_0/bb[31] VSUBS col_512a_512x8m81_0/WL[27] VSUBS VDD col_512a_512x8m81_0/b[14]
+ VDD col_512a_512x8m81_0/bb[25] VDD VDD col_512a_512x8m81_0/WL[29] VDD VSUBS VDD
+ col_512a_512x8m81_0/bb[17] VDD col_512a_512x8m81_0/WL[31] VSUBS col_512a_512x8m81_0/bb[11]
+ col_512a_512x8m81_0/WL[35] ldummy_512x4_512x8m81
Xdcap_103_novia_512x8m81_0[0] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[1] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[2] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[3] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[4] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[5] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[6] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[7] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[8] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[9] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[10] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[11] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[12] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[13] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[14] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[15] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[16] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[17] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[18] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[19] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[20] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[21] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[22] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[23] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[24] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[25] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[26] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[27] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[28] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[29] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[30] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[31] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[32] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[33] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[34] VDD VDD VSUBS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[35] VDD VDD VSUBS dcap_103_novia_512x8m81
Xcol_512a_512x8m81_0 col_512a_512x8m81_0/WL[3] col_512a_512x8m81_0/ypass[0] col_512a_512x8m81_0/ypass[1]
+ col_512a_512x8m81_0/ypass[3] col_512a_512x8m81_0/ypass[4] col_512a_512x8m81_0/ypass[5]
+ col_512a_512x8m81_0/GWE col_512a_512x8m81_0/WL[2] col_512a_512x8m81_0/WL[1] col_512a_512x8m81_0/WL[32]
+ col_512a_512x8m81_0/WL[31] col_512a_512x8m81_0/WL[30] col_512a_512x8m81_0/WL[29]
+ col_512a_512x8m81_0/WL[24] col_512a_512x8m81_0/WL[23] col_512a_512x8m81_0/WL[22]
+ col_512a_512x8m81_0/WL[21] col_512a_512x8m81_0/WL[57] col_512a_512x8m81_0/WL[56]
+ col_512a_512x8m81_0/WL[20] col_512a_512x8m81_0/WL[19] col_512a_512x8m81_0/WL[58]
+ col_512a_512x8m81_0/WL[59] col_512a_512x8m81_0/WL[49] col_512a_512x8m81_0/WL[48]
+ col_512a_512x8m81_0/WL[12] col_512a_512x8m81_0/WL[11] col_512a_512x8m81_0/WL[50]
+ col_512a_512x8m81_0/WL[51] col_512a_512x8m81_0/WL[41] col_512a_512x8m81_0/WL[40]
+ col_512a_512x8m81_0/WL[10] col_512a_512x8m81_0/WL[9] col_512a_512x8m81_0/WL[42]
+ col_512a_512x8m81_0/WL[43] col_512a_512x8m81_0/WL[35] col_512a_512x8m81_0/WL[34]
+ col_512a_512x8m81_0/WL[8] col_512a_512x8m81_0/WL[39] col_512a_512x8m81_0/WL[37]
+ col_512a_512x8m81_0/WL[7] col_512a_512x8m81_0/WL[33] col_512a_512x8m81_0/WL[6] col_512a_512x8m81_0/WL[38]
+ col_512a_512x8m81_0/WL[36] col_512a_512x8m81_0/WL[5] col_512a_512x8m81_0/WL[47]
+ col_512a_512x8m81_0/WL[45] col_512a_512x8m81_0/WL[4] col_512a_512x8m81_0/WL[46]
+ col_512a_512x8m81_0/WL[44] col_512a_512x8m81_0/WL[18] col_512a_512x8m81_0/WL[55]
+ col_512a_512x8m81_0/WL[53] col_512a_512x8m81_0/WL[17] col_512a_512x8m81_0/WL[54]
+ col_512a_512x8m81_0/WL[52] col_512a_512x8m81_0/WL[16] col_512a_512x8m81_0/WL[63]
+ col_512a_512x8m81_0/WL[61] col_512a_512x8m81_0/WL[15] col_512a_512x8m81_0/WL[14]
+ col_512a_512x8m81_0/WL[62] col_512a_512x8m81_0/WL[60] col_512a_512x8m81_0/WL[13]
+ col_512a_512x8m81_0/WL[28] col_512a_512x8m81_0/WL[27] col_512a_512x8m81_0/WL[26]
+ col_512a_512x8m81_0/WL[0] col_512a_512x8m81_0/ypass[2] col_512a_512x8m81_0/WL[25]
+ col_512a_512x8m81_0/b[10] col_512a_512x8m81_0/b[13] col_512a_512x8m81_0/b[16] col_512a_512x8m81_0/b[22]
+ col_512a_512x8m81_0/b[31] col_512a_512x8m81_0/din[1] col_512a_512x8m81_0/din[3]
+ col_512a_512x8m81_0/din[2] col_512a_512x8m81_0/din[0] col_512a_512x8m81_0/q[0] col_512a_512x8m81_0/q[1]
+ col_512a_512x8m81_0/q[2] col_512a_512x8m81_0/q[3] col_512a_512x8m81_0/b[17] col_512a_512x8m81_0/bb[10]
+ col_512a_512x8m81_0/bb[11] col_512a_512x8m81_0/bb[12] col_512a_512x8m81_0/bb[14]
+ col_512a_512x8m81_0/bb[15] col_512a_512x8m81_0/bb[16] col_512a_512x8m81_0/bb[22]
+ col_512a_512x8m81_0/bb[23] col_512a_512x8m81_0/bb[25] col_512a_512x8m81_0/bb[31]
+ col_512a_512x8m81_0/b[27] col_512a_512x8m81_0/b[0] col_512a_512x8m81_0/b[18] col_512a_512x8m81_0/pcb[0]
+ col_512a_512x8m81_0/pcb[1] col_512a_512x8m81_0/pcb[3] col_512a_512x8m81_0/pcb[2]
+ col_512a_512x8m81_0/WEN[3] col_512a_512x8m81_0/WEN[2] col_512a_512x8m81_0/WEN[1]
+ col_512a_512x8m81_0/WEN[0] col_512a_512x8m81_0/a_15501_29383# VSUBS col_512a_512x8m81_0/saout_R_m2_512x8m81_0/wen_wm1_512x8m81_0/wen
+ col_512a_512x8m81_0/a_15261_28608# col_512a_512x8m81_0/saout_m2_512x8m81_1/GWEN
+ col_512a_512x8m81_0/a_4701_29383# col_512a_512x8m81_0/b[8] col_512a_512x8m81_0/b[2]
+ col_512a_512x8m81_0/a_4461_28608# col_512a_512x8m81_0/bb[3] col_512a_512x8m81_0/a_15501_28608#
+ col_512a_512x8m81_0/b[5] col_512a_512x8m81_0/b[4] col_512a_512x8m81_0/ypass[6] col_512a_512x8m81_0/ypass[7]
+ col_512a_512x8m81_0/bb[5] col_512a_512x8m81_0/bb[26] col_512a_512x8m81_0/a_15261_29383#
+ col_512a_512x8m81_0/b[11] col_512a_512x8m81_0/bb[0] col_512a_512x8m81_0/bb[19] col_512a_512x8m81_0/b[1]
+ col_512a_512x8m81_0/saout_m2_512x8m81_1/sa_512x8m81_0/pcb col_512a_512x8m81_0/bb[24]
+ col_512a_512x8m81_0/bb[9] col_512a_512x8m81_0/bb[21] col_512a_512x8m81_0/b[24] col_512a_512x8m81_0/bb[2]
+ col_512a_512x8m81_0/b[6] col_512a_512x8m81_0/a_4701_28608# col_512a_512x8m81_0/b[3]
+ col_512a_512x8m81_0/saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# col_512a_512x8m81_0/bb[18]
+ col_512a_512x8m81_0/b[30] col_512a_512x8m81_0/b[20] col_512a_512x8m81_0/bb[8] col_512a_512x8m81_0/bb[4]
+ col_512a_512x8m81_0/b[19] col_512a_512x8m81_0/bb[29] col_512a_512x8m81_0/saout_m2_512x8m81_0/WEN
+ col_512a_512x8m81_0/b[23] col_512a_512x8m81_0/b[14] col_512a_512x8m81_0/b[5] col_512a_512x8m81_0/bb[20]
+ col_512a_512x8m81_0/b[29] col_512a_512x8m81_0/b[28] col_512a_512x8m81_0/b[25] col_512a_512x8m81_0/saout_m2_512x8m81_0/pcb
+ col_512a_512x8m81_0/bb[13] col_512a_512x8m81_0/men col_512a_512x8m81_0/saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb
+ col_512a_512x8m81_0/saout_R_m2_512x8m81_1/sa_512x8m81_0/pcb col_512a_512x8m81_0/bb[28]
+ col_512a_512x8m81_0/bb[7] col_512a_512x8m81_0/bb[17] col_512a_512x8m81_0/bb[6] col_512a_512x8m81_0/bb[1]
+ col_512a_512x8m81_0/b[21] col_512a_512x8m81_0/b[26] col_512a_512x8m81_0/bb[27] col_512a_512x8m81_0/b[12]
+ col_512a_512x8m81_0/b[9] col_512a_512x8m81_0/a_4461_29383# col_512a_512x8m81_0/b[15]
+ col_512a_512x8m81_0/bb[30] VDD col_512a_512x8m81_0/b[7] VSUBS col_512a_512x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_512x8m81 a_n36_52# a_444_n42# a_246_342# a_126_298#
+ m3_n36_330# a_36_n42# w_n68_622# VSUBS
X0 a_444_206# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_126_298# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_444_206# a_246_342# a_126_298# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_444_206# a_246_342# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt nmos_5p04310591302098_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.38u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.38u l=0.6u
.ends

.subckt ypass_gate_512x8m81_0 vss bb db ypass pcb vdd d m3_n1_4331# m3_n1_1708# m3_n1_1160#
+ m3_n1_2030# m3_n1_3366# m3_n1_2352# b m3_n1_3688# m3_n1_4009# m3_n1_2674# a_66_539#
+ pmos_5p0431059130201_512x8m81_2/D
Xnmos_5p0431059130202_512x8m81_0 nmos_5p0431059130202_512x8m81_0/D a_66_539# vss a_66_539#
+ vss nmos_5p0431059130202_512x8m81
Xnmos_5p0431059130200_512x8m81_0 pmos_5p0431059130201_512x8m81_2/D a_66_539# bb vss
+ nmos_5p0431059130200_512x8m81
Xnmos_5p0431059130200_512x8m81_1 d a_66_539# b vss nmos_5p0431059130200_512x8m81
Xpmos_5p0431059130201_512x8m81_0 vdd d nmos_5p0431059130202_512x8m81_0/D b pmos_5p0431059130201_512x8m81
Xpmos_5p0431059130201_512x8m81_1 vdd b pcb bb pmos_5p0431059130201_512x8m81
Xpmos_5p0431059130201_512x8m81_2 vdd pmos_5p0431059130201_512x8m81_2/D nmos_5p0431059130202_512x8m81_0/D
+ bb pmos_5p0431059130201_512x8m81
X0 nmos_5p0431059130202_512x8m81_0/D a_66_539# vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd a_66_539# nmos_5p0431059130202_512x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt nmos_5p04310591302096_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=8.5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=8.5u l=0.6u
.ends

.subckt pmos_5p04310591302097_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10.64u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.64u l=0.6u
.ends

.subckt pmos_5p04310591302095_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.51u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.51u l=0.6u
.ends

.subckt rdummy_512x4_512x8m81 tblhl pcb 018SRAM_cell1_dummy_512x8m81_39/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_20/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_36/m3_n36_330#
+ 018SRAM_strap1_bndry_512x8m81_21/a_36_52# 018SRAM_cell1_dummy_512x8m81_45/m2_90_n50#
+ m3_22279_n11418# 018SRAM_cell1_dummy_R_512x8m81_62/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_23/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_21/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_37/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_55/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_16/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_52/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_33/a_246_342# 018SRAM_strap1_bndry_512x8m81_37/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_1/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_39/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_22/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_38/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_26/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_0/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_43/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_12/a_36_52# 018SRAM_cell1_dummy_512x8m81_23/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_39/m3_n36_330# 018SRAM_cell1_dummy_R_512x8m81_20/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_31/a_126_298# 018SRAM_cell1_dummy_512x8m81_36/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_53/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_14/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_43/a_36_52# 018SRAM_cell1_dummy_512x8m81_24/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_21/m3_n36_330# 018SRAM_strap1_bndry_512x8m81_28/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_46/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_63/a_246_342#
+ m3_22279_n9439# 018SRAM_cell1_dummy_R_512x8m81_24/a_246_342# m3_22426_n25051# 018SRAM_cell1_dummy_512x8m81_25/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_1/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_22/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_56/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_40/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_17/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_59/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_34/a_246_342# 018SRAM_cell1_dummy_512x8m81_26/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_8/a_36_52# 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_23/m3_n36_330# 018SRAM_cell1_dummy_R_512x8m81_1/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_27/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_34/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_44/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_19/a_36_52# 018SRAM_cell1_dummy_512x8m81_27/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_24/m3_n36_330# 018SRAM_cell1_dummy_R_512x8m81_60/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_37/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_35/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_65/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_54/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_15/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_0/w_n68_622# 018SRAM_cell1_dummy_512x8m81_28/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_25/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_60/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_40/a_36_52# 018SRAM_cell1_dummy_512x8m81_47/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_25/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_64/a_246_342# 018SRAM_cell1_dummy_512x8m81_29/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_25/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_31/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_2/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_26/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_61/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_57/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_64/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_18/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_35/a_246_342# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_56/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_27/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_62/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_58/a_126_298# 018SRAM_cell1_dummy_512x8m81_28/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_8/a_126_298# 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_5/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_45/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_31/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_40/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_28/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_63/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_16/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_61/a_126_298# 018SRAM_cell1_dummy_512x8m81_38/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_60/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_16/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_55/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_29/m3_n36_330#
+ 018SRAM_strap1_bndry_512x8m81_62/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_10/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_48/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_32/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_61/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_47/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_65/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_26/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_60/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_3/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_11/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_19/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_58/m2_90_n50#
+ 018SRAM_strap1_bndry_512x8m81_22/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_62/m3_n36_330#
+ DWL 018SRAM_cell1_dummy_R_512x8m81_36/a_246_342# 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_12/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_6/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_63/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_29/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_53/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_46/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_64/w_n68_622# 018SRAM_cell1_dummy_512x8m81_16/m2_390_n50#
+ 018SRAM_strap1_bndry_512x8m81_2/a_36_52# 018SRAM_strap1_bndry_512x8m81_38/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_13/m3_n36_330# 018SRAM_cell1_dummy_R_512x8m81_62/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_64/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_39/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_56/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_17/a_246_342# 018SRAM_strap1_bndry_512x8m81_13/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_17/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_8/w_n68_622#
+ 018SRAM_cell1_dummy_R_512x8m81_58/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_14/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_65/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_49/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_27/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_61/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_18/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_44/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_4/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_15/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_50/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_59/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_57/a_126_298# 018SRAM_strap1_bndry_512x8m81_29/a_36_52#
+ ypass_gate_512x8m81_0_0/d 018SRAM_cell1_dummy_R_512x8m81_37/a_246_342# m3_22279_n11740#
+ 018SRAM_cell1_dummy_512x8m81_19/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_32/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_16/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_51/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_53/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_2/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_47/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_50/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_17/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_52/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_9/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_63/a_126_298# 018SRAM_strap1_bndry_512x8m81_35/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_18/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_57/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_6/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_18/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_53/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_10/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_34/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_50/m3_n36_330#
+ m3_22279_n9760# 018SRAM_cell1_dummy_R_512x8m81_28/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_62/w_n68_622#
+ 018SRAM_cell1_dummy_R_512x8m81_5/a_246_342# 018SRAM_cell1_dummy_512x8m81_54/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_51/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ 018SRAM_strap1_bndry_512x8m81_41/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_38/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_26/a_36_52# 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_55/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_54/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_20/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_4/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_48/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_57/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_56/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_57/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_53/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_30/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_33/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_58/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_6/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_53/w_n68_622#
+ 018SRAM_cell1_dummy_R_512x8m81_2/w_n68_622# 018SRAM_strap1_bndry_512x8m81_32/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_57/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_54/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_40/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_17/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_29/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_63/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_58/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_6/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_bndry_512x8m81_63/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_55/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_50/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ a_23341_1594# 018SRAM_cell1_dummy_R_512x8m81_39/a_246_342# 018SRAM_strap1_bndry_512x8m81_48/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_34/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_40/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_59/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_56/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_21/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_60/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_7/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_55/a_126_298# 018SRAM_strap1_bndry_512x8m81_23/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_49/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_2/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_41/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_57/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_65/a_126_298# 018SRAM_cell1_dummy_512x8m81_31/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_59/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_54/w_n68_622#
+ 018SRAM_cell1_dummy_R_512x8m81_4/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_3/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_42/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_3/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_58/m3_n36_330# 018SRAM_strap1_bndry_512x8m81_39/a_36_52#
+ w_22685_n22093# 018SRAM_cell1_dummy_512x8m81_41/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_36/a_126_298#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_33/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_4/m3_n36_330#
+ 018SRAM_strap1_bndry_512x8m81_14/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_7/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_43/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_59/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_40/m3_n36_330#
+ m3_22279_n11096# 018SRAM_cell1_dummy_512x8m81_51/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_60/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_35/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_5/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_44/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ 018SRAM_strap1_bndry_512x8m81_45/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_41/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_61/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_56/a_126_298#
+ 018SRAM_cell1_dummy_512x8m81_22/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_5/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_6/m3_n36_330# m3_22279_n10082# 018SRAM_strap1_bndry_512x8m81_20/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_45/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_42/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_32/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_55/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_7/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_7/w_n68_622# 018SRAM_cell1_dummy_512x8m81_46/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_43/m3_n36_330# 018SRAM_strap1_bndry_512x8m81_51/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_42/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_37/a_126_298#
+ 018SRAM_cell1_dummy_R_512x8m81_20/a_246_342# 018SRAM_strap1_bndry_512x8m81_36/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_65/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_8/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_47/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_8/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_44/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_52/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_11/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_30/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_9/m3_n36_330#
+ 018SRAM_cell1_dummy_R_512x8m81_36/w_n68_622# 018SRAM_cell1_dummy_512x8m81_48/m2_390_n50#
+ 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_45/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_23/m2_90_n50# 018SRAM_cell1_dummy_512x8m81_62/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_3/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_40/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_42/a_36_52# 018SRAM_cell1_dummy_512x8m81_49/m2_390_n50#
+ VSS 018SRAM_cell1_dummy_512x8m81_30/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_27/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_46/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_33/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_11/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_50/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_5/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_56/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_31/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_47/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_43/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_38/a_126_298#
+ 018SRAM_strap1_bndry_512x8m81_58/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_60/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_21/a_246_342# 018SRAM_strap1_bndry_512x8m81_7/a_36_52#
+ m3_22279_n10774# pmos_5p04310591302097_512x8m81_0/S 018SRAM_cell1_dummy_R_512x8m81_9/a_246_342#
+ 018SRAM_cell1_dummy_512x8m81_32/m2_390_n50# 018SRAM_strap1_bndry_512x8m81_33/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_48/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_512x8m81_53/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_31/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_18/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_37/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_33/m2_390_n50# 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_49/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_63/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_30/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_24/m2_90_n50#
+ 018SRAM_strap1_bndry_512x8m81_64/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_41/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_49/a_36_52# 018SRAM_cell1_dummy_512x8m81_34/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_31/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_34/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_51/a_246_342# 018SRAM_strap1_bndry_512x8m81_24/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_12/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_3/w_n68_622#
+ 018SRAM_cell1_dummy_512x8m81_35/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_32/m3_n36_330#
+ 018SRAM_cell1_dummy_512x8m81_44/m2_90_n50# 018SRAM_cell1_dummy_R_512x8m81_39/a_126_298#
+ a_n257_52# 018SRAM_cell1_dummy_R_512x8m81_22/a_246_342# 018SRAM_cell1_dummy_R_512x8m81_61/a_246_342#
+ 018SRAM_strap1_bndry_512x8m81_55/a_36_52# 018SRAM_cell1_dummy_512x8m81_36/m2_390_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_33/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_54/m2_90_n50#
+ 018SRAM_strap1_bndry_512x8m81_4/a_36_52# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_R_512x8m81_32/a_246_342# 018SRAM_strap1_bndry_512x8m81_30/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_38/w_n68_622# 018SRAM_cell1_dummy_512x8m81_37/m2_390_n50#
+ a_n257_1594# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50# 018SRAM_strap1_bndry_512x8m81_15/a_36_52#
+ 018SRAM_cell1_dummy_R_512x8m81_34/m3_n36_330# 018SRAM_cell1_dummy_512x8m81_25/m2_90_n50#
+ vdd 018SRAM_cell1_dummy_R_512x8m81_42/a_246_342# 018SRAM_strap1_bndry_512x8m81_61/a_36_52#
+ 018SRAM_cell1_dummy_512x8m81_38/m2_390_n50# 018SRAM_cell1_dummy_R_512x8m81_35/m3_n36_330#
+ m3_22279_n9117# vss 018SRAM_cell1_dummy_512x8m81_35/m2_90_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_strap1_bndry_512x8m81_46/a_36_52# 018SRAM_cell1_dummy_R_512x8m81_13/a_246_342#
X018SRAM_cell1_dummy_512x8m81_13 a_n257_52# 018SRAM_cell1_dummy_512x8m81_13/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_13/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_24 a_n257_52# 018SRAM_cell1_dummy_512x8m81_24/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_24/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_35 DWL 018SRAM_cell1_dummy_512x8m81_35/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_35/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_46 DWL 018SRAM_cell1_dummy_512x8m81_46/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_46/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_57 DWL 018SRAM_cell1_dummy_512x8m81_57/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_57/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_14 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_14/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_2/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_14/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_2/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_25 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_25/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_33/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_25/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_33/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_36 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_36/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_36/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_36/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_36/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_47 DWL ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_47/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_56/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_47/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_56/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_58 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_58/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_58/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_58/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_58/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_58 DWL 018SRAM_cell1_dummy_512x8m81_58/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_58/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_14 a_n257_52# 018SRAM_cell1_dummy_512x8m81_14/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_14/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_25 a_n257_52# 018SRAM_cell1_dummy_512x8m81_25/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_25/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_36 DWL 018SRAM_cell1_dummy_512x8m81_36/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_36/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_47 DWL 018SRAM_cell1_dummy_512x8m81_47/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_47/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_0 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_17/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_10/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_15 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_15/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_4/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_15/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_4/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_26 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_26/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_65/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_26/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_65/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_37 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_37/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_37/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_37/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_37/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_48 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_48/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_61/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_48/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_61/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_59 DWL ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_59/a_246_342#
+ 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_59/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_59 DWL 018SRAM_cell1_dummy_512x8m81_59/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_59/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_15 a_n257_52# 018SRAM_cell1_dummy_512x8m81_15/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_15/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_26 a_n257_52# 018SRAM_cell1_dummy_512x8m81_26/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_26/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_37 DWL 018SRAM_cell1_dummy_512x8m81_37/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_37/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_48 DWL 018SRAM_cell1_dummy_512x8m81_48/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_48/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_1 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_2/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_6/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_16 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_16/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_7/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_16/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_7/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_27 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_27/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_38/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_27/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_38/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_38 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_38/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_38/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_38/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_38/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_49 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_49/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_63/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_49/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_63/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_16 a_n257_52# 018SRAM_cell1_dummy_512x8m81_16/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_16/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_27 a_n257_52# 018SRAM_cell1_dummy_512x8m81_27/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_27/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_38 DWL 018SRAM_cell1_dummy_512x8m81_38/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_38/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_49 DWL 018SRAM_cell1_dummy_512x8m81_49/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_49/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_2 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_18/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_7/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_17 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_17/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_17/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_28 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_28/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_40/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_28/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_40/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_39 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_39/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_39/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_39/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_39/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_17 a_n257_52# 018SRAM_cell1_dummy_512x8m81_17/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_17/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_28 a_n257_52# 018SRAM_cell1_dummy_512x8m81_28/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_28/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_39 DWL 018SRAM_cell1_dummy_512x8m81_39/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_39/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_3 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_5/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_19/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_18 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_18/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_3/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_18/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_3/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_29 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_29/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_34/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_29/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_34/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_18 a_n257_52# 018SRAM_cell1_dummy_512x8m81_18/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_18/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_29 a_n257_52# 018SRAM_cell1_dummy_512x8m81_29/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_29/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_4 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_15/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_9/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_19 a_23341_1594# ypass_gate_512x8m81_0_0/bb vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# ypass_gate_512x8m81_0_0/b 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_19 a_n257_52# 018SRAM_cell1_dummy_512x8m81_19/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_19/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_2x_512x8m81_5 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_12/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_16/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_6 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_1/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_4/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_7 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_14/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_8/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_8 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_11/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_3/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_9 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_24/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_27/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_30 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_64/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_47/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_31 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_13/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_65/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_20 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_62/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_48/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
Xnmos_5p04310591302098_512x8m81_0 pmos_5p04310591302095_512x8m81_0/D ypass_gate_512x8m81_0_0/d
+ vss ypass_gate_512x8m81_0_0/d vss nmos_5p04310591302098_512x8m81
X018SRAM_cell1_2x_512x8m81_10 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_25/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_21/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_21 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_55/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_45/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_0 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_0/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_0/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_0/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_11 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_29/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_20/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_22 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_42/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_52/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_1 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_1/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_1/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_1/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_12 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_32/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_22/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_23 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_56/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_43/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_2 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_2/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_2/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_2/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_2/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_13 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_30/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_40/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_24 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_60/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_44/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_512x8m81_0 a_n257_52# 018SRAM_cell1_dummy_512x8m81_0/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_0/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_3 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_3/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_3/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_3/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_3/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_14 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_34/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_38/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_25 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_61/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_46/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_512x8m81_1 a_n257_52# 018SRAM_cell1_dummy_512x8m81_1/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_1/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_4 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_4/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_4/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_4/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_4/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_15 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_26/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_31/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_26 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_57/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_49/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_512x8m81_2 a_n257_52# 018SRAM_cell1_dummy_512x8m81_2/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_2/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_5 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_5/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
Xypass_gate_512x8m81_0_0 vss ypass_gate_512x8m81_0_0/bb ypass_gate_512x8m81_0_0/db
+ ypass_gate_512x8m81_0_0/ypass ypass_gate_512x8m81_0_0/pcb vdd ypass_gate_512x8m81_0_0/d
+ m3_22279_n9117# m3_22279_n11740# vdd m3_22279_n11418# m3_22279_n10082# m3_22279_n11096#
+ ypass_gate_512x8m81_0_0/b m3_22279_n9760# m3_22279_n9439# m3_22279_n10774# vdd ypass_gate_512x8m81_0_0/bb
+ ypass_gate_512x8m81_0
X018SRAM_cell1_2x_512x8m81_16 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_23/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_35/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_27 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_59/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_53/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_60 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_60/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_60/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_60/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_60/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_3 a_n257_52# 018SRAM_cell1_dummy_512x8m81_3/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_3/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
Xnmos_5p04310591302096_512x8m81_0 tblhl pmos_5p04310591302095_512x8m81_0/D vss pmos_5p04310591302095_512x8m81_0/D
+ vss nmos_5p04310591302096_512x8m81
X018SRAM_cell1_dummy_512x8m81_60 DWL 018SRAM_cell1_dummy_512x8m81_60/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_60/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
Xpmos_5p04310591302097_512x8m81_0 w_22685_n22093# tblhl pmos_5p04310591302095_512x8m81_0/D
+ pmos_5p04310591302097_512x8m81_0/S pmos_5p04310591302095_512x8m81_0/D pmos_5p04310591302097_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_6 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_6/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_6/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_6/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_6/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_17 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_39/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_36/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_28 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_63/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_50/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_50 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_50/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_60/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_50/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_60/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_61 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_61/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_61/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_61/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_61/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_4 a_n257_52# 018SRAM_cell1_dummy_512x8m81_4/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_4/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_61 DWL 018SRAM_cell1_dummy_512x8m81_61/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_61/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_50 DWL 018SRAM_cell1_dummy_512x8m81_50/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_50/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_7 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_7/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_7/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_7/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_7/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_18 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_28/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_33/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_29 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_58/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_51/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_512x8m81_5 a_n257_52# 018SRAM_cell1_dummy_512x8m81_5/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_5/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_40 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_40/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_40/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_40/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_40/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_51 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_51/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_58/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_51/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_58/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_62 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_62/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_62/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_62/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_62/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_62 DWL 018SRAM_cell1_dummy_512x8m81_62/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_62/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_40 DWL 018SRAM_cell1_dummy_512x8m81_40/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_40/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_51 DWL 018SRAM_cell1_dummy_512x8m81_51/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_51/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_8 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_8/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_8/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_8/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_8/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_2x_512x8m81_19 vss 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_strap1_bndry_512x8m81_41/a_36_52#
+ 018SRAM_strap1_bndry_512x8m81_37/a_36_52# 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_1594# 018SRAM_cell1_512x8m81_1/a_36_n42# a_n257_1594# vss vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ 018SRAM_cell1_512x8m81_1/a_444_n42# x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_dummy_512x8m81_6 a_n257_52# 018SRAM_cell1_dummy_512x8m81_6/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_6/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_30 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_30/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_39/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_30/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_39/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_41 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_41/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_64/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_41/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_64/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_52 DWL ypass_gate_512x8m81_0_0/bb vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL ypass_gate_512x8m81_0_0/b 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_63 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_63/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_63/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_63/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_63/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_63 DWL 018SRAM_cell1_dummy_512x8m81_63/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_63/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_30 a_n257_52# 018SRAM_cell1_dummy_512x8m81_30/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_30/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_41 DWL 018SRAM_cell1_dummy_512x8m81_41/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_41/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_52 DWL 018SRAM_cell1_dummy_512x8m81_52/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_52/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_9 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_9/a_246_342#
+ 018SRAM_cell1_512x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_512x8m81_9/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_64 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_64/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_64/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_64/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_64/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_20 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_20/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_31/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_20/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_31/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_31 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_31/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_31/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_31/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_31/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_42 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_42/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_53/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_42/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_53/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_53 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_53/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_53/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_53/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_53/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_7 a_n257_52# 018SRAM_cell1_dummy_512x8m81_7/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_7/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_20 a_n257_52# 018SRAM_cell1_dummy_512x8m81_20/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_20/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_31 a_n257_52# 018SRAM_cell1_dummy_512x8m81_31/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_31/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_42 DWL 018SRAM_cell1_dummy_512x8m81_42/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_42/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_53 DWL 018SRAM_cell1_dummy_512x8m81_53/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_53/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_65 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_65/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_65/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_65/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_65/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_10 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_0/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_10/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_0/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_21 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_21/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_35/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_21/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_35/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_32 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_32/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_32/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_32/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_32/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_43 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_43/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_57/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_43/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_57/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_54 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_54/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_54/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_54/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_54/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_8 a_n257_52# 018SRAM_cell1_dummy_512x8m81_8/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_8/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_10 a_n257_52# 018SRAM_cell1_dummy_512x8m81_10/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_10/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_21 a_n257_52# 018SRAM_cell1_dummy_512x8m81_21/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_21/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_32 DWL 018SRAM_cell1_dummy_512x8m81_32/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_32/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_43 DWL 018SRAM_cell1_dummy_512x8m81_43/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_43/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_54 DWL 018SRAM_cell1_dummy_512x8m81_54/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_54/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_11 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_11/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_1/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_11/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_22 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_22/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_37/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_22/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_37/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_33 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_33/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_33/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_33/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_33/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_44 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_44/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_55/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_44/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_55/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_55 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_55/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_55/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_55/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_55/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_512x8m81_9 a_n257_52# 018SRAM_cell1_dummy_512x8m81_9/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_9/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_11 a_n257_52# 018SRAM_cell1_dummy_512x8m81_11/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_11/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_22 a_n257_52# 018SRAM_cell1_dummy_512x8m81_22/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_22/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_33 DWL 018SRAM_cell1_dummy_512x8m81_33/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_33/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_44 DWL 018SRAM_cell1_dummy_512x8m81_44/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_44/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_55 DWL 018SRAM_cell1_dummy_512x8m81_55/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_55/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_12 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_12/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_8/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_12/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_8/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
Xpmos_5p04310591302095_512x8m81_0 vdd pmos_5p04310591302095_512x8m81_0/D ypass_gate_512x8m81_0_0/d
+ vdd ypass_gate_512x8m81_0_0/d pmos_5p04310591302095_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_23 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_23/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_36/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_23/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_36/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_34 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_34/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_34/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_34/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_34/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_45 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_45/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_62/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_45/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_62/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_56 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_56/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_56/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_56/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_56/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_512x8m81_0 a_n257_52# 018SRAM_cell1_512x8m81_1/a_444_n42# vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_512x8m81
X018SRAM_cell1_dummy_512x8m81_12 a_n257_52# 018SRAM_cell1_dummy_512x8m81_12/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_12/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_23 a_n257_52# 018SRAM_cell1_dummy_512x8m81_23/m2_90_n50#
+ vss 018SRAM_cell1_dummy_512x8m81_23/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_34 DWL 018SRAM_cell1_dummy_512x8m81_34/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_34/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_45 DWL 018SRAM_cell1_dummy_512x8m81_45/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_45/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_512x8m81_56 DWL 018SRAM_cell1_dummy_512x8m81_56/m2_90_n50# vss
+ 018SRAM_cell1_dummy_512x8m81_56/m2_390_n50# 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_13 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_13/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_6/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_13/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_6/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_24 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_24/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_32/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_24/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_32/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_35 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_35/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_35/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_35/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_35/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_46 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_46/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_54/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_46/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_54/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_dummy_R_512x8m81_57 a_23341_1594# ypass_gate_512x8m81_0_0/bb 018SRAM_cell1_dummy_R_512x8m81_57/a_246_342#
+ 018SRAM_cell1_dummy_R_512x8m81_57/a_126_298# 018SRAM_cell1_dummy_R_512x8m81_57/m3_n36_330#
+ ypass_gate_512x8m81_0_0/b 018SRAM_cell1_dummy_R_512x8m81_57/w_n68_622# vss x018SRAM_cell1_dummy_R_512x8m81
X018SRAM_cell1_512x8m81_1 a_n257_1594# 018SRAM_cell1_512x8m81_1/a_444_n42# vss 018SRAM_cell1_512x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_512x8m81_1/a_36_n42# 018SRAM_cell1_512x8m81_1/w_n68_622# vss x018SRAM_cell1_512x8m81
.ends

.subckt rarray4_512_512x8m81 WL[46] WL[35] WL[33] WL[49] WL[45] WL[39] WL[32] WL[54]
+ WL[38] WL[37] WL[44] WL[48] WL[34] WL[36] WL[43] WL[53] WL[50] WL[42] WL[52] WL[51]
+ WL[63] WL[62] WL[59] WL[56] WL[57] WL[60] WL[55] WL[29] WL[19] WL[7] WL[8] WL[25]
+ WL[9] WL[1] WL[22] WL[30] WL[24] WL[18] WL[31] WL[10] WL[14] WL[17] WL[11] WL[15]
+ WL[0] WL[2] WL[28] WL[12] WL[21] WL[4] WL[3] b[3] b[1] b[6] 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ WL[23] WL[5] 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42# WL[58] 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ WL[6] 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42# WL[40] 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ WL[26] bb[7] 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42# WL[47]
+ WL[61] b[7] b[5] 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ WL[20] 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42# WL[41] WL[27]
+ 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42# b[4] BL1B bb[4]
+ WL[13] BL1 BL WL[16] VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# b[0]
X018SRAM_cell1_2x_512x8m81_519 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_508 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_349 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_305 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_327 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_338 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_316 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_894 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_872 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_883 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_861 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_850 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[3] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_168 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_179 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_124 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[1] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_146 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[5] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_102 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[4] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_157 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[6] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_135 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[6] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_113 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[7] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_680 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_691 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_509 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_306 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_328 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_339 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_317 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_895 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_873 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_884 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_862 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_851 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[3] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_840 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[7] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_169 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_0 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_114 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[0] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_125 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[4] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_147 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[5] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_136 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[5] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_103 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[4] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_158 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[6] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_670 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_681 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_692 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_307 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_329 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_318 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_896 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_874 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_885 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_830 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[0] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_863 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_852 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[3] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_841 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[7] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_115 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[0] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_137 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_126 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[4] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_148 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[5] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_104 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[4] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_159 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[7] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_660 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_671 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_682 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_693 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_490 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_308 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_319 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_897 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_875 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_886 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_831 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[0] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_820 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[1] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_864 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_853 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[3] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_842 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[7] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_2 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_116 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[0] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_105 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[4] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_138 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_149 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[5] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_127 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[6] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_661 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_672 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_650 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_683 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_694 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_491 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_480 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_309 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_898 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_876 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_887 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_843 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[0] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_832 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[0] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_810 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[0] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_821 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[1] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_865 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_854 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[3] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_3 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_139 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_117 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[4] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_128 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[6] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_106 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[6] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_673 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_684 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_662 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_695 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_640 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_651 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_492 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_481 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_470 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_899 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_877 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_888 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_833 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[0] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_822 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[1] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_811 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[1] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_866 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_800 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[3] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_855 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[4] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_844 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[5] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_4 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_118 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[0] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_129 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[1] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_107 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[6] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_674 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_685 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_663 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_696 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_630 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_641 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_652 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_493 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_482 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_471 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_460 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_290 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_878 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_889 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_834 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[0] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_823 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[1] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_812 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[1] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_867 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[4] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_856 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[6] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_845 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[6] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_801 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[6] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_5 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_119 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[4] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_108 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[6] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_675 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_664 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_697 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_686 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_620 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_631 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_642 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_653 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_483 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_494 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_472 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_461 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_450 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_291 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_280 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_802 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[6] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_879 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_835 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[0] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_824 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[1] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_857 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[4] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_868 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[4] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_846 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] b[6] WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_813 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[6] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_6 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_109 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[6] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_665 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_676 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_698 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_632 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_687 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_654 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_621 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_610 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_643 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_473 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_462 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_484 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_440 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_451 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_495 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_270 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_281 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_292 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_825 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[1] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_847 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] b[5] WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_869 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[4] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_858 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[4] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_814 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[6] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_803 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[6] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_836 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[7] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_7 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_655 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_666 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_677 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_633 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_600 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_611 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_688 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_622 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_644 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_699 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_485 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_474 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_441 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_463 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_430 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_452 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_496 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_271 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_293 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_282 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_260 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_815 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[1] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_848 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[3] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_804 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[3] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_826 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[5] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_859 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[4] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_837 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[7] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_8 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_656 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_645 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_667 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_678 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_634 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_601 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_612 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_689 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_623 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_486 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_431 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_442 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_420 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_475 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_464 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_453 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_497 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_272 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_294 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_250 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_283 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_261 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_849 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[3] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_805 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[3] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_827 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[6] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_816 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[6] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_838 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[7] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_9 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_646 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_657 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_668 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_679 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_635 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_602 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_624 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_613 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_432 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_443 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_410 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_454 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_421 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_487 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_465 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_476 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_498 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_273 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_240 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_295 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_251 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_284 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_262 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_806 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[3] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_828 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[6] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_817 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[6] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_839 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] b[7] WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_647 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_658 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_669 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_636 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_625 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_603 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_614 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_488 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_400 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_433 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_444 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_466 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_477 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_455 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_411 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_422 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_499 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_230 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_274 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_241 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_252 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_296 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_285 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_263 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_807 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_818 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] b[5] WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_829 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] b[5] WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_637 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_659 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_626 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_604 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_615 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_648 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_489 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_401 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_478 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_434 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_445 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_456 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_467 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_412 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_423 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_990 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_220 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_231 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_264 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_242 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_275 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_253 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_297 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_286 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_819 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[1] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_808 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[4] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_90 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[0] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_605 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_627 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_616 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_638 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_649 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_402 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_479 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_435 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_446 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_468 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_457 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_413 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_424 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_980 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_991 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_221 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_210 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_232 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[6] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_265 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_243 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_276 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_254 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_298 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_287 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_809 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[6] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_91 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[0] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_80 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_606 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_628 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_617 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_639 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_403 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_436 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_458 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_447 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_469 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_414 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_425 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_981 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_970 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_992 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_200 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_222 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_211 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_233 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[6] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_266 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_244 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_277 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_255 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_299 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_288 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_92 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[0] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_70 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[1] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_81 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_607 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_629 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_618 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_404 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_459 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_437 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_448 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_415 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_426 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_982 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_960 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_971 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_993 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_201 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_234 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_223 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_212 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[3] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_267 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_245 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_289 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_278 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_256 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_790 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[7] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_93 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[0] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_71 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[1] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_82 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[5] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_60 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[7] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_608 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_619 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_405 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_427 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_438 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_449 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_416 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_983 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_961 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_950 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[0] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_972 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_994 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_235 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_202 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_213 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[3] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_224 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[5] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_268 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_246 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_279 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_257 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_780 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[4] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_791 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[7] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_50 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_94 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[0] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_83 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[1] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_72 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[5] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_61 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[7] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_609 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_428 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_406 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_417 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_439 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_940 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_984 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_962 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_951 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[0] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_973 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_995 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_203 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_225 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[5] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_214 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[7] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_770 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[1] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_781 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[4] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_236 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[4] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_269 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_247 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_258 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_792 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[4] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_40 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_51 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_84 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[3] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_73 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[5] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_62 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[7] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_95 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[0] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_407 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_429 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_418 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_941 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_985 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_930 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_963 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_952 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[3] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_974 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_996 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_204 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_226 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL1 WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_237 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[4] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_215 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[7] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_248 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_259 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_760 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_782 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[0] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_771 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[1] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_793 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[5] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_590 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_41 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_52 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_30 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_96 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[0] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_85 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[3] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_74 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[5] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_63 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[6] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_408 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_419 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_920 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_942 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_986 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_931 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_953 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[3] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_975 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_997 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_964 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_216 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_205 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_227 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL1 WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_238 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[0] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_249 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_761 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_750 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_783 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[0] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_772 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[3] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_794 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[4] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_580 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_591 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_42 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_53 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_20 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_31 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_97 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[3] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_86 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[3] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_75 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[5] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_64 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[6] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1020 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[7] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_409 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_921 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_910 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_943 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_987 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_954 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_932 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[7] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_976 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_998 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_965 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_217 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_206 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_239 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[0] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_228 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] b[1] WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_762 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_751 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_740 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_784 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[0] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_795 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_773 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[3] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_581 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_592 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_570 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_10 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_43 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_54 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_21 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_32 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_76 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_98 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[3] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_87 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[3] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_65 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[6] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1010 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[0] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1021 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[7] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_900 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_922 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_911 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_944 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_988 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_955 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_933 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[7] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_977 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_999 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_966 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_207 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_229 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] b[1] WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_218 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_763 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_752 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_730 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_741 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_785 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[0] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_796 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_774 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[5] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_560 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_582 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_593 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_571 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_11 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_44 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_55 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_22 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_33 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_66 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[1] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_77 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_88 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] b[3] WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_99 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] b[4] WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_390 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1011 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[0] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1022 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[6] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1000 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_934 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_901 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_923 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_945 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_989 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_912 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_956 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[5] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_978 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_967 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_208 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[14]
+ WL[15] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[14] BL WL[15] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_219 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_764 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_753 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_731 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_742 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_720 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_786 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[0] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_797 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_775 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[5] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_561 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_583 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_550 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_572 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_594 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_12 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_45 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_34 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_23 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_89 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] b[1] WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_78 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_67 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_56 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[7] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_391 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_380 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1012 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[3] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1023 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[6] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1001 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_935 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_902 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_924 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_946 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_913 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_957 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[5] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_979 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_968 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_209 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[16]
+ WL[17] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[16] BL WL[17] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_765 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_743 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_721 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_754 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_732 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_798 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_787 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[4] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_776 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[5] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_710 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_562 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_584 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_540 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_551 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_573 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_595 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_392 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_370 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_381 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_13 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_46 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_35 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_24 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_68 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[1] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_79 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_57 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[7] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1013 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[3] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1002 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_903 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_936 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_925 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_947 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_914 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_958 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[4] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_969 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_766 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_744 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_755 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_733 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_722 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_799 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_777 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] b[5] WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_788 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] b[7] WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_700 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_711 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_552 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_530 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_541 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_563 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_585 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_574 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_596 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_393 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_371 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_360 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_382 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_14 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_47 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_36 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_25 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_69 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[1] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_58 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] b[7] WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_190 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1014 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1003 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_904 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_937 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_926 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_915 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_948 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[1] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_959 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[4] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_745 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_767 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_756 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_734 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_723 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_789 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[7] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_778 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] b[7] WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_712 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_701 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_520 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_553 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_531 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_542 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_586 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_564 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_575 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_597 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_372 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_350 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_394 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_361 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_383 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_15 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_48 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_37 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_26 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_59 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] b[7] WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_191 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_180 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1015 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1004 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_927 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_905 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_916 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_949 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[1] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_938 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] b[6] WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_746 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_724 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_757 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_735 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_768 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] b[1] WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_779 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] b[5] WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_702 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_713 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_510 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_532 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_543 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_587 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_565 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_576 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL1 WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_598 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_554 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_521 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_49 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_38 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_16 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_27 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_351 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_395 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_362 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_340 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_384 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_373 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_192 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_181 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_170 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1016 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[5] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1005 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_906 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_917 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_928 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_939 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] b[6] WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_725 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_758 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_747 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_736 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_769 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] b[7] WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_703 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_714 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_522 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_511 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_599 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_555 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_533 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_544 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_588 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_566 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_577 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL1 WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_500 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_39 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_17 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_28 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_374 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_352 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_396 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_341 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_363 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_330 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_385 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_193 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_182 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_160 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_171 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1017 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[5] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1006 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] BL1 WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_907 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_918 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_929 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_759 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_737 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_748 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_726 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_704 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_715 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_501 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_523 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_973/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_512 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL1 WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_556 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_534 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_578 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_589 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL1 WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_545 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_567 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_375 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_320 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_353 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_397 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_364 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_342 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_386 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_331 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_18 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_29 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_183 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_194 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_161 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_172 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_150 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[3] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1018 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[4] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1007 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] BL1 WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_919 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_908 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_727 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_749 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_738 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_705 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_716 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_502 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_513 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_557 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_546 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_535 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_579 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_568 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_524 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_376 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_310 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_354 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_398 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_365 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_343 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_387 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_321 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_332 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_19 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_184 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_195 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_162 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_173 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_140 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_151 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[3] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1008 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[30]
+ WL[31] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[30] b[1] WL[31] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1019 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[4] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_909 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_23/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_728 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_739 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_706 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_717 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_503 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_514 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_558 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_536 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_547 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_569 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_525 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_377 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_311 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_344 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL1 WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_399 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_300 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_333 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_366 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_388 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_322 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_355 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_185 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_196 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_163 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_174 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_130 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[1] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_141 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_152 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[3] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_1009 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[32]
+ WL[33] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[32] b[1] WL[33] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_729 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_707 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_718 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_504 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL1 WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_515 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_559 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_537 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_548 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[38]
+ WL[39] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[38] BL WL[39] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_526 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_345 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_301 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_334 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_323 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_312 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL1 WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_890 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[62]
+ WL[63] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[62] BL1 WL[63] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_378 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL1 WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_367 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_389 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_356 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_186 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_197 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_164 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_175 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_131 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[1] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_142 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_153 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[3] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_120 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[7] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_708 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_719 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_505 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_977/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_516 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_538 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_549 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_527 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_965/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_346 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] BL WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_717/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_379 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] BL WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_302 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_335 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[12]
+ WL[13] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[12] BL WL[13] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_713/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_368 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_324 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_313 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL1 WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_357 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_891 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_880 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[56]
+ WL[57] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[56] BL1 WL[57] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_187 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_198 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_165 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_176 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_132 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[1] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_154 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] b[3] WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_110 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[5] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_143 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] b[7] WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_121 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[7] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_709 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[48]
+ WL[49] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[48] BL1 WL[49] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_506 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[40]
+ WL[41] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[40] BL1 WL[41] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_517 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_969/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_539 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[42]
+ WL[43] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[42] BL WL[43] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_528 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_347 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] BL WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_303 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL1 WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_336 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_369 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_325 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[8]
+ WL[9] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[8] BL WL[9] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_997/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_314 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL1 WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_358 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] BL1 WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_892 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] BL WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_881 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[58]
+ WL[59] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[58] BL1 WL[59] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_870 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] b[5] WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_100 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[2]
+ WL[3] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[2] b[4] WL[3] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_188 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_199 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_177 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] BL1 WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_166 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_6/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_155 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] b[3] WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_98/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_122 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[4] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_133 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[18]
+ WL[19] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[18] b[4] WL[19] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_111 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[5] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_144 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[7] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[7] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_518 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[44]
+ WL[45] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[44] BL1 WL[45] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_507 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[36]
+ WL[37] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[36] BL1 WL[37] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_529 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[34]
+ WL[35] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[34] BL1 WL[35] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_326 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_348 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[4]
+ WL[5] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[4] BL WL[5] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_993/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_304 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[10]
+ WL[11] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[10] BL1 WL[11] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_337 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_315 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[6]
+ WL[7] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[6] BL1 WL[7] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_359 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[26]
+ WL[27] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[26] BL1 WL[27] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_893 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[54]
+ WL[55] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[54] BL WL[55] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_8/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_882 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[60]
+ WL[61] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[60] BL1 WL[61] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_860 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[50]
+ WL[51] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[50] BL WL[51] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_871 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[52]
+ WL[53] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[52] b[5] WL[53] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_189 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL1 WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_167 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[28]
+ WL[29] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[28] BL WL[29] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_55/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_178 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[22]
+ WL[23] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[22] BL1 WL[23] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_112 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[24]
+ WL[25] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[24] b[0] WL[25] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_134 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[0] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_123 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[1] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_89/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_145 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[5] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_cell1_2x_512x8m81_82/018SRAM_cell1_512x8m81_1/a_444_n42#
+ x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_101 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[0]
+ WL[1] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[0] b[4] WL[1] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# bb[4] x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_156 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[20]
+ WL[21] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[20] b[6] WL[21] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
X018SRAM_cell1_2x_512x8m81_690 VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# WL[46]
+ WL[47] 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# 018SRAM_strap1_bndry_512x8m81_9/w_n68_622#
+ WL[46] BL1 WL[47] VSS VSS 018SRAM_strap1_bndry_512x8m81_9/w_n68_622# BL1B x018SRAM_cell1_2x_512x8m81
.ends

.subckt rcol4_512_512x8m81 WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[42] WL[44]
+ WL[46] WL[48] WL[50] WL[52] WL[54] WL[56] WL[57] WL[59] DWL WL[61] WL[51] WL[29]
+ WL[25] WL[24] WL[23] WL[22] WL[20] WL[27] WL[30] WL[18] WL[41] WL[15] WL[38] WL[45]
+ WL[43] WL[40] WL[39] WL[31] WL[14] WL[16] WL[17] WL[26] WL[19] WL[58] WL[60] WL[62]
+ WL[28] WL[63] WL[21] WL[49] WL[53] WL[47] WL[55] WL[0] WL[2] WL[12] WL[3] WL[4]
+ WL[7] WL[8] WL[9] WL[1] ypass[7] WL[5] ypass[0] WL[10] WL[13] ypass[1] ypass[2]
+ ypass[3] ypass[4] ypass[5] ypass[6] WL[6] tblhl GWEN WL[11] din[4] din[7] q[5] q[6]
+ q[7] din[5] din[6] q[4] pcb[6] pcb[7] pcb[4] vdd WEN[4] WEN[7] pcb[5] WEN[5] WEN[6]
+ rarray4_512_512x8m81_0/WL[39] rarray4_512_512x8m81_0/WL[56] a_17474_27175# rarray4_512_512x8m81_0/WL[57]
+ rarray4_512_512x8m81_0/WL[58] a_17474_27950# rarray4_512_512x8m81_0/WL[59] rarray4_512_512x8m81_0/WL[20]
+ GWE rarray4_512_512x8m81_0/WL[21] saout_R_m2_512x8m81_1/WEN rarray4_512_512x8m81_0/WL[22]
+ rarray4_512_512x8m81_0/WL[23] rarray4_512_512x8m81_0/WL[40] rdummy_512x4_512x8m81_0/VSS
+ rarray4_512_512x8m81_0/WL[24] rarray4_512_512x8m81_0/WL[41] rarray4_512_512x8m81_0/WL[25]
+ rarray4_512_512x8m81_0/WL[0] rarray4_512_512x8m81_0/WL[42] a_6674_27175# rarray4_512_512x8m81_0/WL[26]
+ rarray4_512_512x8m81_0/WL[1] rarray4_512_512x8m81_0/WL[43] rarray4_512_512x8m81_0/WL[60]
+ rarray4_512_512x8m81_0/WL[27] rarray4_512_512x8m81_0/WL[2] rarray4_512_512x8m81_0/WL[44]
+ a_17234_27175# a_6674_27950# rarray4_512_512x8m81_0/WL[61] rarray4_512_512x8m81_0/WL[28]
+ rarray4_512_512x8m81_0/WL[3] rarray4_512_512x8m81_0/WL[45] rarray4_512_512x8m81_0/WL[62]
+ rarray4_512_512x8m81_0/WL[29] rarray4_512_512x8m81_0/WL[4] rarray4_512_512x8m81_0/WL[46]
+ a_17234_27950# rarray4_512_512x8m81_0/WL[63] rdummy_512x4_512x8m81_0/pcb rarray4_512_512x8m81_0/WL[5]
+ rdummy_512x4_512x8m81_0/a_23341_1594# rarray4_512_512x8m81_0/WL[47] rarray4_512_512x8m81_0/WL[6]
+ rarray4_512_512x8m81_0/WL[48] rarray4_512_512x8m81_0/WL[7] rarray4_512_512x8m81_0/WL[49]
+ rarray4_512_512x8m81_0/WL[8] rarray4_512_512x8m81_0/WL[9] rarray4_512_512x8m81_0/WL[10]
+ men rarray4_512_512x8m81_0/WL[11] rarray4_512_512x8m81_0/WL[12] a_6434_27175# saout_m2_512x8m81_1/sa_512x8m81_0/pcb
+ rarray4_512_512x8m81_0/WL[13] rarray4_512_512x8m81_0/WL[30] rarray4_512_512x8m81_0/WL[14]
+ rarray4_512_512x8m81_0/WL[31] a_6434_27950# rarray4_512_512x8m81_0/WL[15] rarray4_512_512x8m81_0/WL[32]
+ saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# rdummy_512x4_512x8m81_0/DWL rarray4_512_512x8m81_0/WL[16]
+ rarray4_512_512x8m81_0/WL[33] rarray4_512_512x8m81_0/WL[50] rarray4_512_512x8m81_0/WL[17]
+ rarray4_512_512x8m81_0/WL[34] rarray4_512_512x8m81_0/WL[51] rarray4_512_512x8m81_0/WL[18]
+ rarray4_512_512x8m81_0/WL[35] rarray4_512_512x8m81_0/WL[52] rarray4_512_512x8m81_0/WL[19]
+ rarray4_512_512x8m81_0/WL[36] saout_m2_512x8m81_0/pcb rarray4_512_512x8m81_0/WL[53]
+ saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb saout_R_m2_512x8m81_1/pcb rarray4_512_512x8m81_0/WL[37]
+ rarray4_512_512x8m81_0/WL[54] rarray4_512_512x8m81_0/WL[38] rarray4_512_512x8m81_0/WL[55]
+ VDD VSS
Xsaout_m2_512x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWEN GWE saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/datain
+ saout_m2_512x8m81_1/q saout_m2_512x8m81_1/pcb saout_m2_512x8m81_1/WEN a_6209_27175#
+ a_6434_27175# a_6209_27950# a_6434_27950# saout_m2_512x8m81_1/bb[5] saout_m2_512x8m81_1/b[6]
+ saout_m2_512x8m81_1/bb[7] saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_1/sacntl_2_512x8m81_0/a_4718_983#
+ ypass[7] saout_m2_512x8m81_1/b[7] saout_m2_512x8m81_1/mux821_512x8m81_0/a_4992_424#
+ saout_m2_512x8m81_1/b[7] men saout_m2_512x8m81_1/b[6] ypass[0] GWEN saout_m2_512x8m81_1/b[7]
+ saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_1/b[6] VDD saout_m2_512x8m81_1/mux821_512x8m81_0/ypass_gate_a_512x8m81_0/b
+ saout_m2_512x8m81_1/bb[3] ypass[1] saout_m2_512x8m81_1/b[7] VDD ypass[4] saout_m2_512x8m81_1/bb[1]
+ saout_m2_512x8m81_1/sa_512x8m81_0/wep saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ VDD ypass[2] saout_m2_512x8m81_1/sacntl_2_512x8m81_0/a_4560_1922# VSS saout_m2_512x8m81_1/sa_512x8m81_0/pcb
+ ypass[3] saout_m2_512x8m81_1/outbuf_oe_512x8m81_0/a_4913_n316# VDD saout_m2_512x8m81_1/bb[6]
+ ypass[5] ypass[6] saout_m2_512x8m81
Xrdummy_512x4_512x8m81_0 tblhl rdummy_512x4_512x8m81_0/pcb saout_m2_512x8m81_1/b[6]
+ saout_R_m2_512x8m81_0/bb[2] rarray4_512_512x8m81_0/WL[35] rarray4_512_512x8m81_0/WL[39]
+ saout_m2_512x8m81_1/bb[6] ypass[1] VSS VSS saout_m2_512x8m81_1/b[6] VSS rarray4_512_512x8m81_0/WL[37]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[55]
+ VSS rarray4_512_512x8m81_0/WL[23] rarray4_512_512x8m81_0/WL[2] VDD saout_m2_512x8m81_0/bb[5]
+ saout_R_m2_512x8m81_0/bb[0] rarray4_512_512x8m81_0/WL[21] saout_m2_512x8m81_1/bb[3]
+ VDD VSS rarray4_512_512x8m81_0/WL[14] saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[25]
+ rarray4_512_512x8m81_0/WL[40] VDD saout_m2_512x8m81_1/bb[7] VSS VSS rarray4_512_512x8m81_0/WL[63]
+ saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[32] rarray4_512_512x8m81_0/WL[30]
+ saout_m2_512x8m81_1/b[7] VSS ypass[6] VSS VSS saout_m2_512x8m81_1/bb[6] VSS rarray4_512_512x8m81_0/WL[38]
+ saout_m2_512x8m81_1/bb[6] VDD saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[52]
+ VSS saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[7] saout_m2_512x8m81_0/b[4]
+ rarray4_512_512x8m81_0/WL[36] VDD saout_m2_512x8m81_1/bb[5] rarray4_512_512x8m81_0/WL[20]
+ saout_m2_512x8m81_0/bb[0] VSS rarray4_512_512x8m81_0/WL[17] saout_m2_512x8m81_1/b[7]
+ rarray4_512_512x8m81_0/WL[34] VDD saout_m2_512x8m81_1/bb[1] VDD saout_m2_512x8m81_0/b[1]
+ rarray4_512_512x8m81_0/WL[19] VSS VSS VDD saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[24]
+ saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[35] saout_m2_512x8m81_1/b[6]
+ saout_m2_512x8m81_1/b[7] VSS VSS saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[38]
+ VDD saout_R_m2_512x8m81_1/bb[4] VSS rarray4_512_512x8m81_0/WL[20] saout_R_m2_512x8m81_1/bb[4]
+ saout_m2_512x8m81_1/b[7] VDD saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_0/b[3]
+ VSS saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[62]
+ rarray4_512_512x8m81_0/WL[22] saout_R_m2_512x8m81_1/bb[0] VDD saout_m2_512x8m81_1/b[6]
+ VDD saout_m2_512x8m81_0/b[5] rarray4_512_512x8m81_0/WL[16] VSS rarray4_512_512x8m81_0/WL[29]
+ VDD saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[30] saout_m2_512x8m81_1/b[6]
+ rarray4_512_512x8m81_0/WL[15] VDD saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[49]
+ saout_m2_512x8m81_0/bb[4] VSS VSS saout_R_m2_512x8m81_1/bb[2] rarray4_512_512x8m81_0/WL[28]
+ rarray4_512_512x8m81_0/WL[46] rarray4_512_512x8m81_0/WL[5] saout_m2_512x8m81_0/bb[5]
+ VDD rarray4_512_512x8m81_0/WL[57] saout_m2_512x8m81_0/bb[6] rarray4_512_512x8m81_0/WL[43]
+ VSS VSS VDD saout_m2_512x8m81_1/b[6] VSS rarray4_512_512x8m81_0/WL[7] saout_m2_512x8m81_1/bb[6]
+ saout_m2_512x8m81_0/b[7] saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[41]
+ rarray4_512_512x8m81_0/WL[45] rdummy_512x4_512x8m81_0/DWL VSS saout_R_m2_512x8m81_1/bb[0]
+ saout_m2_512x8m81_0/bb[7] rarray4_512_512x8m81_0/WL[11] VDD rarray4_512_512x8m81_0/WL[53]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[53]
+ VSS VDD saout_R_m2_512x8m81_0/bb[6] rarray4_512_512x8m81_0/WL[4] rarray4_512_512x8m81_0/WL[21]
+ rarray4_512_512x8m81_0/WL[15] VDD rarray4_512_512x8m81_0/WL[42] saout_R_m2_512x8m81_1/bb[6]
+ saout_m2_512x8m81_1/bb[6] VSS VSS rarray4_512_512x8m81_0/WL[18] saout_R_m2_512x8m81_0/bb[4]
+ VDD VDD rarray4_512_512x8m81_0/WL[3] rarray4_512_512x8m81_0/WL[19] saout_m2_512x8m81_0/bb[1]
+ VSS VDD saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[59] VSS rarray4_512_512x8m81_0/WL[9]
+ saout_m2_512x8m81_0/b[7] saout_m2_512x8m81_1/bb[6] VDD rarray4_512_512x8m81_0/WL[36]
+ rdummy_512x4_512x8m81_0/ypass_gate_512x8m81_0_0/d VSS ypass[0] saout_m2_512x8m81_1/b[6]
+ VDD saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[13] saout_m2_512x8m81_0/bb[6]
+ VDD VDD VSS rarray4_512_512x8m81_0/WL[61] rarray4_512_512x8m81_0/WL[17] saout_m2_512x8m81_0/bb[0]
+ rarray4_512_512x8m81_0/WL[11] VDD rarray4_512_512x8m81_0/WL[25] VSS VSS VDD rarray4_512_512x8m81_0/WL[1]
+ saout_m2_512x8m81_0/bb[4] rarray4_512_512x8m81_0/WL[13] VDD rarray4_512_512x8m81_0/WL[50]
+ ypass[5] VSS VDD VSS saout_m2_512x8m81_0/b[3] rarray4_512_512x8m81_0/WL[48] saout_m2_512x8m81_1/b[7]
+ rarray4_512_512x8m81_0/WL[22] VSS rarray4_512_512x8m81_0/WL[28] saout_m2_512x8m81_1/b[7]
+ saout_m2_512x8m81_1/b[7] VDD saout_m2_512x8m81_1/b[7] VDD VSS VDD saout_m2_512x8m81_1/b[6]
+ rarray4_512_512x8m81_0/WL[48] rarray4_512_512x8m81_0/WL[59] saout_m2_512x8m81_1/bb[7]
+ VDD VSS rarray4_512_512x8m81_0/WL[5] VDD VDD rarray4_512_512x8m81_0/WL[40] saout_R_m2_512x8m81_1/bb[6]
+ rarray4_512_512x8m81_0/WL[43] saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[12]
+ VSS VDD saout_R_m2_512x8m81_1/bb[2] rarray4_512_512x8m81_0/WL[6] VSS VDD rarray4_512_512x8m81_0/WL[60]
+ rarray4_512_512x8m81_0/WL[51] saout_m2_512x8m81_0/bb[7] saout_m2_512x8m81_1/bb[6]
+ rdummy_512x4_512x8m81_0/a_23341_1594# VSS rarray4_512_512x8m81_0/WL[47] VDD rarray4_512_512x8m81_0/WL[8]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[61]
+ saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_1/bb[6] VDD VDD rarray4_512_512x8m81_0/WL[24]
+ VSS rarray4_512_512x8m81_0/WL[4] saout_R_m2_512x8m81_0/bb[0] rarray4_512_512x8m81_0/WL[55]
+ VDD saout_m2_512x8m81_1/bb[6] VSS VDD VDD rarray4_512_512x8m81_0/WL[2] saout_R_m2_512x8m81_0/bb[6]
+ rarray4_512_512x8m81_0/WL[1] rarray4_512_512x8m81_0/WL[47] rarray4_512_512x8m81_0/WL[26]
+ VDD saout_m2_512x8m81_1/b[7] VDD rdummy_512x4_512x8m81_0/ypass_gate_512x8m81_0_0/d
+ VDD rarray4_512_512x8m81_0/WL[10] rarray4_512_512x8m81_0/WL[6] VSS saout_R_m2_512x8m81_0/bb[4]
+ rarray4_512_512x8m81_0/WL[63] saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[29]
+ ypass[2] saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[58] VDD rarray4_512_512x8m81_0/WL[18]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[6] rarray4_512_512x8m81_0/WL[51]
+ rarray4_512_512x8m81_0/WL[41] saout_m2_512x8m81_1/b[7] VDD saout_m2_512x8m81_1/b[7]
+ VDD rarray4_512_512x8m81_0/WL[16] ypass[4] rarray4_512_512x8m81_0/WL[37] saout_m2_512x8m81_1/b[6]
+ rarray4_512_512x8m81_0/WL[60] saout_m2_512x8m81_1/bb[3] VSS VDD rarray4_512_512x8m81_0/WL[14]
+ VDD saout_R_m2_512x8m81_0/bb[2] rarray4_512_512x8m81_0/WL[56] rarray4_512_512x8m81_0/WL[57]
+ saout_m2_512x8m81_1/b[7] VDD VSS rarray4_512_512x8m81_0/WL[27] VDD rarray4_512_512x8m81_0/WL[12]
+ saout_m2_512x8m81_1/bb[6] VSS rarray4_512_512x8m81_0/WL[52] saout_m2_512x8m81_1/b[6]
+ saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[0] VSS rarray4_512_512x8m81_0/WL[0]
+ VDD saout_m2_512x8m81_0/b[5] saout_m2_512x8m81_0/bb[1] rarray4_512_512x8m81_0/WL[46]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_1/b[7] VDD VSS rarray4_512_512x8m81_0/WL[54]
+ saout_m2_512x8m81_0/b[1] rdummy_512x4_512x8m81_0/VSS saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[33]
+ rarray4_512_512x8m81_0/WL[44] saout_m2_512x8m81_1/bb[5] VSS VSS VDD VDD saout_m2_512x8m81_1/b[6]
+ rarray4_512_512x8m81_0/WL[62] saout_m2_512x8m81_1/b[7] VDD rarray4_512_512x8m81_0/WL[56]
+ VSS VSS rarray4_512_512x8m81_0/WL[9] ypass[3] VDD VSS saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[31]
+ rarray4_512_512x8m81_0/WL[58] saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_0/b[4]
+ VSS rarray4_512_512x8m81_0/WL[8] VDD saout_m2_512x8m81_1/b[7] saout_m2_512x8m81_1/b[6]
+ rarray4_512_512x8m81_0/WL[54] saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[26]
+ saout_m2_512x8m81_1/bb[1] rarray4_512_512x8m81_0/WL[42] VSS rarray4_512_512x8m81_0/WL[49]
+ saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[39] saout_m2_512x8m81_1/b[6]
+ VSS rarray4_512_512x8m81_0/WL[32] VSS VDD saout_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[33]
+ saout_m2_512x8m81_1/bb[6] VDD VSS VSS VSS rarray4_512_512x8m81_0/WL[50] saout_m2_512x8m81_1/b[7]
+ rarray4_512_512x8m81_0/WL[23] saout_m2_512x8m81_0/bb[3] rarray4_512_512x8m81_0/WL[3]
+ saout_m2_512x8m81_1/b[7] VSS rarray4_512_512x8m81_0/WL[34] VDD saout_m2_512x8m81_1/b[7]
+ VSS saout_m2_512x8m81_0/bb[3] rarray4_512_512x8m81_0/WL[10] rarray4_512_512x8m81_0/WL[27]
+ saout_m2_512x8m81_1/b[6] VDD VSS rarray4_512_512x8m81_0/WL[44] saout_m2_512x8m81_1/bb[6]
+ rarray4_512_512x8m81_0/WL[31] ypass[7] VSS saout_m2_512x8m81_1/b[6] VDD rarray4_512_512x8m81_0/WL[45]
+ VSS rdummy_512x4_512x8m81
Xdcap_103_novia_512x8m81_0[0] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[1] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[2] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[3] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[4] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[5] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[6] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[7] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[8] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[9] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[10] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[11] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[12] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[13] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[14] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[15] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[16] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[17] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[18] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[19] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[20] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[21] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[22] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[23] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[24] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[25] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[26] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[27] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[28] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[29] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[30] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[31] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[32] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[33] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[34] VDD VDD VSS dcap_103_novia_512x8m81
Xdcap_103_novia_512x8m81_0[35] VDD VDD VSS dcap_103_novia_512x8m81
Xrarray4_512_512x8m81_0 rarray4_512_512x8m81_0/WL[46] rarray4_512_512x8m81_0/WL[35]
+ rarray4_512_512x8m81_0/WL[33] rarray4_512_512x8m81_0/WL[49] rarray4_512_512x8m81_0/WL[45]
+ rarray4_512_512x8m81_0/WL[39] rarray4_512_512x8m81_0/WL[32] rarray4_512_512x8m81_0/WL[54]
+ rarray4_512_512x8m81_0/WL[38] rarray4_512_512x8m81_0/WL[37] rarray4_512_512x8m81_0/WL[44]
+ rarray4_512_512x8m81_0/WL[48] rarray4_512_512x8m81_0/WL[34] rarray4_512_512x8m81_0/WL[36]
+ rarray4_512_512x8m81_0/WL[43] rarray4_512_512x8m81_0/WL[53] rarray4_512_512x8m81_0/WL[50]
+ rarray4_512_512x8m81_0/WL[42] rarray4_512_512x8m81_0/WL[52] rarray4_512_512x8m81_0/WL[51]
+ rarray4_512_512x8m81_0/WL[63] rarray4_512_512x8m81_0/WL[62] rarray4_512_512x8m81_0/WL[59]
+ rarray4_512_512x8m81_0/WL[56] rarray4_512_512x8m81_0/WL[57] rarray4_512_512x8m81_0/WL[60]
+ rarray4_512_512x8m81_0/WL[55] rarray4_512_512x8m81_0/WL[29] rarray4_512_512x8m81_0/WL[19]
+ rarray4_512_512x8m81_0/WL[7] rarray4_512_512x8m81_0/WL[8] rarray4_512_512x8m81_0/WL[25]
+ rarray4_512_512x8m81_0/WL[9] rarray4_512_512x8m81_0/WL[1] rarray4_512_512x8m81_0/WL[22]
+ rarray4_512_512x8m81_0/WL[30] rarray4_512_512x8m81_0/WL[24] rarray4_512_512x8m81_0/WL[18]
+ rarray4_512_512x8m81_0/WL[31] rarray4_512_512x8m81_0/WL[10] rarray4_512_512x8m81_0/WL[14]
+ rarray4_512_512x8m81_0/WL[17] rarray4_512_512x8m81_0/WL[11] rarray4_512_512x8m81_0/WL[15]
+ rarray4_512_512x8m81_0/WL[0] rarray4_512_512x8m81_0/WL[2] rarray4_512_512x8m81_0/WL[28]
+ rarray4_512_512x8m81_0/WL[12] rarray4_512_512x8m81_0/WL[21] rarray4_512_512x8m81_0/WL[4]
+ rarray4_512_512x8m81_0/WL[3] saout_m2_512x8m81_0/b[3] saout_m2_512x8m81_0/b[1] saout_m2_512x8m81_0/bb[6]
+ saout_m2_512x8m81_1/bb[1] rarray4_512_512x8m81_0/WL[23] rarray4_512_512x8m81_0/WL[5]
+ saout_R_m2_512x8m81_0/bb[4] saout_R_m2_512x8m81_0/bb[2] saout_R_m2_512x8m81_1/bb[0]
+ rarray4_512_512x8m81_0/WL[58] saout_m2_512x8m81_0/bb[5] saout_m2_512x8m81_1/bb[5]
+ saout_R_m2_512x8m81_1/bb[6] rarray4_512_512x8m81_0/WL[6] saout_R_m2_512x8m81_0/bb[0]
+ rarray4_512_512x8m81_0/WL[40] saout_m2_512x8m81_1/bb[7] rarray4_512_512x8m81_0/WL[26]
+ saout_m2_512x8m81_0/bb[7] saout_m2_512x8m81_1/bb[3] rarray4_512_512x8m81_0/WL[47]
+ rarray4_512_512x8m81_0/WL[61] saout_m2_512x8m81_0/b[7] saout_m2_512x8m81_0/b[5]
+ saout_m2_512x8m81_0/bb[3] rarray4_512_512x8m81_0/WL[20] saout_R_m2_512x8m81_1/bb[2]
+ rarray4_512_512x8m81_0/WL[41] rarray4_512_512x8m81_0/WL[27] saout_m2_512x8m81_0/bb[1]
+ saout_R_m2_512x8m81_1/bb[4] saout_R_m2_512x8m81_0/bb[6] saout_m2_512x8m81_0/bb[4]
+ saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_0/b[4] rarray4_512_512x8m81_0/WL[13]
+ saout_m2_512x8m81_1/bb[6] saout_m2_512x8m81_1/b[7] rarray4_512_512x8m81_0/WL[16]
+ VSS VDD saout_m2_512x8m81_0/bb[0] rarray4_512_512x8m81
Xsaout_R_m2_512x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWE GWEN saout_R_m2_512x8m81_0/datain saout_m2_512x8m81_1/b[7] saout_R_m2_512x8m81_0/q
+ saout_m2_512x8m81_1/bb[6] saout_R_m2_512x8m81_0/pcb saout_R_m2_512x8m81_0/WEN saout_R_m2_512x8m81_0/wen_wm1_512x8m81_0/wen
+ saout_R_m2_512x8m81_0/mux821_512x8m81_0/ypass_gate_512x8m81_4/b saout_R_m2_512x8m81_0/bb[2]
+ saout_m2_512x8m81_1/b[6] ypass[7] saout_R_m2_512x8m81_0/bb[0] saout_m2_512x8m81_1/bb[6]
+ saout_R_m2_512x8m81_0/sacntl_2_512x8m81_0/a_4718_983# men saout_m2_512x8m81_1/b[6]
+ a_6900_27175# a_6674_27175# a_6900_27950# a_6674_27950# saout_m2_512x8m81_1/b[7]
+ saout_m2_512x8m81_1/b[6] GWEN saout_m2_512x8m81_1/b[7] saout_m2_512x8m81_1/bb[6]
+ saout_m2_512x8m81_1/b[6] ypass[0] VDD saout_R_m2_512x8m81_0/bb[4] saout_m2_512x8m81_1/b[7]
+ ypass[1] VDD ypass[4] saout_R_m2_512x8m81_0/bb[6] saout_R_m2_512x8m81_0/sa_512x8m81_0/wep
+ saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# VDD ypass[2] ypass[5] saout_R_m2_512x8m81_0/sacntl_2_512x8m81_0/a_4560_1922#
+ ypass[6] VSS saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb ypass[3] VSS VDD saout_m2_512x8m81_1/bb[6]
+ saout_R_m2_512x8m81
Xsaout_R_m2_512x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWE GWEN saout_R_m2_512x8m81_1/datain saout_m2_512x8m81_1/b[7] saout_R_m2_512x8m81_1/q
+ saout_m2_512x8m81_1/bb[6] saout_R_m2_512x8m81_1/pcb saout_R_m2_512x8m81_1/WEN saout_R_m2_512x8m81_1/wen_wm1_512x8m81_0/wen
+ saout_R_m2_512x8m81_1/mux821_512x8m81_0/ypass_gate_512x8m81_4/b saout_R_m2_512x8m81_1/bb[2]
+ saout_m2_512x8m81_1/b[6] ypass[7] saout_R_m2_512x8m81_1/bb[0] saout_m2_512x8m81_1/bb[6]
+ saout_R_m2_512x8m81_1/sacntl_2_512x8m81_0/a_4718_983# men saout_m2_512x8m81_1/b[6]
+ a_17700_27175# a_17474_27175# a_17700_27950# a_17474_27950# saout_m2_512x8m81_1/b[7]
+ saout_m2_512x8m81_1/b[6] GWEN saout_m2_512x8m81_1/b[7] saout_m2_512x8m81_1/bb[6]
+ saout_m2_512x8m81_1/b[6] ypass[0] VDD saout_R_m2_512x8m81_1/bb[4] saout_m2_512x8m81_1/b[7]
+ ypass[1] VDD ypass[4] saout_R_m2_512x8m81_1/bb[6] saout_R_m2_512x8m81_1/sa_512x8m81_0/wep
+ saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735# VDD ypass[2] ypass[5] saout_R_m2_512x8m81_1/sacntl_2_512x8m81_0/a_4560_1922#
+ ypass[6] VSS saout_R_m2_512x8m81_1/pcb ypass[3] saout_R_m2_512x8m81_1/outbuf_oe_512x8m81_0/a_4913_n316#
+ VDD saout_m2_512x8m81_1/b[7] saout_R_m2_512x8m81
Xsaout_m2_512x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ ypass[0] GWEN GWE saout_m2_512x8m81_0/bb[6] saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_0/datain
+ saout_m2_512x8m81_0/q saout_m2_512x8m81_0/pcb saout_m2_512x8m81_0/WEN a_17009_27175#
+ a_17234_27175# a_17009_27950# a_17234_27950# saout_m2_512x8m81_0/bb[5] saout_m2_512x8m81_0/b[4]
+ saout_m2_512x8m81_0/bb[7] saout_m2_512x8m81_1/b[7] VSS ypass[7] saout_m2_512x8m81_0/b[7]
+ saout_m2_512x8m81_0/mux821_512x8m81_0/a_4992_424# saout_m2_512x8m81_0/b[5] men saout_m2_512x8m81_1/b[6]
+ ypass[0] GWEN saout_m2_512x8m81_0/b[1] saout_m2_512x8m81_0/bb[4] saout_m2_512x8m81_1/b[6]
+ VDD saout_m2_512x8m81_1/b[6] saout_m2_512x8m81_0/bb[3] ypass[1] saout_m2_512x8m81_0/b[3]
+ VDD ypass[4] saout_m2_512x8m81_0/bb[1] saout_m2_512x8m81_0/sa_512x8m81_0/wep saout_m2_512x8m81_1/mux821_512x8m81_0/a_656_7735#
+ VDD ypass[2] VSS VSS saout_m2_512x8m81_0/pcb ypass[3] VSS VDD saout_m2_512x8m81_0/bb[0]
+ ypass[5] ypass[6] saout_m2_512x8m81
.ends

.subckt pmoscap_R270_512x8m81 m3_489_n1# m3_1409_n1# w_n60_n407# a_81_507#
X0 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
X1 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_5p043105913020100_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.63u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.63u l=0.6u
.ends

.subckt pmos_1p2_02_R90_512x8m81 pmos_5p043105913020100_512x8m81_0/S a_193_n71# a_n31_n71#
+ pmos_5p043105913020100_512x8m81_0/D w_n296_n137#
Xpmos_5p043105913020100_512x8m81_0 w_n296_n137# pmos_5p043105913020100_512x8m81_0/D
+ a_n31_n71# pmos_5p043105913020100_512x8m81_0/S a_193_n71# pmos_5p043105913020100_512x8m81
.ends

.subckt nmos_5p043105913020111_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.64u l=0.6u
.ends

.subckt pmoscap_L1_W2_R270_512x8m81 w_n60_n407# a_81_507# m3_509_n1#
X0 a_81_507# M3_M2$01_R270_512x8m81_0/VSUBS a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmos_5p043105913020101_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.59u l=0.6u
.ends

.subckt pmos_1p2_01_R90_512x8m81 w_n295_n137# pmos_5p043105913020101_512x8m81_0/S
+ pmos_5p043105913020101_512x8m81_0/D a_n31_n71#
Xpmos_5p043105913020101_512x8m81_0 w_n295_n137# pmos_5p043105913020101_512x8m81_0/D
+ a_n31_n71# pmos_5p043105913020101_512x8m81_0/S pmos_5p043105913020101_512x8m81
.ends

.subckt nmos_5p04310591302099_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=10.11u l=0.6u
.ends

.subckt nmos_5p043105913020102_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.59u l=0.6u
.ends

.subckt nmos_1p2_01_R270_512x8m81 nmos_5p043105913020102_512x8m81_0/S nmos_5p043105913020102_512x8m81_0/D
+ a_n31_n71# VSUBS
Xnmos_5p043105913020102_512x8m81_0 nmos_5p043105913020102_512x8m81_0/D a_n31_n71#
+ nmos_5p043105913020102_512x8m81_0/S VSUBS nmos_5p043105913020102_512x8m81
.ends

.subckt nmos_1p2_02_R90_512x8m81 nmos_5p04310591302099_512x8m81_0/D a_n31_n71# nmos_5p04310591302099_512x8m81_0/S
+ VSUBS
Xnmos_5p04310591302099_512x8m81_0 nmos_5p04310591302099_512x8m81_0/D a_n31_n71# nmos_5p04310591302099_512x8m81_0/S
+ VSUBS nmos_5p04310591302099_512x8m81
.ends

.subckt pmos_5p043105913020108_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.5u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.5u l=0.6u
.ends

.subckt pmos_1p2_01_R270_512x8m81 w_n296_n137# pmos_5p043105913020108_512x8m81_0/D
+ a_n31_n71# a_193_n71# pmos_5p043105913020108_512x8m81_0/S
Xpmos_5p043105913020108_512x8m81_0 w_n296_n137# pmos_5p043105913020108_512x8m81_0/D
+ a_n31_n71# pmos_5p043105913020108_512x8m81_0/S a_193_n71# pmos_5p043105913020108_512x8m81
.ends

.subckt pmos_5p043105913020104_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_1p2_02_R270_512x8m81 w_n296_n137# pmos_5p043105913020104_512x8m81_0/D
+ a_193_n71# pmos_5p043105913020104_512x8m81_0/S a_n31_n71#
Xpmos_5p043105913020104_512x8m81_0 w_n296_n137# pmos_5p043105913020104_512x8m81_0/D
+ a_n31_n71# pmos_5p043105913020104_512x8m81_0/S a_193_n71# pmos_5p043105913020104_512x8m81
.ends

.subckt pmos_5p043105913020105_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.62u l=0.6u
.ends

.subckt nmos_5p043105913020109_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_5p043105913020103_512x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
.ends

.subckt pmos_1p2_03_R270_512x8m81 w_n296_n137# pmos_5p043105913020103_512x8m81_0/D
+ a_193_n71# a_n31_n71# a_417_n71# pmos_5p043105913020103_512x8m81_0/S
Xpmos_5p043105913020103_512x8m81_0 w_n296_n137# pmos_5p043105913020103_512x8m81_0/D
+ a_n31_n71# pmos_5p043105913020103_512x8m81_0/S a_417_n71# a_193_n71# pmos_5p043105913020103_512x8m81
.ends

.subckt nmos_5p043105913020107_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=5u l=0.6u
.ends

.subckt nmos_5p043105913020106_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.66u l=0.6u
.ends

.subckt pmos_5p043105913020110_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.59u l=0.6u
.ends

.subckt nmos_1p2_02_R270_512x8m81 nmos_5p04310591302044_512x8m81_0/S a_n31_n71# nmos_5p04310591302044_512x8m81_0/D
+ VSUBS
Xnmos_5p04310591302044_512x8m81_0 nmos_5p04310591302044_512x8m81_0/D a_n31_n71# nmos_5p04310591302044_512x8m81_0/S
+ VSUBS nmos_5p04310591302044_512x8m81
.ends

.subckt xdec_512x8m81 RWL xc xb xa m2_16621_n223# m2_17754_n223# m2_11825_n223# m2_12202_n223#
+ m2_12958_n223# m2_15487_n223# m2_12580_n223# m2_15110_n223# m2_11069_n223# m2_15865_n223#
+ m2_16243_n223# m2_10314_n223# m2_16998_n223# m2_17376_n223# men m2_11447_n223# vdd
+ vss LWL m2_10691_n223#
Xpmos_1p2_01_R270_512x8m81_0 vdd pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D
+ nmos_5p043105913020109_512x8m81_0/S nmos_5p043105913020109_512x8m81_0/S vdd pmos_1p2_01_R270_512x8m81
Xpmos_1p2_01_R270_512x8m81_1 vdd pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D
+ nmos_5p043105913020109_512x8m81_0/S nmos_5p043105913020109_512x8m81_0/S vdd pmos_1p2_01_R270_512x8m81
Xpmos_1p2_02_R270_512x8m81_0 vdd men pmos_5p043105913020105_512x8m81_2/S nmos_5p043105913020109_512x8m81_0/S
+ pmos_5p043105913020105_512x8m81_2/S pmos_1p2_02_R270_512x8m81
Xpmos_5p043105913020105_512x8m81_0 vdd pmos_5p043105913020105_512x8m81_2/S xb vdd
+ pmos_5p043105913020105_512x8m81
Xpmos_5p043105913020105_512x8m81_1 vdd vdd xc pmos_5p043105913020105_512x8m81_2/S
+ pmos_5p043105913020105_512x8m81
Xpmos_5p043105913020105_512x8m81_2 vdd vdd xa pmos_5p043105913020105_512x8m81_2/S
+ pmos_5p043105913020105_512x8m81
Xnmos_5p043105913020109_512x8m81_0 men pmos_5p043105913020110_512x8m81_0/S nmos_5p043105913020109_512x8m81_0/S
+ pmos_5p043105913020110_512x8m81_0/S vss nmos_5p043105913020109_512x8m81
Xpmos_1p2_03_R270_512x8m81_0 vdd vdd pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D
+ pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D
+ LWL pmos_1p2_03_R270_512x8m81
Xpmos_5p043105913020103_512x8m81_0 vdd vdd pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D
+ RWL pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D
+ pmos_5p043105913020103_512x8m81
Xnmos_5p043105913020107_512x8m81_0 LWL pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D
+ vss pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D vss nmos_5p043105913020107_512x8m81
Xnmos_5p043105913020107_512x8m81_1 RWL pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D
+ vss pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D vss nmos_5p043105913020107_512x8m81
Xnmos_5p043105913020106_512x8m81_0 vss pmos_5p043105913020105_512x8m81_2/S pmos_5p043105913020110_512x8m81_0/S
+ vss nmos_5p043105913020106_512x8m81
Xpmos_5p043105913020110_512x8m81_0 vdd vdd pmos_5p043105913020105_512x8m81_2/S pmos_5p043105913020110_512x8m81_0/S
+ pmos_5p043105913020110_512x8m81
Xnmos_1p2_02_R270_512x8m81_0 nmos_5p043105913020109_512x8m81_0/S pmos_5p043105913020105_512x8m81_2/S
+ vss vss nmos_1p2_02_R270_512x8m81
X0 a_13291_624# xb a_13291_400# vss nmos_3p3 w=3.15u l=0.6u
X1 vss xc a_13291_624# vss nmos_3p3 w=3.15u l=0.6u
X2 a_13291_400# xa pmos_5p043105913020105_512x8m81_2/S vss nmos_3p3 w=3.15u l=0.6u
X3 vss nmos_5p043105913020109_512x8m81_0/S pmos_1p2_01_R270_512x8m81_0/pmos_5p043105913020108_512x8m81_0/D vss nmos_3p3 w=5u l=0.6u
X4 vss nmos_5p043105913020109_512x8m81_0/S pmos_1p2_01_R270_512x8m81_1/pmos_5p043105913020108_512x8m81_0/D vss nmos_3p3 w=5u l=0.6u
.ends

.subckt xdec8_512x8m81 RWL[0] LWL[4] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0] xa[4]
+ xa[7] xa[1] xa[3] xdec_512x8m81_3/RWL xa[0] xa[6] RWL[1] xc xdec_512x8m81_7/m2_10314_n223#
+ RWL[7] xb xa[5] xa[2] LWL[5] RWL[5] xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_16621_n223#
+ RWL[4] xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_12958_n223# xdec_512x8m81_7/m2_17376_n223#
+ xdec_512x8m81_7/m2_15110_n223# LWL[2] xdec_512x8m81_7/m2_11447_n223# LWL[3] xdec_512x8m81_7/m2_15487_n223#
+ xdec_512x8m81_7/m2_15865_n223# vdd xdec_512x8m81_7/m2_17754_n223# RWL[3] men xdec_512x8m81_7/m2_11825_n223#
+ xdec_512x8m81_7/m2_10691_n223# xdec_512x8m81_7/m2_16243_n223# xdec_512x8m81_7/m2_12202_n223#
+ xdec_512x8m81_7/m2_12580_n223# vss
Xxdec_512x8m81_0 RWL[6] xc xb xa[6] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[6] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_1 RWL[4] xc xb xa[4] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[4] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_2 RWL[2] xc xb xa[2] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[2] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_3 xdec_512x8m81_3/RWL xc xb xa[0] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[0] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_5 RWL[5] xc xb xa[5] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[5] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_4 RWL[7] xc xb xa[7] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[7] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_6 RWL[3] xc xb xa[3] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[3] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
Xxdec_512x8m81_7 RWL[1] xc xb xa[1] xdec_512x8m81_7/m2_16621_n223# xdec_512x8m81_7/m2_17754_n223#
+ xdec_512x8m81_7/m2_11825_n223# xdec_512x8m81_7/m2_12202_n223# xdec_512x8m81_7/m2_12958_n223#
+ xdec_512x8m81_7/m2_15487_n223# xdec_512x8m81_7/m2_12580_n223# xdec_512x8m81_7/m2_15110_n223#
+ xdec_512x8m81_7/m2_11069_n223# xdec_512x8m81_7/m2_15865_n223# xdec_512x8m81_7/m2_16243_n223#
+ xdec_512x8m81_7/m2_10314_n223# xdec_512x8m81_7/m2_16998_n223# xdec_512x8m81_7/m2_17376_n223#
+ men xdec_512x8m81_7/m2_11447_n223# vdd vss LWL[1] xdec_512x8m81_7/m2_10691_n223#
+ xdec_512x8m81
.ends

.subckt xdec32_468_512x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[16] RWL[15] RWL[14]
+ RWL[12] LWL[9] LWL[0] LWL[1] LWL[4] LWL[5] RWL[11] RWL[9] RWL[8] RWL[7] RWL[3] RWL[0]
+ LWL[18] LWL[15] LWL[13] LWL[12] RWL[6] LWL[27] LWL[22] LWL[21] LWL[20] LWL[19] RWL[22]
+ RWL[24] RWL[26] RWL[29] RWL[30] LWL[30] xa[2] xa[0] xa[3] xa[4] xa[5] xa[7] xb[3]
+ xb[2] xb[1] xb[0] xc xa[1] xdec8_512x8m81_2/xdec_512x8m81_3/RWL LWL[24] RWL[23]
+ xdec8_512x8m81_1/xdec_512x8m81_3/RWL RWL[20] xa[6] RWL[27] LWL[25] xdec8_512x8m81_0/xdec_512x8m81_3/RWL
+ LWL[31] RWL[1] LWL[10] RWL[21] LWL[28] LWL[16] RWL[4] RWL[25] LWL[2] RWL[13] LWL[11]
+ RWL[31] RWL[10] LWL[29] LWL[8] RWL[19] RWL[28] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11447_n223#
+ LWL[17] LWL[26] RWL[5] men LWL[14] xdec8_512x8m81_3/xdec_512x8m81_3/RWL LWL[3] LWL[23]
+ xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223# RWL[2] vdd vss xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223#
Xxdec8_512x8m81_3 RWL[16] LWL[20] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22] LWL[16]
+ xa[4] xa[7] xa[1] xa[3] xdec8_512x8m81_3/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[17]
+ xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223# RWL[23] xb[2] xa[5] xa[2] LWL[21]
+ RWL[21] xa[2] xa[3] RWL[20] xc xb[0] xa[1] xa[7] LWL[18] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11447_n223#
+ LWL[19] xa[6] xa[5] vdd xa[0] RWL[19] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
Xxdec8_512x8m81_0 RWL[24] LWL[28] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30] LWL[24]
+ xa[4] xa[7] xa[1] xa[3] xdec8_512x8m81_0/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[25]
+ xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223# RWL[31] xb[3] xa[5] xa[2] LWL[29]
+ RWL[29] xa[2] xa[3] RWL[28] xc xb[0] xa[1] xa[7] LWL[26] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11447_n223#
+ LWL[27] xa[6] xa[5] vdd xa[0] RWL[27] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
Xxdec8_512x8m81_1 RWL[0] LWL[4] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0] xa[4] xa[7]
+ xa[1] xa[3] xdec8_512x8m81_1/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[1] xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223#
+ RWL[7] xb[0] xa[5] xa[2] LWL[5] RWL[5] xa[2] xa[3] RWL[4] xc xb[0] xa[1] xa[7] LWL[2]
+ xdec8_512x8m81_3/xdec_512x8m81_7/m2_11447_n223# LWL[3] xa[6] xa[5] vdd xa[0] RWL[3]
+ men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223# xa[4] xb[2] xb[1] vss
+ xdec8_512x8m81
Xxdec8_512x8m81_2 RWL[8] LWL[12] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14] LWL[8] xa[4]
+ xa[7] xa[1] xa[3] xdec8_512x8m81_2/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[9] xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223#
+ RWL[15] xb[1] xa[5] xa[2] LWL[13] RWL[13] xa[2] xa[3] RWL[12] xc xb[0] xa[1] xa[7]
+ LWL[10] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11447_n223# LWL[11] xa[6] xa[5] vdd
+ xa[0] RWL[11] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223# xa[4] xb[2]
+ xb[1] vss xdec8_512x8m81
.ends

.subckt xdec32_512x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[16] RWL[15] RWL[14] RWL[12]
+ LWL[9] LWL[0] LWL[1] LWL[4] LWL[5] RWL[11] RWL[9] RWL[8] RWL[7] RWL[3] RWL[0] LWL[18]
+ LWL[15] LWL[13] LWL[12] RWL[6] LWL[22] LWL[21] LWL[20] LWL[19] RWL[22] RWL[24] RWL[26]
+ RWL[29] RWL[30] LWL[30] xa[2] xb[3] xb[2] xb[1] xb[0] xc xdec8_512x8m81_2/xdec_512x8m81_3/RWL
+ LWL[24] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223# RWL[23] xa[3] xdec8_512x8m81_1/xdec_512x8m81_3/RWL
+ RWL[20] xa[0] LWL[25] RWL[27] xdec8_512x8m81_0/xdec_512x8m81_3/RWL LWL[31] RWL[1]
+ LWL[10] RWL[21] LWL[28] LWL[27] LWL[16] RWL[4] RWL[25] LWL[2] RWL[13] LWL[11] RWL[31]
+ RWL[10] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11069_n223# LWL[29] xa[1] LWL[8] RWL[19]
+ RWL[28] LWL[17] LWL[26] RWL[5] xa[5] men LWL[14] xdec8_512x8m81_3/xdec_512x8m81_3/RWL
+ LWL[3] xa[6] xa[4] LWL[23] vdd RWL[2] xa[7] vss xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223#
Xxdec8_512x8m81_3 RWL[16] LWL[20] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22] LWL[16]
+ xa[4] xa[7] xa[1] xa[3] xdec8_512x8m81_3/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[17]
+ xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223# RWL[23] xb[2] xa[5] xa[2] LWL[21]
+ RWL[21] xa[2] xa[3] RWL[20] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11069_n223# xb[0]
+ xa[1] xa[7] LWL[18] xc LWL[19] xa[6] xa[5] vdd xa[0] RWL[19] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
Xxdec8_512x8m81_0 RWL[24] LWL[28] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30] LWL[24]
+ xa[4] xa[7] xa[1] xa[3] xdec8_512x8m81_0/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[25]
+ xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223# RWL[31] xb[3] xa[5] xa[2] LWL[29]
+ RWL[29] xa[2] xa[3] RWL[28] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11069_n223# xb[0]
+ xa[1] xa[7] LWL[26] xc LWL[27] xa[6] xa[5] vdd xa[0] RWL[27] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
Xxdec8_512x8m81_1 xdec8_512x8m81_1/RWL[0] LWL[4] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6]
+ LWL[0] xa[4] xa[7] xa[1] xa[3] xdec8_512x8m81_1/xdec_512x8m81_3/RWL xa[0] xa[6]
+ RWL[1] xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223# RWL[7] xb[0] xa[5] xa[2]
+ LWL[5] RWL[5] xa[2] xa[3] RWL[4] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11069_n223#
+ xb[0] xa[1] xa[7] LWL[2] xc LWL[3] xa[6] xa[5] vdd xa[0] RWL[3] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
Xxdec8_512x8m81_2 RWL[8] LWL[12] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14] LWL[8] xa[4]
+ xa[7] xa[1] xa[3] xdec8_512x8m81_2/xdec_512x8m81_3/RWL xa[0] xa[6] RWL[9] xc xdec8_512x8m81_3/xdec_512x8m81_7/m2_10314_n223#
+ RWL[15] xb[1] xa[5] xa[2] LWL[13] RWL[13] xa[2] xa[3] RWL[12] xdec8_512x8m81_3/xdec_512x8m81_7/m2_11069_n223#
+ xb[0] xa[1] xa[7] LWL[10] xc LWL[11] xa[6] xa[5] vdd xa[0] RWL[11] men xb[3] xdec8_512x8m81_3/xdec_512x8m81_7/m2_10691_n223#
+ xa[4] xb[2] xb[1] vss xdec8_512x8m81
.ends

.subckt xdec64_512x8m81 DRWL RWL[34] RWL[35] RWL[36] RWL[37] RWL[38] RWL[39] RWL[40]
+ RWL[42] RWL[43] RWL[44] RWL[45] RWL[46] RWL[48] RWL[50] RWL[53] RWL[55] RWL[57]
+ RWL[58] RWL[61] RWL[62] RWL[63] LWL[58] LWL[56] LWL[55] LWL[54] LWL[53] LWL[52]
+ LWL[51] LWL[50] LWL[46] LWL[38] LWL[36] LWL[35] LWL[34] DLWL LWL[19] LWL[20] LWL[21]
+ LWL[22] LWL[27] LWL[11] LWL[13] LWL[15] LWL[18] LWL[5] LWL[4] LWL[2] LWL[8] LWL[9]
+ LWL[6] LWL[7] LWL[29] RWL[31] RWL[30] RWL[6] RWL[4] RWL[2] RWL[0] RWL[1] RWL[3]
+ RWL[5] RWL[7] RWL[8] RWL[10] RWL[12] RWL[14] RWL[15] RWL[16] RWL[17] xb[0] xb[1]
+ xb[2] xb[3] xa[7] xa[6] xa[5] xa[4] xa[0] xa[3] xa[2] xc[0] xc[1] LWL[44] LWL[42]
+ LWL[25] LWL[40] RWL[41] LWL[23] LWL[49] RWL[60] RWL[59] LWL[62] LWL[60] RWL[29]
+ LWL[47] RWL[27] LWL[48] LWL[45] RWL[25] LWL[0] LWL[30] LWL[63] LWL[28] LWL[43] LWL[26]
+ RWL[23] LWL[24] LWL[33] LWL[3] RWL[28] LWL[61] RWL[13] RWL[26] LWL[41] LWL[32] RWL[24]
+ RWL[51] RWL[21] RWL[32] RWL[22] LWL[1] RWL[33] RWL[20] LWL[59] RWL[11] RWL[18] LWL[39]
+ xa[1] LWL[16] RWL[49] RWL[19] LWL[14] LWL[31] LWL[12] RWL[56] LWL[57] men LWL[10]
+ RWL[9] vdd LWL[37] RWL[54] vss LWL[17] RWL[52] RWL[47]
Xpmoscap_R270_512x8m81_23 LWL[3] LWL[2] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_12 RWL[25] RWL[24] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_45 LWL[37] LWL[36] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_56 RWL[45] RWL[44] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_34 LWL[59] LWL[58] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_24 LWL[1] LWL[0] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_13 RWL[23] RWL[22] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_46 LWL[35] LWL[34] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_57 RWL[43] RWL[42] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_35 LWL[57] LWL[56] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_14 RWL[21] RWL[20] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_25 LWL[31] LWL[30] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_58 RWL[41] RWL[40] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_36 LWL[55] LWL[54] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_47 RWL[63] RWL[62] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_15 RWL[19] RWL[18] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_26 LWL[29] LWL[28] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_59 RWL[39] RWL[38] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_37 LWL[53] LWL[52] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_48 RWL[61] RWL[60] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_16 LWL[17] LWL[16] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_27 LWL[27] LWL[26] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_38 LWL[51] LWL[50] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_49 RWL[59] RWL[58] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_17 LWL[15] LWL[14] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_28 LWL[25] LWL[24] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_39 LWL[49] LWL[48] vdd vdd pmoscap_R270_512x8m81
Xpmos_1p2_02_R90_512x8m81_0 vdd nmos_5p043105913020111_512x8m81_0/S nmos_5p043105913020111_512x8m81_0/S
+ DLWL vdd pmos_1p2_02_R90_512x8m81
Xnmos_5p043105913020111_512x8m81_0 vss pmos_5p043105913020101_512x8m81_1/D nmos_5p043105913020111_512x8m81_0/S
+ vss nmos_5p043105913020111_512x8m81
Xpmoscap_R270_512x8m81_18 LWL[13] LWL[12] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_29 LWL[23] LWL[22] vdd vdd pmoscap_R270_512x8m81
Xnmos_5p043105913020111_512x8m81_1 vss pmos_5p043105913020101_512x8m81_1/D pmos_5p043105913020101_512x8m81_0/S
+ vss nmos_5p043105913020111_512x8m81
Xpmos_1p2_02_R90_512x8m81_1 vdd pmos_5p043105913020101_512x8m81_0/S pmos_5p043105913020101_512x8m81_0/S
+ DRWL vdd pmos_1p2_02_R90_512x8m81
Xpmoscap_R270_512x8m81_19 LWL[11] LWL[10] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_L1_W2_R270_512x8m81_0 vdd vdd DLWL pmoscap_L1_W2_R270_512x8m81
Xpmoscap_L1_W2_R270_512x8m81_1 vdd vdd DRWL pmoscap_L1_W2_R270_512x8m81
Xpmoscap_R270_512x8m81_0 RWL[17] RWL[16] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_1 RWL[15] RWL[14] vdd vdd pmoscap_R270_512x8m81
Xpmos_1p2_01_R90_512x8m81_0 vdd nmos_5p043105913020111_512x8m81_0/S vdd pmos_5p043105913020101_512x8m81_1/D
+ pmos_1p2_01_R90_512x8m81
Xpmoscap_R270_512x8m81_2 RWL[13] RWL[12] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_3 RWL[11] RWL[10] vdd vdd pmoscap_R270_512x8m81
Xnmos_5p04310591302099_512x8m81_0 vss pmos_5p043105913020101_512x8m81_0/S DRWL vss
+ nmos_5p04310591302099_512x8m81
Xpmoscap_R270_512x8m81_4 RWL[9] RWL[8] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_5 RWL[7] RWL[6] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_6 RWL[5] RWL[4] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_7 RWL[3] RWL[2] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_8 RWL[1] RWL[0] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_9 RWL[31] RWL[30] vdd vdd pmoscap_R270_512x8m81
Xnmos_1p2_01_R270_512x8m81_0 pmos_5p043105913020101_512x8m81_1/D men vdd vss nmos_1p2_01_R270_512x8m81
Xpmos_5p043105913020101_512x8m81_0 vdd vdd pmos_5p043105913020101_512x8m81_1/D pmos_5p043105913020101_512x8m81_0/S
+ pmos_5p043105913020101_512x8m81
Xnmos_1p2_02_R90_512x8m81_0 vss nmos_5p043105913020111_512x8m81_0/S DLWL vss nmos_1p2_02_R90_512x8m81
Xpmos_5p043105913020101_512x8m81_1 vdd pmos_5p043105913020101_512x8m81_1/D vss men
+ pmos_5p043105913020101_512x8m81
Xpmoscap_R270_512x8m81_60 RWL[37] RWL[36] vdd vdd pmoscap_R270_512x8m81
Xxdec32_468_512x8m81_0 LWL[38] LWL[39] RWL[50] RWL[49] RWL[48] RWL[47] RWL[46] RWL[44]
+ LWL[41] LWL[32] LWL[33] LWL[36] LWL[37] RWL[43] RWL[41] RWL[40] RWL[39] RWL[35]
+ RWL[32] LWL[50] LWL[47] LWL[45] LWL[44] RWL[38] LWL[59] LWL[54] LWL[53] LWL[52]
+ LWL[51] RWL[54] RWL[56] RWL[58] RWL[61] RWL[62] LWL[62] xa[2] xa[0] xa[3] xa[4]
+ xa[5] xa[7] xb[3] xb[2] xb[1] xb[0] xc[1] xa[1] RWL[40] LWL[56] RWL[55] RWL[32]
+ RWL[52] xa[6] RWL[59] LWL[57] RWL[56] LWL[63] RWL[33] LWL[42] RWL[53] LWL[60] LWL[48]
+ RWL[36] RWL[57] LWL[34] RWL[45] LWL[43] RWL[63] RWL[42] LWL[61] LWL[40] RWL[51]
+ RWL[60] xc[0] LWL[49] LWL[58] RWL[37] men LWL[46] RWL[48] LWL[35] LWL[55] vdd RWL[34]
+ vdd vss vdd xdec32_468_512x8m81
Xpmoscap_R270_512x8m81_61 RWL[35] RWL[34] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_50 RWL[57] RWL[56] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_62 LWL[33] LWL[32] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_40 LWL[47] LWL[46] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_51 RWL[55] RWL[54] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_30 LWL[21] LWL[20] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_63 RWL[33] RWL[32] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_41 LWL[45] LWL[44] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_52 RWL[53] RWL[52] vdd vdd pmoscap_R270_512x8m81
Xxdec32_512x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[16] RWL[15] RWL[14] RWL[12] LWL[9]
+ LWL[0] LWL[1] LWL[4] LWL[5] RWL[11] RWL[9] RWL[8] RWL[7] RWL[3] RWL[0] LWL[18] LWL[15]
+ LWL[13] LWL[12] RWL[6] LWL[22] LWL[21] LWL[20] LWL[19] RWL[22] RWL[24] RWL[26] RWL[29]
+ RWL[30] LWL[30] xa[2] xb[3] xb[2] xb[1] xb[0] xc[0] RWL[8] LWL[24] vdd RWL[23] xa[3]
+ RWL[0] RWL[20] xa[0] LWL[25] RWL[27] RWL[24] LWL[31] RWL[1] LWL[10] RWL[21] LWL[28]
+ LWL[27] LWL[16] RWL[4] RWL[25] LWL[2] RWL[13] LWL[11] RWL[31] RWL[10] xc[1] LWL[29]
+ xa[1] LWL[8] RWL[19] RWL[28] LWL[17] LWL[26] RWL[5] xa[5] men LWL[14] RWL[16] LWL[3]
+ xa[6] xa[4] LWL[23] vdd RWL[2] xa[7] vss vdd xdec32_512x8m81
Xpmoscap_R270_512x8m81_20 LWL[9] LWL[8] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_31 LWL[19] LWL[18] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_42 LWL[43] LWL[42] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_53 RWL[51] RWL[50] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_21 LWL[7] LWL[6] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_10 RWL[29] RWL[28] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_43 LWL[41] LWL[40] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_54 RWL[49] RWL[48] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_32 LWL[63] LWL[62] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_22 LWL[5] LWL[4] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_11 RWL[27] RWL[26] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_44 LWL[39] LWL[38] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_55 RWL[47] RWL[46] vdd vdd pmoscap_R270_512x8m81
Xpmoscap_R270_512x8m81_33 LWL[61] LWL[60] vdd vdd pmoscap_R270_512x8m81
.ends

.subckt pmos_5p04310591302087_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=22.68u l=0.6u
.ends

.subckt pmos_1p2$$47815724_512x8m81 pmos_5p04310591302087_512x8m81_0/S w_n286_n141#
+ a_n31_n74# pmos_5p04310591302087_512x8m81_0/D
Xpmos_5p04310591302087_512x8m81_0 w_n286_n141# pmos_5p04310591302087_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302087_512x8m81_0/S pmos_5p04310591302087_512x8m81
.ends

.subckt nmos_5p04310591302093_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1.2u
.ends

.subckt pmos_5p04310591302094_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.89u l=0.6u
.ends

.subckt nmos_5p04310591302083_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.75u l=0.6u
.ends

.subckt nmos_5p04310591302086_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.02u l=0.6u
.ends

.subckt nmos_1p2$$48302124_512x8m81 a_n31_n74# nmos_5p04310591302086_512x8m81_0/S
+ nmos_5p04310591302086_512x8m81_0/D VSUBS
Xnmos_5p04310591302086_512x8m81_0 nmos_5p04310591302086_512x8m81_0/D a_n31_n74# nmos_5p04310591302086_512x8m81_0/S
+ VSUBS nmos_5p04310591302086_512x8m81
.ends

.subckt pmos_5p04310591302074_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1.2u
.ends

.subckt nmos_5p04310591302085_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
.ends

.subckt nmos_1p2$$48306220_512x8m81 nmos_5p04310591302085_512x8m81_0/S a_865_n74#
+ nmos_5p04310591302085_512x8m81_0/D a_641_n74# a_417_n74# a_193_n74# a_n31_n74# VSUBS
Xnmos_5p04310591302085_512x8m81_0 nmos_5p04310591302085_512x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310591302085_512x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310591302085_512x8m81
.ends

.subckt pmos_5p04310591302092_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1u
.ends

.subckt nmos_5p04310591302090_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1u
.ends

.subckt pmos_5p04310591302073_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.77u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.77u l=0.6u
.ends

.subckt pmos_1p2$$48623660_512x8m81 pmos_5p04310591302073_512x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310591302073_512x8m81_0/S
Xpmos_5p04310591302073_512x8m81_0 w_n286_n142# pmos_5p04310591302073_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302073_512x8m81_0/S a_193_n74# pmos_5p04310591302073_512x8m81
.ends

.subckt nmos_5p04310591302053_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.36u l=0.6u
.ends

.subckt nmos_1p2$$47342636_512x8m81 nmos_5p04310591302053_512x8m81_0/D nmos_5p04310591302053_512x8m81_0/S
+ a_n31_n73# VSUBS
Xnmos_5p04310591302053_512x8m81_0 nmos_5p04310591302053_512x8m81_0/D a_n31_n73# nmos_5p04310591302053_512x8m81_0/S
+ VSUBS nmos_5p04310591302053_512x8m81
.ends

.subckt pmos_5p04310591302091_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=19.5u l=0.6u
.ends

.subckt pmos_1p2$$48624684_512x8m81 pmos_5p04310591302091_512x8m81_0/S pmos_5p04310591302091_512x8m81_0/D
+ w_n286_n141# a_n31_n74#
Xpmos_5p04310591302091_512x8m81_0 w_n286_n141# pmos_5p04310591302091_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302091_512x8m81_0/S pmos_5p04310591302091_512x8m81
.ends

.subckt nmos_5p04310591302084_512x8m81 a_2464_n44# D a_2240_n44# a_3584_n44# a_2016_n44#
+ a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44# a_3808_n44#
+ a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44#
+ a_1120_n44# a_2688_n44# VSUBS
X0 S a_4256_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X1 S a_224_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X2 D a_448_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X3 D a_0_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X4 S a_2912_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X5 D a_3136_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X6 S a_672_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X7 D a_896_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X8 S a_3360_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X9 S a_2016_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X10 D a_3584_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X11 D a_2240_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X12 S a_2464_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X13 D a_2688_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X14 S a_1120_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X15 D a_1344_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X16 S a_1568_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X17 D a_1792_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X18 S a_3808_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X19 D a_4032_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
.ends

.subckt nmos_1p2$$48308268_512x8m81 nmos_5p04310591302084_512x8m81_0/a_1120_n44# nmos_5p04310591302084_512x8m81_0/a_2688_n44#
+ nmos_5p04310591302084_512x8m81_0/a_0_n44# nmos_5p04310591302084_512x8m81_0/a_2464_n44#
+ nmos_5p04310591302084_512x8m81_0/a_2240_n44# nmos_5p04310591302084_512x8m81_0/a_2016_n44#
+ nmos_5p04310591302084_512x8m81_0/a_3584_n44# nmos_5p04310591302084_512x8m81_0/a_3360_n44#
+ nmos_5p04310591302084_512x8m81_0/a_3136_n44# nmos_5p04310591302084_512x8m81_0/a_2912_n44#
+ nmos_5p04310591302084_512x8m81_0/a_896_n44# nmos_5p04310591302084_512x8m81_0/S nmos_5p04310591302084_512x8m81_0/a_672_n44#
+ nmos_5p04310591302084_512x8m81_0/a_4256_n44# nmos_5p04310591302084_512x8m81_0/a_4032_n44#
+ nmos_5p04310591302084_512x8m81_0/a_448_n44# nmos_5p04310591302084_512x8m81_0/a_3808_n44#
+ nmos_5p04310591302084_512x8m81_0/a_224_n44# nmos_5p04310591302084_512x8m81_0/a_1792_n44#
+ nmos_5p04310591302084_512x8m81_0/a_1568_n44# nmos_5p04310591302084_512x8m81_0/D
+ VSUBS nmos_5p04310591302084_512x8m81_0/a_1344_n44#
Xnmos_5p04310591302084_512x8m81_0 nmos_5p04310591302084_512x8m81_0/a_2464_n44# nmos_5p04310591302084_512x8m81_0/D
+ nmos_5p04310591302084_512x8m81_0/a_2240_n44# nmos_5p04310591302084_512x8m81_0/a_3584_n44#
+ nmos_5p04310591302084_512x8m81_0/a_2016_n44# nmos_5p04310591302084_512x8m81_0/a_3360_n44#
+ nmos_5p04310591302084_512x8m81_0/a_3136_n44# nmos_5p04310591302084_512x8m81_0/a_2912_n44#
+ nmos_5p04310591302084_512x8m81_0/a_0_n44# nmos_5p04310591302084_512x8m81_0/a_4256_n44#
+ nmos_5p04310591302084_512x8m81_0/a_4032_n44# nmos_5p04310591302084_512x8m81_0/a_3808_n44#
+ nmos_5p04310591302084_512x8m81_0/a_896_n44# nmos_5p04310591302084_512x8m81_0/a_672_n44#
+ nmos_5p04310591302084_512x8m81_0/S nmos_5p04310591302084_512x8m81_0/a_1792_n44#
+ nmos_5p04310591302084_512x8m81_0/a_448_n44# nmos_5p04310591302084_512x8m81_0/a_224_n44#
+ nmos_5p04310591302084_512x8m81_0/a_1568_n44# nmos_5p04310591302084_512x8m81_0/a_1344_n44#
+ nmos_5p04310591302084_512x8m81_0/a_1120_n44# nmos_5p04310591302084_512x8m81_0/a_2688_n44#
+ VSUBS nmos_5p04310591302084_512x8m81
.ends

.subckt pmos_5p04310591302089_512x8m81 a_2464_n44# w_n208_n120# D a_2240_n44# a_3584_n44#
+ a_2016_n44# a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44#
+ a_3808_n44# a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44#
+ a_1344_n44# a_1120_n44# a_2688_n44#
X0 D a_4032_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X1 S a_4256_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X2 S a_224_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X3 D a_448_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X4 D a_0_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X5 S a_2912_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X6 D a_3136_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X7 S a_672_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X8 D a_896_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X9 S a_3360_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X10 S a_2016_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X11 D a_3584_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X12 D a_2240_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X13 S a_2464_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X14 D a_2688_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X15 S a_1120_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X16 D a_1344_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X17 S a_1568_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X18 D a_1792_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X19 S a_3808_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
.ends

.subckt pmos_5p04310591302088_512x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
.ends

.subckt nmos_5p04310591302081_512x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
.ends

.subckt pmos_5p04310591302082_512x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
.ends

.subckt pmos_5p04310591302080_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310591302078_512x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_5p04310591302079_512x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X6 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310591302076_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310591302077_512x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
.ends

.subckt nmos_5p04310591302075_512x8m81 D a_2016_n44# a_0_n44# a_896_n44# a_672_n44#
+ S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X5 S a_2016_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X6 S a_1120_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X7 D a_1344_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X8 S a_1568_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X9 D a_1792_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
.ends

.subckt wen_v2_512x8m81 IGWEN clk wen GWE vss vdd
Xpmos_1p2$$202586156_512x8m81_0 pmos_5p04310591302041_512x8m81_1/D vdd pmos_5p04310591302014_512x8m81_2/S
+ vdd pmos_1p2$$202586156_512x8m81
Xpmos_5p04310591302014_512x8m81_0 vdd vdd pmos_5p04310591302079_512x8m81_0/D nmos_5p0431059130208_512x8m81_1/D
+ pmos_5p04310591302014_512x8m81
Xnmos_5p04310591302081_512x8m81_0 pmos_5p04310591302079_512x8m81_0/D nmos_5p0431059130208_512x8m81_1/S
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S vss nmos_5p0431059130208_512x8m81_1/S
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S
+ vss nmos_5p04310591302081_512x8m81
Xpmos_5p04310591302082_512x8m81_0 vdd pmos_5p04310591302082_512x8m81_0/D wen wen wen
+ vdd wen wen wen pmos_5p04310591302082_512x8m81
Xpmos_5p04310591302014_512x8m81_1 vdd nmos_5p0431059130208_512x8m81_3/D clk vdd pmos_5p04310591302014_512x8m81
Xpmos_1p2$$202587180_512x8m81_0 nmos_5p0431059130208_512x8m81_2/S vdd nmos_5p0431059130208_512x8m81_4/D
+ pmos_5p04310591302041_512x8m81_1/S pmos_1p2$$202587180_512x8m81
Xpmos_5p04310591302014_512x8m81_2 vdd vdd pmos_5p04310591302041_512x8m81_1/S pmos_5p04310591302014_512x8m81_2/S
+ pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302014_512x8m81_3 vdd vdd wen nmos_5p0431059130208_512x8m81_2/S pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302014_512x8m81_4 vdd nmos_5p0431059130208_512x8m81_4/D nmos_5p0431059130208_512x8m81_3/D
+ vdd pmos_5p04310591302014_512x8m81
Xpmos_5p04310591302041_512x8m81_0 vdd nmos_5p0431059130208_512x8m81_1/D nmos_5p0431059130208_512x8m81_4/D
+ nmos_5p0431059130208_512x8m81_1/S pmos_5p04310591302041_512x8m81
Xpmos_5p04310591302080_512x8m81_0 vdd pmos_5p04310591302080_512x8m81_0/D pmos_5p04310591302014_512x8m81_2/S
+ vdd pmos_5p04310591302014_512x8m81_2/S pmos_5p04310591302080_512x8m81
Xpmos_5p04310591302041_512x8m81_1 vdd pmos_5p04310591302041_512x8m81_1/D nmos_5p0431059130208_512x8m81_3/D
+ pmos_5p04310591302041_512x8m81_1/S pmos_5p04310591302041_512x8m81
Xnmos_5p0431059130208_512x8m81_0 vss pmos_5p04310591302079_512x8m81_0/D nmos_5p0431059130208_512x8m81_1/D
+ vss nmos_5p0431059130208_512x8m81
Xnmos_5p04310591302010_512x8m81_0 pmos_5p04310591302041_512x8m81_1/S nmos_5p0431059130208_512x8m81_3/D
+ nmos_5p0431059130208_512x8m81_2/S vss nmos_5p04310591302010_512x8m81
Xnmos_5p0431059130208_512x8m81_1 nmos_5p0431059130208_512x8m81_1/D nmos_5p0431059130208_512x8m81_3/D
+ nmos_5p0431059130208_512x8m81_1/S vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_2 vss wen nmos_5p0431059130208_512x8m81_2/S vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_3 nmos_5p0431059130208_512x8m81_3/D clk vss vss nmos_5p0431059130208_512x8m81
Xnmos_5p0431059130208_512x8m81_4 nmos_5p0431059130208_512x8m81_4/D nmos_5p0431059130208_512x8m81_3/D
+ vss vss nmos_5p0431059130208_512x8m81
Xpmos_5p04310591302020_512x8m81_0 vdd pmos_5p04310591302080_512x8m81_0/D nmos_5p0431059130208_512x8m81_3/D
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_3/D pmos_5p04310591302020_512x8m81
Xnmos_1p2$$202595372_512x8m81_0 vss pmos_5p04310591302041_512x8m81_1/S pmos_5p04310591302014_512x8m81_2/S
+ vss nmos_1p2$$202595372_512x8m81
Xnmos_1p2$$202595372_512x8m81_1 pmos_5p04310591302041_512x8m81_1/D nmos_5p0431059130208_512x8m81_4/D
+ pmos_5p04310591302041_512x8m81_1/S vss nmos_1p2$$202595372_512x8m81
Xnmos_5p04310591302078_512x8m81_0 pmos_5p04310591302082_512x8m81_0/D wen vss wen wen
+ vss nmos_5p04310591302078_512x8m81
Xnmos_5p04310591302039_512x8m81_0 pmos_5p04310591302080_512x8m81_0/D nmos_5p0431059130208_512x8m81_4/D
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_4/D vss nmos_5p04310591302039_512x8m81
Xpmos_5p04310591302079_512x8m81_0 vdd pmos_5p04310591302079_512x8m81_0/D nmos_5p0431059130208_512x8m81_1/S
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S vdd nmos_5p0431059130208_512x8m81_1/S
+ nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S nmos_5p0431059130208_512x8m81_1/S
+ pmos_5p04310591302079_512x8m81
Xnmos_1p2$$202596396_512x8m81_0 vss pmos_5p04310591302014_512x8m81_2/S pmos_5p04310591302041_512x8m81_1/D
+ vss nmos_1p2$$202596396_512x8m81
Xnmos_5p04310591302076_512x8m81_0 pmos_5p04310591302080_512x8m81_0/D pmos_5p04310591302014_512x8m81_2/S
+ vss pmos_5p04310591302014_512x8m81_2/S vss nmos_5p04310591302076_512x8m81
Xpmos_5p04310591302077_512x8m81_0 vdd GWE pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D vdd pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302077_512x8m81
Xpmos_5p04310591302077_512x8m81_1 vdd IGWEN pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D vdd pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302077_512x8m81
Xnmos_5p04310591302075_512x8m81_0 GWE pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D vss pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D
+ pmos_5p04310591302079_512x8m81_0/D pmos_5p04310591302079_512x8m81_0/D vss nmos_5p04310591302075_512x8m81
Xnmos_5p04310591302075_512x8m81_1 IGWEN pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D vss pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D
+ pmos_5p04310591302082_512x8m81_0/D pmos_5p04310591302082_512x8m81_0/D vss nmos_5p04310591302075_512x8m81
.ends

.subckt pmos_1p2$$47330348_512x8m81 pmos_5p04310591302041_512x8m81_0/S a_n31_n73#
+ pmos_5p04310591302041_512x8m81_0/D w_n286_n141#
Xpmos_5p04310591302041_512x8m81_0 w_n286_n141# pmos_5p04310591302041_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302041_512x8m81_0/S pmos_5p04310591302041_512x8m81
.ends

.subckt nmos_1p2$$48629804_512x8m81 nmos_5p04310591302039_512x8m81_0/D a_193_n73#
+ a_n31_n73# nmos_5p04310591302039_512x8m81_0/S VSUBS
Xnmos_5p04310591302039_512x8m81_0 nmos_5p04310591302039_512x8m81_0/D a_n31_n73# nmos_5p04310591302039_512x8m81_0/S
+ a_193_n73# VSUBS nmos_5p04310591302039_512x8m81
.ends

.subckt gen_512x8_512x8m81 tblhl IGWEN clk WEN GWE pmos_5p04310591302088_512x8m81_0/D
+ cen men VDD VSS
Xpmos_1p2$$47815724_512x8m81_7 pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ VDD pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S VDD pmos_1p2$$47815724_512x8m81
Xnmos_5p04310591302093_512x8m81_0 pmos_5p04310591302074_512x8m81_0/D clk VSS VSS nmos_5p04310591302093_512x8m81
Xpmos_5p04310591302094_512x8m81_0 VDD pmos_5p04310591302094_512x8m81_0/D pmos_5p04310591302092_512x8m81_0/D
+ VDD pmos_5p04310591302094_512x8m81
Xnmos_5p04310591302083_512x8m81_0 pmos_5p04310591302094_512x8m81_0/D pmos_5p04310591302092_512x8m81_0/D
+ VSS VSS nmos_5p04310591302083_512x8m81
Xnmos_1p2$$48302124_512x8m81_0 pmos_5p04310591302094_512x8m81_0/D VSS pmos_1p2$$48623660_512x8m81_0/pmos_5p04310591302073_512x8m81_0/D
+ VSS nmos_1p2$$48302124_512x8m81
Xnmos_5p04310591302093_512x8m81_1 pmos_5p04310591302074_512x8m81_1/D pmos_5p04310591302074_512x8m81_0/D
+ VSS VSS nmos_5p04310591302093_512x8m81
Xpmos_5p04310591302074_512x8m81_0 VDD pmos_5p04310591302074_512x8m81_0/D clk VDD pmos_5p04310591302074_512x8m81
Xpmos_5p04310591302074_512x8m81_1 VDD pmos_5p04310591302074_512x8m81_1/D pmos_5p04310591302074_512x8m81_0/D
+ VDD pmos_5p04310591302074_512x8m81
Xpmos_1p2$$46285868_512x8m81_0 VDD VDD nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S
+ nmos_1p2$$46563372_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D pmos_1p2$$46285868_512x8m81
Xnmos_1p2$$48306220_512x8m81_0 VSS pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_5p04310591302088_512x8m81_0/D pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S VSS nmos_1p2$$48306220_512x8m81
Xnmos_1p2$$46563372_512x8m81_0 nmos_1p2$$46563372_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D
+ nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S VSS VSS nmos_1p2$$46563372_512x8m81
Xpmos_1p2$$46285868_512x8m81_1 nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S
+ VDD nmos_1p2$$46563372_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D cen pmos_1p2$$46285868_512x8m81
Xnmos_1p2$$46563372_512x8m81_1 VSS pmos_5p04310591302051_512x8m81_0/D pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ VSS nmos_1p2$$46563372_512x8m81
Xnmos_1p2$$46563372_512x8m81_2 pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ nmos_1p2$$46563372_512x8m81_0/nmos_5p0431059130208_512x8m81_0/D nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S
+ VSS nmos_1p2$$46563372_512x8m81
Xpmos_5p04310591302092_512x8m81_0 VDD pmos_5p04310591302092_512x8m81_0/D pmos_5p04310591302074_512x8m81_1/D
+ VDD pmos_5p04310591302092_512x8m81
Xpmos_1p2$$46273580_512x8m81_0 VDD pmos_5p04310591302051_512x8m81_0/D pmos_5p04310591302051_512x8m81_0/D
+ pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D VDD pmos_1p2$$46273580_512x8m81
Xnmos_5p04310591302090_512x8m81_0 pmos_5p04310591302092_512x8m81_0/D pmos_5p04310591302074_512x8m81_1/D
+ VSS VSS nmos_5p04310591302090_512x8m81
Xnmos_1p2$$46551084_512x8m81_0 cen nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S
+ nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S VSS nmos_1p2$$46551084_512x8m81
Xpmos_1p2$$48623660_512x8m81_0 pmos_1p2$$48623660_512x8m81_0/pmos_5p04310591302073_512x8m81_0/D
+ pmos_5p04310591302094_512x8m81_0/D VDD pmos_5p04310591302094_512x8m81_0/D VDD pmos_1p2$$48623660_512x8m81
Xpmos_5p04310591302051_512x8m81_0 VDD pmos_5p04310591302051_512x8m81_0/D nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S
+ VDD nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S pmos_5p04310591302051_512x8m81
Xnmos_1p2$$47342636_512x8m81_0 nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S
+ VSS clk VSS nmos_1p2$$47342636_512x8m81
Xnmos_1p2$$47342636_512x8m81_1 VSS nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S
+ men VSS nmos_1p2$$47342636_512x8m81
Xpmos_1p2$$48624684_512x8m81_0 VDD pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S
+ VDD pmos_5p04310591302051_512x8m81_0/D pmos_1p2$$48624684_512x8m81
Xnmos_1p2$$48308268_512x8m81_0 pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ VSS pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D men VSS pmos_5p04310591302088_512x8m81_0/D
+ nmos_1p2$$48308268_512x8m81
Xpmos_5p04310591302089_512x8m81_0 pmos_5p04310591302088_512x8m81_0/D VDD men pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D VDD pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D pmos_5p04310591302088_512x8m81_0/D
+ pmos_5p04310591302089_512x8m81
Xpmos_1p2$$48624684_512x8m81_1 VDD pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S
+ VDD pmos_1p2$$48623660_512x8m81_0/pmos_5p04310591302073_512x8m81_0/D pmos_1p2$$48624684_512x8m81
Xpmos_1p2$$48624684_512x8m81_2 pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S
+ VDD VDD clk pmos_1p2$$48624684_512x8m81
Xpmos_5p04310591302088_512x8m81_0 VDD pmos_5p04310591302088_512x8m81_0/D pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S VDD pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_5p04310591302088_512x8m81
Xpmos_1p2$$47815724_512x8m81_0 pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S
+ VDD tblhl VDD pmos_1p2$$47815724_512x8m81
Xwen_v2_512x8m81_0 wen_v2_512x8m81_0/IGWEN clk wen_v2_512x8m81_0/wen wen_v2_512x8m81_0/GWE
+ VSS VDD wen_v2_512x8m81
Xpmos_1p2$$47815724_512x8m81_1 VDD VDD pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81
Xpmos_1p2$$47815724_512x8m81_2 VDD VDD tblhl pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81
Xpmos_1p2$$47815724_512x8m81_3 pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S
+ VDD pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S VDD pmos_1p2$$47815724_512x8m81
Xpmos_1p2$$47815724_512x8m81_4 VDD VDD pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81
Xpmos_1p2$$47815724_512x8m81_5 VDD VDD pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S
+ pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$47815724_512x8m81
Xpmos_1p2$$47330348_512x8m81_0 nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S
+ nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S pmos_1p2$$46273580_512x8m81_0/pmos_5p0431059130203_512x8m81_0/D
+ VDD pmos_1p2$$47330348_512x8m81
Xpmos_1p2$$47815724_512x8m81_6 pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S
+ VDD pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S VDD pmos_1p2$$47815724_512x8m81
Xnmos_1p2$$48629804_512x8m81_0 pmos_5p04310591302051_512x8m81_0/D nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S
+ nmos_1p2$$46563372_512x8m81_2/nmos_5p0431059130208_512x8m81_0/S VSS VSS nmos_1p2$$48629804_512x8m81
X0 VSS pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S a_11293_484# VSS nmos_6p0 w=18.145u l=0.6u
X1 a_9646_262# pmos_1p2$$48623660_512x8m81_0/pmos_5p04310591302073_512x8m81_0/D VSS VSS nmos_6p0 w=22.68u l=0.6u
X2 pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S a_10845_484# VSS nmos_6p0 w=18.145u l=0.6u
X3 a_12578_3205# tblhl pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S VSS nmos_6p0 w=4.54u l=0.6u
X4 pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S pmos_5p04310591302051_512x8m81_0/D a_9870_262# VSS nmos_6p0 w=22.68u l=0.6u
X5 a_11293_484# pmos_1p2$$48624684_512x8m81_2/pmos_5p04310591302091_512x8m81_0/S pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S VSS nmos_6p0 w=18.145u l=0.6u
X6 a_12130_3205# pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S VSS VSS nmos_6p0 w=4.54u l=0.6u
X7 a_10845_484# pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S VSS VSS nmos_6p0 w=18.145u l=0.6u
X8 pmos_1p2$$47815724_512x8m81_3/pmos_5p04310591302087_512x8m81_0/S tblhl a_12130_3205# VSS nmos_6p0 w=4.54u l=0.6u
X9 nmos_1p2$$47342636_512x8m81_1/nmos_5p04310591302053_512x8m81_0/S clk a_5174_6131# VDD pmos_6p0 w=2.28u l=0.595u
X10 VSS pmos_1p2$$47815724_512x8m81_7/pmos_5p04310591302087_512x8m81_0/S a_12578_3205# VSS nmos_6p0 w=4.54u l=0.6u
X11 a_9870_262# clk a_9646_262# VSS nmos_6p0 w=22.68u l=0.6u
X12 a_5174_6131# men VDD VDD pmos_6p0 w=2.28u l=0.595u
.ends

.subckt nmos_5p04310591302054_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=9.08u l=0.6u
.ends

.subckt pmos_5p04310591302055_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=20u l=0.6u
.ends

.subckt ypredec1_ys_512x8m81 a_254_2184# nmos_5p04310591302054_512x8m81_1/D nmos_5p04310591302054_512x8m81_3/D
+ nmos_5p04310591302054_512x8m81_2/S pmos_5p04310591302055_512x8m81_3/S pmos_5p04310591302055_512x8m81_3/D
+ VSUBS pmos_5p04310591302055_512x8m81_1/S
Xnmos_5p04310591302054_512x8m81_0 pmos_5p04310591302055_512x8m81_3/S pmos_5p04310591302055_512x8m81_0/D
+ nmos_5p04310591302054_512x8m81_1/D VSUBS nmos_5p04310591302054_512x8m81
Xpmos_5p04310591302055_512x8m81_0 pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81_0/D
+ a_254_2184# pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81
Xnmos_5p04310591302054_512x8m81_1 nmos_5p04310591302054_512x8m81_1/D pmos_5p04310591302055_512x8m81_0/D
+ pmos_5p04310591302055_512x8m81_1/S VSUBS nmos_5p04310591302054_512x8m81
Xpmos_5p04310591302055_512x8m81_1 pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81_3/D
+ pmos_5p04310591302055_512x8m81_0/D pmos_5p04310591302055_512x8m81_1/S pmos_5p04310591302055_512x8m81
Xnmos_5p04310591302054_512x8m81_2 pmos_5p04310591302055_512x8m81_0/D a_254_2184# nmos_5p04310591302054_512x8m81_2/S
+ VSUBS nmos_5p04310591302054_512x8m81
Xpmos_5p04310591302055_512x8m81_2 pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81_3/S
+ pmos_5p04310591302055_512x8m81_0/D pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81
Xnmos_5p04310591302054_512x8m81_3 nmos_5p04310591302054_512x8m81_3/D pmos_5p04310591302055_512x8m81_0/D
+ pmos_5p04310591302055_512x8m81_3/S VSUBS nmos_5p04310591302054_512x8m81
Xpmos_5p04310591302055_512x8m81_3 pmos_5p04310591302055_512x8m81_3/D pmos_5p04310591302055_512x8m81_3/D
+ pmos_5p04310591302055_512x8m81_0/D pmos_5p04310591302055_512x8m81_3/S pmos_5p04310591302055_512x8m81
.ends

.subckt pmos_5p04310591302058_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$47331372_512x8m81 pmos_5p04310591302058_512x8m81_0/S a_n30_n74#
+ pmos_5p04310591302058_512x8m81_0/D w_n286_n142# a_194_n74#
Xpmos_5p04310591302058_512x8m81_0 w_n286_n142# pmos_5p04310591302058_512x8m81_0/D
+ a_n30_n74# pmos_5p04310591302058_512x8m81_0/S a_194_n74# pmos_5p04310591302058_512x8m81
.ends

.subckt nmos_1p2_157_512x8m81 nmos_5p04310591302010_512x8m81_0/D a_n31_n74# nmos_5p04310591302010_512x8m81_0/S
+ VSUBS
Xnmos_5p04310591302010_512x8m81_0 nmos_5p04310591302010_512x8m81_0/D a_n31_n74# nmos_5p04310591302010_512x8m81_0/S
+ VSUBS nmos_5p04310591302010_512x8m81
.ends

.subckt pmos_1p2_161_512x8m81 pmos_5p04310591302041_512x8m81_0/S a_n31_191# pmos_5p04310591302041_512x8m81_0/D
+ w_n286_n141#
Xpmos_5p04310591302041_512x8m81_0 w_n286_n141# pmos_5p04310591302041_512x8m81_0/D
+ a_n31_191# pmos_5p04310591302041_512x8m81_0/S pmos_5p04310591302041_512x8m81
.ends

.subckt pmos_1p2_160_512x8m81 a_n31_n74# pmos_5p04310591302014_512x8m81_0/S w_n286_n142#
+ pmos_5p04310591302014_512x8m81_0/D
Xpmos_5p04310591302014_512x8m81_0 w_n286_n142# pmos_5p04310591302014_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302014_512x8m81_0/S pmos_5p04310591302014_512x8m81
.ends

.subckt nmos_5p04310591302059_512x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.82u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.82u l=0.6u
.ends

.subckt nmos_1p2$$47329324_512x8m81 a_194_n74# nmos_5p04310591302059_512x8m81_0/S
+ nmos_5p04310591302059_512x8m81_0/D a_n30_n74# VSUBS
Xnmos_5p04310591302059_512x8m81_0 nmos_5p04310591302059_512x8m81_0/D a_n30_n74# nmos_5p04310591302059_512x8m81_0/S
+ a_194_n74# VSUBS nmos_5p04310591302059_512x8m81
.ends

.subckt alatch_512x8m81 enb en ab a vss vdd
Xpmos_1p2$$47331372_512x8m81_0 vdd nmos_5p0431059130208_512x8m81_1/S ab vdd nmos_5p0431059130208_512x8m81_1/S
+ pmos_1p2$$47331372_512x8m81
Xnmos_1p2_157_512x8m81_0 a en nmos_5p0431059130208_512x8m81_1/S vss nmos_1p2_157_512x8m81
Xpmos_1p2_161_512x8m81_0 nmos_5p0431059130208_512x8m81_1/S en nmos_5p0431059130208_512x8m81_1/D
+ vdd pmos_1p2_161_512x8m81
Xnmos_5p0431059130208_512x8m81_0 vss ab nmos_5p0431059130208_512x8m81_1/D vss nmos_5p0431059130208_512x8m81
Xpmos_1p2_161_512x8m81_1 nmos_5p0431059130208_512x8m81_1/D ab vdd vdd pmos_1p2_161_512x8m81
Xnmos_5p0431059130208_512x8m81_1 nmos_5p0431059130208_512x8m81_1/D enb nmos_5p0431059130208_512x8m81_1/S
+ vss nmos_5p0431059130208_512x8m81
Xpmos_1p2_160_512x8m81_0 enb nmos_5p0431059130208_512x8m81_1/S vdd a pmos_1p2_160_512x8m81
Xnmos_1p2$$47329324_512x8m81_0 nmos_5p0431059130208_512x8m81_1/S vss ab nmos_5p0431059130208_512x8m81_1/S
+ vss nmos_1p2$$47329324_512x8m81
.ends

.subckt nmos_5p04310591302057_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=4.54u l=0.6u
.ends

.subckt nmos_1p2$$47514668_512x8m81 nmos_5p04310591302057_512x8m81_0/D a_n30_n73#
+ nmos_5p04310591302057_512x8m81_0/S VSUBS
Xnmos_5p04310591302057_512x8m81_0 nmos_5p04310591302057_512x8m81_0/D a_n30_n73# nmos_5p04310591302057_512x8m81_0/S
+ VSUBS nmos_5p04310591302057_512x8m81
.ends

.subckt ypredec1_bot_512x8m81 m1_n14_3279# m1_n14_2674# alatch_512x8m81_0/a m1_n14_2876#
+ alatch_512x8m81_0/en m1_n14_3078# m1_n14_3481# pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ alatch_512x8m81_0/vdd m1_n14_2472# pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ alatch_512x8m81_0/enb pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ alatch_512x8m81_0/vss
Xalatch_512x8m81_0 alatch_512x8m81_0/enb alatch_512x8m81_0/en alatch_512x8m81_0/ab
+ alatch_512x8m81_0/a alatch_512x8m81_0/vss alatch_512x8m81_0/vdd alatch_512x8m81
Xpmos_1p2$$46887980_512x8m81_0 pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S pmos_1p2$$46887980_512x8m81
Xpmos_1p2$$46887980_512x8m81_1 pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ alatch_512x8m81_0/ab pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S pmos_1p2$$46887980_512x8m81
Xnmos_1p2$$47514668_512x8m81_0 pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D alatch_512x8m81_0/vss
+ alatch_512x8m81_0/vss nmos_1p2$$47514668_512x8m81
Xnmos_1p2$$47514668_512x8m81_1 pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ alatch_512x8m81_0/ab alatch_512x8m81_0/vss alatch_512x8m81_0/vss nmos_1p2$$47514668_512x8m81
.ends

.subckt pmos_5p04310591302061_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.77u l=0.6u
.ends

.subckt pmos_1p2$$47820844_512x8m81 pmos_5p04310591302061_512x8m81_0/D w_n286_n141#
+ a_n30_n74# pmos_5p04310591302061_512x8m81_0/S
Xpmos_5p04310591302061_512x8m81_0 w_n286_n141# pmos_5p04310591302061_512x8m81_0/D
+ a_n30_n74# pmos_5p04310591302061_512x8m81_0/S pmos_5p04310591302061_512x8m81
.ends

.subckt pmos_5p04310591302060_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$47821868_512x8m81 pmos_5p04310591302060_512x8m81_0/S pmos_5p04310591302060_512x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310591302060_512x8m81_0 w_n286_n142# pmos_5p04310591302060_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302060_512x8m81_0/S pmos_5p04310591302060_512x8m81
.ends

.subckt ypredec1_xa_512x8m81 m1_n58_n4290# m1_n58_n4895# m1_n58_n5097# m3_n1_n7124#
+ a_644_n6680# m1_n58_n4492# m1_n58_n4088# a_421_n4311# a_n1_81# a_197_n5120# m1_n58_n4694#
+ M3_M2$$47819820_512x8m81_0/VSUBS pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
Xnmos_1p2$$46551084_512x8m81_0 pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D M3_M2$$47819820_512x8m81_0/VSUBS
+ M3_M2$$47819820_512x8m81_0/VSUBS nmos_1p2$$46551084_512x8m81
Xnmos_1p2$$46551084_512x8m81_2 pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D M3_M2$$47819820_512x8m81_0/VSUBS
+ M3_M2$$47819820_512x8m81_0/VSUBS nmos_1p2$$46551084_512x8m81
Xnmos_1p2$$46551084_512x8m81_1 M3_M2$$47819820_512x8m81_0/VSUBS pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D
+ pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S M3_M2$$47819820_512x8m81_0/VSUBS
+ nmos_1p2$$46551084_512x8m81
Xpmos_1p2$$47820844_512x8m81_0 pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47820844_512x8m81
Xpmos_1p2$$47820844_512x8m81_1 pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47820844_512x8m81
Xpmos_1p2$$47820844_512x8m81_2 pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D
+ pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S pmos_1p2$$47820844_512x8m81
Xpmos_1p2$$47821868_512x8m81_0 pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ a_197_n5120# pmos_1p2$$47821868_512x8m81
Xpmos_1p2$$47821868_512x8m81_1 pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ a_421_n4311# pmos_1p2$$47821868_512x8m81
Xpmos_1p2$$47821868_512x8m81_2 pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ a_644_n6680# pmos_1p2$$47821868_512x8m81
X0 pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/D a_644_n6680# a_542_n6607# M3_M2$$47819820_512x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X1 a_318_n6607# a_197_n5120# M3_M2$$47819820_512x8m81_0/VSUBS M3_M2$$47819820_512x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X2 a_542_n6607# a_421_n4311# a_318_n6607# M3_M2$$47819820_512x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
.ends

.subckt ypredec1_xax8_512x8m81 ypredec1_xa_512x8m81_4/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_3/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_7/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_2/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ a_527_2758# ypredec1_xa_512x8m81_6/a_n1_81# a_6100_2150# ypredec1_xa_512x8m81_6/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_1/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ a_975_1949# ypredec1_xa_512x8m81_3/a_n1_81# a_6324_2352# ypredec1_xa_512x8m81_0/a_n1_81#
+ ypredec1_xa_512x8m81_5/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_0/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81_7/a_n1_81# a_751_2554# a_303_2957# VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
Xypredec1_xa_512x8m81_0 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_512x8m81_0/a_n1_81# a_751_2554# a_6324_2352#
+ VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_0/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_1 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS a_751_2554# a_6324_2352# VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_1/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_2 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS a_751_2554# a_6324_2352# VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_2/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_3 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_512x8m81_3/a_n1_81# a_751_2554# a_6324_2352#
+ VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_3/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_4 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_512x8m81_4/a_n1_81# a_975_1949# a_6324_2352#
+ VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_4/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_5 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_6324_2352# a_751_2554#
+ a_303_2957# a_6100_2150# VSUBS a_975_1949# a_6324_2352# VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_5/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_6 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_6100_2150# ypredec1_xa_512x8m81_6/a_n1_81# a_975_1949# a_6324_2352#
+ VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_6/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
Xypredec1_xa_512x8m81_7 a_527_2758# a_6100_2150# a_975_1949# VSUBS a_303_2957# a_751_2554#
+ a_303_2957# a_527_2758# ypredec1_xa_512x8m81_7/a_n1_81# a_975_1949# a_6324_2352#
+ VSUBS ypredec1_xa_512x8m81_7/pmos_1p2$$47821868_512x8m81_2/pmos_5p04310591302060_512x8m81_0/S
+ ypredec1_xa_512x8m81_7/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xa_512x8m81
.ends

.subckt nmos_5p04310591302056_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.91u l=0.6u
.ends

.subckt pmos_5p04310591302062_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$47109164_512x8m81 a_n31_341# pmos_5p04310591302062_512x8m81_0/D
+ pmos_5p04310591302062_512x8m81_0/w_n208_n120# pmos_5p04310591302062_512x8m81_0/S
+ a_193_341#
Xpmos_5p04310591302062_512x8m81_0 pmos_5p04310591302062_512x8m81_0/w_n208_n120# pmos_5p04310591302062_512x8m81_0/D
+ a_n31_341# pmos_5p04310591302062_512x8m81_0/S a_193_341# pmos_5p04310591302062_512x8m81
.ends

.subckt ypredec1_512x8m81 ly[5] ly[4] ly[7] ly[3] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120#
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS
Xypredec1_ys_512x8m81_4 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_5/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[0] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[0] ypredec1_ys_512x8m81
Xypredec1_bot_512x8m81_2 ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ A[1] ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/enb ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81
Xypredec1_ys_512x8m81_5 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_1/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[1] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[1] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_6 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_4/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[2] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[2] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_7 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_2/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[5] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[5] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_8 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_7/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[6] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[6] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_10 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_1/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[1] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[1] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_9 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_3/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[7] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[7] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_11 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_4/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[2] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[2] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_12 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_0/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[3] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[3] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_13 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_6/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[4] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[4] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_14 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_5/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ry[0] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ry[0] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_15 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_3/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[7] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[7] ypredec1_ys_512x8m81
Xnmos_1p2$$47342636_512x8m81_0 M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81_2/alatch_512x8m81_0/enb
+ nmos_5p04310591302056_512x8m81_1/D M1_NWELL13_512x8m81_0/VSUBS nmos_1p2$$47342636_512x8m81
Xypredec1_xax8_512x8m81_0 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_4/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_3/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_7/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_2/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_6/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_1/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_5/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_0/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ ypredec1_xax8_512x8m81
Xnmos_5p04310591302056_512x8m81_0 M1_NWELL13_512x8m81_0/VSUBS clk nmos_5p04310591302056_512x8m81_1/D
+ M1_NWELL13_512x8m81_0/VSUBS nmos_5p04310591302056_512x8m81
Xnmos_5p04310591302056_512x8m81_1 nmos_5p04310591302056_512x8m81_1/D men M1_NWELL13_512x8m81_0/VSUBS
+ M1_NWELL13_512x8m81_0/VSUBS nmos_5p04310591302056_512x8m81
Xypredec1_ys_512x8m81_0 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_0/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[3] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[3] ypredec1_ys_512x8m81
Xypredec1_ys_512x8m81_1 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_6/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[4] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[4] ypredec1_ys_512x8m81
Xypredec1_bot_512x8m81_0 ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ A[0] ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/enb ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81
Xypredec1_ys_512x8m81_2 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_2/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[5] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[5] ypredec1_ys_512x8m81
Xpmos_1p2$$47109164_512x8m81_0 nmos_5p04310591302056_512x8m81_1/D ypredec1_bot_512x8m81_2/alatch_512x8m81_0/enb
+ pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120# pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S
+ nmos_5p04310591302056_512x8m81_1/D pmos_1p2$$47109164_512x8m81
Xypredec1_bot_512x8m81_1 ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ A[2] ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd ypredec1_bot_512x8m81_0/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_1/pmos_1p2$$46887980_512x8m81_0/pmos_5p0431059130204_512x8m81_0/D
+ ypredec1_bot_512x8m81_2/alatch_512x8m81_0/enb ypredec1_bot_512x8m81_2/pmos_1p2$$46887980_512x8m81_1/pmos_5p0431059130204_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS ypredec1_bot_512x8m81
Xypredec1_ys_512x8m81_3 ypredec1_xax8_512x8m81_0/ypredec1_xa_512x8m81_7/pmos_1p2$$47820844_512x8m81_2/pmos_5p04310591302061_512x8m81_0/S
+ M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS M1_NWELL13_512x8m81_0/VSUBS
+ ly[6] ypredec1_ys_512x8m81_9/pmos_5p04310591302055_512x8m81_3/D M1_NWELL13_512x8m81_0/VSUBS
+ ly[6] ypredec1_ys_512x8m81
X0 a_7843_267# clk nmos_5p04310591302056_512x8m81_1/D pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X1 nmos_5p04310591302056_512x8m81_1/D clk a_7395_267# pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X2 a_7395_267# men pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X3 pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S men a_7843_267# pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/S pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310591302072_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.43u l=0.6u
.ends

.subckt pmos_1p2$$47512620_512x8m81 pmos_5p04310591302072_512x8m81_0/S a_n30_n74#
+ pmos_5p04310591302072_512x8m81_0/D w_n286_n142#
Xpmos_5p04310591302072_512x8m81_0 w_n286_n142# pmos_5p04310591302072_512x8m81_0/D
+ a_n30_n74# pmos_5p04310591302072_512x8m81_0/S pmos_5p04310591302072_512x8m81
.ends

.subckt pmos_5p04310591302068_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt pmos_1p2$$47513644_512x8m81 a_n30_n74# pmos_5p04310591302068_512x8m81_0/S
+ w_n286_n141# pmos_5p04310591302068_512x8m81_0/D
Xpmos_5p04310591302068_512x8m81_0 w_n286_n141# pmos_5p04310591302068_512x8m81_0/D
+ a_n30_n74# pmos_5p04310591302068_512x8m81_0/S pmos_5p04310591302068_512x8m81
.ends

.subckt xpredec1_xa_512x8m81 a_197_n10255# m1_n58_n7539# a_421_n10255# m1_n58_n6933#
+ a_645_n10255# m1_n58_n7135# m1_n58_n6530# pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D
+ m1_n58_n7337# a_n1_81# m1_n58_n6732# pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ M3_M2$$47333420_512x8m81_1/VSUBS
Xpmos_1p2$$47512620_512x8m81_0 pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ a_645_n10255# pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47512620_512x8m81
Xpmos_1p2$$47512620_512x8m81_1 pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D
+ a_421_n10255# pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47512620_512x8m81
Xpmos_1p2$$47512620_512x8m81_2 pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ a_197_n10255# pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47512620_512x8m81
Xnmos_1p2$$47514668_512x8m81_0 pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D
+ pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D M3_M2$$47333420_512x8m81_1/VSUBS
+ M3_M2$$47333420_512x8m81_1/VSUBS nmos_1p2$$47514668_512x8m81
Xnmos_1p2$$47514668_512x8m81_1 M3_M2$$47333420_512x8m81_1/VSUBS pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D M3_M2$$47333420_512x8m81_1/VSUBS
+ nmos_1p2$$47514668_512x8m81
Xnmos_1p2$$47514668_512x8m81_2 pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D
+ pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D M3_M2$$47333420_512x8m81_1/VSUBS
+ M3_M2$$47333420_512x8m81_1/VSUBS nmos_1p2$$47514668_512x8m81
Xpmos_1p2$$47513644_512x8m81_0 pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81
Xpmos_1p2$$47513644_512x8m81_1 pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47513644_512x8m81
Xpmos_1p2$$47513644_512x8m81_2 pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_2/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47513644_512x8m81
X0 pmos_1p2$$47512620_512x8m81_2/pmos_5p04310591302072_512x8m81_0/D a_645_n10255# a_541_n10182# M3_M2$$47333420_512x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X1 a_317_n10182# a_197_n10255# M3_M2$$47333420_512x8m81_1/VSUBS M3_M2$$47333420_512x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X2 a_541_n10182# a_421_n10255# a_317_n10182# M3_M2$$47333420_512x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
.ends

.subckt nmos_5p04310591302071_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.58u l=0.6u
.ends

.subckt nmos_1p2$$47336492_512x8m81 nmos_5p04310591302071_512x8m81_0/D nmos_5p04310591302071_512x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310591302071_512x8m81_0 nmos_5p04310591302071_512x8m81_0/D a_n31_n74# nmos_5p04310591302071_512x8m81_0/S
+ VSUBS nmos_5p04310591302071_512x8m81
.ends

.subckt pmos_5p04310591302070_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=16.33u l=0.6u
.ends

.subckt pmos_1p2$$47337516_512x8m81 pmos_5p04310591302070_512x8m81_0/S a_n31_n73#
+ w_n286_n141# pmos_5p04310591302070_512x8m81_0/D
Xpmos_5p04310591302070_512x8m81_0 w_n286_n141# pmos_5p04310591302070_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302070_512x8m81_0/S pmos_5p04310591302070_512x8m81
.ends

.subckt xpredec1_bot_512x8m81 m1_n106_2472# pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ m1_n106_3279# alatch_512x8m81_0/a m1_n106_2674# alatch_512x8m81_0/en alatch_512x8m81_0/vdd
+ pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/S
+ alatch_512x8m81_0/enb m1_n106_2876# m1_n106_3078# m1_n106_3481# VSUBS
Xnmos_1p2$$47336492_512x8m81_0 pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ VSUBS pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D VSUBS nmos_1p2$$47336492_512x8m81
Xpmos_1p2$$47337516_512x8m81_0 pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/S
+ pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/S
+ pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D pmos_1p2$$47337516_512x8m81
Xnmos_1p2$$47336492_512x8m81_1 pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ VSUBS alatch_512x8m81_0/ab VSUBS nmos_1p2$$47336492_512x8m81
Xpmos_1p2$$47337516_512x8m81_1 pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/S
+ alatch_512x8m81_0/ab pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/S
+ pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D pmos_1p2$$47337516_512x8m81
Xalatch_512x8m81_0 alatch_512x8m81_0/enb alatch_512x8m81_0/en alatch_512x8m81_0/ab
+ alatch_512x8m81_0/a VSUBS alatch_512x8m81_0/vdd alatch_512x8m81
.ends

.subckt xpredec1_512x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1] A[0]
+ clk w_7178_9364# pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120#
+ vss vdd
Xxpredec1_xa_512x8m81_0 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[3] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_xa_512x8m81_1 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[1] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_xa_512x8m81_1/a_n1_81# xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_xa_512x8m81_2 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[5] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_bot_512x8m81_0 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ A[0] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D vdd xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd xpredec1_bot_512x8m81_2/alatch_512x8m81_0/enb xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81
Xxpredec1_xa_512x8m81_3 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[7] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_xa_512x8m81_3/a_n1_81# xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_bot_512x8m81_1 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ A[2] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D vdd xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd xpredec1_bot_512x8m81_2/alatch_512x8m81_0/enb xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81
Xxpredec1_xa_512x8m81_4 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[2] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_bot_512x8m81_2 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ A[1] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ nmos_5p04310591302056_512x8m81_1/D vdd xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd xpredec1_bot_512x8m81_2/alatch_512x8m81_0/enb xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81
Xxpredec1_xa_512x8m81_5 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[0] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_xa_512x8m81_6 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[4] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ vss xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xxpredec1_xa_512x8m81_7 xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_0/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_bot_512x8m81_1/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ x[6] xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_0/pmos_5p04310591302070_512x8m81_0/D
+ xpredec1_xa_512x8m81_7/a_n1_81# xpredec1_bot_512x8m81_2/pmos_1p2$$47337516_512x8m81_1/pmos_5p04310591302070_512x8m81_0/D
+ vdd vss xpredec1_xa_512x8m81
Xnmos_1p2$$47342636_512x8m81_0 vss xpredec1_bot_512x8m81_2/alatch_512x8m81_0/enb nmos_5p04310591302056_512x8m81_1/D
+ vss nmos_1p2$$47342636_512x8m81
Xnmos_5p04310591302056_512x8m81_0 vss clk nmos_5p04310591302056_512x8m81_1/D vss nmos_5p04310591302056_512x8m81
Xnmos_5p04310591302056_512x8m81_1 nmos_5p04310591302056_512x8m81_1/D men vss vss nmos_5p04310591302056_512x8m81
Xpmos_1p2$$47109164_512x8m81_0 nmos_5p04310591302056_512x8m81_1/D xpredec1_bot_512x8m81_2/alatch_512x8m81_0/enb
+ pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120# vdd
+ nmos_5p04310591302056_512x8m81_1/D pmos_1p2$$47109164_512x8m81
X0 nmos_5p04310591302056_512x8m81_1/D clk a_7553_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X1 a_7553_9505# men vdd w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X2 a_8001_9505# clk nmos_5p04310591302056_512x8m81_1/D w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X3 vdd men a_8001_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
.ends

.subckt nmos_5p04310591302065_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=5.22u l=0.6u
.ends

.subckt nmos_1p2$$47502380_512x8m81 nmos_5p04310591302065_512x8m81_0/D nmos_5p04310591302065_512x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310591302065_512x8m81_0 nmos_5p04310591302065_512x8m81_0/D a_n31_n74# nmos_5p04310591302065_512x8m81_0/S
+ VSUBS nmos_5p04310591302065_512x8m81
.ends

.subckt pmos_5p04310591302064_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=17.69u l=0.6u
.ends

.subckt pmos_1p2$$47503404_512x8m81 a_n31_n73# pmos_5p04310591302064_512x8m81_0/S
+ w_n286_n141# pmos_5p04310591302064_512x8m81_0/D
Xpmos_5p04310591302064_512x8m81_0 w_n286_n141# pmos_5p04310591302064_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302064_512x8m81_0/S pmos_5p04310591302064_512x8m81
.ends

.subckt nmos_5p04310591302066_512x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=7.04u l=0.6u
.ends

.subckt pmos_5p04310591302063_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.16u l=0.6u
.ends

.subckt pmos_1p2$$47504428_512x8m81 pmos_5p04310591302063_512x8m81_0/S w_n286_n142#
+ pmos_5p04310591302063_512x8m81_0/w_n208_n120# pmos_5p04310591302063_512x8m81_0/D
+ a_n31_n73#
Xpmos_5p04310591302063_512x8m81_0 pmos_5p04310591302063_512x8m81_0/w_n208_n120# pmos_5p04310591302063_512x8m81_0/D
+ a_n31_n73# pmos_5p04310591302063_512x8m81_0/S pmos_5p04310591302063_512x8m81
.ends

.subckt xpredec0_bot_512x8m81 m1_n106_2472# alatch_512x8m81_0/a m1_n106_2674# alatch_512x8m81_0/en
+ alatch_512x8m81_0/vdd pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ alatch_512x8m81_0/enb m1_n106_2876# nmos_5p04310591302066_512x8m81_0/D m1_n106_3078#
+ VSUBS pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S
Xalatch_512x8m81_0 alatch_512x8m81_0/enb alatch_512x8m81_0/en alatch_512x8m81_0/ab
+ alatch_512x8m81_0/a VSUBS alatch_512x8m81_0/vdd alatch_512x8m81
Xnmos_1p2$$47502380_512x8m81_0 pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ VSUBS nmos_5p04310591302066_512x8m81_0/D VSUBS nmos_1p2$$47502380_512x8m81
Xpmos_1p2$$47503404_512x8m81_0 alatch_512x8m81_0/ab pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S
+ pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S nmos_5p04310591302066_512x8m81_0/D
+ pmos_1p2$$47503404_512x8m81
Xnmos_5p04310591302066_512x8m81_0 nmos_5p04310591302066_512x8m81_0/D alatch_512x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310591302066_512x8m81
Xpmos_1p2$$47504428_512x8m81_0 pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S
+ pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/S
+ pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D nmos_5p04310591302066_512x8m81_0/D
+ pmos_1p2$$47504428_512x8m81
.ends

.subckt pmos_5p04310591302067_512x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=15.2u l=0.6u
.ends

.subckt pmos_1p2$$47642668_512x8m81 pmos_5p04310591302067_512x8m81_0/D w_n546_n142#
+ pmos_5p04310591302067_512x8m81_0/S a_n31_n74#
Xpmos_5p04310591302067_512x8m81_0 w_n546_n142# pmos_5p04310591302067_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302067_512x8m81_0/S pmos_5p04310591302067_512x8m81
.ends

.subckt pmos_1p2$$47643692_512x8m81 pmos_5p04310591302067_512x8m81_0/D w_n286_n142#
+ pmos_5p04310591302067_512x8m81_0/S a_n31_n74#
Xpmos_5p04310591302067_512x8m81_0 w_n286_n142# pmos_5p04310591302067_512x8m81_0/D
+ a_n31_n74# pmos_5p04310591302067_512x8m81_0/S pmos_5p04310591302067_512x8m81
.ends

.subckt nmos_1p2$$47641644_512x8m81 a_n31_n73# nmos_5p04310591302057_512x8m81_0/D
+ nmos_5p04310591302057_512x8m81_0/S VSUBS
Xnmos_5p04310591302057_512x8m81_0 nmos_5p04310591302057_512x8m81_0/D a_n31_n73# nmos_5p04310591302057_512x8m81_0/S
+ VSUBS nmos_5p04310591302057_512x8m81
.ends

.subckt xpredec0_xa_512x8m81 m1_342_3273# a_875_414# m3_855_1044# a_651_414# nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D m1_342_3474# m3_153_8117#
+ m1_342_3071# pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/S m1_342_3676#
+ M3_M2$$47644716_512x8m81_2/VSUBS pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ nmos_1p2$$47641644_512x8m81_3/nmos_5p04310591302057_512x8m81_0/D
Xpmos_1p2$$47642668_512x8m81_0 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ a_875_414# pmos_1p2$$47642668_512x8m81
Xpmos_1p2$$47643692_512x8m81_0 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ a_651_414# pmos_1p2$$47643692_512x8m81
Xnmos_1p2$$47641644_512x8m81_0 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ M3_M2$$47644716_512x8m81_2/VSUBS nmos_1p2$$47641644_512x8m81
Xnmos_1p2$$47641644_512x8m81_1 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D nmos_1p2$$47641644_512x8m81_3/nmos_5p04310591302057_512x8m81_0/D
+ M3_M2$$47644716_512x8m81_2/VSUBS nmos_1p2$$47641644_512x8m81
Xnmos_1p2$$47641644_512x8m81_2 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ nmos_1p2$$47641644_512x8m81_3/nmos_5p04310591302057_512x8m81_0/D pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D
+ M3_M2$$47644716_512x8m81_2/VSUBS nmos_1p2$$47641644_512x8m81
Xnmos_1p2$$47641644_512x8m81_3 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ nmos_1p2$$47641644_512x8m81_3/nmos_5p04310591302057_512x8m81_0/D pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D
+ M3_M2$$47644716_512x8m81_2/VSUBS nmos_1p2$$47641644_512x8m81
Xpmos_1p2$$47513644_512x8m81_0 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81
Xpmos_1p2$$47513644_512x8m81_1 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47513644_512x8m81
Xpmos_1p2$$47513644_512x8m81_2 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47513644_512x8m81
Xpmos_1p2$$47513644_512x8m81_3 pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/S pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/D
+ pmos_1p2$$47513644_512x8m81_3/pmos_5p04310591302068_512x8m81_0/D pmos_1p2$$47513644_512x8m81
X0 a_771_486# a_651_414# pmos_1p2$$47643692_512x8m81_0/pmos_5p04310591302067_512x8m81_0/S M3_M2$$47644716_512x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
X1 M3_M2$$47644716_512x8m81_2/VSUBS a_875_414# a_771_486# M3_M2$$47644716_512x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
.ends

.subckt pmos_5p04310591302069_512x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt xpredec0_512x8m81 A[0] men x[0] x[1] x[2] x[3] A[1] clk xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ vdd vss
Xnmos_1p2$$46563372_512x8m81_0 vss nmos_5p04310591302040_512x8m81_1/S pmos_5p04310591302069_512x8m81_0/D
+ vss nmos_1p2$$46563372_512x8m81
Xxpredec0_bot_512x8m81_0 xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ A[0] xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D nmos_5p04310591302040_512x8m81_1/S
+ vdd xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ pmos_5p04310591302069_512x8m81_0/D xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D
+ vss vdd xpredec0_bot_512x8m81
Xxpredec0_bot_512x8m81_1 xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ A[1] xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D nmos_5p04310591302040_512x8m81_1/S
+ vdd xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ pmos_5p04310591302069_512x8m81_0/D xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D
+ vss vdd xpredec0_bot_512x8m81
Xnmos_5p04310591302040_512x8m81_0 nmos_5p04310591302040_512x8m81_1/S men vss vss nmos_5p04310591302040_512x8m81
Xxpredec0_xa_512x8m81_0 xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D
+ xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ x[0] xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vss xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D vss vdd vss xpredec0_xa_512x8m81
Xnmos_5p04310591302040_512x8m81_1 vss clk nmos_5p04310591302040_512x8m81_1/S vss nmos_5p04310591302040_512x8m81
Xxpredec0_xa_512x8m81_1 xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D
+ xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ x[2] xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vss xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D vss vdd vss xpredec0_xa_512x8m81
Xxpredec0_xa_512x8m81_2 xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D
+ xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D vdd xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ x[1] xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vss xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D vss vdd vss xpredec0_xa_512x8m81
Xxpredec0_xa_512x8m81_3 xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D
+ xpredec0_bot_512x8m81_0/nmos_5p04310591302066_512x8m81_0/D vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D
+ xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ x[3] xpredec0_bot_512x8m81_1/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vss xpredec0_bot_512x8m81_0/pmos_1p2$$47504428_512x8m81_0/pmos_5p04310591302063_512x8m81_0/D
+ vdd xpredec0_bot_512x8m81_1/nmos_5p04310591302066_512x8m81_0/D vss vdd vss xpredec0_xa_512x8m81
Xpmos_5p04310591302069_512x8m81_0 vdd pmos_5p04310591302069_512x8m81_0/D nmos_5p04310591302040_512x8m81_1/S
+ vdd nmos_5p04310591302040_512x8m81_1/S pmos_5p04310591302069_512x8m81
X0 vdd men a_4894_9505# vdd pmos_3p3 w=1.705u l=0.6u
X1 a_4446_9505# men vdd vdd pmos_3p3 w=1.705u l=0.6u
X2 a_4894_9505# clk nmos_5p04310591302040_512x8m81_1/S vdd pmos_3p3 w=1.705u l=0.6u
X3 nmos_5p04310591302040_512x8m81_1/S clk a_4446_9505# vdd pmos_3p3 w=1.705u l=0.6u
.ends

.subckt prexdec_top_512x8m81 clk A[2] A[6] A[4] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1]
+ xb[2] xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1] xpredec1_512x8m81_0/w_7178_9364#
+ xpredec1_512x8m81_0/pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120#
+ xpredec0_512x8m81_0/xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_512x8m81_0/xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_512x8m81_1/xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_512x8m81_1/xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xc[0] men xpredec1_512x8m81_0/vdd VSUBS
Xxpredec1_512x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] clk xpredec1_512x8m81_0/w_7178_9364# xpredec1_512x8m81_0/pmos_1p2$$47109164_512x8m81_0/pmos_5p04310591302062_512x8m81_0/w_n208_n120#
+ VSUBS xpredec1_512x8m81_0/vdd xpredec1_512x8m81
Xxpredec0_512x8m81_0 A[3] men xb[0] xb[1] xb[2] xb[3] A[4] clk xpredec0_512x8m81_0/xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_512x8m81_0/xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec1_512x8m81_0/vdd VSUBS xpredec0_512x8m81
Xxpredec0_512x8m81_1 A[5] men xc[0] xc[1] xc[2] xc[3] A[6] clk xpredec0_512x8m81_1/xpredec0_xa_512x8m81_3/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec0_512x8m81_1/xpredec0_xa_512x8m81_2/nmos_1p2$$47641644_512x8m81_0/nmos_5p04310591302057_512x8m81_0/S
+ xpredec1_512x8m81_0/vdd VSUBS xpredec0_512x8m81
.ends

.subckt control_512x8_512x8m81 VSS VDD RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xb[1] xc[3] xc[1] xc[2] xc[0] xa[0]
+ xa[1] A[9] A[7] CLK A[6] A[3] A[4] A[5] A[8] GWE GWEN ypredec1_512x8m81_0/ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd
+ ypredec1_512x8m81_0/ly[2] CEN A[0] A[1] A[2] men VSUBS gen_512x8_512x8m81_0/VDD
+ prexdec_top_512x8m81_0/xpredec1_512x8m81_0/vdd gen_512x8_512x8m81_0/tblhl
Xgen_512x8_512x8m81_0 gen_512x8_512x8m81_0/tblhl IGWEN CLK GWEN GWE gen_512x8_512x8m81_0/pmos_5p04310591302088_512x8m81_0/D
+ CEN men gen_512x8_512x8m81_0/VDD VSUBS gen_512x8_512x8m81
Xypredec1_512x8m81_0 ypredec1_512x8m81_0/ly[5] ypredec1_512x8m81_0/ly[4] ypredec1_512x8m81_0/ly[7]
+ ypredec1_512x8m81_0/ly[3] ypredec1_512x8m81_0/ly[2] ypredec1_512x8m81_0/ly[1] ypredec1_512x8m81_0/ly[0]
+ RYS[0] RYS[1] RYS[2] RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_512x8m81_0/ly[6]
+ men A[0] A[1] A[2] CLK gen_512x8_512x8m81_0/VDD ypredec1_512x8m81_0/ypredec1_bot_512x8m81_2/alatch_512x8m81_0/vdd
+ gen_512x8_512x8m81_0/VDD gen_512x8_512x8m81_0/VDD gen_512x8_512x8m81_0/VDD VSUBS
+ ypredec1_512x8m81
Xprexdec_top_512x8m81_0 CLK A[5] A[9] A[7] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1] xb[2]
+ xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] prexdec_top_512x8m81_0/xpredec1_512x8m81_0/vdd
+ prexdec_top_512x8m81_0/xpredec1_512x8m81_0/vdd VSUBS VSUBS VSUBS VSUBS xc[0] men
+ prexdec_top_512x8m81_0/xpredec1_512x8m81_0/vdd VSUBS prexdec_top_512x8m81
.ends

.subckt gf180mcu_fd_ip_sram__sram512x8m8wm1 VSS CLK D[0] A[8] A[7] A[2] A[1] A[0]
+ Q[2] Q[3] CEN A[5] A[6] A[4] WEN[3] D[7] Q[7] D[3] D[1] D[2] A[3] Q[1] Q[6] D[5]
+ Q[4] WEN[5] WEN[2] WEN[1] WEN[4] WEN[7] WEN[6] D[4] D[6] Q[5] Q[0] GWEN WEN[0]
Xlcol4_512_512x8m81_0 lcol4_512_512x8m81_0/WL[32] lcol4_512_512x8m81_0/WL[33] lcol4_512_512x8m81_0/WL[34]
+ lcol4_512_512x8m81_0/WL[38] lcol4_512_512x8m81_0/WL[39] lcol4_512_512x8m81_0/WL[35]
+ lcol4_512_512x8m81_0/WL[36] lcol4_512_512x8m81_0/WL[37] lcol4_512_512x8m81_0/WL[40]
+ lcol4_512_512x8m81_0/WL[41] lcol4_512_512x8m81_0/WL[42] lcol4_512_512x8m81_0/WL[43]
+ lcol4_512_512x8m81_0/WL[44] lcol4_512_512x8m81_0/WL[45] lcol4_512_512x8m81_0/WL[46]
+ lcol4_512_512x8m81_0/WL[47] lcol4_512_512x8m81_0/WL[48] lcol4_512_512x8m81_0/WL[49]
+ lcol4_512_512x8m81_0/WL[50] lcol4_512_512x8m81_0/WL[51] lcol4_512_512x8m81_0/WL[52]
+ lcol4_512_512x8m81_0/WL[53] lcol4_512_512x8m81_0/WL[54] lcol4_512_512x8m81_0/WL[55]
+ lcol4_512_512x8m81_0/WL[56] lcol4_512_512x8m81_0/WL[57] lcol4_512_512x8m81_0/WL[58]
+ lcol4_512_512x8m81_0/WL[59] lcol4_512_512x8m81_0/WL[60] lcol4_512_512x8m81_0/WL[61]
+ lcol4_512_512x8m81_0/WL[62] lcol4_512_512x8m81_0/WL[63] lcol4_512_512x8m81_0/WL[25]
+ lcol4_512_512x8m81_0/WL[24] lcol4_512_512x8m81_0/WL[23] lcol4_512_512x8m81_0/WL[22]
+ lcol4_512_512x8m81_0/WL[21] lcol4_512_512x8m81_0/WL[20] lcol4_512_512x8m81_0/WL[19]
+ lcol4_512_512x8m81_0/WL[18] lcol4_512_512x8m81_0/WL[17] lcol4_512_512x8m81_0/WL[16]
+ lcol4_512_512x8m81_0/WL[15] lcol4_512_512x8m81_0/WL[14] lcol4_512_512x8m81_0/WL[13]
+ lcol4_512_512x8m81_0/WL[12] lcol4_512_512x8m81_0/WL[11] lcol4_512_512x8m81_0/WL[10]
+ lcol4_512_512x8m81_0/WL[9] lcol4_512_512x8m81_0/WL[8] lcol4_512_512x8m81_0/WL[7]
+ lcol4_512_512x8m81_0/WL[6] lcol4_512_512x8m81_0/WL[5] lcol4_512_512x8m81_0/WL[4]
+ lcol4_512_512x8m81_0/WL[3] lcol4_512_512x8m81_0/WL[2] lcol4_512_512x8m81_0/WL[1]
+ lcol4_512_512x8m81_0/WL[0] lcol4_512_512x8m81_0/WL[31] lcol4_512_512x8m81_0/WL[30]
+ lcol4_512_512x8m81_0/WL[29] lcol4_512_512x8m81_0/WL[28] lcol4_512_512x8m81_0/WL[27]
+ lcol4_512_512x8m81_0/WL[26] lcol4_512_512x8m81_0/men lcol4_512_512x8m81_0/ypass[0]
+ lcol4_512_512x8m81_0/ypass[1] lcol4_512_512x8m81_0/ypass[2] lcol4_512_512x8m81_0/ypass[3]
+ lcol4_512_512x8m81_0/ypass[4] lcol4_512_512x8m81_0/ypass[5] lcol4_512_512x8m81_0/ypass[6]
+ lcol4_512_512x8m81_0/ypass[7] VSS lcol4_512_512x8m81_0/GWEN lcol4_512_512x8m81_0/GWE
+ D[0] D[1] D[3] D[2] Q[0] Q[1] Q[2] Q[3] lcol4_512_512x8m81_0/pcb[2] lcol4_512_512x8m81_0/pcb[3]
+ lcol4_512_512x8m81_0/pcb[0] lcol4_512_512x8m81_0/pcb[1] VSS WEN[0] WEN[1] WEN[2]
+ WEN[3] xdec64_512x8m81_0/LWL[62] xdec64_512x8m81_0/LWL[29] xdec64_512x8m81_0/LWL[46]
+ xdec64_512x8m81_0/LWL[63] VSS xdec64_512x8m81_0/LWL[47] xdec64_512x8m81_0/LWL[48]
+ WEN[3] xdec64_512x8m81_0/LWL[49] xdec64_512x8m81_0/LWL[10] xdec64_512x8m81_0/LWL[11]
+ xdec64_512x8m81_0/LWL[12] xdec64_512x8m81_0/LWL[13] xdec64_512x8m81_0/LWL[30] xdec64_512x8m81_0/LWL[14]
+ xdec64_512x8m81_0/LWL[31] VSS xdec64_512x8m81_0/LWL[15] xdec64_512x8m81_0/LWL[32]
+ xdec64_512x8m81_0/LWL[0] xdec64_512x8m81_0/LWL[16] xdec64_512x8m81_0/LWL[33] xdec64_512x8m81_0/LWL[1]
+ xdec64_512x8m81_0/LWL[50] VSS xdec64_512x8m81_0/LWL[17] xdec64_512x8m81_0/LWL[34]
+ xdec64_512x8m81_0/LWL[2] xdec64_512x8m81_0/LWL[51] xdec64_512x8m81_0/LWL[18] xdec64_512x8m81_0/LWL[35]
+ VSS xdec64_512x8m81_0/LWL[3] xdec64_512x8m81_0/LWL[52] xdec64_512x8m81_0/LWL[19]
+ xdec64_512x8m81_0/LWL[36] xdec64_512x8m81_0/LWL[53] xdec64_512x8m81_0/LWL[4] xdec64_512x8m81_0/LWL[37]
+ xdec64_512x8m81_0/LWL[54] xdec64_512x8m81_0/LWL[5] xdec64_512x8m81_0/LWL[38] xdec64_512x8m81_0/LWL[6]
+ xdec64_512x8m81_0/LWL[55] xdec64_512x8m81_0/LWL[39] xdec64_512x8m81_0/LWL[7] xdec64_512x8m81_0/LWL[56]
+ VSS xdec64_512x8m81_0/LWL[8] xdec64_512x8m81_0/LWL[57] xdec64_512x8m81_0/LWL[58]
+ xdec64_512x8m81_0/LWL[9] xdec64_512x8m81_0/LWL[59] WEN[0] xdec64_512x8m81_0/men
+ lcol4_512_512x8m81_0/col_512a_512x8m81_0/saout_m2_512x8m81_1/sa_512x8m81_0/pcb xdec64_512x8m81_0/LWL[20]
+ xdec64_512x8m81_0/LWL[21] control_512x8_512x8m81_0/LYS[0] rcol4_512_512x8m81_0/GWE
+ VSS xdec64_512x8m81_0/LWL[22] control_512x8_512x8m81_0/LYS[1] xdec64_512x8m81_0/LWL[23]
+ xdec64_512x8m81_0/LWL[40] control_512x8_512x8m81_0/LYS[2] rcol4_512_512x8m81_0/GWEN
+ xdec64_512x8m81_0/LWL[24] xdec64_512x8m81_0/LWL[41] control_512x8_512x8m81_0/LYS[3]
+ xdec64_512x8m81_0/LWL[25] VSS lcol4_512_512x8m81_0/col_512a_512x8m81_0/saout_m2_512x8m81_0/pcb
+ xdec64_512x8m81_0/LWL[42] control_512x8_512x8m81_0/LYS[4] xdec64_512x8m81_0/LWL[26]
+ control_512x8_512x8m81_0/LYS[5] xdec64_512x8m81_0/LWL[43] xdec64_512x8m81_0/LWL[60]
+ VSS VSS lcol4_512_512x8m81_0/col_512a_512x8m81_0/saout_R_m2_512x8m81_1/sa_512x8m81_0/pcb
+ lcol4_512_512x8m81_0/col_512a_512x8m81_0/saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb
+ xdec64_512x8m81_0/LWL[27] control_512x8_512x8m81_0/LYS[6] xdec64_512x8m81_0/LWL[44]
+ xdec64_512x8m81_0/LWL[61] xdec64_512x8m81_0/LWL[28] VSS control_512x8_512x8m81_0/LYS[7]
+ xdec64_512x8m81_0/LWL[45] VSS VSS lcol4_512_512x8m81
Xrcol4_512_512x8m81_0 xdec64_512x8m81_0/RWL[32] xdec64_512x8m81_0/RWL[33] xdec64_512x8m81_0/RWL[34]
+ xdec64_512x8m81_0/RWL[35] xdec64_512x8m81_0/RWL[36] xdec64_512x8m81_0/RWL[37] xdec64_512x8m81_0/RWL[42]
+ xdec64_512x8m81_0/RWL[44] xdec64_512x8m81_0/RWL[46] xdec64_512x8m81_0/RWL[48] xdec64_512x8m81_0/RWL[50]
+ xdec64_512x8m81_0/RWL[52] xdec64_512x8m81_0/RWL[54] xdec64_512x8m81_0/RWL[56] xdec64_512x8m81_0/RWL[57]
+ xdec64_512x8m81_0/RWL[59] xdec64_512x8m81_0/DRWL xdec64_512x8m81_0/RWL[61] xdec64_512x8m81_0/RWL[51]
+ xdec64_512x8m81_0/RWL[29] xdec64_512x8m81_0/RWL[25] xdec64_512x8m81_0/RWL[24] xdec64_512x8m81_0/RWL[23]
+ xdec64_512x8m81_0/RWL[22] xdec64_512x8m81_0/RWL[20] xdec64_512x8m81_0/RWL[27] xdec64_512x8m81_0/RWL[30]
+ xdec64_512x8m81_0/RWL[18] xdec64_512x8m81_0/RWL[41] xdec64_512x8m81_0/RWL[15] xdec64_512x8m81_0/RWL[38]
+ xdec64_512x8m81_0/RWL[45] xdec64_512x8m81_0/RWL[43] xdec64_512x8m81_0/RWL[40] xdec64_512x8m81_0/RWL[39]
+ xdec64_512x8m81_0/RWL[31] xdec64_512x8m81_0/RWL[14] xdec64_512x8m81_0/RWL[16] xdec64_512x8m81_0/RWL[17]
+ xdec64_512x8m81_0/RWL[26] xdec64_512x8m81_0/RWL[19] xdec64_512x8m81_0/RWL[58] xdec64_512x8m81_0/RWL[60]
+ xdec64_512x8m81_0/RWL[62] xdec64_512x8m81_0/RWL[28] xdec64_512x8m81_0/RWL[63] xdec64_512x8m81_0/RWL[21]
+ xdec64_512x8m81_0/RWL[49] xdec64_512x8m81_0/RWL[53] xdec64_512x8m81_0/RWL[47] xdec64_512x8m81_0/RWL[55]
+ xdec64_512x8m81_0/RWL[0] xdec64_512x8m81_0/RWL[2] xdec64_512x8m81_0/RWL[12] xdec64_512x8m81_0/RWL[3]
+ xdec64_512x8m81_0/RWL[4] xdec64_512x8m81_0/RWL[7] xdec64_512x8m81_0/RWL[8] xdec64_512x8m81_0/RWL[9]
+ xdec64_512x8m81_0/RWL[1] rcol4_512_512x8m81_0/ypass[7] xdec64_512x8m81_0/RWL[5]
+ rcol4_512_512x8m81_0/ypass[0] xdec64_512x8m81_0/RWL[10] xdec64_512x8m81_0/RWL[13]
+ rcol4_512_512x8m81_0/ypass[1] rcol4_512_512x8m81_0/ypass[2] rcol4_512_512x8m81_0/ypass[3]
+ rcol4_512_512x8m81_0/ypass[4] rcol4_512_512x8m81_0/ypass[5] rcol4_512_512x8m81_0/ypass[6]
+ xdec64_512x8m81_0/RWL[6] rcol4_512_512x8m81_0/tblhl rcol4_512_512x8m81_0/GWEN xdec64_512x8m81_0/RWL[11]
+ D[4] D[7] Q[5] Q[6] Q[7] D[5] D[6] Q[4] rcol4_512_512x8m81_0/pcb[6] rcol4_512_512x8m81_0/pcb[7]
+ rcol4_512_512x8m81_0/pcb[4] rcol4_512_512x8m81_0/vdd WEN[7] WEN[4] rcol4_512_512x8m81_0/pcb[5]
+ WEN[6] WEN[5] xdec64_512x8m81_0/RWL[39] xdec64_512x8m81_0/RWL[56] VSS xdec64_512x8m81_0/RWL[57]
+ xdec64_512x8m81_0/RWL[58] VSS xdec64_512x8m81_0/RWL[59] xdec64_512x8m81_0/RWL[20]
+ rcol4_512_512x8m81_0/GWE xdec64_512x8m81_0/RWL[21] WEN[7] xdec64_512x8m81_0/RWL[22]
+ xdec64_512x8m81_0/RWL[23] xdec64_512x8m81_0/RWL[40] VSS xdec64_512x8m81_0/RWL[24]
+ xdec64_512x8m81_0/RWL[41] xdec64_512x8m81_0/RWL[25] xdec64_512x8m81_0/RWL[0] xdec64_512x8m81_0/RWL[42]
+ VSS xdec64_512x8m81_0/RWL[26] xdec64_512x8m81_0/RWL[1] xdec64_512x8m81_0/RWL[43]
+ xdec64_512x8m81_0/RWL[60] xdec64_512x8m81_0/RWL[27] xdec64_512x8m81_0/RWL[2] xdec64_512x8m81_0/RWL[44]
+ VSS VSS xdec64_512x8m81_0/RWL[61] xdec64_512x8m81_0/RWL[28] xdec64_512x8m81_0/RWL[3]
+ xdec64_512x8m81_0/RWL[45] xdec64_512x8m81_0/RWL[62] xdec64_512x8m81_0/RWL[29] xdec64_512x8m81_0/RWL[4]
+ xdec64_512x8m81_0/RWL[46] VSS xdec64_512x8m81_0/RWL[63] rcol4_512_512x8m81_0/saout_R_m2_512x8m81_1/pcb
+ xdec64_512x8m81_0/RWL[5] VSS xdec64_512x8m81_0/RWL[47] xdec64_512x8m81_0/RWL[6]
+ xdec64_512x8m81_0/RWL[48] xdec64_512x8m81_0/RWL[7] xdec64_512x8m81_0/RWL[49] xdec64_512x8m81_0/RWL[8]
+ xdec64_512x8m81_0/RWL[9] xdec64_512x8m81_0/RWL[10] xdec64_512x8m81_0/men xdec64_512x8m81_0/RWL[11]
+ xdec64_512x8m81_0/RWL[12] VSS rcol4_512_512x8m81_0/saout_m2_512x8m81_1/sa_512x8m81_0/pcb
+ xdec64_512x8m81_0/RWL[13] xdec64_512x8m81_0/RWL[30] xdec64_512x8m81_0/RWL[14] xdec64_512x8m81_0/RWL[31]
+ VSS xdec64_512x8m81_0/RWL[15] xdec64_512x8m81_0/RWL[32] VSS xdec64_512x8m81_0/DRWL
+ xdec64_512x8m81_0/RWL[16] xdec64_512x8m81_0/RWL[33] xdec64_512x8m81_0/RWL[50] xdec64_512x8m81_0/RWL[17]
+ xdec64_512x8m81_0/RWL[34] xdec64_512x8m81_0/RWL[51] xdec64_512x8m81_0/RWL[18] xdec64_512x8m81_0/RWL[35]
+ xdec64_512x8m81_0/RWL[52] xdec64_512x8m81_0/RWL[19] xdec64_512x8m81_0/RWL[36] rcol4_512_512x8m81_0/saout_m2_512x8m81_0/pcb
+ xdec64_512x8m81_0/RWL[53] rcol4_512_512x8m81_0/saout_R_m2_512x8m81_0/sa_512x8m81_0/pcb
+ rcol4_512_512x8m81_0/saout_R_m2_512x8m81_1/pcb xdec64_512x8m81_0/RWL[37] xdec64_512x8m81_0/RWL[54]
+ xdec64_512x8m81_0/RWL[38] xdec64_512x8m81_0/RWL[55] VSS VSS rcol4_512_512x8m81
Xxdec64_512x8m81_0 xdec64_512x8m81_0/DRWL xdec64_512x8m81_0/RWL[34] xdec64_512x8m81_0/RWL[35]
+ xdec64_512x8m81_0/RWL[36] xdec64_512x8m81_0/RWL[37] xdec64_512x8m81_0/RWL[38] xdec64_512x8m81_0/RWL[39]
+ xdec64_512x8m81_0/RWL[40] xdec64_512x8m81_0/RWL[42] xdec64_512x8m81_0/RWL[43] xdec64_512x8m81_0/RWL[44]
+ xdec64_512x8m81_0/RWL[45] xdec64_512x8m81_0/RWL[46] xdec64_512x8m81_0/RWL[48] xdec64_512x8m81_0/RWL[50]
+ xdec64_512x8m81_0/RWL[53] xdec64_512x8m81_0/RWL[55] xdec64_512x8m81_0/RWL[57] xdec64_512x8m81_0/RWL[58]
+ xdec64_512x8m81_0/RWL[61] xdec64_512x8m81_0/RWL[62] xdec64_512x8m81_0/RWL[63] xdec64_512x8m81_0/LWL[58]
+ xdec64_512x8m81_0/LWL[56] xdec64_512x8m81_0/LWL[55] xdec64_512x8m81_0/LWL[54] xdec64_512x8m81_0/LWL[53]
+ xdec64_512x8m81_0/LWL[52] xdec64_512x8m81_0/LWL[51] xdec64_512x8m81_0/LWL[50] xdec64_512x8m81_0/LWL[46]
+ xdec64_512x8m81_0/LWL[38] xdec64_512x8m81_0/LWL[36] xdec64_512x8m81_0/LWL[35] xdec64_512x8m81_0/LWL[34]
+ xdec64_512x8m81_0/DLWL xdec64_512x8m81_0/LWL[19] xdec64_512x8m81_0/LWL[20] xdec64_512x8m81_0/LWL[21]
+ xdec64_512x8m81_0/LWL[22] xdec64_512x8m81_0/LWL[27] xdec64_512x8m81_0/LWL[11] xdec64_512x8m81_0/LWL[13]
+ xdec64_512x8m81_0/LWL[15] xdec64_512x8m81_0/LWL[18] xdec64_512x8m81_0/LWL[5] xdec64_512x8m81_0/LWL[4]
+ xdec64_512x8m81_0/LWL[2] xdec64_512x8m81_0/LWL[8] xdec64_512x8m81_0/LWL[9] xdec64_512x8m81_0/LWL[6]
+ xdec64_512x8m81_0/LWL[7] xdec64_512x8m81_0/LWL[29] xdec64_512x8m81_0/RWL[31] xdec64_512x8m81_0/RWL[30]
+ xdec64_512x8m81_0/RWL[6] xdec64_512x8m81_0/RWL[4] xdec64_512x8m81_0/RWL[2] xdec64_512x8m81_0/RWL[0]
+ xdec64_512x8m81_0/RWL[1] xdec64_512x8m81_0/RWL[3] xdec64_512x8m81_0/RWL[5] xdec64_512x8m81_0/RWL[7]
+ xdec64_512x8m81_0/RWL[8] xdec64_512x8m81_0/RWL[10] xdec64_512x8m81_0/RWL[12] xdec64_512x8m81_0/RWL[14]
+ xdec64_512x8m81_0/RWL[15] xdec64_512x8m81_0/RWL[16] xdec64_512x8m81_0/RWL[17] xdec64_512x8m81_0/xb[0]
+ xdec64_512x8m81_0/xb[1] xdec64_512x8m81_0/xb[2] xdec64_512x8m81_0/xb[3] xdec64_512x8m81_0/xa[7]
+ xdec64_512x8m81_0/xa[6] xdec64_512x8m81_0/xa[5] xdec64_512x8m81_0/xa[4] xdec64_512x8m81_0/xa[0]
+ xdec64_512x8m81_0/xa[3] xdec64_512x8m81_0/xa[2] xdec64_512x8m81_0/xc[0] xdec64_512x8m81_0/xc[1]
+ xdec64_512x8m81_0/LWL[44] xdec64_512x8m81_0/LWL[42] xdec64_512x8m81_0/LWL[25] xdec64_512x8m81_0/LWL[40]
+ xdec64_512x8m81_0/RWL[41] xdec64_512x8m81_0/LWL[23] xdec64_512x8m81_0/LWL[49] xdec64_512x8m81_0/RWL[60]
+ xdec64_512x8m81_0/RWL[59] xdec64_512x8m81_0/LWL[62] xdec64_512x8m81_0/LWL[60] xdec64_512x8m81_0/RWL[29]
+ xdec64_512x8m81_0/LWL[47] xdec64_512x8m81_0/RWL[27] xdec64_512x8m81_0/LWL[48] xdec64_512x8m81_0/LWL[45]
+ xdec64_512x8m81_0/RWL[25] xdec64_512x8m81_0/LWL[0] xdec64_512x8m81_0/LWL[30] xdec64_512x8m81_0/LWL[63]
+ xdec64_512x8m81_0/LWL[28] xdec64_512x8m81_0/LWL[43] xdec64_512x8m81_0/LWL[26] xdec64_512x8m81_0/RWL[23]
+ xdec64_512x8m81_0/LWL[24] xdec64_512x8m81_0/LWL[33] xdec64_512x8m81_0/LWL[3] xdec64_512x8m81_0/RWL[28]
+ xdec64_512x8m81_0/LWL[61] xdec64_512x8m81_0/RWL[13] xdec64_512x8m81_0/RWL[26] xdec64_512x8m81_0/LWL[41]
+ xdec64_512x8m81_0/LWL[32] xdec64_512x8m81_0/RWL[24] xdec64_512x8m81_0/RWL[51] xdec64_512x8m81_0/RWL[21]
+ xdec64_512x8m81_0/RWL[32] xdec64_512x8m81_0/RWL[22] xdec64_512x8m81_0/LWL[1] xdec64_512x8m81_0/RWL[33]
+ xdec64_512x8m81_0/RWL[20] xdec64_512x8m81_0/LWL[59] xdec64_512x8m81_0/RWL[11] xdec64_512x8m81_0/RWL[18]
+ xdec64_512x8m81_0/LWL[39] xdec64_512x8m81_0/xa[1] xdec64_512x8m81_0/LWL[16] xdec64_512x8m81_0/RWL[49]
+ xdec64_512x8m81_0/RWL[19] xdec64_512x8m81_0/LWL[14] xdec64_512x8m81_0/LWL[31] xdec64_512x8m81_0/LWL[12]
+ xdec64_512x8m81_0/RWL[56] xdec64_512x8m81_0/LWL[57] xdec64_512x8m81_0/men xdec64_512x8m81_0/LWL[10]
+ xdec64_512x8m81_0/RWL[9] VSS xdec64_512x8m81_0/LWL[37] xdec64_512x8m81_0/RWL[54]
+ VSS xdec64_512x8m81_0/LWL[17] xdec64_512x8m81_0/RWL[52] xdec64_512x8m81_0/RWL[47]
+ xdec64_512x8m81
Xcontrol_512x8_512x8m81_0 VSS VSS rcol4_512_512x8m81_0/ypass[7] rcol4_512_512x8m81_0/ypass[6]
+ rcol4_512_512x8m81_0/ypass[5] rcol4_512_512x8m81_0/ypass[4] rcol4_512_512x8m81_0/ypass[3]
+ rcol4_512_512x8m81_0/ypass[2] rcol4_512_512x8m81_0/ypass[1] rcol4_512_512x8m81_0/ypass[0]
+ control_512x8_512x8m81_0/LYS[0] control_512x8_512x8m81_0/LYS[1] control_512x8_512x8m81_0/LYS[2]
+ control_512x8_512x8m81_0/LYS[3] control_512x8_512x8m81_0/LYS[6] control_512x8_512x8m81_0/LYS[5]
+ control_512x8_512x8m81_0/LYS[4] control_512x8_512x8m81_0/LYS[7] rcol4_512_512x8m81_0/tblhl
+ rcol4_512_512x8m81_0/GWEN xdec64_512x8m81_0/xb[3] xdec64_512x8m81_0/xb[2] xdec64_512x8m81_0/xb[0]
+ xdec64_512x8m81_0/xa[7] xdec64_512x8m81_0/xa[6] xdec64_512x8m81_0/xa[5] xdec64_512x8m81_0/xa[4]
+ xdec64_512x8m81_0/xa[3] xdec64_512x8m81_0/xa[2] xdec64_512x8m81_0/xb[1] control_512x8_512x8m81_0/xc[3]
+ xdec64_512x8m81_0/xc[1] control_512x8_512x8m81_0/xc[2] xdec64_512x8m81_0/xc[0] xdec64_512x8m81_0/xa[0]
+ xdec64_512x8m81_0/xa[1] VSS A[7] CLK A[6] A[3] A[4] A[5] A[8] rcol4_512_512x8m81_0/GWE
+ GWEN VSS control_512x8_512x8m81_0/LYS[2] CEN A[0] A[1] A[2] xdec64_512x8m81_0/men
+ VSS VSS VSS rcol4_512_512x8m81_0/tblhl control_512x8_512x8m81
.ends

