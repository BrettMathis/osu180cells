magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1008 844
rect 80 636 126 724
rect 252 589 330 678
rect 488 636 534 724
rect 692 590 754 678
rect 896 636 942 724
rect 692 589 982 590
rect 252 543 982 589
rect 132 378 280 438
rect 132 242 204 378
rect 80 60 126 196
rect 360 122 428 438
rect 580 122 648 438
rect 804 242 874 438
rect 920 196 982 543
rect 755 106 982 196
rect 0 -60 1008 60
<< labels >>
rlabel metal1 s 804 242 874 438 6 A1
port 1 nsew default input
rlabel metal1 s 580 122 648 438 6 A2
port 2 nsew default input
rlabel metal1 s 360 122 428 438 6 A3
port 3 nsew default input
rlabel metal1 s 132 378 280 438 6 A4
port 4 nsew default input
rlabel metal1 s 132 242 204 378 6 A4
port 4 nsew default input
rlabel metal1 s 692 590 754 678 6 ZN
port 5 nsew default output
rlabel metal1 s 252 590 330 678 6 ZN
port 5 nsew default output
rlabel metal1 s 692 589 982 590 6 ZN
port 5 nsew default output
rlabel metal1 s 252 589 330 590 6 ZN
port 5 nsew default output
rlabel metal1 s 252 543 982 589 6 ZN
port 5 nsew default output
rlabel metal1 s 920 196 982 543 6 ZN
port 5 nsew default output
rlabel metal1 s 755 106 982 196 6 ZN
port 5 nsew default output
rlabel metal1 s 0 724 1008 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 896 636 942 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 488 636 534 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 80 636 126 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 80 60 126 196 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1008 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1008 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 711982
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 708912
<< end >>
