magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 918 224 1098
rect 30 263 95 643
rect 0 -90 224 90
<< labels >>
rlabel metal1 s 30 263 95 643 6 I
port 1 nsew default input
rlabel metal1 s 0 918 224 1098 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -90 224 90 8 VSS
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 1008
string LEFclass core gf180mcu_fd_sc_mcu9t5v0__antennaCELL
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1144494
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1143014
<< end >>
