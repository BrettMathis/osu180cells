magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect 85432 578 85816 67902
<< metal1 >>
rect 0 403 1000 67894
rect 84808 403 85808 67894
<< metal2 >>
rect 424 403 1424 67376
rect 84384 403 85384 67376
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_0
timestamp 1669390400
transform 1 0 85474 0 1 1140
box -42 -42 342 66242
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_1
timestamp 1669390400
transform 1 0 27139 0 1 1140
box -42 -42 342 66242
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_2
timestamp 1669390400
transform 1 0 57047 0 1 1140
box -42 -42 342 66242
use M1_PSUB43105908781105_256x8m81  M1_PSUB43105908781105_256x8m81_3
timestamp 1669390400
transform 1 0 112 0 1 1140
box -42 -42 342 66242
use M1_PSUB43105908781106_256x8m81  M1_PSUB43105908781106_256x8m81_0
timestamp 1669390400
transform 1 0 27587 0 1 34265
box -42 -42 29342 342
use M1_PSUB43105908781107_256x8m81  M1_PSUB43105908781107_256x8m81_0
timestamp 1669390400
transform 1 0 56133 0 1 36019
box -42 -42 842 31342
use M1_PSUB43105908781107_256x8m81  M1_PSUB43105908781107_256x8m81_1
timestamp 1669390400
transform 1 0 27587 0 1 36019
box -42 -42 842 31342
use M1_PSUB43105908781108_256x8m81  M1_PSUB43105908781108_256x8m81_0
timestamp 1669390400
transform 1 0 112 0 1 67488
box -42 -42 85602 414
use M1_PSUB43105908781108_256x8m81  M1_PSUB43105908781108_256x8m81_1
timestamp 1669390400
transform 1 0 112 0 1 620
box -42 -42 85602 414
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2141308
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2140054
string path 4.620 11.160 4.620 0.000 
<< end >>
