magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 2021 89 2091
rect -31 -71 89 -1
use nmos_5p04310590548799_128x8m81  nmos_5p04310590548799_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 2066
<< properties >>
string GDS_END 1700688
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1700438
<< end >>
