magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -817 23 817 79
rect -817 -23 -758 23
rect -712 -23 -595 23
rect -549 -23 -431 23
rect -385 -23 -268 23
rect -222 -23 -105 23
rect -59 -23 59 23
rect 105 -23 222 23
rect 268 -23 385 23
rect 431 -23 549 23
rect 595 -23 712 23
rect 758 -23 817 23
rect -817 -80 817 -23
<< psubdiffcont >>
rect -758 -23 -712 23
rect -595 -23 -549 23
rect -431 -23 -385 23
rect -268 -23 -222 23
rect -105 -23 -59 23
rect 59 -23 105 23
rect 222 -23 268 23
rect 385 -23 431 23
rect 549 -23 595 23
rect 712 -23 758 23
<< metal1 >>
rect -808 23 808 70
rect -808 -23 -758 23
rect -712 -23 -595 23
rect -549 -23 -431 23
rect -385 -23 -268 23
rect -222 -23 -105 23
rect -59 -23 59 23
rect 105 -23 222 23
rect 268 -23 385 23
rect 431 -23 549 23
rect 595 -23 712 23
rect 758 -23 808 23
rect -808 -71 808 -23
<< properties >>
string GDS_END 228818
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 227950
<< end >>
