magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 1361 89 1434
rect -31 -74 89 -1
use nmos_5p0431059087812_256x8m81  nmos_5p0431059087812_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 1406
<< properties >>
string GDS_END 46672
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 46422
<< end >>
