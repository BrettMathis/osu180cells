magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1008 844
rect 49 528 95 724
rect 244 536 316 676
rect 457 617 503 724
rect 661 536 707 676
rect 865 617 911 724
rect 244 472 898 536
rect 124 360 806 424
rect 124 248 632 312
rect 852 307 898 472
rect 692 253 898 307
rect 692 200 764 253
rect 49 60 95 181
rect 430 136 764 200
rect 852 60 924 127
rect 0 -60 1008 60
<< labels >>
rlabel metal1 s 124 248 632 312 6 A1
port 1 nsew default input
rlabel metal1 s 124 360 806 424 6 A2
port 2 nsew default input
rlabel metal1 s 661 536 707 676 6 ZN
port 3 nsew default output
rlabel metal1 s 244 536 316 676 6 ZN
port 3 nsew default output
rlabel metal1 s 244 472 898 536 6 ZN
port 3 nsew default output
rlabel metal1 s 852 307 898 472 6 ZN
port 3 nsew default output
rlabel metal1 s 692 253 898 307 6 ZN
port 3 nsew default output
rlabel metal1 s 692 200 764 253 6 ZN
port 3 nsew default output
rlabel metal1 s 430 136 764 200 6 ZN
port 3 nsew default output
rlabel metal1 s 0 724 1008 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 865 617 911 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 457 617 503 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 49 617 95 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 49 528 95 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 49 127 95 181 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 852 60 924 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1008 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1008 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 691406
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 688316
<< end >>
