magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -5784 1125 5784 1144
rect -5784 1079 -5765 1125
rect -5719 1079 -5649 1125
rect -5603 1079 -5533 1125
rect -5487 1079 -5417 1125
rect -5371 1079 -5301 1125
rect -5255 1079 -5185 1125
rect -5139 1079 -5069 1125
rect -5023 1079 -4953 1125
rect -4907 1079 -4837 1125
rect -4791 1079 -4721 1125
rect -4675 1079 -4605 1125
rect -4559 1079 -4489 1125
rect -4443 1079 -4373 1125
rect -4327 1079 -4257 1125
rect -4211 1079 -4141 1125
rect -4095 1079 -4025 1125
rect -3979 1079 -3909 1125
rect -3863 1079 -3793 1125
rect -3747 1079 -3677 1125
rect -3631 1079 -3561 1125
rect -3515 1079 -3445 1125
rect -3399 1079 -3329 1125
rect -3283 1079 -3213 1125
rect -3167 1079 -3097 1125
rect -3051 1079 -2981 1125
rect -2935 1079 -2865 1125
rect -2819 1079 -2749 1125
rect -2703 1079 -2633 1125
rect -2587 1079 -2517 1125
rect -2471 1079 -2401 1125
rect -2355 1079 -2285 1125
rect -2239 1079 -2169 1125
rect -2123 1079 -2053 1125
rect -2007 1079 -1937 1125
rect -1891 1079 -1821 1125
rect -1775 1079 -1705 1125
rect -1659 1079 -1589 1125
rect -1543 1079 -1473 1125
rect -1427 1079 -1357 1125
rect -1311 1079 -1241 1125
rect -1195 1079 -1125 1125
rect -1079 1079 -1009 1125
rect -963 1079 -893 1125
rect -847 1079 -777 1125
rect -731 1079 -661 1125
rect -615 1079 -545 1125
rect -499 1079 -429 1125
rect -383 1079 -313 1125
rect -267 1079 -197 1125
rect -151 1079 -81 1125
rect -35 1079 35 1125
rect 81 1079 151 1125
rect 197 1079 267 1125
rect 313 1079 383 1125
rect 429 1079 499 1125
rect 545 1079 615 1125
rect 661 1079 731 1125
rect 777 1079 847 1125
rect 893 1079 963 1125
rect 1009 1079 1079 1125
rect 1125 1079 1195 1125
rect 1241 1079 1311 1125
rect 1357 1079 1427 1125
rect 1473 1079 1543 1125
rect 1589 1079 1659 1125
rect 1705 1079 1775 1125
rect 1821 1079 1891 1125
rect 1937 1079 2007 1125
rect 2053 1079 2123 1125
rect 2169 1079 2239 1125
rect 2285 1079 2355 1125
rect 2401 1079 2471 1125
rect 2517 1079 2587 1125
rect 2633 1079 2703 1125
rect 2749 1079 2819 1125
rect 2865 1079 2935 1125
rect 2981 1079 3051 1125
rect 3097 1079 3167 1125
rect 3213 1079 3283 1125
rect 3329 1079 3399 1125
rect 3445 1079 3515 1125
rect 3561 1079 3631 1125
rect 3677 1079 3747 1125
rect 3793 1079 3863 1125
rect 3909 1079 3979 1125
rect 4025 1079 4095 1125
rect 4141 1079 4211 1125
rect 4257 1079 4327 1125
rect 4373 1079 4443 1125
rect 4489 1079 4559 1125
rect 4605 1079 4675 1125
rect 4721 1079 4791 1125
rect 4837 1079 4907 1125
rect 4953 1079 5023 1125
rect 5069 1079 5139 1125
rect 5185 1079 5255 1125
rect 5301 1079 5371 1125
rect 5417 1079 5487 1125
rect 5533 1079 5603 1125
rect 5649 1079 5719 1125
rect 5765 1079 5784 1125
rect -5784 1009 5784 1079
rect -5784 963 -5765 1009
rect -5719 963 -5649 1009
rect -5603 963 -5533 1009
rect -5487 963 -5417 1009
rect -5371 963 -5301 1009
rect -5255 963 -5185 1009
rect -5139 963 -5069 1009
rect -5023 963 -4953 1009
rect -4907 963 -4837 1009
rect -4791 963 -4721 1009
rect -4675 963 -4605 1009
rect -4559 963 -4489 1009
rect -4443 963 -4373 1009
rect -4327 963 -4257 1009
rect -4211 963 -4141 1009
rect -4095 963 -4025 1009
rect -3979 963 -3909 1009
rect -3863 963 -3793 1009
rect -3747 963 -3677 1009
rect -3631 963 -3561 1009
rect -3515 963 -3445 1009
rect -3399 963 -3329 1009
rect -3283 963 -3213 1009
rect -3167 963 -3097 1009
rect -3051 963 -2981 1009
rect -2935 963 -2865 1009
rect -2819 963 -2749 1009
rect -2703 963 -2633 1009
rect -2587 963 -2517 1009
rect -2471 963 -2401 1009
rect -2355 963 -2285 1009
rect -2239 963 -2169 1009
rect -2123 963 -2053 1009
rect -2007 963 -1937 1009
rect -1891 963 -1821 1009
rect -1775 963 -1705 1009
rect -1659 963 -1589 1009
rect -1543 963 -1473 1009
rect -1427 963 -1357 1009
rect -1311 963 -1241 1009
rect -1195 963 -1125 1009
rect -1079 963 -1009 1009
rect -963 963 -893 1009
rect -847 963 -777 1009
rect -731 963 -661 1009
rect -615 963 -545 1009
rect -499 963 -429 1009
rect -383 963 -313 1009
rect -267 963 -197 1009
rect -151 963 -81 1009
rect -35 963 35 1009
rect 81 963 151 1009
rect 197 963 267 1009
rect 313 963 383 1009
rect 429 963 499 1009
rect 545 963 615 1009
rect 661 963 731 1009
rect 777 963 847 1009
rect 893 963 963 1009
rect 1009 963 1079 1009
rect 1125 963 1195 1009
rect 1241 963 1311 1009
rect 1357 963 1427 1009
rect 1473 963 1543 1009
rect 1589 963 1659 1009
rect 1705 963 1775 1009
rect 1821 963 1891 1009
rect 1937 963 2007 1009
rect 2053 963 2123 1009
rect 2169 963 2239 1009
rect 2285 963 2355 1009
rect 2401 963 2471 1009
rect 2517 963 2587 1009
rect 2633 963 2703 1009
rect 2749 963 2819 1009
rect 2865 963 2935 1009
rect 2981 963 3051 1009
rect 3097 963 3167 1009
rect 3213 963 3283 1009
rect 3329 963 3399 1009
rect 3445 963 3515 1009
rect 3561 963 3631 1009
rect 3677 963 3747 1009
rect 3793 963 3863 1009
rect 3909 963 3979 1009
rect 4025 963 4095 1009
rect 4141 963 4211 1009
rect 4257 963 4327 1009
rect 4373 963 4443 1009
rect 4489 963 4559 1009
rect 4605 963 4675 1009
rect 4721 963 4791 1009
rect 4837 963 4907 1009
rect 4953 963 5023 1009
rect 5069 963 5139 1009
rect 5185 963 5255 1009
rect 5301 963 5371 1009
rect 5417 963 5487 1009
rect 5533 963 5603 1009
rect 5649 963 5719 1009
rect 5765 963 5784 1009
rect -5784 893 5784 963
rect -5784 847 -5765 893
rect -5719 847 -5649 893
rect -5603 847 -5533 893
rect -5487 847 -5417 893
rect -5371 847 -5301 893
rect -5255 847 -5185 893
rect -5139 847 -5069 893
rect -5023 847 -4953 893
rect -4907 847 -4837 893
rect -4791 847 -4721 893
rect -4675 847 -4605 893
rect -4559 847 -4489 893
rect -4443 847 -4373 893
rect -4327 847 -4257 893
rect -4211 847 -4141 893
rect -4095 847 -4025 893
rect -3979 847 -3909 893
rect -3863 847 -3793 893
rect -3747 847 -3677 893
rect -3631 847 -3561 893
rect -3515 847 -3445 893
rect -3399 847 -3329 893
rect -3283 847 -3213 893
rect -3167 847 -3097 893
rect -3051 847 -2981 893
rect -2935 847 -2865 893
rect -2819 847 -2749 893
rect -2703 847 -2633 893
rect -2587 847 -2517 893
rect -2471 847 -2401 893
rect -2355 847 -2285 893
rect -2239 847 -2169 893
rect -2123 847 -2053 893
rect -2007 847 -1937 893
rect -1891 847 -1821 893
rect -1775 847 -1705 893
rect -1659 847 -1589 893
rect -1543 847 -1473 893
rect -1427 847 -1357 893
rect -1311 847 -1241 893
rect -1195 847 -1125 893
rect -1079 847 -1009 893
rect -963 847 -893 893
rect -847 847 -777 893
rect -731 847 -661 893
rect -615 847 -545 893
rect -499 847 -429 893
rect -383 847 -313 893
rect -267 847 -197 893
rect -151 847 -81 893
rect -35 847 35 893
rect 81 847 151 893
rect 197 847 267 893
rect 313 847 383 893
rect 429 847 499 893
rect 545 847 615 893
rect 661 847 731 893
rect 777 847 847 893
rect 893 847 963 893
rect 1009 847 1079 893
rect 1125 847 1195 893
rect 1241 847 1311 893
rect 1357 847 1427 893
rect 1473 847 1543 893
rect 1589 847 1659 893
rect 1705 847 1775 893
rect 1821 847 1891 893
rect 1937 847 2007 893
rect 2053 847 2123 893
rect 2169 847 2239 893
rect 2285 847 2355 893
rect 2401 847 2471 893
rect 2517 847 2587 893
rect 2633 847 2703 893
rect 2749 847 2819 893
rect 2865 847 2935 893
rect 2981 847 3051 893
rect 3097 847 3167 893
rect 3213 847 3283 893
rect 3329 847 3399 893
rect 3445 847 3515 893
rect 3561 847 3631 893
rect 3677 847 3747 893
rect 3793 847 3863 893
rect 3909 847 3979 893
rect 4025 847 4095 893
rect 4141 847 4211 893
rect 4257 847 4327 893
rect 4373 847 4443 893
rect 4489 847 4559 893
rect 4605 847 4675 893
rect 4721 847 4791 893
rect 4837 847 4907 893
rect 4953 847 5023 893
rect 5069 847 5139 893
rect 5185 847 5255 893
rect 5301 847 5371 893
rect 5417 847 5487 893
rect 5533 847 5603 893
rect 5649 847 5719 893
rect 5765 847 5784 893
rect -5784 777 5784 847
rect -5784 731 -5765 777
rect -5719 731 -5649 777
rect -5603 731 -5533 777
rect -5487 731 -5417 777
rect -5371 731 -5301 777
rect -5255 731 -5185 777
rect -5139 731 -5069 777
rect -5023 731 -4953 777
rect -4907 731 -4837 777
rect -4791 731 -4721 777
rect -4675 731 -4605 777
rect -4559 731 -4489 777
rect -4443 731 -4373 777
rect -4327 731 -4257 777
rect -4211 731 -4141 777
rect -4095 731 -4025 777
rect -3979 731 -3909 777
rect -3863 731 -3793 777
rect -3747 731 -3677 777
rect -3631 731 -3561 777
rect -3515 731 -3445 777
rect -3399 731 -3329 777
rect -3283 731 -3213 777
rect -3167 731 -3097 777
rect -3051 731 -2981 777
rect -2935 731 -2865 777
rect -2819 731 -2749 777
rect -2703 731 -2633 777
rect -2587 731 -2517 777
rect -2471 731 -2401 777
rect -2355 731 -2285 777
rect -2239 731 -2169 777
rect -2123 731 -2053 777
rect -2007 731 -1937 777
rect -1891 731 -1821 777
rect -1775 731 -1705 777
rect -1659 731 -1589 777
rect -1543 731 -1473 777
rect -1427 731 -1357 777
rect -1311 731 -1241 777
rect -1195 731 -1125 777
rect -1079 731 -1009 777
rect -963 731 -893 777
rect -847 731 -777 777
rect -731 731 -661 777
rect -615 731 -545 777
rect -499 731 -429 777
rect -383 731 -313 777
rect -267 731 -197 777
rect -151 731 -81 777
rect -35 731 35 777
rect 81 731 151 777
rect 197 731 267 777
rect 313 731 383 777
rect 429 731 499 777
rect 545 731 615 777
rect 661 731 731 777
rect 777 731 847 777
rect 893 731 963 777
rect 1009 731 1079 777
rect 1125 731 1195 777
rect 1241 731 1311 777
rect 1357 731 1427 777
rect 1473 731 1543 777
rect 1589 731 1659 777
rect 1705 731 1775 777
rect 1821 731 1891 777
rect 1937 731 2007 777
rect 2053 731 2123 777
rect 2169 731 2239 777
rect 2285 731 2355 777
rect 2401 731 2471 777
rect 2517 731 2587 777
rect 2633 731 2703 777
rect 2749 731 2819 777
rect 2865 731 2935 777
rect 2981 731 3051 777
rect 3097 731 3167 777
rect 3213 731 3283 777
rect 3329 731 3399 777
rect 3445 731 3515 777
rect 3561 731 3631 777
rect 3677 731 3747 777
rect 3793 731 3863 777
rect 3909 731 3979 777
rect 4025 731 4095 777
rect 4141 731 4211 777
rect 4257 731 4327 777
rect 4373 731 4443 777
rect 4489 731 4559 777
rect 4605 731 4675 777
rect 4721 731 4791 777
rect 4837 731 4907 777
rect 4953 731 5023 777
rect 5069 731 5139 777
rect 5185 731 5255 777
rect 5301 731 5371 777
rect 5417 731 5487 777
rect 5533 731 5603 777
rect 5649 731 5719 777
rect 5765 731 5784 777
rect -5784 661 5784 731
rect -5784 615 -5765 661
rect -5719 615 -5649 661
rect -5603 615 -5533 661
rect -5487 615 -5417 661
rect -5371 615 -5301 661
rect -5255 615 -5185 661
rect -5139 615 -5069 661
rect -5023 615 -4953 661
rect -4907 615 -4837 661
rect -4791 615 -4721 661
rect -4675 615 -4605 661
rect -4559 615 -4489 661
rect -4443 615 -4373 661
rect -4327 615 -4257 661
rect -4211 615 -4141 661
rect -4095 615 -4025 661
rect -3979 615 -3909 661
rect -3863 615 -3793 661
rect -3747 615 -3677 661
rect -3631 615 -3561 661
rect -3515 615 -3445 661
rect -3399 615 -3329 661
rect -3283 615 -3213 661
rect -3167 615 -3097 661
rect -3051 615 -2981 661
rect -2935 615 -2865 661
rect -2819 615 -2749 661
rect -2703 615 -2633 661
rect -2587 615 -2517 661
rect -2471 615 -2401 661
rect -2355 615 -2285 661
rect -2239 615 -2169 661
rect -2123 615 -2053 661
rect -2007 615 -1937 661
rect -1891 615 -1821 661
rect -1775 615 -1705 661
rect -1659 615 -1589 661
rect -1543 615 -1473 661
rect -1427 615 -1357 661
rect -1311 615 -1241 661
rect -1195 615 -1125 661
rect -1079 615 -1009 661
rect -963 615 -893 661
rect -847 615 -777 661
rect -731 615 -661 661
rect -615 615 -545 661
rect -499 615 -429 661
rect -383 615 -313 661
rect -267 615 -197 661
rect -151 615 -81 661
rect -35 615 35 661
rect 81 615 151 661
rect 197 615 267 661
rect 313 615 383 661
rect 429 615 499 661
rect 545 615 615 661
rect 661 615 731 661
rect 777 615 847 661
rect 893 615 963 661
rect 1009 615 1079 661
rect 1125 615 1195 661
rect 1241 615 1311 661
rect 1357 615 1427 661
rect 1473 615 1543 661
rect 1589 615 1659 661
rect 1705 615 1775 661
rect 1821 615 1891 661
rect 1937 615 2007 661
rect 2053 615 2123 661
rect 2169 615 2239 661
rect 2285 615 2355 661
rect 2401 615 2471 661
rect 2517 615 2587 661
rect 2633 615 2703 661
rect 2749 615 2819 661
rect 2865 615 2935 661
rect 2981 615 3051 661
rect 3097 615 3167 661
rect 3213 615 3283 661
rect 3329 615 3399 661
rect 3445 615 3515 661
rect 3561 615 3631 661
rect 3677 615 3747 661
rect 3793 615 3863 661
rect 3909 615 3979 661
rect 4025 615 4095 661
rect 4141 615 4211 661
rect 4257 615 4327 661
rect 4373 615 4443 661
rect 4489 615 4559 661
rect 4605 615 4675 661
rect 4721 615 4791 661
rect 4837 615 4907 661
rect 4953 615 5023 661
rect 5069 615 5139 661
rect 5185 615 5255 661
rect 5301 615 5371 661
rect 5417 615 5487 661
rect 5533 615 5603 661
rect 5649 615 5719 661
rect 5765 615 5784 661
rect -5784 545 5784 615
rect -5784 499 -5765 545
rect -5719 499 -5649 545
rect -5603 499 -5533 545
rect -5487 499 -5417 545
rect -5371 499 -5301 545
rect -5255 499 -5185 545
rect -5139 499 -5069 545
rect -5023 499 -4953 545
rect -4907 499 -4837 545
rect -4791 499 -4721 545
rect -4675 499 -4605 545
rect -4559 499 -4489 545
rect -4443 499 -4373 545
rect -4327 499 -4257 545
rect -4211 499 -4141 545
rect -4095 499 -4025 545
rect -3979 499 -3909 545
rect -3863 499 -3793 545
rect -3747 499 -3677 545
rect -3631 499 -3561 545
rect -3515 499 -3445 545
rect -3399 499 -3329 545
rect -3283 499 -3213 545
rect -3167 499 -3097 545
rect -3051 499 -2981 545
rect -2935 499 -2865 545
rect -2819 499 -2749 545
rect -2703 499 -2633 545
rect -2587 499 -2517 545
rect -2471 499 -2401 545
rect -2355 499 -2285 545
rect -2239 499 -2169 545
rect -2123 499 -2053 545
rect -2007 499 -1937 545
rect -1891 499 -1821 545
rect -1775 499 -1705 545
rect -1659 499 -1589 545
rect -1543 499 -1473 545
rect -1427 499 -1357 545
rect -1311 499 -1241 545
rect -1195 499 -1125 545
rect -1079 499 -1009 545
rect -963 499 -893 545
rect -847 499 -777 545
rect -731 499 -661 545
rect -615 499 -545 545
rect -499 499 -429 545
rect -383 499 -313 545
rect -267 499 -197 545
rect -151 499 -81 545
rect -35 499 35 545
rect 81 499 151 545
rect 197 499 267 545
rect 313 499 383 545
rect 429 499 499 545
rect 545 499 615 545
rect 661 499 731 545
rect 777 499 847 545
rect 893 499 963 545
rect 1009 499 1079 545
rect 1125 499 1195 545
rect 1241 499 1311 545
rect 1357 499 1427 545
rect 1473 499 1543 545
rect 1589 499 1659 545
rect 1705 499 1775 545
rect 1821 499 1891 545
rect 1937 499 2007 545
rect 2053 499 2123 545
rect 2169 499 2239 545
rect 2285 499 2355 545
rect 2401 499 2471 545
rect 2517 499 2587 545
rect 2633 499 2703 545
rect 2749 499 2819 545
rect 2865 499 2935 545
rect 2981 499 3051 545
rect 3097 499 3167 545
rect 3213 499 3283 545
rect 3329 499 3399 545
rect 3445 499 3515 545
rect 3561 499 3631 545
rect 3677 499 3747 545
rect 3793 499 3863 545
rect 3909 499 3979 545
rect 4025 499 4095 545
rect 4141 499 4211 545
rect 4257 499 4327 545
rect 4373 499 4443 545
rect 4489 499 4559 545
rect 4605 499 4675 545
rect 4721 499 4791 545
rect 4837 499 4907 545
rect 4953 499 5023 545
rect 5069 499 5139 545
rect 5185 499 5255 545
rect 5301 499 5371 545
rect 5417 499 5487 545
rect 5533 499 5603 545
rect 5649 499 5719 545
rect 5765 499 5784 545
rect -5784 429 5784 499
rect -5784 383 -5765 429
rect -5719 383 -5649 429
rect -5603 383 -5533 429
rect -5487 383 -5417 429
rect -5371 383 -5301 429
rect -5255 383 -5185 429
rect -5139 383 -5069 429
rect -5023 383 -4953 429
rect -4907 383 -4837 429
rect -4791 383 -4721 429
rect -4675 383 -4605 429
rect -4559 383 -4489 429
rect -4443 383 -4373 429
rect -4327 383 -4257 429
rect -4211 383 -4141 429
rect -4095 383 -4025 429
rect -3979 383 -3909 429
rect -3863 383 -3793 429
rect -3747 383 -3677 429
rect -3631 383 -3561 429
rect -3515 383 -3445 429
rect -3399 383 -3329 429
rect -3283 383 -3213 429
rect -3167 383 -3097 429
rect -3051 383 -2981 429
rect -2935 383 -2865 429
rect -2819 383 -2749 429
rect -2703 383 -2633 429
rect -2587 383 -2517 429
rect -2471 383 -2401 429
rect -2355 383 -2285 429
rect -2239 383 -2169 429
rect -2123 383 -2053 429
rect -2007 383 -1937 429
rect -1891 383 -1821 429
rect -1775 383 -1705 429
rect -1659 383 -1589 429
rect -1543 383 -1473 429
rect -1427 383 -1357 429
rect -1311 383 -1241 429
rect -1195 383 -1125 429
rect -1079 383 -1009 429
rect -963 383 -893 429
rect -847 383 -777 429
rect -731 383 -661 429
rect -615 383 -545 429
rect -499 383 -429 429
rect -383 383 -313 429
rect -267 383 -197 429
rect -151 383 -81 429
rect -35 383 35 429
rect 81 383 151 429
rect 197 383 267 429
rect 313 383 383 429
rect 429 383 499 429
rect 545 383 615 429
rect 661 383 731 429
rect 777 383 847 429
rect 893 383 963 429
rect 1009 383 1079 429
rect 1125 383 1195 429
rect 1241 383 1311 429
rect 1357 383 1427 429
rect 1473 383 1543 429
rect 1589 383 1659 429
rect 1705 383 1775 429
rect 1821 383 1891 429
rect 1937 383 2007 429
rect 2053 383 2123 429
rect 2169 383 2239 429
rect 2285 383 2355 429
rect 2401 383 2471 429
rect 2517 383 2587 429
rect 2633 383 2703 429
rect 2749 383 2819 429
rect 2865 383 2935 429
rect 2981 383 3051 429
rect 3097 383 3167 429
rect 3213 383 3283 429
rect 3329 383 3399 429
rect 3445 383 3515 429
rect 3561 383 3631 429
rect 3677 383 3747 429
rect 3793 383 3863 429
rect 3909 383 3979 429
rect 4025 383 4095 429
rect 4141 383 4211 429
rect 4257 383 4327 429
rect 4373 383 4443 429
rect 4489 383 4559 429
rect 4605 383 4675 429
rect 4721 383 4791 429
rect 4837 383 4907 429
rect 4953 383 5023 429
rect 5069 383 5139 429
rect 5185 383 5255 429
rect 5301 383 5371 429
rect 5417 383 5487 429
rect 5533 383 5603 429
rect 5649 383 5719 429
rect 5765 383 5784 429
rect -5784 313 5784 383
rect -5784 267 -5765 313
rect -5719 267 -5649 313
rect -5603 267 -5533 313
rect -5487 267 -5417 313
rect -5371 267 -5301 313
rect -5255 267 -5185 313
rect -5139 267 -5069 313
rect -5023 267 -4953 313
rect -4907 267 -4837 313
rect -4791 267 -4721 313
rect -4675 267 -4605 313
rect -4559 267 -4489 313
rect -4443 267 -4373 313
rect -4327 267 -4257 313
rect -4211 267 -4141 313
rect -4095 267 -4025 313
rect -3979 267 -3909 313
rect -3863 267 -3793 313
rect -3747 267 -3677 313
rect -3631 267 -3561 313
rect -3515 267 -3445 313
rect -3399 267 -3329 313
rect -3283 267 -3213 313
rect -3167 267 -3097 313
rect -3051 267 -2981 313
rect -2935 267 -2865 313
rect -2819 267 -2749 313
rect -2703 267 -2633 313
rect -2587 267 -2517 313
rect -2471 267 -2401 313
rect -2355 267 -2285 313
rect -2239 267 -2169 313
rect -2123 267 -2053 313
rect -2007 267 -1937 313
rect -1891 267 -1821 313
rect -1775 267 -1705 313
rect -1659 267 -1589 313
rect -1543 267 -1473 313
rect -1427 267 -1357 313
rect -1311 267 -1241 313
rect -1195 267 -1125 313
rect -1079 267 -1009 313
rect -963 267 -893 313
rect -847 267 -777 313
rect -731 267 -661 313
rect -615 267 -545 313
rect -499 267 -429 313
rect -383 267 -313 313
rect -267 267 -197 313
rect -151 267 -81 313
rect -35 267 35 313
rect 81 267 151 313
rect 197 267 267 313
rect 313 267 383 313
rect 429 267 499 313
rect 545 267 615 313
rect 661 267 731 313
rect 777 267 847 313
rect 893 267 963 313
rect 1009 267 1079 313
rect 1125 267 1195 313
rect 1241 267 1311 313
rect 1357 267 1427 313
rect 1473 267 1543 313
rect 1589 267 1659 313
rect 1705 267 1775 313
rect 1821 267 1891 313
rect 1937 267 2007 313
rect 2053 267 2123 313
rect 2169 267 2239 313
rect 2285 267 2355 313
rect 2401 267 2471 313
rect 2517 267 2587 313
rect 2633 267 2703 313
rect 2749 267 2819 313
rect 2865 267 2935 313
rect 2981 267 3051 313
rect 3097 267 3167 313
rect 3213 267 3283 313
rect 3329 267 3399 313
rect 3445 267 3515 313
rect 3561 267 3631 313
rect 3677 267 3747 313
rect 3793 267 3863 313
rect 3909 267 3979 313
rect 4025 267 4095 313
rect 4141 267 4211 313
rect 4257 267 4327 313
rect 4373 267 4443 313
rect 4489 267 4559 313
rect 4605 267 4675 313
rect 4721 267 4791 313
rect 4837 267 4907 313
rect 4953 267 5023 313
rect 5069 267 5139 313
rect 5185 267 5255 313
rect 5301 267 5371 313
rect 5417 267 5487 313
rect 5533 267 5603 313
rect 5649 267 5719 313
rect 5765 267 5784 313
rect -5784 197 5784 267
rect -5784 151 -5765 197
rect -5719 151 -5649 197
rect -5603 151 -5533 197
rect -5487 151 -5417 197
rect -5371 151 -5301 197
rect -5255 151 -5185 197
rect -5139 151 -5069 197
rect -5023 151 -4953 197
rect -4907 151 -4837 197
rect -4791 151 -4721 197
rect -4675 151 -4605 197
rect -4559 151 -4489 197
rect -4443 151 -4373 197
rect -4327 151 -4257 197
rect -4211 151 -4141 197
rect -4095 151 -4025 197
rect -3979 151 -3909 197
rect -3863 151 -3793 197
rect -3747 151 -3677 197
rect -3631 151 -3561 197
rect -3515 151 -3445 197
rect -3399 151 -3329 197
rect -3283 151 -3213 197
rect -3167 151 -3097 197
rect -3051 151 -2981 197
rect -2935 151 -2865 197
rect -2819 151 -2749 197
rect -2703 151 -2633 197
rect -2587 151 -2517 197
rect -2471 151 -2401 197
rect -2355 151 -2285 197
rect -2239 151 -2169 197
rect -2123 151 -2053 197
rect -2007 151 -1937 197
rect -1891 151 -1821 197
rect -1775 151 -1705 197
rect -1659 151 -1589 197
rect -1543 151 -1473 197
rect -1427 151 -1357 197
rect -1311 151 -1241 197
rect -1195 151 -1125 197
rect -1079 151 -1009 197
rect -963 151 -893 197
rect -847 151 -777 197
rect -731 151 -661 197
rect -615 151 -545 197
rect -499 151 -429 197
rect -383 151 -313 197
rect -267 151 -197 197
rect -151 151 -81 197
rect -35 151 35 197
rect 81 151 151 197
rect 197 151 267 197
rect 313 151 383 197
rect 429 151 499 197
rect 545 151 615 197
rect 661 151 731 197
rect 777 151 847 197
rect 893 151 963 197
rect 1009 151 1079 197
rect 1125 151 1195 197
rect 1241 151 1311 197
rect 1357 151 1427 197
rect 1473 151 1543 197
rect 1589 151 1659 197
rect 1705 151 1775 197
rect 1821 151 1891 197
rect 1937 151 2007 197
rect 2053 151 2123 197
rect 2169 151 2239 197
rect 2285 151 2355 197
rect 2401 151 2471 197
rect 2517 151 2587 197
rect 2633 151 2703 197
rect 2749 151 2819 197
rect 2865 151 2935 197
rect 2981 151 3051 197
rect 3097 151 3167 197
rect 3213 151 3283 197
rect 3329 151 3399 197
rect 3445 151 3515 197
rect 3561 151 3631 197
rect 3677 151 3747 197
rect 3793 151 3863 197
rect 3909 151 3979 197
rect 4025 151 4095 197
rect 4141 151 4211 197
rect 4257 151 4327 197
rect 4373 151 4443 197
rect 4489 151 4559 197
rect 4605 151 4675 197
rect 4721 151 4791 197
rect 4837 151 4907 197
rect 4953 151 5023 197
rect 5069 151 5139 197
rect 5185 151 5255 197
rect 5301 151 5371 197
rect 5417 151 5487 197
rect 5533 151 5603 197
rect 5649 151 5719 197
rect 5765 151 5784 197
rect -5784 81 5784 151
rect -5784 35 -5765 81
rect -5719 35 -5649 81
rect -5603 35 -5533 81
rect -5487 35 -5417 81
rect -5371 35 -5301 81
rect -5255 35 -5185 81
rect -5139 35 -5069 81
rect -5023 35 -4953 81
rect -4907 35 -4837 81
rect -4791 35 -4721 81
rect -4675 35 -4605 81
rect -4559 35 -4489 81
rect -4443 35 -4373 81
rect -4327 35 -4257 81
rect -4211 35 -4141 81
rect -4095 35 -4025 81
rect -3979 35 -3909 81
rect -3863 35 -3793 81
rect -3747 35 -3677 81
rect -3631 35 -3561 81
rect -3515 35 -3445 81
rect -3399 35 -3329 81
rect -3283 35 -3213 81
rect -3167 35 -3097 81
rect -3051 35 -2981 81
rect -2935 35 -2865 81
rect -2819 35 -2749 81
rect -2703 35 -2633 81
rect -2587 35 -2517 81
rect -2471 35 -2401 81
rect -2355 35 -2285 81
rect -2239 35 -2169 81
rect -2123 35 -2053 81
rect -2007 35 -1937 81
rect -1891 35 -1821 81
rect -1775 35 -1705 81
rect -1659 35 -1589 81
rect -1543 35 -1473 81
rect -1427 35 -1357 81
rect -1311 35 -1241 81
rect -1195 35 -1125 81
rect -1079 35 -1009 81
rect -963 35 -893 81
rect -847 35 -777 81
rect -731 35 -661 81
rect -615 35 -545 81
rect -499 35 -429 81
rect -383 35 -313 81
rect -267 35 -197 81
rect -151 35 -81 81
rect -35 35 35 81
rect 81 35 151 81
rect 197 35 267 81
rect 313 35 383 81
rect 429 35 499 81
rect 545 35 615 81
rect 661 35 731 81
rect 777 35 847 81
rect 893 35 963 81
rect 1009 35 1079 81
rect 1125 35 1195 81
rect 1241 35 1311 81
rect 1357 35 1427 81
rect 1473 35 1543 81
rect 1589 35 1659 81
rect 1705 35 1775 81
rect 1821 35 1891 81
rect 1937 35 2007 81
rect 2053 35 2123 81
rect 2169 35 2239 81
rect 2285 35 2355 81
rect 2401 35 2471 81
rect 2517 35 2587 81
rect 2633 35 2703 81
rect 2749 35 2819 81
rect 2865 35 2935 81
rect 2981 35 3051 81
rect 3097 35 3167 81
rect 3213 35 3283 81
rect 3329 35 3399 81
rect 3445 35 3515 81
rect 3561 35 3631 81
rect 3677 35 3747 81
rect 3793 35 3863 81
rect 3909 35 3979 81
rect 4025 35 4095 81
rect 4141 35 4211 81
rect 4257 35 4327 81
rect 4373 35 4443 81
rect 4489 35 4559 81
rect 4605 35 4675 81
rect 4721 35 4791 81
rect 4837 35 4907 81
rect 4953 35 5023 81
rect 5069 35 5139 81
rect 5185 35 5255 81
rect 5301 35 5371 81
rect 5417 35 5487 81
rect 5533 35 5603 81
rect 5649 35 5719 81
rect 5765 35 5784 81
rect -5784 -35 5784 35
rect -5784 -81 -5765 -35
rect -5719 -81 -5649 -35
rect -5603 -81 -5533 -35
rect -5487 -81 -5417 -35
rect -5371 -81 -5301 -35
rect -5255 -81 -5185 -35
rect -5139 -81 -5069 -35
rect -5023 -81 -4953 -35
rect -4907 -81 -4837 -35
rect -4791 -81 -4721 -35
rect -4675 -81 -4605 -35
rect -4559 -81 -4489 -35
rect -4443 -81 -4373 -35
rect -4327 -81 -4257 -35
rect -4211 -81 -4141 -35
rect -4095 -81 -4025 -35
rect -3979 -81 -3909 -35
rect -3863 -81 -3793 -35
rect -3747 -81 -3677 -35
rect -3631 -81 -3561 -35
rect -3515 -81 -3445 -35
rect -3399 -81 -3329 -35
rect -3283 -81 -3213 -35
rect -3167 -81 -3097 -35
rect -3051 -81 -2981 -35
rect -2935 -81 -2865 -35
rect -2819 -81 -2749 -35
rect -2703 -81 -2633 -35
rect -2587 -81 -2517 -35
rect -2471 -81 -2401 -35
rect -2355 -81 -2285 -35
rect -2239 -81 -2169 -35
rect -2123 -81 -2053 -35
rect -2007 -81 -1937 -35
rect -1891 -81 -1821 -35
rect -1775 -81 -1705 -35
rect -1659 -81 -1589 -35
rect -1543 -81 -1473 -35
rect -1427 -81 -1357 -35
rect -1311 -81 -1241 -35
rect -1195 -81 -1125 -35
rect -1079 -81 -1009 -35
rect -963 -81 -893 -35
rect -847 -81 -777 -35
rect -731 -81 -661 -35
rect -615 -81 -545 -35
rect -499 -81 -429 -35
rect -383 -81 -313 -35
rect -267 -81 -197 -35
rect -151 -81 -81 -35
rect -35 -81 35 -35
rect 81 -81 151 -35
rect 197 -81 267 -35
rect 313 -81 383 -35
rect 429 -81 499 -35
rect 545 -81 615 -35
rect 661 -81 731 -35
rect 777 -81 847 -35
rect 893 -81 963 -35
rect 1009 -81 1079 -35
rect 1125 -81 1195 -35
rect 1241 -81 1311 -35
rect 1357 -81 1427 -35
rect 1473 -81 1543 -35
rect 1589 -81 1659 -35
rect 1705 -81 1775 -35
rect 1821 -81 1891 -35
rect 1937 -81 2007 -35
rect 2053 -81 2123 -35
rect 2169 -81 2239 -35
rect 2285 -81 2355 -35
rect 2401 -81 2471 -35
rect 2517 -81 2587 -35
rect 2633 -81 2703 -35
rect 2749 -81 2819 -35
rect 2865 -81 2935 -35
rect 2981 -81 3051 -35
rect 3097 -81 3167 -35
rect 3213 -81 3283 -35
rect 3329 -81 3399 -35
rect 3445 -81 3515 -35
rect 3561 -81 3631 -35
rect 3677 -81 3747 -35
rect 3793 -81 3863 -35
rect 3909 -81 3979 -35
rect 4025 -81 4095 -35
rect 4141 -81 4211 -35
rect 4257 -81 4327 -35
rect 4373 -81 4443 -35
rect 4489 -81 4559 -35
rect 4605 -81 4675 -35
rect 4721 -81 4791 -35
rect 4837 -81 4907 -35
rect 4953 -81 5023 -35
rect 5069 -81 5139 -35
rect 5185 -81 5255 -35
rect 5301 -81 5371 -35
rect 5417 -81 5487 -35
rect 5533 -81 5603 -35
rect 5649 -81 5719 -35
rect 5765 -81 5784 -35
rect -5784 -151 5784 -81
rect -5784 -197 -5765 -151
rect -5719 -197 -5649 -151
rect -5603 -197 -5533 -151
rect -5487 -197 -5417 -151
rect -5371 -197 -5301 -151
rect -5255 -197 -5185 -151
rect -5139 -197 -5069 -151
rect -5023 -197 -4953 -151
rect -4907 -197 -4837 -151
rect -4791 -197 -4721 -151
rect -4675 -197 -4605 -151
rect -4559 -197 -4489 -151
rect -4443 -197 -4373 -151
rect -4327 -197 -4257 -151
rect -4211 -197 -4141 -151
rect -4095 -197 -4025 -151
rect -3979 -197 -3909 -151
rect -3863 -197 -3793 -151
rect -3747 -197 -3677 -151
rect -3631 -197 -3561 -151
rect -3515 -197 -3445 -151
rect -3399 -197 -3329 -151
rect -3283 -197 -3213 -151
rect -3167 -197 -3097 -151
rect -3051 -197 -2981 -151
rect -2935 -197 -2865 -151
rect -2819 -197 -2749 -151
rect -2703 -197 -2633 -151
rect -2587 -197 -2517 -151
rect -2471 -197 -2401 -151
rect -2355 -197 -2285 -151
rect -2239 -197 -2169 -151
rect -2123 -197 -2053 -151
rect -2007 -197 -1937 -151
rect -1891 -197 -1821 -151
rect -1775 -197 -1705 -151
rect -1659 -197 -1589 -151
rect -1543 -197 -1473 -151
rect -1427 -197 -1357 -151
rect -1311 -197 -1241 -151
rect -1195 -197 -1125 -151
rect -1079 -197 -1009 -151
rect -963 -197 -893 -151
rect -847 -197 -777 -151
rect -731 -197 -661 -151
rect -615 -197 -545 -151
rect -499 -197 -429 -151
rect -383 -197 -313 -151
rect -267 -197 -197 -151
rect -151 -197 -81 -151
rect -35 -197 35 -151
rect 81 -197 151 -151
rect 197 -197 267 -151
rect 313 -197 383 -151
rect 429 -197 499 -151
rect 545 -197 615 -151
rect 661 -197 731 -151
rect 777 -197 847 -151
rect 893 -197 963 -151
rect 1009 -197 1079 -151
rect 1125 -197 1195 -151
rect 1241 -197 1311 -151
rect 1357 -197 1427 -151
rect 1473 -197 1543 -151
rect 1589 -197 1659 -151
rect 1705 -197 1775 -151
rect 1821 -197 1891 -151
rect 1937 -197 2007 -151
rect 2053 -197 2123 -151
rect 2169 -197 2239 -151
rect 2285 -197 2355 -151
rect 2401 -197 2471 -151
rect 2517 -197 2587 -151
rect 2633 -197 2703 -151
rect 2749 -197 2819 -151
rect 2865 -197 2935 -151
rect 2981 -197 3051 -151
rect 3097 -197 3167 -151
rect 3213 -197 3283 -151
rect 3329 -197 3399 -151
rect 3445 -197 3515 -151
rect 3561 -197 3631 -151
rect 3677 -197 3747 -151
rect 3793 -197 3863 -151
rect 3909 -197 3979 -151
rect 4025 -197 4095 -151
rect 4141 -197 4211 -151
rect 4257 -197 4327 -151
rect 4373 -197 4443 -151
rect 4489 -197 4559 -151
rect 4605 -197 4675 -151
rect 4721 -197 4791 -151
rect 4837 -197 4907 -151
rect 4953 -197 5023 -151
rect 5069 -197 5139 -151
rect 5185 -197 5255 -151
rect 5301 -197 5371 -151
rect 5417 -197 5487 -151
rect 5533 -197 5603 -151
rect 5649 -197 5719 -151
rect 5765 -197 5784 -151
rect -5784 -267 5784 -197
rect -5784 -313 -5765 -267
rect -5719 -313 -5649 -267
rect -5603 -313 -5533 -267
rect -5487 -313 -5417 -267
rect -5371 -313 -5301 -267
rect -5255 -313 -5185 -267
rect -5139 -313 -5069 -267
rect -5023 -313 -4953 -267
rect -4907 -313 -4837 -267
rect -4791 -313 -4721 -267
rect -4675 -313 -4605 -267
rect -4559 -313 -4489 -267
rect -4443 -313 -4373 -267
rect -4327 -313 -4257 -267
rect -4211 -313 -4141 -267
rect -4095 -313 -4025 -267
rect -3979 -313 -3909 -267
rect -3863 -313 -3793 -267
rect -3747 -313 -3677 -267
rect -3631 -313 -3561 -267
rect -3515 -313 -3445 -267
rect -3399 -313 -3329 -267
rect -3283 -313 -3213 -267
rect -3167 -313 -3097 -267
rect -3051 -313 -2981 -267
rect -2935 -313 -2865 -267
rect -2819 -313 -2749 -267
rect -2703 -313 -2633 -267
rect -2587 -313 -2517 -267
rect -2471 -313 -2401 -267
rect -2355 -313 -2285 -267
rect -2239 -313 -2169 -267
rect -2123 -313 -2053 -267
rect -2007 -313 -1937 -267
rect -1891 -313 -1821 -267
rect -1775 -313 -1705 -267
rect -1659 -313 -1589 -267
rect -1543 -313 -1473 -267
rect -1427 -313 -1357 -267
rect -1311 -313 -1241 -267
rect -1195 -313 -1125 -267
rect -1079 -313 -1009 -267
rect -963 -313 -893 -267
rect -847 -313 -777 -267
rect -731 -313 -661 -267
rect -615 -313 -545 -267
rect -499 -313 -429 -267
rect -383 -313 -313 -267
rect -267 -313 -197 -267
rect -151 -313 -81 -267
rect -35 -313 35 -267
rect 81 -313 151 -267
rect 197 -313 267 -267
rect 313 -313 383 -267
rect 429 -313 499 -267
rect 545 -313 615 -267
rect 661 -313 731 -267
rect 777 -313 847 -267
rect 893 -313 963 -267
rect 1009 -313 1079 -267
rect 1125 -313 1195 -267
rect 1241 -313 1311 -267
rect 1357 -313 1427 -267
rect 1473 -313 1543 -267
rect 1589 -313 1659 -267
rect 1705 -313 1775 -267
rect 1821 -313 1891 -267
rect 1937 -313 2007 -267
rect 2053 -313 2123 -267
rect 2169 -313 2239 -267
rect 2285 -313 2355 -267
rect 2401 -313 2471 -267
rect 2517 -313 2587 -267
rect 2633 -313 2703 -267
rect 2749 -313 2819 -267
rect 2865 -313 2935 -267
rect 2981 -313 3051 -267
rect 3097 -313 3167 -267
rect 3213 -313 3283 -267
rect 3329 -313 3399 -267
rect 3445 -313 3515 -267
rect 3561 -313 3631 -267
rect 3677 -313 3747 -267
rect 3793 -313 3863 -267
rect 3909 -313 3979 -267
rect 4025 -313 4095 -267
rect 4141 -313 4211 -267
rect 4257 -313 4327 -267
rect 4373 -313 4443 -267
rect 4489 -313 4559 -267
rect 4605 -313 4675 -267
rect 4721 -313 4791 -267
rect 4837 -313 4907 -267
rect 4953 -313 5023 -267
rect 5069 -313 5139 -267
rect 5185 -313 5255 -267
rect 5301 -313 5371 -267
rect 5417 -313 5487 -267
rect 5533 -313 5603 -267
rect 5649 -313 5719 -267
rect 5765 -313 5784 -267
rect -5784 -383 5784 -313
rect -5784 -429 -5765 -383
rect -5719 -429 -5649 -383
rect -5603 -429 -5533 -383
rect -5487 -429 -5417 -383
rect -5371 -429 -5301 -383
rect -5255 -429 -5185 -383
rect -5139 -429 -5069 -383
rect -5023 -429 -4953 -383
rect -4907 -429 -4837 -383
rect -4791 -429 -4721 -383
rect -4675 -429 -4605 -383
rect -4559 -429 -4489 -383
rect -4443 -429 -4373 -383
rect -4327 -429 -4257 -383
rect -4211 -429 -4141 -383
rect -4095 -429 -4025 -383
rect -3979 -429 -3909 -383
rect -3863 -429 -3793 -383
rect -3747 -429 -3677 -383
rect -3631 -429 -3561 -383
rect -3515 -429 -3445 -383
rect -3399 -429 -3329 -383
rect -3283 -429 -3213 -383
rect -3167 -429 -3097 -383
rect -3051 -429 -2981 -383
rect -2935 -429 -2865 -383
rect -2819 -429 -2749 -383
rect -2703 -429 -2633 -383
rect -2587 -429 -2517 -383
rect -2471 -429 -2401 -383
rect -2355 -429 -2285 -383
rect -2239 -429 -2169 -383
rect -2123 -429 -2053 -383
rect -2007 -429 -1937 -383
rect -1891 -429 -1821 -383
rect -1775 -429 -1705 -383
rect -1659 -429 -1589 -383
rect -1543 -429 -1473 -383
rect -1427 -429 -1357 -383
rect -1311 -429 -1241 -383
rect -1195 -429 -1125 -383
rect -1079 -429 -1009 -383
rect -963 -429 -893 -383
rect -847 -429 -777 -383
rect -731 -429 -661 -383
rect -615 -429 -545 -383
rect -499 -429 -429 -383
rect -383 -429 -313 -383
rect -267 -429 -197 -383
rect -151 -429 -81 -383
rect -35 -429 35 -383
rect 81 -429 151 -383
rect 197 -429 267 -383
rect 313 -429 383 -383
rect 429 -429 499 -383
rect 545 -429 615 -383
rect 661 -429 731 -383
rect 777 -429 847 -383
rect 893 -429 963 -383
rect 1009 -429 1079 -383
rect 1125 -429 1195 -383
rect 1241 -429 1311 -383
rect 1357 -429 1427 -383
rect 1473 -429 1543 -383
rect 1589 -429 1659 -383
rect 1705 -429 1775 -383
rect 1821 -429 1891 -383
rect 1937 -429 2007 -383
rect 2053 -429 2123 -383
rect 2169 -429 2239 -383
rect 2285 -429 2355 -383
rect 2401 -429 2471 -383
rect 2517 -429 2587 -383
rect 2633 -429 2703 -383
rect 2749 -429 2819 -383
rect 2865 -429 2935 -383
rect 2981 -429 3051 -383
rect 3097 -429 3167 -383
rect 3213 -429 3283 -383
rect 3329 -429 3399 -383
rect 3445 -429 3515 -383
rect 3561 -429 3631 -383
rect 3677 -429 3747 -383
rect 3793 -429 3863 -383
rect 3909 -429 3979 -383
rect 4025 -429 4095 -383
rect 4141 -429 4211 -383
rect 4257 -429 4327 -383
rect 4373 -429 4443 -383
rect 4489 -429 4559 -383
rect 4605 -429 4675 -383
rect 4721 -429 4791 -383
rect 4837 -429 4907 -383
rect 4953 -429 5023 -383
rect 5069 -429 5139 -383
rect 5185 -429 5255 -383
rect 5301 -429 5371 -383
rect 5417 -429 5487 -383
rect 5533 -429 5603 -383
rect 5649 -429 5719 -383
rect 5765 -429 5784 -383
rect -5784 -499 5784 -429
rect -5784 -545 -5765 -499
rect -5719 -545 -5649 -499
rect -5603 -545 -5533 -499
rect -5487 -545 -5417 -499
rect -5371 -545 -5301 -499
rect -5255 -545 -5185 -499
rect -5139 -545 -5069 -499
rect -5023 -545 -4953 -499
rect -4907 -545 -4837 -499
rect -4791 -545 -4721 -499
rect -4675 -545 -4605 -499
rect -4559 -545 -4489 -499
rect -4443 -545 -4373 -499
rect -4327 -545 -4257 -499
rect -4211 -545 -4141 -499
rect -4095 -545 -4025 -499
rect -3979 -545 -3909 -499
rect -3863 -545 -3793 -499
rect -3747 -545 -3677 -499
rect -3631 -545 -3561 -499
rect -3515 -545 -3445 -499
rect -3399 -545 -3329 -499
rect -3283 -545 -3213 -499
rect -3167 -545 -3097 -499
rect -3051 -545 -2981 -499
rect -2935 -545 -2865 -499
rect -2819 -545 -2749 -499
rect -2703 -545 -2633 -499
rect -2587 -545 -2517 -499
rect -2471 -545 -2401 -499
rect -2355 -545 -2285 -499
rect -2239 -545 -2169 -499
rect -2123 -545 -2053 -499
rect -2007 -545 -1937 -499
rect -1891 -545 -1821 -499
rect -1775 -545 -1705 -499
rect -1659 -545 -1589 -499
rect -1543 -545 -1473 -499
rect -1427 -545 -1357 -499
rect -1311 -545 -1241 -499
rect -1195 -545 -1125 -499
rect -1079 -545 -1009 -499
rect -963 -545 -893 -499
rect -847 -545 -777 -499
rect -731 -545 -661 -499
rect -615 -545 -545 -499
rect -499 -545 -429 -499
rect -383 -545 -313 -499
rect -267 -545 -197 -499
rect -151 -545 -81 -499
rect -35 -545 35 -499
rect 81 -545 151 -499
rect 197 -545 267 -499
rect 313 -545 383 -499
rect 429 -545 499 -499
rect 545 -545 615 -499
rect 661 -545 731 -499
rect 777 -545 847 -499
rect 893 -545 963 -499
rect 1009 -545 1079 -499
rect 1125 -545 1195 -499
rect 1241 -545 1311 -499
rect 1357 -545 1427 -499
rect 1473 -545 1543 -499
rect 1589 -545 1659 -499
rect 1705 -545 1775 -499
rect 1821 -545 1891 -499
rect 1937 -545 2007 -499
rect 2053 -545 2123 -499
rect 2169 -545 2239 -499
rect 2285 -545 2355 -499
rect 2401 -545 2471 -499
rect 2517 -545 2587 -499
rect 2633 -545 2703 -499
rect 2749 -545 2819 -499
rect 2865 -545 2935 -499
rect 2981 -545 3051 -499
rect 3097 -545 3167 -499
rect 3213 -545 3283 -499
rect 3329 -545 3399 -499
rect 3445 -545 3515 -499
rect 3561 -545 3631 -499
rect 3677 -545 3747 -499
rect 3793 -545 3863 -499
rect 3909 -545 3979 -499
rect 4025 -545 4095 -499
rect 4141 -545 4211 -499
rect 4257 -545 4327 -499
rect 4373 -545 4443 -499
rect 4489 -545 4559 -499
rect 4605 -545 4675 -499
rect 4721 -545 4791 -499
rect 4837 -545 4907 -499
rect 4953 -545 5023 -499
rect 5069 -545 5139 -499
rect 5185 -545 5255 -499
rect 5301 -545 5371 -499
rect 5417 -545 5487 -499
rect 5533 -545 5603 -499
rect 5649 -545 5719 -499
rect 5765 -545 5784 -499
rect -5784 -615 5784 -545
rect -5784 -661 -5765 -615
rect -5719 -661 -5649 -615
rect -5603 -661 -5533 -615
rect -5487 -661 -5417 -615
rect -5371 -661 -5301 -615
rect -5255 -661 -5185 -615
rect -5139 -661 -5069 -615
rect -5023 -661 -4953 -615
rect -4907 -661 -4837 -615
rect -4791 -661 -4721 -615
rect -4675 -661 -4605 -615
rect -4559 -661 -4489 -615
rect -4443 -661 -4373 -615
rect -4327 -661 -4257 -615
rect -4211 -661 -4141 -615
rect -4095 -661 -4025 -615
rect -3979 -661 -3909 -615
rect -3863 -661 -3793 -615
rect -3747 -661 -3677 -615
rect -3631 -661 -3561 -615
rect -3515 -661 -3445 -615
rect -3399 -661 -3329 -615
rect -3283 -661 -3213 -615
rect -3167 -661 -3097 -615
rect -3051 -661 -2981 -615
rect -2935 -661 -2865 -615
rect -2819 -661 -2749 -615
rect -2703 -661 -2633 -615
rect -2587 -661 -2517 -615
rect -2471 -661 -2401 -615
rect -2355 -661 -2285 -615
rect -2239 -661 -2169 -615
rect -2123 -661 -2053 -615
rect -2007 -661 -1937 -615
rect -1891 -661 -1821 -615
rect -1775 -661 -1705 -615
rect -1659 -661 -1589 -615
rect -1543 -661 -1473 -615
rect -1427 -661 -1357 -615
rect -1311 -661 -1241 -615
rect -1195 -661 -1125 -615
rect -1079 -661 -1009 -615
rect -963 -661 -893 -615
rect -847 -661 -777 -615
rect -731 -661 -661 -615
rect -615 -661 -545 -615
rect -499 -661 -429 -615
rect -383 -661 -313 -615
rect -267 -661 -197 -615
rect -151 -661 -81 -615
rect -35 -661 35 -615
rect 81 -661 151 -615
rect 197 -661 267 -615
rect 313 -661 383 -615
rect 429 -661 499 -615
rect 545 -661 615 -615
rect 661 -661 731 -615
rect 777 -661 847 -615
rect 893 -661 963 -615
rect 1009 -661 1079 -615
rect 1125 -661 1195 -615
rect 1241 -661 1311 -615
rect 1357 -661 1427 -615
rect 1473 -661 1543 -615
rect 1589 -661 1659 -615
rect 1705 -661 1775 -615
rect 1821 -661 1891 -615
rect 1937 -661 2007 -615
rect 2053 -661 2123 -615
rect 2169 -661 2239 -615
rect 2285 -661 2355 -615
rect 2401 -661 2471 -615
rect 2517 -661 2587 -615
rect 2633 -661 2703 -615
rect 2749 -661 2819 -615
rect 2865 -661 2935 -615
rect 2981 -661 3051 -615
rect 3097 -661 3167 -615
rect 3213 -661 3283 -615
rect 3329 -661 3399 -615
rect 3445 -661 3515 -615
rect 3561 -661 3631 -615
rect 3677 -661 3747 -615
rect 3793 -661 3863 -615
rect 3909 -661 3979 -615
rect 4025 -661 4095 -615
rect 4141 -661 4211 -615
rect 4257 -661 4327 -615
rect 4373 -661 4443 -615
rect 4489 -661 4559 -615
rect 4605 -661 4675 -615
rect 4721 -661 4791 -615
rect 4837 -661 4907 -615
rect 4953 -661 5023 -615
rect 5069 -661 5139 -615
rect 5185 -661 5255 -615
rect 5301 -661 5371 -615
rect 5417 -661 5487 -615
rect 5533 -661 5603 -615
rect 5649 -661 5719 -615
rect 5765 -661 5784 -615
rect -5784 -731 5784 -661
rect -5784 -777 -5765 -731
rect -5719 -777 -5649 -731
rect -5603 -777 -5533 -731
rect -5487 -777 -5417 -731
rect -5371 -777 -5301 -731
rect -5255 -777 -5185 -731
rect -5139 -777 -5069 -731
rect -5023 -777 -4953 -731
rect -4907 -777 -4837 -731
rect -4791 -777 -4721 -731
rect -4675 -777 -4605 -731
rect -4559 -777 -4489 -731
rect -4443 -777 -4373 -731
rect -4327 -777 -4257 -731
rect -4211 -777 -4141 -731
rect -4095 -777 -4025 -731
rect -3979 -777 -3909 -731
rect -3863 -777 -3793 -731
rect -3747 -777 -3677 -731
rect -3631 -777 -3561 -731
rect -3515 -777 -3445 -731
rect -3399 -777 -3329 -731
rect -3283 -777 -3213 -731
rect -3167 -777 -3097 -731
rect -3051 -777 -2981 -731
rect -2935 -777 -2865 -731
rect -2819 -777 -2749 -731
rect -2703 -777 -2633 -731
rect -2587 -777 -2517 -731
rect -2471 -777 -2401 -731
rect -2355 -777 -2285 -731
rect -2239 -777 -2169 -731
rect -2123 -777 -2053 -731
rect -2007 -777 -1937 -731
rect -1891 -777 -1821 -731
rect -1775 -777 -1705 -731
rect -1659 -777 -1589 -731
rect -1543 -777 -1473 -731
rect -1427 -777 -1357 -731
rect -1311 -777 -1241 -731
rect -1195 -777 -1125 -731
rect -1079 -777 -1009 -731
rect -963 -777 -893 -731
rect -847 -777 -777 -731
rect -731 -777 -661 -731
rect -615 -777 -545 -731
rect -499 -777 -429 -731
rect -383 -777 -313 -731
rect -267 -777 -197 -731
rect -151 -777 -81 -731
rect -35 -777 35 -731
rect 81 -777 151 -731
rect 197 -777 267 -731
rect 313 -777 383 -731
rect 429 -777 499 -731
rect 545 -777 615 -731
rect 661 -777 731 -731
rect 777 -777 847 -731
rect 893 -777 963 -731
rect 1009 -777 1079 -731
rect 1125 -777 1195 -731
rect 1241 -777 1311 -731
rect 1357 -777 1427 -731
rect 1473 -777 1543 -731
rect 1589 -777 1659 -731
rect 1705 -777 1775 -731
rect 1821 -777 1891 -731
rect 1937 -777 2007 -731
rect 2053 -777 2123 -731
rect 2169 -777 2239 -731
rect 2285 -777 2355 -731
rect 2401 -777 2471 -731
rect 2517 -777 2587 -731
rect 2633 -777 2703 -731
rect 2749 -777 2819 -731
rect 2865 -777 2935 -731
rect 2981 -777 3051 -731
rect 3097 -777 3167 -731
rect 3213 -777 3283 -731
rect 3329 -777 3399 -731
rect 3445 -777 3515 -731
rect 3561 -777 3631 -731
rect 3677 -777 3747 -731
rect 3793 -777 3863 -731
rect 3909 -777 3979 -731
rect 4025 -777 4095 -731
rect 4141 -777 4211 -731
rect 4257 -777 4327 -731
rect 4373 -777 4443 -731
rect 4489 -777 4559 -731
rect 4605 -777 4675 -731
rect 4721 -777 4791 -731
rect 4837 -777 4907 -731
rect 4953 -777 5023 -731
rect 5069 -777 5139 -731
rect 5185 -777 5255 -731
rect 5301 -777 5371 -731
rect 5417 -777 5487 -731
rect 5533 -777 5603 -731
rect 5649 -777 5719 -731
rect 5765 -777 5784 -731
rect -5784 -847 5784 -777
rect -5784 -893 -5765 -847
rect -5719 -893 -5649 -847
rect -5603 -893 -5533 -847
rect -5487 -893 -5417 -847
rect -5371 -893 -5301 -847
rect -5255 -893 -5185 -847
rect -5139 -893 -5069 -847
rect -5023 -893 -4953 -847
rect -4907 -893 -4837 -847
rect -4791 -893 -4721 -847
rect -4675 -893 -4605 -847
rect -4559 -893 -4489 -847
rect -4443 -893 -4373 -847
rect -4327 -893 -4257 -847
rect -4211 -893 -4141 -847
rect -4095 -893 -4025 -847
rect -3979 -893 -3909 -847
rect -3863 -893 -3793 -847
rect -3747 -893 -3677 -847
rect -3631 -893 -3561 -847
rect -3515 -893 -3445 -847
rect -3399 -893 -3329 -847
rect -3283 -893 -3213 -847
rect -3167 -893 -3097 -847
rect -3051 -893 -2981 -847
rect -2935 -893 -2865 -847
rect -2819 -893 -2749 -847
rect -2703 -893 -2633 -847
rect -2587 -893 -2517 -847
rect -2471 -893 -2401 -847
rect -2355 -893 -2285 -847
rect -2239 -893 -2169 -847
rect -2123 -893 -2053 -847
rect -2007 -893 -1937 -847
rect -1891 -893 -1821 -847
rect -1775 -893 -1705 -847
rect -1659 -893 -1589 -847
rect -1543 -893 -1473 -847
rect -1427 -893 -1357 -847
rect -1311 -893 -1241 -847
rect -1195 -893 -1125 -847
rect -1079 -893 -1009 -847
rect -963 -893 -893 -847
rect -847 -893 -777 -847
rect -731 -893 -661 -847
rect -615 -893 -545 -847
rect -499 -893 -429 -847
rect -383 -893 -313 -847
rect -267 -893 -197 -847
rect -151 -893 -81 -847
rect -35 -893 35 -847
rect 81 -893 151 -847
rect 197 -893 267 -847
rect 313 -893 383 -847
rect 429 -893 499 -847
rect 545 -893 615 -847
rect 661 -893 731 -847
rect 777 -893 847 -847
rect 893 -893 963 -847
rect 1009 -893 1079 -847
rect 1125 -893 1195 -847
rect 1241 -893 1311 -847
rect 1357 -893 1427 -847
rect 1473 -893 1543 -847
rect 1589 -893 1659 -847
rect 1705 -893 1775 -847
rect 1821 -893 1891 -847
rect 1937 -893 2007 -847
rect 2053 -893 2123 -847
rect 2169 -893 2239 -847
rect 2285 -893 2355 -847
rect 2401 -893 2471 -847
rect 2517 -893 2587 -847
rect 2633 -893 2703 -847
rect 2749 -893 2819 -847
rect 2865 -893 2935 -847
rect 2981 -893 3051 -847
rect 3097 -893 3167 -847
rect 3213 -893 3283 -847
rect 3329 -893 3399 -847
rect 3445 -893 3515 -847
rect 3561 -893 3631 -847
rect 3677 -893 3747 -847
rect 3793 -893 3863 -847
rect 3909 -893 3979 -847
rect 4025 -893 4095 -847
rect 4141 -893 4211 -847
rect 4257 -893 4327 -847
rect 4373 -893 4443 -847
rect 4489 -893 4559 -847
rect 4605 -893 4675 -847
rect 4721 -893 4791 -847
rect 4837 -893 4907 -847
rect 4953 -893 5023 -847
rect 5069 -893 5139 -847
rect 5185 -893 5255 -847
rect 5301 -893 5371 -847
rect 5417 -893 5487 -847
rect 5533 -893 5603 -847
rect 5649 -893 5719 -847
rect 5765 -893 5784 -847
rect -5784 -963 5784 -893
rect -5784 -1009 -5765 -963
rect -5719 -1009 -5649 -963
rect -5603 -1009 -5533 -963
rect -5487 -1009 -5417 -963
rect -5371 -1009 -5301 -963
rect -5255 -1009 -5185 -963
rect -5139 -1009 -5069 -963
rect -5023 -1009 -4953 -963
rect -4907 -1009 -4837 -963
rect -4791 -1009 -4721 -963
rect -4675 -1009 -4605 -963
rect -4559 -1009 -4489 -963
rect -4443 -1009 -4373 -963
rect -4327 -1009 -4257 -963
rect -4211 -1009 -4141 -963
rect -4095 -1009 -4025 -963
rect -3979 -1009 -3909 -963
rect -3863 -1009 -3793 -963
rect -3747 -1009 -3677 -963
rect -3631 -1009 -3561 -963
rect -3515 -1009 -3445 -963
rect -3399 -1009 -3329 -963
rect -3283 -1009 -3213 -963
rect -3167 -1009 -3097 -963
rect -3051 -1009 -2981 -963
rect -2935 -1009 -2865 -963
rect -2819 -1009 -2749 -963
rect -2703 -1009 -2633 -963
rect -2587 -1009 -2517 -963
rect -2471 -1009 -2401 -963
rect -2355 -1009 -2285 -963
rect -2239 -1009 -2169 -963
rect -2123 -1009 -2053 -963
rect -2007 -1009 -1937 -963
rect -1891 -1009 -1821 -963
rect -1775 -1009 -1705 -963
rect -1659 -1009 -1589 -963
rect -1543 -1009 -1473 -963
rect -1427 -1009 -1357 -963
rect -1311 -1009 -1241 -963
rect -1195 -1009 -1125 -963
rect -1079 -1009 -1009 -963
rect -963 -1009 -893 -963
rect -847 -1009 -777 -963
rect -731 -1009 -661 -963
rect -615 -1009 -545 -963
rect -499 -1009 -429 -963
rect -383 -1009 -313 -963
rect -267 -1009 -197 -963
rect -151 -1009 -81 -963
rect -35 -1009 35 -963
rect 81 -1009 151 -963
rect 197 -1009 267 -963
rect 313 -1009 383 -963
rect 429 -1009 499 -963
rect 545 -1009 615 -963
rect 661 -1009 731 -963
rect 777 -1009 847 -963
rect 893 -1009 963 -963
rect 1009 -1009 1079 -963
rect 1125 -1009 1195 -963
rect 1241 -1009 1311 -963
rect 1357 -1009 1427 -963
rect 1473 -1009 1543 -963
rect 1589 -1009 1659 -963
rect 1705 -1009 1775 -963
rect 1821 -1009 1891 -963
rect 1937 -1009 2007 -963
rect 2053 -1009 2123 -963
rect 2169 -1009 2239 -963
rect 2285 -1009 2355 -963
rect 2401 -1009 2471 -963
rect 2517 -1009 2587 -963
rect 2633 -1009 2703 -963
rect 2749 -1009 2819 -963
rect 2865 -1009 2935 -963
rect 2981 -1009 3051 -963
rect 3097 -1009 3167 -963
rect 3213 -1009 3283 -963
rect 3329 -1009 3399 -963
rect 3445 -1009 3515 -963
rect 3561 -1009 3631 -963
rect 3677 -1009 3747 -963
rect 3793 -1009 3863 -963
rect 3909 -1009 3979 -963
rect 4025 -1009 4095 -963
rect 4141 -1009 4211 -963
rect 4257 -1009 4327 -963
rect 4373 -1009 4443 -963
rect 4489 -1009 4559 -963
rect 4605 -1009 4675 -963
rect 4721 -1009 4791 -963
rect 4837 -1009 4907 -963
rect 4953 -1009 5023 -963
rect 5069 -1009 5139 -963
rect 5185 -1009 5255 -963
rect 5301 -1009 5371 -963
rect 5417 -1009 5487 -963
rect 5533 -1009 5603 -963
rect 5649 -1009 5719 -963
rect 5765 -1009 5784 -963
rect -5784 -1079 5784 -1009
rect -5784 -1125 -5765 -1079
rect -5719 -1125 -5649 -1079
rect -5603 -1125 -5533 -1079
rect -5487 -1125 -5417 -1079
rect -5371 -1125 -5301 -1079
rect -5255 -1125 -5185 -1079
rect -5139 -1125 -5069 -1079
rect -5023 -1125 -4953 -1079
rect -4907 -1125 -4837 -1079
rect -4791 -1125 -4721 -1079
rect -4675 -1125 -4605 -1079
rect -4559 -1125 -4489 -1079
rect -4443 -1125 -4373 -1079
rect -4327 -1125 -4257 -1079
rect -4211 -1125 -4141 -1079
rect -4095 -1125 -4025 -1079
rect -3979 -1125 -3909 -1079
rect -3863 -1125 -3793 -1079
rect -3747 -1125 -3677 -1079
rect -3631 -1125 -3561 -1079
rect -3515 -1125 -3445 -1079
rect -3399 -1125 -3329 -1079
rect -3283 -1125 -3213 -1079
rect -3167 -1125 -3097 -1079
rect -3051 -1125 -2981 -1079
rect -2935 -1125 -2865 -1079
rect -2819 -1125 -2749 -1079
rect -2703 -1125 -2633 -1079
rect -2587 -1125 -2517 -1079
rect -2471 -1125 -2401 -1079
rect -2355 -1125 -2285 -1079
rect -2239 -1125 -2169 -1079
rect -2123 -1125 -2053 -1079
rect -2007 -1125 -1937 -1079
rect -1891 -1125 -1821 -1079
rect -1775 -1125 -1705 -1079
rect -1659 -1125 -1589 -1079
rect -1543 -1125 -1473 -1079
rect -1427 -1125 -1357 -1079
rect -1311 -1125 -1241 -1079
rect -1195 -1125 -1125 -1079
rect -1079 -1125 -1009 -1079
rect -963 -1125 -893 -1079
rect -847 -1125 -777 -1079
rect -731 -1125 -661 -1079
rect -615 -1125 -545 -1079
rect -499 -1125 -429 -1079
rect -383 -1125 -313 -1079
rect -267 -1125 -197 -1079
rect -151 -1125 -81 -1079
rect -35 -1125 35 -1079
rect 81 -1125 151 -1079
rect 197 -1125 267 -1079
rect 313 -1125 383 -1079
rect 429 -1125 499 -1079
rect 545 -1125 615 -1079
rect 661 -1125 731 -1079
rect 777 -1125 847 -1079
rect 893 -1125 963 -1079
rect 1009 -1125 1079 -1079
rect 1125 -1125 1195 -1079
rect 1241 -1125 1311 -1079
rect 1357 -1125 1427 -1079
rect 1473 -1125 1543 -1079
rect 1589 -1125 1659 -1079
rect 1705 -1125 1775 -1079
rect 1821 -1125 1891 -1079
rect 1937 -1125 2007 -1079
rect 2053 -1125 2123 -1079
rect 2169 -1125 2239 -1079
rect 2285 -1125 2355 -1079
rect 2401 -1125 2471 -1079
rect 2517 -1125 2587 -1079
rect 2633 -1125 2703 -1079
rect 2749 -1125 2819 -1079
rect 2865 -1125 2935 -1079
rect 2981 -1125 3051 -1079
rect 3097 -1125 3167 -1079
rect 3213 -1125 3283 -1079
rect 3329 -1125 3399 -1079
rect 3445 -1125 3515 -1079
rect 3561 -1125 3631 -1079
rect 3677 -1125 3747 -1079
rect 3793 -1125 3863 -1079
rect 3909 -1125 3979 -1079
rect 4025 -1125 4095 -1079
rect 4141 -1125 4211 -1079
rect 4257 -1125 4327 -1079
rect 4373 -1125 4443 -1079
rect 4489 -1125 4559 -1079
rect 4605 -1125 4675 -1079
rect 4721 -1125 4791 -1079
rect 4837 -1125 4907 -1079
rect 4953 -1125 5023 -1079
rect 5069 -1125 5139 -1079
rect 5185 -1125 5255 -1079
rect 5301 -1125 5371 -1079
rect 5417 -1125 5487 -1079
rect 5533 -1125 5603 -1079
rect 5649 -1125 5719 -1079
rect 5765 -1125 5784 -1079
rect -5784 -1144 5784 -1125
<< psubdiffcont >>
rect -5765 1079 -5719 1125
rect -5649 1079 -5603 1125
rect -5533 1079 -5487 1125
rect -5417 1079 -5371 1125
rect -5301 1079 -5255 1125
rect -5185 1079 -5139 1125
rect -5069 1079 -5023 1125
rect -4953 1079 -4907 1125
rect -4837 1079 -4791 1125
rect -4721 1079 -4675 1125
rect -4605 1079 -4559 1125
rect -4489 1079 -4443 1125
rect -4373 1079 -4327 1125
rect -4257 1079 -4211 1125
rect -4141 1079 -4095 1125
rect -4025 1079 -3979 1125
rect -3909 1079 -3863 1125
rect -3793 1079 -3747 1125
rect -3677 1079 -3631 1125
rect -3561 1079 -3515 1125
rect -3445 1079 -3399 1125
rect -3329 1079 -3283 1125
rect -3213 1079 -3167 1125
rect -3097 1079 -3051 1125
rect -2981 1079 -2935 1125
rect -2865 1079 -2819 1125
rect -2749 1079 -2703 1125
rect -2633 1079 -2587 1125
rect -2517 1079 -2471 1125
rect -2401 1079 -2355 1125
rect -2285 1079 -2239 1125
rect -2169 1079 -2123 1125
rect -2053 1079 -2007 1125
rect -1937 1079 -1891 1125
rect -1821 1079 -1775 1125
rect -1705 1079 -1659 1125
rect -1589 1079 -1543 1125
rect -1473 1079 -1427 1125
rect -1357 1079 -1311 1125
rect -1241 1079 -1195 1125
rect -1125 1079 -1079 1125
rect -1009 1079 -963 1125
rect -893 1079 -847 1125
rect -777 1079 -731 1125
rect -661 1079 -615 1125
rect -545 1079 -499 1125
rect -429 1079 -383 1125
rect -313 1079 -267 1125
rect -197 1079 -151 1125
rect -81 1079 -35 1125
rect 35 1079 81 1125
rect 151 1079 197 1125
rect 267 1079 313 1125
rect 383 1079 429 1125
rect 499 1079 545 1125
rect 615 1079 661 1125
rect 731 1079 777 1125
rect 847 1079 893 1125
rect 963 1079 1009 1125
rect 1079 1079 1125 1125
rect 1195 1079 1241 1125
rect 1311 1079 1357 1125
rect 1427 1079 1473 1125
rect 1543 1079 1589 1125
rect 1659 1079 1705 1125
rect 1775 1079 1821 1125
rect 1891 1079 1937 1125
rect 2007 1079 2053 1125
rect 2123 1079 2169 1125
rect 2239 1079 2285 1125
rect 2355 1079 2401 1125
rect 2471 1079 2517 1125
rect 2587 1079 2633 1125
rect 2703 1079 2749 1125
rect 2819 1079 2865 1125
rect 2935 1079 2981 1125
rect 3051 1079 3097 1125
rect 3167 1079 3213 1125
rect 3283 1079 3329 1125
rect 3399 1079 3445 1125
rect 3515 1079 3561 1125
rect 3631 1079 3677 1125
rect 3747 1079 3793 1125
rect 3863 1079 3909 1125
rect 3979 1079 4025 1125
rect 4095 1079 4141 1125
rect 4211 1079 4257 1125
rect 4327 1079 4373 1125
rect 4443 1079 4489 1125
rect 4559 1079 4605 1125
rect 4675 1079 4721 1125
rect 4791 1079 4837 1125
rect 4907 1079 4953 1125
rect 5023 1079 5069 1125
rect 5139 1079 5185 1125
rect 5255 1079 5301 1125
rect 5371 1079 5417 1125
rect 5487 1079 5533 1125
rect 5603 1079 5649 1125
rect 5719 1079 5765 1125
rect -5765 963 -5719 1009
rect -5649 963 -5603 1009
rect -5533 963 -5487 1009
rect -5417 963 -5371 1009
rect -5301 963 -5255 1009
rect -5185 963 -5139 1009
rect -5069 963 -5023 1009
rect -4953 963 -4907 1009
rect -4837 963 -4791 1009
rect -4721 963 -4675 1009
rect -4605 963 -4559 1009
rect -4489 963 -4443 1009
rect -4373 963 -4327 1009
rect -4257 963 -4211 1009
rect -4141 963 -4095 1009
rect -4025 963 -3979 1009
rect -3909 963 -3863 1009
rect -3793 963 -3747 1009
rect -3677 963 -3631 1009
rect -3561 963 -3515 1009
rect -3445 963 -3399 1009
rect -3329 963 -3283 1009
rect -3213 963 -3167 1009
rect -3097 963 -3051 1009
rect -2981 963 -2935 1009
rect -2865 963 -2819 1009
rect -2749 963 -2703 1009
rect -2633 963 -2587 1009
rect -2517 963 -2471 1009
rect -2401 963 -2355 1009
rect -2285 963 -2239 1009
rect -2169 963 -2123 1009
rect -2053 963 -2007 1009
rect -1937 963 -1891 1009
rect -1821 963 -1775 1009
rect -1705 963 -1659 1009
rect -1589 963 -1543 1009
rect -1473 963 -1427 1009
rect -1357 963 -1311 1009
rect -1241 963 -1195 1009
rect -1125 963 -1079 1009
rect -1009 963 -963 1009
rect -893 963 -847 1009
rect -777 963 -731 1009
rect -661 963 -615 1009
rect -545 963 -499 1009
rect -429 963 -383 1009
rect -313 963 -267 1009
rect -197 963 -151 1009
rect -81 963 -35 1009
rect 35 963 81 1009
rect 151 963 197 1009
rect 267 963 313 1009
rect 383 963 429 1009
rect 499 963 545 1009
rect 615 963 661 1009
rect 731 963 777 1009
rect 847 963 893 1009
rect 963 963 1009 1009
rect 1079 963 1125 1009
rect 1195 963 1241 1009
rect 1311 963 1357 1009
rect 1427 963 1473 1009
rect 1543 963 1589 1009
rect 1659 963 1705 1009
rect 1775 963 1821 1009
rect 1891 963 1937 1009
rect 2007 963 2053 1009
rect 2123 963 2169 1009
rect 2239 963 2285 1009
rect 2355 963 2401 1009
rect 2471 963 2517 1009
rect 2587 963 2633 1009
rect 2703 963 2749 1009
rect 2819 963 2865 1009
rect 2935 963 2981 1009
rect 3051 963 3097 1009
rect 3167 963 3213 1009
rect 3283 963 3329 1009
rect 3399 963 3445 1009
rect 3515 963 3561 1009
rect 3631 963 3677 1009
rect 3747 963 3793 1009
rect 3863 963 3909 1009
rect 3979 963 4025 1009
rect 4095 963 4141 1009
rect 4211 963 4257 1009
rect 4327 963 4373 1009
rect 4443 963 4489 1009
rect 4559 963 4605 1009
rect 4675 963 4721 1009
rect 4791 963 4837 1009
rect 4907 963 4953 1009
rect 5023 963 5069 1009
rect 5139 963 5185 1009
rect 5255 963 5301 1009
rect 5371 963 5417 1009
rect 5487 963 5533 1009
rect 5603 963 5649 1009
rect 5719 963 5765 1009
rect -5765 847 -5719 893
rect -5649 847 -5603 893
rect -5533 847 -5487 893
rect -5417 847 -5371 893
rect -5301 847 -5255 893
rect -5185 847 -5139 893
rect -5069 847 -5023 893
rect -4953 847 -4907 893
rect -4837 847 -4791 893
rect -4721 847 -4675 893
rect -4605 847 -4559 893
rect -4489 847 -4443 893
rect -4373 847 -4327 893
rect -4257 847 -4211 893
rect -4141 847 -4095 893
rect -4025 847 -3979 893
rect -3909 847 -3863 893
rect -3793 847 -3747 893
rect -3677 847 -3631 893
rect -3561 847 -3515 893
rect -3445 847 -3399 893
rect -3329 847 -3283 893
rect -3213 847 -3167 893
rect -3097 847 -3051 893
rect -2981 847 -2935 893
rect -2865 847 -2819 893
rect -2749 847 -2703 893
rect -2633 847 -2587 893
rect -2517 847 -2471 893
rect -2401 847 -2355 893
rect -2285 847 -2239 893
rect -2169 847 -2123 893
rect -2053 847 -2007 893
rect -1937 847 -1891 893
rect -1821 847 -1775 893
rect -1705 847 -1659 893
rect -1589 847 -1543 893
rect -1473 847 -1427 893
rect -1357 847 -1311 893
rect -1241 847 -1195 893
rect -1125 847 -1079 893
rect -1009 847 -963 893
rect -893 847 -847 893
rect -777 847 -731 893
rect -661 847 -615 893
rect -545 847 -499 893
rect -429 847 -383 893
rect -313 847 -267 893
rect -197 847 -151 893
rect -81 847 -35 893
rect 35 847 81 893
rect 151 847 197 893
rect 267 847 313 893
rect 383 847 429 893
rect 499 847 545 893
rect 615 847 661 893
rect 731 847 777 893
rect 847 847 893 893
rect 963 847 1009 893
rect 1079 847 1125 893
rect 1195 847 1241 893
rect 1311 847 1357 893
rect 1427 847 1473 893
rect 1543 847 1589 893
rect 1659 847 1705 893
rect 1775 847 1821 893
rect 1891 847 1937 893
rect 2007 847 2053 893
rect 2123 847 2169 893
rect 2239 847 2285 893
rect 2355 847 2401 893
rect 2471 847 2517 893
rect 2587 847 2633 893
rect 2703 847 2749 893
rect 2819 847 2865 893
rect 2935 847 2981 893
rect 3051 847 3097 893
rect 3167 847 3213 893
rect 3283 847 3329 893
rect 3399 847 3445 893
rect 3515 847 3561 893
rect 3631 847 3677 893
rect 3747 847 3793 893
rect 3863 847 3909 893
rect 3979 847 4025 893
rect 4095 847 4141 893
rect 4211 847 4257 893
rect 4327 847 4373 893
rect 4443 847 4489 893
rect 4559 847 4605 893
rect 4675 847 4721 893
rect 4791 847 4837 893
rect 4907 847 4953 893
rect 5023 847 5069 893
rect 5139 847 5185 893
rect 5255 847 5301 893
rect 5371 847 5417 893
rect 5487 847 5533 893
rect 5603 847 5649 893
rect 5719 847 5765 893
rect -5765 731 -5719 777
rect -5649 731 -5603 777
rect -5533 731 -5487 777
rect -5417 731 -5371 777
rect -5301 731 -5255 777
rect -5185 731 -5139 777
rect -5069 731 -5023 777
rect -4953 731 -4907 777
rect -4837 731 -4791 777
rect -4721 731 -4675 777
rect -4605 731 -4559 777
rect -4489 731 -4443 777
rect -4373 731 -4327 777
rect -4257 731 -4211 777
rect -4141 731 -4095 777
rect -4025 731 -3979 777
rect -3909 731 -3863 777
rect -3793 731 -3747 777
rect -3677 731 -3631 777
rect -3561 731 -3515 777
rect -3445 731 -3399 777
rect -3329 731 -3283 777
rect -3213 731 -3167 777
rect -3097 731 -3051 777
rect -2981 731 -2935 777
rect -2865 731 -2819 777
rect -2749 731 -2703 777
rect -2633 731 -2587 777
rect -2517 731 -2471 777
rect -2401 731 -2355 777
rect -2285 731 -2239 777
rect -2169 731 -2123 777
rect -2053 731 -2007 777
rect -1937 731 -1891 777
rect -1821 731 -1775 777
rect -1705 731 -1659 777
rect -1589 731 -1543 777
rect -1473 731 -1427 777
rect -1357 731 -1311 777
rect -1241 731 -1195 777
rect -1125 731 -1079 777
rect -1009 731 -963 777
rect -893 731 -847 777
rect -777 731 -731 777
rect -661 731 -615 777
rect -545 731 -499 777
rect -429 731 -383 777
rect -313 731 -267 777
rect -197 731 -151 777
rect -81 731 -35 777
rect 35 731 81 777
rect 151 731 197 777
rect 267 731 313 777
rect 383 731 429 777
rect 499 731 545 777
rect 615 731 661 777
rect 731 731 777 777
rect 847 731 893 777
rect 963 731 1009 777
rect 1079 731 1125 777
rect 1195 731 1241 777
rect 1311 731 1357 777
rect 1427 731 1473 777
rect 1543 731 1589 777
rect 1659 731 1705 777
rect 1775 731 1821 777
rect 1891 731 1937 777
rect 2007 731 2053 777
rect 2123 731 2169 777
rect 2239 731 2285 777
rect 2355 731 2401 777
rect 2471 731 2517 777
rect 2587 731 2633 777
rect 2703 731 2749 777
rect 2819 731 2865 777
rect 2935 731 2981 777
rect 3051 731 3097 777
rect 3167 731 3213 777
rect 3283 731 3329 777
rect 3399 731 3445 777
rect 3515 731 3561 777
rect 3631 731 3677 777
rect 3747 731 3793 777
rect 3863 731 3909 777
rect 3979 731 4025 777
rect 4095 731 4141 777
rect 4211 731 4257 777
rect 4327 731 4373 777
rect 4443 731 4489 777
rect 4559 731 4605 777
rect 4675 731 4721 777
rect 4791 731 4837 777
rect 4907 731 4953 777
rect 5023 731 5069 777
rect 5139 731 5185 777
rect 5255 731 5301 777
rect 5371 731 5417 777
rect 5487 731 5533 777
rect 5603 731 5649 777
rect 5719 731 5765 777
rect -5765 615 -5719 661
rect -5649 615 -5603 661
rect -5533 615 -5487 661
rect -5417 615 -5371 661
rect -5301 615 -5255 661
rect -5185 615 -5139 661
rect -5069 615 -5023 661
rect -4953 615 -4907 661
rect -4837 615 -4791 661
rect -4721 615 -4675 661
rect -4605 615 -4559 661
rect -4489 615 -4443 661
rect -4373 615 -4327 661
rect -4257 615 -4211 661
rect -4141 615 -4095 661
rect -4025 615 -3979 661
rect -3909 615 -3863 661
rect -3793 615 -3747 661
rect -3677 615 -3631 661
rect -3561 615 -3515 661
rect -3445 615 -3399 661
rect -3329 615 -3283 661
rect -3213 615 -3167 661
rect -3097 615 -3051 661
rect -2981 615 -2935 661
rect -2865 615 -2819 661
rect -2749 615 -2703 661
rect -2633 615 -2587 661
rect -2517 615 -2471 661
rect -2401 615 -2355 661
rect -2285 615 -2239 661
rect -2169 615 -2123 661
rect -2053 615 -2007 661
rect -1937 615 -1891 661
rect -1821 615 -1775 661
rect -1705 615 -1659 661
rect -1589 615 -1543 661
rect -1473 615 -1427 661
rect -1357 615 -1311 661
rect -1241 615 -1195 661
rect -1125 615 -1079 661
rect -1009 615 -963 661
rect -893 615 -847 661
rect -777 615 -731 661
rect -661 615 -615 661
rect -545 615 -499 661
rect -429 615 -383 661
rect -313 615 -267 661
rect -197 615 -151 661
rect -81 615 -35 661
rect 35 615 81 661
rect 151 615 197 661
rect 267 615 313 661
rect 383 615 429 661
rect 499 615 545 661
rect 615 615 661 661
rect 731 615 777 661
rect 847 615 893 661
rect 963 615 1009 661
rect 1079 615 1125 661
rect 1195 615 1241 661
rect 1311 615 1357 661
rect 1427 615 1473 661
rect 1543 615 1589 661
rect 1659 615 1705 661
rect 1775 615 1821 661
rect 1891 615 1937 661
rect 2007 615 2053 661
rect 2123 615 2169 661
rect 2239 615 2285 661
rect 2355 615 2401 661
rect 2471 615 2517 661
rect 2587 615 2633 661
rect 2703 615 2749 661
rect 2819 615 2865 661
rect 2935 615 2981 661
rect 3051 615 3097 661
rect 3167 615 3213 661
rect 3283 615 3329 661
rect 3399 615 3445 661
rect 3515 615 3561 661
rect 3631 615 3677 661
rect 3747 615 3793 661
rect 3863 615 3909 661
rect 3979 615 4025 661
rect 4095 615 4141 661
rect 4211 615 4257 661
rect 4327 615 4373 661
rect 4443 615 4489 661
rect 4559 615 4605 661
rect 4675 615 4721 661
rect 4791 615 4837 661
rect 4907 615 4953 661
rect 5023 615 5069 661
rect 5139 615 5185 661
rect 5255 615 5301 661
rect 5371 615 5417 661
rect 5487 615 5533 661
rect 5603 615 5649 661
rect 5719 615 5765 661
rect -5765 499 -5719 545
rect -5649 499 -5603 545
rect -5533 499 -5487 545
rect -5417 499 -5371 545
rect -5301 499 -5255 545
rect -5185 499 -5139 545
rect -5069 499 -5023 545
rect -4953 499 -4907 545
rect -4837 499 -4791 545
rect -4721 499 -4675 545
rect -4605 499 -4559 545
rect -4489 499 -4443 545
rect -4373 499 -4327 545
rect -4257 499 -4211 545
rect -4141 499 -4095 545
rect -4025 499 -3979 545
rect -3909 499 -3863 545
rect -3793 499 -3747 545
rect -3677 499 -3631 545
rect -3561 499 -3515 545
rect -3445 499 -3399 545
rect -3329 499 -3283 545
rect -3213 499 -3167 545
rect -3097 499 -3051 545
rect -2981 499 -2935 545
rect -2865 499 -2819 545
rect -2749 499 -2703 545
rect -2633 499 -2587 545
rect -2517 499 -2471 545
rect -2401 499 -2355 545
rect -2285 499 -2239 545
rect -2169 499 -2123 545
rect -2053 499 -2007 545
rect -1937 499 -1891 545
rect -1821 499 -1775 545
rect -1705 499 -1659 545
rect -1589 499 -1543 545
rect -1473 499 -1427 545
rect -1357 499 -1311 545
rect -1241 499 -1195 545
rect -1125 499 -1079 545
rect -1009 499 -963 545
rect -893 499 -847 545
rect -777 499 -731 545
rect -661 499 -615 545
rect -545 499 -499 545
rect -429 499 -383 545
rect -313 499 -267 545
rect -197 499 -151 545
rect -81 499 -35 545
rect 35 499 81 545
rect 151 499 197 545
rect 267 499 313 545
rect 383 499 429 545
rect 499 499 545 545
rect 615 499 661 545
rect 731 499 777 545
rect 847 499 893 545
rect 963 499 1009 545
rect 1079 499 1125 545
rect 1195 499 1241 545
rect 1311 499 1357 545
rect 1427 499 1473 545
rect 1543 499 1589 545
rect 1659 499 1705 545
rect 1775 499 1821 545
rect 1891 499 1937 545
rect 2007 499 2053 545
rect 2123 499 2169 545
rect 2239 499 2285 545
rect 2355 499 2401 545
rect 2471 499 2517 545
rect 2587 499 2633 545
rect 2703 499 2749 545
rect 2819 499 2865 545
rect 2935 499 2981 545
rect 3051 499 3097 545
rect 3167 499 3213 545
rect 3283 499 3329 545
rect 3399 499 3445 545
rect 3515 499 3561 545
rect 3631 499 3677 545
rect 3747 499 3793 545
rect 3863 499 3909 545
rect 3979 499 4025 545
rect 4095 499 4141 545
rect 4211 499 4257 545
rect 4327 499 4373 545
rect 4443 499 4489 545
rect 4559 499 4605 545
rect 4675 499 4721 545
rect 4791 499 4837 545
rect 4907 499 4953 545
rect 5023 499 5069 545
rect 5139 499 5185 545
rect 5255 499 5301 545
rect 5371 499 5417 545
rect 5487 499 5533 545
rect 5603 499 5649 545
rect 5719 499 5765 545
rect -5765 383 -5719 429
rect -5649 383 -5603 429
rect -5533 383 -5487 429
rect -5417 383 -5371 429
rect -5301 383 -5255 429
rect -5185 383 -5139 429
rect -5069 383 -5023 429
rect -4953 383 -4907 429
rect -4837 383 -4791 429
rect -4721 383 -4675 429
rect -4605 383 -4559 429
rect -4489 383 -4443 429
rect -4373 383 -4327 429
rect -4257 383 -4211 429
rect -4141 383 -4095 429
rect -4025 383 -3979 429
rect -3909 383 -3863 429
rect -3793 383 -3747 429
rect -3677 383 -3631 429
rect -3561 383 -3515 429
rect -3445 383 -3399 429
rect -3329 383 -3283 429
rect -3213 383 -3167 429
rect -3097 383 -3051 429
rect -2981 383 -2935 429
rect -2865 383 -2819 429
rect -2749 383 -2703 429
rect -2633 383 -2587 429
rect -2517 383 -2471 429
rect -2401 383 -2355 429
rect -2285 383 -2239 429
rect -2169 383 -2123 429
rect -2053 383 -2007 429
rect -1937 383 -1891 429
rect -1821 383 -1775 429
rect -1705 383 -1659 429
rect -1589 383 -1543 429
rect -1473 383 -1427 429
rect -1357 383 -1311 429
rect -1241 383 -1195 429
rect -1125 383 -1079 429
rect -1009 383 -963 429
rect -893 383 -847 429
rect -777 383 -731 429
rect -661 383 -615 429
rect -545 383 -499 429
rect -429 383 -383 429
rect -313 383 -267 429
rect -197 383 -151 429
rect -81 383 -35 429
rect 35 383 81 429
rect 151 383 197 429
rect 267 383 313 429
rect 383 383 429 429
rect 499 383 545 429
rect 615 383 661 429
rect 731 383 777 429
rect 847 383 893 429
rect 963 383 1009 429
rect 1079 383 1125 429
rect 1195 383 1241 429
rect 1311 383 1357 429
rect 1427 383 1473 429
rect 1543 383 1589 429
rect 1659 383 1705 429
rect 1775 383 1821 429
rect 1891 383 1937 429
rect 2007 383 2053 429
rect 2123 383 2169 429
rect 2239 383 2285 429
rect 2355 383 2401 429
rect 2471 383 2517 429
rect 2587 383 2633 429
rect 2703 383 2749 429
rect 2819 383 2865 429
rect 2935 383 2981 429
rect 3051 383 3097 429
rect 3167 383 3213 429
rect 3283 383 3329 429
rect 3399 383 3445 429
rect 3515 383 3561 429
rect 3631 383 3677 429
rect 3747 383 3793 429
rect 3863 383 3909 429
rect 3979 383 4025 429
rect 4095 383 4141 429
rect 4211 383 4257 429
rect 4327 383 4373 429
rect 4443 383 4489 429
rect 4559 383 4605 429
rect 4675 383 4721 429
rect 4791 383 4837 429
rect 4907 383 4953 429
rect 5023 383 5069 429
rect 5139 383 5185 429
rect 5255 383 5301 429
rect 5371 383 5417 429
rect 5487 383 5533 429
rect 5603 383 5649 429
rect 5719 383 5765 429
rect -5765 267 -5719 313
rect -5649 267 -5603 313
rect -5533 267 -5487 313
rect -5417 267 -5371 313
rect -5301 267 -5255 313
rect -5185 267 -5139 313
rect -5069 267 -5023 313
rect -4953 267 -4907 313
rect -4837 267 -4791 313
rect -4721 267 -4675 313
rect -4605 267 -4559 313
rect -4489 267 -4443 313
rect -4373 267 -4327 313
rect -4257 267 -4211 313
rect -4141 267 -4095 313
rect -4025 267 -3979 313
rect -3909 267 -3863 313
rect -3793 267 -3747 313
rect -3677 267 -3631 313
rect -3561 267 -3515 313
rect -3445 267 -3399 313
rect -3329 267 -3283 313
rect -3213 267 -3167 313
rect -3097 267 -3051 313
rect -2981 267 -2935 313
rect -2865 267 -2819 313
rect -2749 267 -2703 313
rect -2633 267 -2587 313
rect -2517 267 -2471 313
rect -2401 267 -2355 313
rect -2285 267 -2239 313
rect -2169 267 -2123 313
rect -2053 267 -2007 313
rect -1937 267 -1891 313
rect -1821 267 -1775 313
rect -1705 267 -1659 313
rect -1589 267 -1543 313
rect -1473 267 -1427 313
rect -1357 267 -1311 313
rect -1241 267 -1195 313
rect -1125 267 -1079 313
rect -1009 267 -963 313
rect -893 267 -847 313
rect -777 267 -731 313
rect -661 267 -615 313
rect -545 267 -499 313
rect -429 267 -383 313
rect -313 267 -267 313
rect -197 267 -151 313
rect -81 267 -35 313
rect 35 267 81 313
rect 151 267 197 313
rect 267 267 313 313
rect 383 267 429 313
rect 499 267 545 313
rect 615 267 661 313
rect 731 267 777 313
rect 847 267 893 313
rect 963 267 1009 313
rect 1079 267 1125 313
rect 1195 267 1241 313
rect 1311 267 1357 313
rect 1427 267 1473 313
rect 1543 267 1589 313
rect 1659 267 1705 313
rect 1775 267 1821 313
rect 1891 267 1937 313
rect 2007 267 2053 313
rect 2123 267 2169 313
rect 2239 267 2285 313
rect 2355 267 2401 313
rect 2471 267 2517 313
rect 2587 267 2633 313
rect 2703 267 2749 313
rect 2819 267 2865 313
rect 2935 267 2981 313
rect 3051 267 3097 313
rect 3167 267 3213 313
rect 3283 267 3329 313
rect 3399 267 3445 313
rect 3515 267 3561 313
rect 3631 267 3677 313
rect 3747 267 3793 313
rect 3863 267 3909 313
rect 3979 267 4025 313
rect 4095 267 4141 313
rect 4211 267 4257 313
rect 4327 267 4373 313
rect 4443 267 4489 313
rect 4559 267 4605 313
rect 4675 267 4721 313
rect 4791 267 4837 313
rect 4907 267 4953 313
rect 5023 267 5069 313
rect 5139 267 5185 313
rect 5255 267 5301 313
rect 5371 267 5417 313
rect 5487 267 5533 313
rect 5603 267 5649 313
rect 5719 267 5765 313
rect -5765 151 -5719 197
rect -5649 151 -5603 197
rect -5533 151 -5487 197
rect -5417 151 -5371 197
rect -5301 151 -5255 197
rect -5185 151 -5139 197
rect -5069 151 -5023 197
rect -4953 151 -4907 197
rect -4837 151 -4791 197
rect -4721 151 -4675 197
rect -4605 151 -4559 197
rect -4489 151 -4443 197
rect -4373 151 -4327 197
rect -4257 151 -4211 197
rect -4141 151 -4095 197
rect -4025 151 -3979 197
rect -3909 151 -3863 197
rect -3793 151 -3747 197
rect -3677 151 -3631 197
rect -3561 151 -3515 197
rect -3445 151 -3399 197
rect -3329 151 -3283 197
rect -3213 151 -3167 197
rect -3097 151 -3051 197
rect -2981 151 -2935 197
rect -2865 151 -2819 197
rect -2749 151 -2703 197
rect -2633 151 -2587 197
rect -2517 151 -2471 197
rect -2401 151 -2355 197
rect -2285 151 -2239 197
rect -2169 151 -2123 197
rect -2053 151 -2007 197
rect -1937 151 -1891 197
rect -1821 151 -1775 197
rect -1705 151 -1659 197
rect -1589 151 -1543 197
rect -1473 151 -1427 197
rect -1357 151 -1311 197
rect -1241 151 -1195 197
rect -1125 151 -1079 197
rect -1009 151 -963 197
rect -893 151 -847 197
rect -777 151 -731 197
rect -661 151 -615 197
rect -545 151 -499 197
rect -429 151 -383 197
rect -313 151 -267 197
rect -197 151 -151 197
rect -81 151 -35 197
rect 35 151 81 197
rect 151 151 197 197
rect 267 151 313 197
rect 383 151 429 197
rect 499 151 545 197
rect 615 151 661 197
rect 731 151 777 197
rect 847 151 893 197
rect 963 151 1009 197
rect 1079 151 1125 197
rect 1195 151 1241 197
rect 1311 151 1357 197
rect 1427 151 1473 197
rect 1543 151 1589 197
rect 1659 151 1705 197
rect 1775 151 1821 197
rect 1891 151 1937 197
rect 2007 151 2053 197
rect 2123 151 2169 197
rect 2239 151 2285 197
rect 2355 151 2401 197
rect 2471 151 2517 197
rect 2587 151 2633 197
rect 2703 151 2749 197
rect 2819 151 2865 197
rect 2935 151 2981 197
rect 3051 151 3097 197
rect 3167 151 3213 197
rect 3283 151 3329 197
rect 3399 151 3445 197
rect 3515 151 3561 197
rect 3631 151 3677 197
rect 3747 151 3793 197
rect 3863 151 3909 197
rect 3979 151 4025 197
rect 4095 151 4141 197
rect 4211 151 4257 197
rect 4327 151 4373 197
rect 4443 151 4489 197
rect 4559 151 4605 197
rect 4675 151 4721 197
rect 4791 151 4837 197
rect 4907 151 4953 197
rect 5023 151 5069 197
rect 5139 151 5185 197
rect 5255 151 5301 197
rect 5371 151 5417 197
rect 5487 151 5533 197
rect 5603 151 5649 197
rect 5719 151 5765 197
rect -5765 35 -5719 81
rect -5649 35 -5603 81
rect -5533 35 -5487 81
rect -5417 35 -5371 81
rect -5301 35 -5255 81
rect -5185 35 -5139 81
rect -5069 35 -5023 81
rect -4953 35 -4907 81
rect -4837 35 -4791 81
rect -4721 35 -4675 81
rect -4605 35 -4559 81
rect -4489 35 -4443 81
rect -4373 35 -4327 81
rect -4257 35 -4211 81
rect -4141 35 -4095 81
rect -4025 35 -3979 81
rect -3909 35 -3863 81
rect -3793 35 -3747 81
rect -3677 35 -3631 81
rect -3561 35 -3515 81
rect -3445 35 -3399 81
rect -3329 35 -3283 81
rect -3213 35 -3167 81
rect -3097 35 -3051 81
rect -2981 35 -2935 81
rect -2865 35 -2819 81
rect -2749 35 -2703 81
rect -2633 35 -2587 81
rect -2517 35 -2471 81
rect -2401 35 -2355 81
rect -2285 35 -2239 81
rect -2169 35 -2123 81
rect -2053 35 -2007 81
rect -1937 35 -1891 81
rect -1821 35 -1775 81
rect -1705 35 -1659 81
rect -1589 35 -1543 81
rect -1473 35 -1427 81
rect -1357 35 -1311 81
rect -1241 35 -1195 81
rect -1125 35 -1079 81
rect -1009 35 -963 81
rect -893 35 -847 81
rect -777 35 -731 81
rect -661 35 -615 81
rect -545 35 -499 81
rect -429 35 -383 81
rect -313 35 -267 81
rect -197 35 -151 81
rect -81 35 -35 81
rect 35 35 81 81
rect 151 35 197 81
rect 267 35 313 81
rect 383 35 429 81
rect 499 35 545 81
rect 615 35 661 81
rect 731 35 777 81
rect 847 35 893 81
rect 963 35 1009 81
rect 1079 35 1125 81
rect 1195 35 1241 81
rect 1311 35 1357 81
rect 1427 35 1473 81
rect 1543 35 1589 81
rect 1659 35 1705 81
rect 1775 35 1821 81
rect 1891 35 1937 81
rect 2007 35 2053 81
rect 2123 35 2169 81
rect 2239 35 2285 81
rect 2355 35 2401 81
rect 2471 35 2517 81
rect 2587 35 2633 81
rect 2703 35 2749 81
rect 2819 35 2865 81
rect 2935 35 2981 81
rect 3051 35 3097 81
rect 3167 35 3213 81
rect 3283 35 3329 81
rect 3399 35 3445 81
rect 3515 35 3561 81
rect 3631 35 3677 81
rect 3747 35 3793 81
rect 3863 35 3909 81
rect 3979 35 4025 81
rect 4095 35 4141 81
rect 4211 35 4257 81
rect 4327 35 4373 81
rect 4443 35 4489 81
rect 4559 35 4605 81
rect 4675 35 4721 81
rect 4791 35 4837 81
rect 4907 35 4953 81
rect 5023 35 5069 81
rect 5139 35 5185 81
rect 5255 35 5301 81
rect 5371 35 5417 81
rect 5487 35 5533 81
rect 5603 35 5649 81
rect 5719 35 5765 81
rect -5765 -81 -5719 -35
rect -5649 -81 -5603 -35
rect -5533 -81 -5487 -35
rect -5417 -81 -5371 -35
rect -5301 -81 -5255 -35
rect -5185 -81 -5139 -35
rect -5069 -81 -5023 -35
rect -4953 -81 -4907 -35
rect -4837 -81 -4791 -35
rect -4721 -81 -4675 -35
rect -4605 -81 -4559 -35
rect -4489 -81 -4443 -35
rect -4373 -81 -4327 -35
rect -4257 -81 -4211 -35
rect -4141 -81 -4095 -35
rect -4025 -81 -3979 -35
rect -3909 -81 -3863 -35
rect -3793 -81 -3747 -35
rect -3677 -81 -3631 -35
rect -3561 -81 -3515 -35
rect -3445 -81 -3399 -35
rect -3329 -81 -3283 -35
rect -3213 -81 -3167 -35
rect -3097 -81 -3051 -35
rect -2981 -81 -2935 -35
rect -2865 -81 -2819 -35
rect -2749 -81 -2703 -35
rect -2633 -81 -2587 -35
rect -2517 -81 -2471 -35
rect -2401 -81 -2355 -35
rect -2285 -81 -2239 -35
rect -2169 -81 -2123 -35
rect -2053 -81 -2007 -35
rect -1937 -81 -1891 -35
rect -1821 -81 -1775 -35
rect -1705 -81 -1659 -35
rect -1589 -81 -1543 -35
rect -1473 -81 -1427 -35
rect -1357 -81 -1311 -35
rect -1241 -81 -1195 -35
rect -1125 -81 -1079 -35
rect -1009 -81 -963 -35
rect -893 -81 -847 -35
rect -777 -81 -731 -35
rect -661 -81 -615 -35
rect -545 -81 -499 -35
rect -429 -81 -383 -35
rect -313 -81 -267 -35
rect -197 -81 -151 -35
rect -81 -81 -35 -35
rect 35 -81 81 -35
rect 151 -81 197 -35
rect 267 -81 313 -35
rect 383 -81 429 -35
rect 499 -81 545 -35
rect 615 -81 661 -35
rect 731 -81 777 -35
rect 847 -81 893 -35
rect 963 -81 1009 -35
rect 1079 -81 1125 -35
rect 1195 -81 1241 -35
rect 1311 -81 1357 -35
rect 1427 -81 1473 -35
rect 1543 -81 1589 -35
rect 1659 -81 1705 -35
rect 1775 -81 1821 -35
rect 1891 -81 1937 -35
rect 2007 -81 2053 -35
rect 2123 -81 2169 -35
rect 2239 -81 2285 -35
rect 2355 -81 2401 -35
rect 2471 -81 2517 -35
rect 2587 -81 2633 -35
rect 2703 -81 2749 -35
rect 2819 -81 2865 -35
rect 2935 -81 2981 -35
rect 3051 -81 3097 -35
rect 3167 -81 3213 -35
rect 3283 -81 3329 -35
rect 3399 -81 3445 -35
rect 3515 -81 3561 -35
rect 3631 -81 3677 -35
rect 3747 -81 3793 -35
rect 3863 -81 3909 -35
rect 3979 -81 4025 -35
rect 4095 -81 4141 -35
rect 4211 -81 4257 -35
rect 4327 -81 4373 -35
rect 4443 -81 4489 -35
rect 4559 -81 4605 -35
rect 4675 -81 4721 -35
rect 4791 -81 4837 -35
rect 4907 -81 4953 -35
rect 5023 -81 5069 -35
rect 5139 -81 5185 -35
rect 5255 -81 5301 -35
rect 5371 -81 5417 -35
rect 5487 -81 5533 -35
rect 5603 -81 5649 -35
rect 5719 -81 5765 -35
rect -5765 -197 -5719 -151
rect -5649 -197 -5603 -151
rect -5533 -197 -5487 -151
rect -5417 -197 -5371 -151
rect -5301 -197 -5255 -151
rect -5185 -197 -5139 -151
rect -5069 -197 -5023 -151
rect -4953 -197 -4907 -151
rect -4837 -197 -4791 -151
rect -4721 -197 -4675 -151
rect -4605 -197 -4559 -151
rect -4489 -197 -4443 -151
rect -4373 -197 -4327 -151
rect -4257 -197 -4211 -151
rect -4141 -197 -4095 -151
rect -4025 -197 -3979 -151
rect -3909 -197 -3863 -151
rect -3793 -197 -3747 -151
rect -3677 -197 -3631 -151
rect -3561 -197 -3515 -151
rect -3445 -197 -3399 -151
rect -3329 -197 -3283 -151
rect -3213 -197 -3167 -151
rect -3097 -197 -3051 -151
rect -2981 -197 -2935 -151
rect -2865 -197 -2819 -151
rect -2749 -197 -2703 -151
rect -2633 -197 -2587 -151
rect -2517 -197 -2471 -151
rect -2401 -197 -2355 -151
rect -2285 -197 -2239 -151
rect -2169 -197 -2123 -151
rect -2053 -197 -2007 -151
rect -1937 -197 -1891 -151
rect -1821 -197 -1775 -151
rect -1705 -197 -1659 -151
rect -1589 -197 -1543 -151
rect -1473 -197 -1427 -151
rect -1357 -197 -1311 -151
rect -1241 -197 -1195 -151
rect -1125 -197 -1079 -151
rect -1009 -197 -963 -151
rect -893 -197 -847 -151
rect -777 -197 -731 -151
rect -661 -197 -615 -151
rect -545 -197 -499 -151
rect -429 -197 -383 -151
rect -313 -197 -267 -151
rect -197 -197 -151 -151
rect -81 -197 -35 -151
rect 35 -197 81 -151
rect 151 -197 197 -151
rect 267 -197 313 -151
rect 383 -197 429 -151
rect 499 -197 545 -151
rect 615 -197 661 -151
rect 731 -197 777 -151
rect 847 -197 893 -151
rect 963 -197 1009 -151
rect 1079 -197 1125 -151
rect 1195 -197 1241 -151
rect 1311 -197 1357 -151
rect 1427 -197 1473 -151
rect 1543 -197 1589 -151
rect 1659 -197 1705 -151
rect 1775 -197 1821 -151
rect 1891 -197 1937 -151
rect 2007 -197 2053 -151
rect 2123 -197 2169 -151
rect 2239 -197 2285 -151
rect 2355 -197 2401 -151
rect 2471 -197 2517 -151
rect 2587 -197 2633 -151
rect 2703 -197 2749 -151
rect 2819 -197 2865 -151
rect 2935 -197 2981 -151
rect 3051 -197 3097 -151
rect 3167 -197 3213 -151
rect 3283 -197 3329 -151
rect 3399 -197 3445 -151
rect 3515 -197 3561 -151
rect 3631 -197 3677 -151
rect 3747 -197 3793 -151
rect 3863 -197 3909 -151
rect 3979 -197 4025 -151
rect 4095 -197 4141 -151
rect 4211 -197 4257 -151
rect 4327 -197 4373 -151
rect 4443 -197 4489 -151
rect 4559 -197 4605 -151
rect 4675 -197 4721 -151
rect 4791 -197 4837 -151
rect 4907 -197 4953 -151
rect 5023 -197 5069 -151
rect 5139 -197 5185 -151
rect 5255 -197 5301 -151
rect 5371 -197 5417 -151
rect 5487 -197 5533 -151
rect 5603 -197 5649 -151
rect 5719 -197 5765 -151
rect -5765 -313 -5719 -267
rect -5649 -313 -5603 -267
rect -5533 -313 -5487 -267
rect -5417 -313 -5371 -267
rect -5301 -313 -5255 -267
rect -5185 -313 -5139 -267
rect -5069 -313 -5023 -267
rect -4953 -313 -4907 -267
rect -4837 -313 -4791 -267
rect -4721 -313 -4675 -267
rect -4605 -313 -4559 -267
rect -4489 -313 -4443 -267
rect -4373 -313 -4327 -267
rect -4257 -313 -4211 -267
rect -4141 -313 -4095 -267
rect -4025 -313 -3979 -267
rect -3909 -313 -3863 -267
rect -3793 -313 -3747 -267
rect -3677 -313 -3631 -267
rect -3561 -313 -3515 -267
rect -3445 -313 -3399 -267
rect -3329 -313 -3283 -267
rect -3213 -313 -3167 -267
rect -3097 -313 -3051 -267
rect -2981 -313 -2935 -267
rect -2865 -313 -2819 -267
rect -2749 -313 -2703 -267
rect -2633 -313 -2587 -267
rect -2517 -313 -2471 -267
rect -2401 -313 -2355 -267
rect -2285 -313 -2239 -267
rect -2169 -313 -2123 -267
rect -2053 -313 -2007 -267
rect -1937 -313 -1891 -267
rect -1821 -313 -1775 -267
rect -1705 -313 -1659 -267
rect -1589 -313 -1543 -267
rect -1473 -313 -1427 -267
rect -1357 -313 -1311 -267
rect -1241 -313 -1195 -267
rect -1125 -313 -1079 -267
rect -1009 -313 -963 -267
rect -893 -313 -847 -267
rect -777 -313 -731 -267
rect -661 -313 -615 -267
rect -545 -313 -499 -267
rect -429 -313 -383 -267
rect -313 -313 -267 -267
rect -197 -313 -151 -267
rect -81 -313 -35 -267
rect 35 -313 81 -267
rect 151 -313 197 -267
rect 267 -313 313 -267
rect 383 -313 429 -267
rect 499 -313 545 -267
rect 615 -313 661 -267
rect 731 -313 777 -267
rect 847 -313 893 -267
rect 963 -313 1009 -267
rect 1079 -313 1125 -267
rect 1195 -313 1241 -267
rect 1311 -313 1357 -267
rect 1427 -313 1473 -267
rect 1543 -313 1589 -267
rect 1659 -313 1705 -267
rect 1775 -313 1821 -267
rect 1891 -313 1937 -267
rect 2007 -313 2053 -267
rect 2123 -313 2169 -267
rect 2239 -313 2285 -267
rect 2355 -313 2401 -267
rect 2471 -313 2517 -267
rect 2587 -313 2633 -267
rect 2703 -313 2749 -267
rect 2819 -313 2865 -267
rect 2935 -313 2981 -267
rect 3051 -313 3097 -267
rect 3167 -313 3213 -267
rect 3283 -313 3329 -267
rect 3399 -313 3445 -267
rect 3515 -313 3561 -267
rect 3631 -313 3677 -267
rect 3747 -313 3793 -267
rect 3863 -313 3909 -267
rect 3979 -313 4025 -267
rect 4095 -313 4141 -267
rect 4211 -313 4257 -267
rect 4327 -313 4373 -267
rect 4443 -313 4489 -267
rect 4559 -313 4605 -267
rect 4675 -313 4721 -267
rect 4791 -313 4837 -267
rect 4907 -313 4953 -267
rect 5023 -313 5069 -267
rect 5139 -313 5185 -267
rect 5255 -313 5301 -267
rect 5371 -313 5417 -267
rect 5487 -313 5533 -267
rect 5603 -313 5649 -267
rect 5719 -313 5765 -267
rect -5765 -429 -5719 -383
rect -5649 -429 -5603 -383
rect -5533 -429 -5487 -383
rect -5417 -429 -5371 -383
rect -5301 -429 -5255 -383
rect -5185 -429 -5139 -383
rect -5069 -429 -5023 -383
rect -4953 -429 -4907 -383
rect -4837 -429 -4791 -383
rect -4721 -429 -4675 -383
rect -4605 -429 -4559 -383
rect -4489 -429 -4443 -383
rect -4373 -429 -4327 -383
rect -4257 -429 -4211 -383
rect -4141 -429 -4095 -383
rect -4025 -429 -3979 -383
rect -3909 -429 -3863 -383
rect -3793 -429 -3747 -383
rect -3677 -429 -3631 -383
rect -3561 -429 -3515 -383
rect -3445 -429 -3399 -383
rect -3329 -429 -3283 -383
rect -3213 -429 -3167 -383
rect -3097 -429 -3051 -383
rect -2981 -429 -2935 -383
rect -2865 -429 -2819 -383
rect -2749 -429 -2703 -383
rect -2633 -429 -2587 -383
rect -2517 -429 -2471 -383
rect -2401 -429 -2355 -383
rect -2285 -429 -2239 -383
rect -2169 -429 -2123 -383
rect -2053 -429 -2007 -383
rect -1937 -429 -1891 -383
rect -1821 -429 -1775 -383
rect -1705 -429 -1659 -383
rect -1589 -429 -1543 -383
rect -1473 -429 -1427 -383
rect -1357 -429 -1311 -383
rect -1241 -429 -1195 -383
rect -1125 -429 -1079 -383
rect -1009 -429 -963 -383
rect -893 -429 -847 -383
rect -777 -429 -731 -383
rect -661 -429 -615 -383
rect -545 -429 -499 -383
rect -429 -429 -383 -383
rect -313 -429 -267 -383
rect -197 -429 -151 -383
rect -81 -429 -35 -383
rect 35 -429 81 -383
rect 151 -429 197 -383
rect 267 -429 313 -383
rect 383 -429 429 -383
rect 499 -429 545 -383
rect 615 -429 661 -383
rect 731 -429 777 -383
rect 847 -429 893 -383
rect 963 -429 1009 -383
rect 1079 -429 1125 -383
rect 1195 -429 1241 -383
rect 1311 -429 1357 -383
rect 1427 -429 1473 -383
rect 1543 -429 1589 -383
rect 1659 -429 1705 -383
rect 1775 -429 1821 -383
rect 1891 -429 1937 -383
rect 2007 -429 2053 -383
rect 2123 -429 2169 -383
rect 2239 -429 2285 -383
rect 2355 -429 2401 -383
rect 2471 -429 2517 -383
rect 2587 -429 2633 -383
rect 2703 -429 2749 -383
rect 2819 -429 2865 -383
rect 2935 -429 2981 -383
rect 3051 -429 3097 -383
rect 3167 -429 3213 -383
rect 3283 -429 3329 -383
rect 3399 -429 3445 -383
rect 3515 -429 3561 -383
rect 3631 -429 3677 -383
rect 3747 -429 3793 -383
rect 3863 -429 3909 -383
rect 3979 -429 4025 -383
rect 4095 -429 4141 -383
rect 4211 -429 4257 -383
rect 4327 -429 4373 -383
rect 4443 -429 4489 -383
rect 4559 -429 4605 -383
rect 4675 -429 4721 -383
rect 4791 -429 4837 -383
rect 4907 -429 4953 -383
rect 5023 -429 5069 -383
rect 5139 -429 5185 -383
rect 5255 -429 5301 -383
rect 5371 -429 5417 -383
rect 5487 -429 5533 -383
rect 5603 -429 5649 -383
rect 5719 -429 5765 -383
rect -5765 -545 -5719 -499
rect -5649 -545 -5603 -499
rect -5533 -545 -5487 -499
rect -5417 -545 -5371 -499
rect -5301 -545 -5255 -499
rect -5185 -545 -5139 -499
rect -5069 -545 -5023 -499
rect -4953 -545 -4907 -499
rect -4837 -545 -4791 -499
rect -4721 -545 -4675 -499
rect -4605 -545 -4559 -499
rect -4489 -545 -4443 -499
rect -4373 -545 -4327 -499
rect -4257 -545 -4211 -499
rect -4141 -545 -4095 -499
rect -4025 -545 -3979 -499
rect -3909 -545 -3863 -499
rect -3793 -545 -3747 -499
rect -3677 -545 -3631 -499
rect -3561 -545 -3515 -499
rect -3445 -545 -3399 -499
rect -3329 -545 -3283 -499
rect -3213 -545 -3167 -499
rect -3097 -545 -3051 -499
rect -2981 -545 -2935 -499
rect -2865 -545 -2819 -499
rect -2749 -545 -2703 -499
rect -2633 -545 -2587 -499
rect -2517 -545 -2471 -499
rect -2401 -545 -2355 -499
rect -2285 -545 -2239 -499
rect -2169 -545 -2123 -499
rect -2053 -545 -2007 -499
rect -1937 -545 -1891 -499
rect -1821 -545 -1775 -499
rect -1705 -545 -1659 -499
rect -1589 -545 -1543 -499
rect -1473 -545 -1427 -499
rect -1357 -545 -1311 -499
rect -1241 -545 -1195 -499
rect -1125 -545 -1079 -499
rect -1009 -545 -963 -499
rect -893 -545 -847 -499
rect -777 -545 -731 -499
rect -661 -545 -615 -499
rect -545 -545 -499 -499
rect -429 -545 -383 -499
rect -313 -545 -267 -499
rect -197 -545 -151 -499
rect -81 -545 -35 -499
rect 35 -545 81 -499
rect 151 -545 197 -499
rect 267 -545 313 -499
rect 383 -545 429 -499
rect 499 -545 545 -499
rect 615 -545 661 -499
rect 731 -545 777 -499
rect 847 -545 893 -499
rect 963 -545 1009 -499
rect 1079 -545 1125 -499
rect 1195 -545 1241 -499
rect 1311 -545 1357 -499
rect 1427 -545 1473 -499
rect 1543 -545 1589 -499
rect 1659 -545 1705 -499
rect 1775 -545 1821 -499
rect 1891 -545 1937 -499
rect 2007 -545 2053 -499
rect 2123 -545 2169 -499
rect 2239 -545 2285 -499
rect 2355 -545 2401 -499
rect 2471 -545 2517 -499
rect 2587 -545 2633 -499
rect 2703 -545 2749 -499
rect 2819 -545 2865 -499
rect 2935 -545 2981 -499
rect 3051 -545 3097 -499
rect 3167 -545 3213 -499
rect 3283 -545 3329 -499
rect 3399 -545 3445 -499
rect 3515 -545 3561 -499
rect 3631 -545 3677 -499
rect 3747 -545 3793 -499
rect 3863 -545 3909 -499
rect 3979 -545 4025 -499
rect 4095 -545 4141 -499
rect 4211 -545 4257 -499
rect 4327 -545 4373 -499
rect 4443 -545 4489 -499
rect 4559 -545 4605 -499
rect 4675 -545 4721 -499
rect 4791 -545 4837 -499
rect 4907 -545 4953 -499
rect 5023 -545 5069 -499
rect 5139 -545 5185 -499
rect 5255 -545 5301 -499
rect 5371 -545 5417 -499
rect 5487 -545 5533 -499
rect 5603 -545 5649 -499
rect 5719 -545 5765 -499
rect -5765 -661 -5719 -615
rect -5649 -661 -5603 -615
rect -5533 -661 -5487 -615
rect -5417 -661 -5371 -615
rect -5301 -661 -5255 -615
rect -5185 -661 -5139 -615
rect -5069 -661 -5023 -615
rect -4953 -661 -4907 -615
rect -4837 -661 -4791 -615
rect -4721 -661 -4675 -615
rect -4605 -661 -4559 -615
rect -4489 -661 -4443 -615
rect -4373 -661 -4327 -615
rect -4257 -661 -4211 -615
rect -4141 -661 -4095 -615
rect -4025 -661 -3979 -615
rect -3909 -661 -3863 -615
rect -3793 -661 -3747 -615
rect -3677 -661 -3631 -615
rect -3561 -661 -3515 -615
rect -3445 -661 -3399 -615
rect -3329 -661 -3283 -615
rect -3213 -661 -3167 -615
rect -3097 -661 -3051 -615
rect -2981 -661 -2935 -615
rect -2865 -661 -2819 -615
rect -2749 -661 -2703 -615
rect -2633 -661 -2587 -615
rect -2517 -661 -2471 -615
rect -2401 -661 -2355 -615
rect -2285 -661 -2239 -615
rect -2169 -661 -2123 -615
rect -2053 -661 -2007 -615
rect -1937 -661 -1891 -615
rect -1821 -661 -1775 -615
rect -1705 -661 -1659 -615
rect -1589 -661 -1543 -615
rect -1473 -661 -1427 -615
rect -1357 -661 -1311 -615
rect -1241 -661 -1195 -615
rect -1125 -661 -1079 -615
rect -1009 -661 -963 -615
rect -893 -661 -847 -615
rect -777 -661 -731 -615
rect -661 -661 -615 -615
rect -545 -661 -499 -615
rect -429 -661 -383 -615
rect -313 -661 -267 -615
rect -197 -661 -151 -615
rect -81 -661 -35 -615
rect 35 -661 81 -615
rect 151 -661 197 -615
rect 267 -661 313 -615
rect 383 -661 429 -615
rect 499 -661 545 -615
rect 615 -661 661 -615
rect 731 -661 777 -615
rect 847 -661 893 -615
rect 963 -661 1009 -615
rect 1079 -661 1125 -615
rect 1195 -661 1241 -615
rect 1311 -661 1357 -615
rect 1427 -661 1473 -615
rect 1543 -661 1589 -615
rect 1659 -661 1705 -615
rect 1775 -661 1821 -615
rect 1891 -661 1937 -615
rect 2007 -661 2053 -615
rect 2123 -661 2169 -615
rect 2239 -661 2285 -615
rect 2355 -661 2401 -615
rect 2471 -661 2517 -615
rect 2587 -661 2633 -615
rect 2703 -661 2749 -615
rect 2819 -661 2865 -615
rect 2935 -661 2981 -615
rect 3051 -661 3097 -615
rect 3167 -661 3213 -615
rect 3283 -661 3329 -615
rect 3399 -661 3445 -615
rect 3515 -661 3561 -615
rect 3631 -661 3677 -615
rect 3747 -661 3793 -615
rect 3863 -661 3909 -615
rect 3979 -661 4025 -615
rect 4095 -661 4141 -615
rect 4211 -661 4257 -615
rect 4327 -661 4373 -615
rect 4443 -661 4489 -615
rect 4559 -661 4605 -615
rect 4675 -661 4721 -615
rect 4791 -661 4837 -615
rect 4907 -661 4953 -615
rect 5023 -661 5069 -615
rect 5139 -661 5185 -615
rect 5255 -661 5301 -615
rect 5371 -661 5417 -615
rect 5487 -661 5533 -615
rect 5603 -661 5649 -615
rect 5719 -661 5765 -615
rect -5765 -777 -5719 -731
rect -5649 -777 -5603 -731
rect -5533 -777 -5487 -731
rect -5417 -777 -5371 -731
rect -5301 -777 -5255 -731
rect -5185 -777 -5139 -731
rect -5069 -777 -5023 -731
rect -4953 -777 -4907 -731
rect -4837 -777 -4791 -731
rect -4721 -777 -4675 -731
rect -4605 -777 -4559 -731
rect -4489 -777 -4443 -731
rect -4373 -777 -4327 -731
rect -4257 -777 -4211 -731
rect -4141 -777 -4095 -731
rect -4025 -777 -3979 -731
rect -3909 -777 -3863 -731
rect -3793 -777 -3747 -731
rect -3677 -777 -3631 -731
rect -3561 -777 -3515 -731
rect -3445 -777 -3399 -731
rect -3329 -777 -3283 -731
rect -3213 -777 -3167 -731
rect -3097 -777 -3051 -731
rect -2981 -777 -2935 -731
rect -2865 -777 -2819 -731
rect -2749 -777 -2703 -731
rect -2633 -777 -2587 -731
rect -2517 -777 -2471 -731
rect -2401 -777 -2355 -731
rect -2285 -777 -2239 -731
rect -2169 -777 -2123 -731
rect -2053 -777 -2007 -731
rect -1937 -777 -1891 -731
rect -1821 -777 -1775 -731
rect -1705 -777 -1659 -731
rect -1589 -777 -1543 -731
rect -1473 -777 -1427 -731
rect -1357 -777 -1311 -731
rect -1241 -777 -1195 -731
rect -1125 -777 -1079 -731
rect -1009 -777 -963 -731
rect -893 -777 -847 -731
rect -777 -777 -731 -731
rect -661 -777 -615 -731
rect -545 -777 -499 -731
rect -429 -777 -383 -731
rect -313 -777 -267 -731
rect -197 -777 -151 -731
rect -81 -777 -35 -731
rect 35 -777 81 -731
rect 151 -777 197 -731
rect 267 -777 313 -731
rect 383 -777 429 -731
rect 499 -777 545 -731
rect 615 -777 661 -731
rect 731 -777 777 -731
rect 847 -777 893 -731
rect 963 -777 1009 -731
rect 1079 -777 1125 -731
rect 1195 -777 1241 -731
rect 1311 -777 1357 -731
rect 1427 -777 1473 -731
rect 1543 -777 1589 -731
rect 1659 -777 1705 -731
rect 1775 -777 1821 -731
rect 1891 -777 1937 -731
rect 2007 -777 2053 -731
rect 2123 -777 2169 -731
rect 2239 -777 2285 -731
rect 2355 -777 2401 -731
rect 2471 -777 2517 -731
rect 2587 -777 2633 -731
rect 2703 -777 2749 -731
rect 2819 -777 2865 -731
rect 2935 -777 2981 -731
rect 3051 -777 3097 -731
rect 3167 -777 3213 -731
rect 3283 -777 3329 -731
rect 3399 -777 3445 -731
rect 3515 -777 3561 -731
rect 3631 -777 3677 -731
rect 3747 -777 3793 -731
rect 3863 -777 3909 -731
rect 3979 -777 4025 -731
rect 4095 -777 4141 -731
rect 4211 -777 4257 -731
rect 4327 -777 4373 -731
rect 4443 -777 4489 -731
rect 4559 -777 4605 -731
rect 4675 -777 4721 -731
rect 4791 -777 4837 -731
rect 4907 -777 4953 -731
rect 5023 -777 5069 -731
rect 5139 -777 5185 -731
rect 5255 -777 5301 -731
rect 5371 -777 5417 -731
rect 5487 -777 5533 -731
rect 5603 -777 5649 -731
rect 5719 -777 5765 -731
rect -5765 -893 -5719 -847
rect -5649 -893 -5603 -847
rect -5533 -893 -5487 -847
rect -5417 -893 -5371 -847
rect -5301 -893 -5255 -847
rect -5185 -893 -5139 -847
rect -5069 -893 -5023 -847
rect -4953 -893 -4907 -847
rect -4837 -893 -4791 -847
rect -4721 -893 -4675 -847
rect -4605 -893 -4559 -847
rect -4489 -893 -4443 -847
rect -4373 -893 -4327 -847
rect -4257 -893 -4211 -847
rect -4141 -893 -4095 -847
rect -4025 -893 -3979 -847
rect -3909 -893 -3863 -847
rect -3793 -893 -3747 -847
rect -3677 -893 -3631 -847
rect -3561 -893 -3515 -847
rect -3445 -893 -3399 -847
rect -3329 -893 -3283 -847
rect -3213 -893 -3167 -847
rect -3097 -893 -3051 -847
rect -2981 -893 -2935 -847
rect -2865 -893 -2819 -847
rect -2749 -893 -2703 -847
rect -2633 -893 -2587 -847
rect -2517 -893 -2471 -847
rect -2401 -893 -2355 -847
rect -2285 -893 -2239 -847
rect -2169 -893 -2123 -847
rect -2053 -893 -2007 -847
rect -1937 -893 -1891 -847
rect -1821 -893 -1775 -847
rect -1705 -893 -1659 -847
rect -1589 -893 -1543 -847
rect -1473 -893 -1427 -847
rect -1357 -893 -1311 -847
rect -1241 -893 -1195 -847
rect -1125 -893 -1079 -847
rect -1009 -893 -963 -847
rect -893 -893 -847 -847
rect -777 -893 -731 -847
rect -661 -893 -615 -847
rect -545 -893 -499 -847
rect -429 -893 -383 -847
rect -313 -893 -267 -847
rect -197 -893 -151 -847
rect -81 -893 -35 -847
rect 35 -893 81 -847
rect 151 -893 197 -847
rect 267 -893 313 -847
rect 383 -893 429 -847
rect 499 -893 545 -847
rect 615 -893 661 -847
rect 731 -893 777 -847
rect 847 -893 893 -847
rect 963 -893 1009 -847
rect 1079 -893 1125 -847
rect 1195 -893 1241 -847
rect 1311 -893 1357 -847
rect 1427 -893 1473 -847
rect 1543 -893 1589 -847
rect 1659 -893 1705 -847
rect 1775 -893 1821 -847
rect 1891 -893 1937 -847
rect 2007 -893 2053 -847
rect 2123 -893 2169 -847
rect 2239 -893 2285 -847
rect 2355 -893 2401 -847
rect 2471 -893 2517 -847
rect 2587 -893 2633 -847
rect 2703 -893 2749 -847
rect 2819 -893 2865 -847
rect 2935 -893 2981 -847
rect 3051 -893 3097 -847
rect 3167 -893 3213 -847
rect 3283 -893 3329 -847
rect 3399 -893 3445 -847
rect 3515 -893 3561 -847
rect 3631 -893 3677 -847
rect 3747 -893 3793 -847
rect 3863 -893 3909 -847
rect 3979 -893 4025 -847
rect 4095 -893 4141 -847
rect 4211 -893 4257 -847
rect 4327 -893 4373 -847
rect 4443 -893 4489 -847
rect 4559 -893 4605 -847
rect 4675 -893 4721 -847
rect 4791 -893 4837 -847
rect 4907 -893 4953 -847
rect 5023 -893 5069 -847
rect 5139 -893 5185 -847
rect 5255 -893 5301 -847
rect 5371 -893 5417 -847
rect 5487 -893 5533 -847
rect 5603 -893 5649 -847
rect 5719 -893 5765 -847
rect -5765 -1009 -5719 -963
rect -5649 -1009 -5603 -963
rect -5533 -1009 -5487 -963
rect -5417 -1009 -5371 -963
rect -5301 -1009 -5255 -963
rect -5185 -1009 -5139 -963
rect -5069 -1009 -5023 -963
rect -4953 -1009 -4907 -963
rect -4837 -1009 -4791 -963
rect -4721 -1009 -4675 -963
rect -4605 -1009 -4559 -963
rect -4489 -1009 -4443 -963
rect -4373 -1009 -4327 -963
rect -4257 -1009 -4211 -963
rect -4141 -1009 -4095 -963
rect -4025 -1009 -3979 -963
rect -3909 -1009 -3863 -963
rect -3793 -1009 -3747 -963
rect -3677 -1009 -3631 -963
rect -3561 -1009 -3515 -963
rect -3445 -1009 -3399 -963
rect -3329 -1009 -3283 -963
rect -3213 -1009 -3167 -963
rect -3097 -1009 -3051 -963
rect -2981 -1009 -2935 -963
rect -2865 -1009 -2819 -963
rect -2749 -1009 -2703 -963
rect -2633 -1009 -2587 -963
rect -2517 -1009 -2471 -963
rect -2401 -1009 -2355 -963
rect -2285 -1009 -2239 -963
rect -2169 -1009 -2123 -963
rect -2053 -1009 -2007 -963
rect -1937 -1009 -1891 -963
rect -1821 -1009 -1775 -963
rect -1705 -1009 -1659 -963
rect -1589 -1009 -1543 -963
rect -1473 -1009 -1427 -963
rect -1357 -1009 -1311 -963
rect -1241 -1009 -1195 -963
rect -1125 -1009 -1079 -963
rect -1009 -1009 -963 -963
rect -893 -1009 -847 -963
rect -777 -1009 -731 -963
rect -661 -1009 -615 -963
rect -545 -1009 -499 -963
rect -429 -1009 -383 -963
rect -313 -1009 -267 -963
rect -197 -1009 -151 -963
rect -81 -1009 -35 -963
rect 35 -1009 81 -963
rect 151 -1009 197 -963
rect 267 -1009 313 -963
rect 383 -1009 429 -963
rect 499 -1009 545 -963
rect 615 -1009 661 -963
rect 731 -1009 777 -963
rect 847 -1009 893 -963
rect 963 -1009 1009 -963
rect 1079 -1009 1125 -963
rect 1195 -1009 1241 -963
rect 1311 -1009 1357 -963
rect 1427 -1009 1473 -963
rect 1543 -1009 1589 -963
rect 1659 -1009 1705 -963
rect 1775 -1009 1821 -963
rect 1891 -1009 1937 -963
rect 2007 -1009 2053 -963
rect 2123 -1009 2169 -963
rect 2239 -1009 2285 -963
rect 2355 -1009 2401 -963
rect 2471 -1009 2517 -963
rect 2587 -1009 2633 -963
rect 2703 -1009 2749 -963
rect 2819 -1009 2865 -963
rect 2935 -1009 2981 -963
rect 3051 -1009 3097 -963
rect 3167 -1009 3213 -963
rect 3283 -1009 3329 -963
rect 3399 -1009 3445 -963
rect 3515 -1009 3561 -963
rect 3631 -1009 3677 -963
rect 3747 -1009 3793 -963
rect 3863 -1009 3909 -963
rect 3979 -1009 4025 -963
rect 4095 -1009 4141 -963
rect 4211 -1009 4257 -963
rect 4327 -1009 4373 -963
rect 4443 -1009 4489 -963
rect 4559 -1009 4605 -963
rect 4675 -1009 4721 -963
rect 4791 -1009 4837 -963
rect 4907 -1009 4953 -963
rect 5023 -1009 5069 -963
rect 5139 -1009 5185 -963
rect 5255 -1009 5301 -963
rect 5371 -1009 5417 -963
rect 5487 -1009 5533 -963
rect 5603 -1009 5649 -963
rect 5719 -1009 5765 -963
rect -5765 -1125 -5719 -1079
rect -5649 -1125 -5603 -1079
rect -5533 -1125 -5487 -1079
rect -5417 -1125 -5371 -1079
rect -5301 -1125 -5255 -1079
rect -5185 -1125 -5139 -1079
rect -5069 -1125 -5023 -1079
rect -4953 -1125 -4907 -1079
rect -4837 -1125 -4791 -1079
rect -4721 -1125 -4675 -1079
rect -4605 -1125 -4559 -1079
rect -4489 -1125 -4443 -1079
rect -4373 -1125 -4327 -1079
rect -4257 -1125 -4211 -1079
rect -4141 -1125 -4095 -1079
rect -4025 -1125 -3979 -1079
rect -3909 -1125 -3863 -1079
rect -3793 -1125 -3747 -1079
rect -3677 -1125 -3631 -1079
rect -3561 -1125 -3515 -1079
rect -3445 -1125 -3399 -1079
rect -3329 -1125 -3283 -1079
rect -3213 -1125 -3167 -1079
rect -3097 -1125 -3051 -1079
rect -2981 -1125 -2935 -1079
rect -2865 -1125 -2819 -1079
rect -2749 -1125 -2703 -1079
rect -2633 -1125 -2587 -1079
rect -2517 -1125 -2471 -1079
rect -2401 -1125 -2355 -1079
rect -2285 -1125 -2239 -1079
rect -2169 -1125 -2123 -1079
rect -2053 -1125 -2007 -1079
rect -1937 -1125 -1891 -1079
rect -1821 -1125 -1775 -1079
rect -1705 -1125 -1659 -1079
rect -1589 -1125 -1543 -1079
rect -1473 -1125 -1427 -1079
rect -1357 -1125 -1311 -1079
rect -1241 -1125 -1195 -1079
rect -1125 -1125 -1079 -1079
rect -1009 -1125 -963 -1079
rect -893 -1125 -847 -1079
rect -777 -1125 -731 -1079
rect -661 -1125 -615 -1079
rect -545 -1125 -499 -1079
rect -429 -1125 -383 -1079
rect -313 -1125 -267 -1079
rect -197 -1125 -151 -1079
rect -81 -1125 -35 -1079
rect 35 -1125 81 -1079
rect 151 -1125 197 -1079
rect 267 -1125 313 -1079
rect 383 -1125 429 -1079
rect 499 -1125 545 -1079
rect 615 -1125 661 -1079
rect 731 -1125 777 -1079
rect 847 -1125 893 -1079
rect 963 -1125 1009 -1079
rect 1079 -1125 1125 -1079
rect 1195 -1125 1241 -1079
rect 1311 -1125 1357 -1079
rect 1427 -1125 1473 -1079
rect 1543 -1125 1589 -1079
rect 1659 -1125 1705 -1079
rect 1775 -1125 1821 -1079
rect 1891 -1125 1937 -1079
rect 2007 -1125 2053 -1079
rect 2123 -1125 2169 -1079
rect 2239 -1125 2285 -1079
rect 2355 -1125 2401 -1079
rect 2471 -1125 2517 -1079
rect 2587 -1125 2633 -1079
rect 2703 -1125 2749 -1079
rect 2819 -1125 2865 -1079
rect 2935 -1125 2981 -1079
rect 3051 -1125 3097 -1079
rect 3167 -1125 3213 -1079
rect 3283 -1125 3329 -1079
rect 3399 -1125 3445 -1079
rect 3515 -1125 3561 -1079
rect 3631 -1125 3677 -1079
rect 3747 -1125 3793 -1079
rect 3863 -1125 3909 -1079
rect 3979 -1125 4025 -1079
rect 4095 -1125 4141 -1079
rect 4211 -1125 4257 -1079
rect 4327 -1125 4373 -1079
rect 4443 -1125 4489 -1079
rect 4559 -1125 4605 -1079
rect 4675 -1125 4721 -1079
rect 4791 -1125 4837 -1079
rect 4907 -1125 4953 -1079
rect 5023 -1125 5069 -1079
rect 5139 -1125 5185 -1079
rect 5255 -1125 5301 -1079
rect 5371 -1125 5417 -1079
rect 5487 -1125 5533 -1079
rect 5603 -1125 5649 -1079
rect 5719 -1125 5765 -1079
<< metal1 >>
rect -5776 1125 5776 1136
rect -5776 1079 -5765 1125
rect -5719 1079 -5649 1125
rect -5603 1079 -5533 1125
rect -5487 1079 -5417 1125
rect -5371 1079 -5301 1125
rect -5255 1079 -5185 1125
rect -5139 1079 -5069 1125
rect -5023 1079 -4953 1125
rect -4907 1079 -4837 1125
rect -4791 1079 -4721 1125
rect -4675 1079 -4605 1125
rect -4559 1079 -4489 1125
rect -4443 1079 -4373 1125
rect -4327 1079 -4257 1125
rect -4211 1079 -4141 1125
rect -4095 1079 -4025 1125
rect -3979 1079 -3909 1125
rect -3863 1079 -3793 1125
rect -3747 1079 -3677 1125
rect -3631 1079 -3561 1125
rect -3515 1079 -3445 1125
rect -3399 1079 -3329 1125
rect -3283 1079 -3213 1125
rect -3167 1079 -3097 1125
rect -3051 1079 -2981 1125
rect -2935 1079 -2865 1125
rect -2819 1079 -2749 1125
rect -2703 1079 -2633 1125
rect -2587 1079 -2517 1125
rect -2471 1079 -2401 1125
rect -2355 1079 -2285 1125
rect -2239 1079 -2169 1125
rect -2123 1079 -2053 1125
rect -2007 1079 -1937 1125
rect -1891 1079 -1821 1125
rect -1775 1079 -1705 1125
rect -1659 1079 -1589 1125
rect -1543 1079 -1473 1125
rect -1427 1079 -1357 1125
rect -1311 1079 -1241 1125
rect -1195 1079 -1125 1125
rect -1079 1079 -1009 1125
rect -963 1079 -893 1125
rect -847 1079 -777 1125
rect -731 1079 -661 1125
rect -615 1079 -545 1125
rect -499 1079 -429 1125
rect -383 1079 -313 1125
rect -267 1079 -197 1125
rect -151 1079 -81 1125
rect -35 1079 35 1125
rect 81 1079 151 1125
rect 197 1079 267 1125
rect 313 1079 383 1125
rect 429 1079 499 1125
rect 545 1079 615 1125
rect 661 1079 731 1125
rect 777 1079 847 1125
rect 893 1079 963 1125
rect 1009 1079 1079 1125
rect 1125 1079 1195 1125
rect 1241 1079 1311 1125
rect 1357 1079 1427 1125
rect 1473 1079 1543 1125
rect 1589 1079 1659 1125
rect 1705 1079 1775 1125
rect 1821 1079 1891 1125
rect 1937 1079 2007 1125
rect 2053 1079 2123 1125
rect 2169 1079 2239 1125
rect 2285 1079 2355 1125
rect 2401 1079 2471 1125
rect 2517 1079 2587 1125
rect 2633 1079 2703 1125
rect 2749 1079 2819 1125
rect 2865 1079 2935 1125
rect 2981 1079 3051 1125
rect 3097 1079 3167 1125
rect 3213 1079 3283 1125
rect 3329 1079 3399 1125
rect 3445 1079 3515 1125
rect 3561 1079 3631 1125
rect 3677 1079 3747 1125
rect 3793 1079 3863 1125
rect 3909 1079 3979 1125
rect 4025 1079 4095 1125
rect 4141 1079 4211 1125
rect 4257 1079 4327 1125
rect 4373 1079 4443 1125
rect 4489 1079 4559 1125
rect 4605 1079 4675 1125
rect 4721 1079 4791 1125
rect 4837 1079 4907 1125
rect 4953 1079 5023 1125
rect 5069 1079 5139 1125
rect 5185 1079 5255 1125
rect 5301 1079 5371 1125
rect 5417 1079 5487 1125
rect 5533 1079 5603 1125
rect 5649 1079 5719 1125
rect 5765 1079 5776 1125
rect -5776 1009 5776 1079
rect -5776 963 -5765 1009
rect -5719 963 -5649 1009
rect -5603 963 -5533 1009
rect -5487 963 -5417 1009
rect -5371 963 -5301 1009
rect -5255 963 -5185 1009
rect -5139 963 -5069 1009
rect -5023 963 -4953 1009
rect -4907 963 -4837 1009
rect -4791 963 -4721 1009
rect -4675 963 -4605 1009
rect -4559 963 -4489 1009
rect -4443 963 -4373 1009
rect -4327 963 -4257 1009
rect -4211 963 -4141 1009
rect -4095 963 -4025 1009
rect -3979 963 -3909 1009
rect -3863 963 -3793 1009
rect -3747 963 -3677 1009
rect -3631 963 -3561 1009
rect -3515 963 -3445 1009
rect -3399 963 -3329 1009
rect -3283 963 -3213 1009
rect -3167 963 -3097 1009
rect -3051 963 -2981 1009
rect -2935 963 -2865 1009
rect -2819 963 -2749 1009
rect -2703 963 -2633 1009
rect -2587 963 -2517 1009
rect -2471 963 -2401 1009
rect -2355 963 -2285 1009
rect -2239 963 -2169 1009
rect -2123 963 -2053 1009
rect -2007 963 -1937 1009
rect -1891 963 -1821 1009
rect -1775 963 -1705 1009
rect -1659 963 -1589 1009
rect -1543 963 -1473 1009
rect -1427 963 -1357 1009
rect -1311 963 -1241 1009
rect -1195 963 -1125 1009
rect -1079 963 -1009 1009
rect -963 963 -893 1009
rect -847 963 -777 1009
rect -731 963 -661 1009
rect -615 963 -545 1009
rect -499 963 -429 1009
rect -383 963 -313 1009
rect -267 963 -197 1009
rect -151 963 -81 1009
rect -35 963 35 1009
rect 81 963 151 1009
rect 197 963 267 1009
rect 313 963 383 1009
rect 429 963 499 1009
rect 545 963 615 1009
rect 661 963 731 1009
rect 777 963 847 1009
rect 893 963 963 1009
rect 1009 963 1079 1009
rect 1125 963 1195 1009
rect 1241 963 1311 1009
rect 1357 963 1427 1009
rect 1473 963 1543 1009
rect 1589 963 1659 1009
rect 1705 963 1775 1009
rect 1821 963 1891 1009
rect 1937 963 2007 1009
rect 2053 963 2123 1009
rect 2169 963 2239 1009
rect 2285 963 2355 1009
rect 2401 963 2471 1009
rect 2517 963 2587 1009
rect 2633 963 2703 1009
rect 2749 963 2819 1009
rect 2865 963 2935 1009
rect 2981 963 3051 1009
rect 3097 963 3167 1009
rect 3213 963 3283 1009
rect 3329 963 3399 1009
rect 3445 963 3515 1009
rect 3561 963 3631 1009
rect 3677 963 3747 1009
rect 3793 963 3863 1009
rect 3909 963 3979 1009
rect 4025 963 4095 1009
rect 4141 963 4211 1009
rect 4257 963 4327 1009
rect 4373 963 4443 1009
rect 4489 963 4559 1009
rect 4605 963 4675 1009
rect 4721 963 4791 1009
rect 4837 963 4907 1009
rect 4953 963 5023 1009
rect 5069 963 5139 1009
rect 5185 963 5255 1009
rect 5301 963 5371 1009
rect 5417 963 5487 1009
rect 5533 963 5603 1009
rect 5649 963 5719 1009
rect 5765 963 5776 1009
rect -5776 893 5776 963
rect -5776 847 -5765 893
rect -5719 847 -5649 893
rect -5603 847 -5533 893
rect -5487 847 -5417 893
rect -5371 847 -5301 893
rect -5255 847 -5185 893
rect -5139 847 -5069 893
rect -5023 847 -4953 893
rect -4907 847 -4837 893
rect -4791 847 -4721 893
rect -4675 847 -4605 893
rect -4559 847 -4489 893
rect -4443 847 -4373 893
rect -4327 847 -4257 893
rect -4211 847 -4141 893
rect -4095 847 -4025 893
rect -3979 847 -3909 893
rect -3863 847 -3793 893
rect -3747 847 -3677 893
rect -3631 847 -3561 893
rect -3515 847 -3445 893
rect -3399 847 -3329 893
rect -3283 847 -3213 893
rect -3167 847 -3097 893
rect -3051 847 -2981 893
rect -2935 847 -2865 893
rect -2819 847 -2749 893
rect -2703 847 -2633 893
rect -2587 847 -2517 893
rect -2471 847 -2401 893
rect -2355 847 -2285 893
rect -2239 847 -2169 893
rect -2123 847 -2053 893
rect -2007 847 -1937 893
rect -1891 847 -1821 893
rect -1775 847 -1705 893
rect -1659 847 -1589 893
rect -1543 847 -1473 893
rect -1427 847 -1357 893
rect -1311 847 -1241 893
rect -1195 847 -1125 893
rect -1079 847 -1009 893
rect -963 847 -893 893
rect -847 847 -777 893
rect -731 847 -661 893
rect -615 847 -545 893
rect -499 847 -429 893
rect -383 847 -313 893
rect -267 847 -197 893
rect -151 847 -81 893
rect -35 847 35 893
rect 81 847 151 893
rect 197 847 267 893
rect 313 847 383 893
rect 429 847 499 893
rect 545 847 615 893
rect 661 847 731 893
rect 777 847 847 893
rect 893 847 963 893
rect 1009 847 1079 893
rect 1125 847 1195 893
rect 1241 847 1311 893
rect 1357 847 1427 893
rect 1473 847 1543 893
rect 1589 847 1659 893
rect 1705 847 1775 893
rect 1821 847 1891 893
rect 1937 847 2007 893
rect 2053 847 2123 893
rect 2169 847 2239 893
rect 2285 847 2355 893
rect 2401 847 2471 893
rect 2517 847 2587 893
rect 2633 847 2703 893
rect 2749 847 2819 893
rect 2865 847 2935 893
rect 2981 847 3051 893
rect 3097 847 3167 893
rect 3213 847 3283 893
rect 3329 847 3399 893
rect 3445 847 3515 893
rect 3561 847 3631 893
rect 3677 847 3747 893
rect 3793 847 3863 893
rect 3909 847 3979 893
rect 4025 847 4095 893
rect 4141 847 4211 893
rect 4257 847 4327 893
rect 4373 847 4443 893
rect 4489 847 4559 893
rect 4605 847 4675 893
rect 4721 847 4791 893
rect 4837 847 4907 893
rect 4953 847 5023 893
rect 5069 847 5139 893
rect 5185 847 5255 893
rect 5301 847 5371 893
rect 5417 847 5487 893
rect 5533 847 5603 893
rect 5649 847 5719 893
rect 5765 847 5776 893
rect -5776 777 5776 847
rect -5776 731 -5765 777
rect -5719 731 -5649 777
rect -5603 731 -5533 777
rect -5487 731 -5417 777
rect -5371 731 -5301 777
rect -5255 731 -5185 777
rect -5139 731 -5069 777
rect -5023 731 -4953 777
rect -4907 731 -4837 777
rect -4791 731 -4721 777
rect -4675 731 -4605 777
rect -4559 731 -4489 777
rect -4443 731 -4373 777
rect -4327 731 -4257 777
rect -4211 731 -4141 777
rect -4095 731 -4025 777
rect -3979 731 -3909 777
rect -3863 731 -3793 777
rect -3747 731 -3677 777
rect -3631 731 -3561 777
rect -3515 731 -3445 777
rect -3399 731 -3329 777
rect -3283 731 -3213 777
rect -3167 731 -3097 777
rect -3051 731 -2981 777
rect -2935 731 -2865 777
rect -2819 731 -2749 777
rect -2703 731 -2633 777
rect -2587 731 -2517 777
rect -2471 731 -2401 777
rect -2355 731 -2285 777
rect -2239 731 -2169 777
rect -2123 731 -2053 777
rect -2007 731 -1937 777
rect -1891 731 -1821 777
rect -1775 731 -1705 777
rect -1659 731 -1589 777
rect -1543 731 -1473 777
rect -1427 731 -1357 777
rect -1311 731 -1241 777
rect -1195 731 -1125 777
rect -1079 731 -1009 777
rect -963 731 -893 777
rect -847 731 -777 777
rect -731 731 -661 777
rect -615 731 -545 777
rect -499 731 -429 777
rect -383 731 -313 777
rect -267 731 -197 777
rect -151 731 -81 777
rect -35 731 35 777
rect 81 731 151 777
rect 197 731 267 777
rect 313 731 383 777
rect 429 731 499 777
rect 545 731 615 777
rect 661 731 731 777
rect 777 731 847 777
rect 893 731 963 777
rect 1009 731 1079 777
rect 1125 731 1195 777
rect 1241 731 1311 777
rect 1357 731 1427 777
rect 1473 731 1543 777
rect 1589 731 1659 777
rect 1705 731 1775 777
rect 1821 731 1891 777
rect 1937 731 2007 777
rect 2053 731 2123 777
rect 2169 731 2239 777
rect 2285 731 2355 777
rect 2401 731 2471 777
rect 2517 731 2587 777
rect 2633 731 2703 777
rect 2749 731 2819 777
rect 2865 731 2935 777
rect 2981 731 3051 777
rect 3097 731 3167 777
rect 3213 731 3283 777
rect 3329 731 3399 777
rect 3445 731 3515 777
rect 3561 731 3631 777
rect 3677 731 3747 777
rect 3793 731 3863 777
rect 3909 731 3979 777
rect 4025 731 4095 777
rect 4141 731 4211 777
rect 4257 731 4327 777
rect 4373 731 4443 777
rect 4489 731 4559 777
rect 4605 731 4675 777
rect 4721 731 4791 777
rect 4837 731 4907 777
rect 4953 731 5023 777
rect 5069 731 5139 777
rect 5185 731 5255 777
rect 5301 731 5371 777
rect 5417 731 5487 777
rect 5533 731 5603 777
rect 5649 731 5719 777
rect 5765 731 5776 777
rect -5776 661 5776 731
rect -5776 615 -5765 661
rect -5719 615 -5649 661
rect -5603 615 -5533 661
rect -5487 615 -5417 661
rect -5371 615 -5301 661
rect -5255 615 -5185 661
rect -5139 615 -5069 661
rect -5023 615 -4953 661
rect -4907 615 -4837 661
rect -4791 615 -4721 661
rect -4675 615 -4605 661
rect -4559 615 -4489 661
rect -4443 615 -4373 661
rect -4327 615 -4257 661
rect -4211 615 -4141 661
rect -4095 615 -4025 661
rect -3979 615 -3909 661
rect -3863 615 -3793 661
rect -3747 615 -3677 661
rect -3631 615 -3561 661
rect -3515 615 -3445 661
rect -3399 615 -3329 661
rect -3283 615 -3213 661
rect -3167 615 -3097 661
rect -3051 615 -2981 661
rect -2935 615 -2865 661
rect -2819 615 -2749 661
rect -2703 615 -2633 661
rect -2587 615 -2517 661
rect -2471 615 -2401 661
rect -2355 615 -2285 661
rect -2239 615 -2169 661
rect -2123 615 -2053 661
rect -2007 615 -1937 661
rect -1891 615 -1821 661
rect -1775 615 -1705 661
rect -1659 615 -1589 661
rect -1543 615 -1473 661
rect -1427 615 -1357 661
rect -1311 615 -1241 661
rect -1195 615 -1125 661
rect -1079 615 -1009 661
rect -963 615 -893 661
rect -847 615 -777 661
rect -731 615 -661 661
rect -615 615 -545 661
rect -499 615 -429 661
rect -383 615 -313 661
rect -267 615 -197 661
rect -151 615 -81 661
rect -35 615 35 661
rect 81 615 151 661
rect 197 615 267 661
rect 313 615 383 661
rect 429 615 499 661
rect 545 615 615 661
rect 661 615 731 661
rect 777 615 847 661
rect 893 615 963 661
rect 1009 615 1079 661
rect 1125 615 1195 661
rect 1241 615 1311 661
rect 1357 615 1427 661
rect 1473 615 1543 661
rect 1589 615 1659 661
rect 1705 615 1775 661
rect 1821 615 1891 661
rect 1937 615 2007 661
rect 2053 615 2123 661
rect 2169 615 2239 661
rect 2285 615 2355 661
rect 2401 615 2471 661
rect 2517 615 2587 661
rect 2633 615 2703 661
rect 2749 615 2819 661
rect 2865 615 2935 661
rect 2981 615 3051 661
rect 3097 615 3167 661
rect 3213 615 3283 661
rect 3329 615 3399 661
rect 3445 615 3515 661
rect 3561 615 3631 661
rect 3677 615 3747 661
rect 3793 615 3863 661
rect 3909 615 3979 661
rect 4025 615 4095 661
rect 4141 615 4211 661
rect 4257 615 4327 661
rect 4373 615 4443 661
rect 4489 615 4559 661
rect 4605 615 4675 661
rect 4721 615 4791 661
rect 4837 615 4907 661
rect 4953 615 5023 661
rect 5069 615 5139 661
rect 5185 615 5255 661
rect 5301 615 5371 661
rect 5417 615 5487 661
rect 5533 615 5603 661
rect 5649 615 5719 661
rect 5765 615 5776 661
rect -5776 545 5776 615
rect -5776 499 -5765 545
rect -5719 499 -5649 545
rect -5603 499 -5533 545
rect -5487 499 -5417 545
rect -5371 499 -5301 545
rect -5255 499 -5185 545
rect -5139 499 -5069 545
rect -5023 499 -4953 545
rect -4907 499 -4837 545
rect -4791 499 -4721 545
rect -4675 499 -4605 545
rect -4559 499 -4489 545
rect -4443 499 -4373 545
rect -4327 499 -4257 545
rect -4211 499 -4141 545
rect -4095 499 -4025 545
rect -3979 499 -3909 545
rect -3863 499 -3793 545
rect -3747 499 -3677 545
rect -3631 499 -3561 545
rect -3515 499 -3445 545
rect -3399 499 -3329 545
rect -3283 499 -3213 545
rect -3167 499 -3097 545
rect -3051 499 -2981 545
rect -2935 499 -2865 545
rect -2819 499 -2749 545
rect -2703 499 -2633 545
rect -2587 499 -2517 545
rect -2471 499 -2401 545
rect -2355 499 -2285 545
rect -2239 499 -2169 545
rect -2123 499 -2053 545
rect -2007 499 -1937 545
rect -1891 499 -1821 545
rect -1775 499 -1705 545
rect -1659 499 -1589 545
rect -1543 499 -1473 545
rect -1427 499 -1357 545
rect -1311 499 -1241 545
rect -1195 499 -1125 545
rect -1079 499 -1009 545
rect -963 499 -893 545
rect -847 499 -777 545
rect -731 499 -661 545
rect -615 499 -545 545
rect -499 499 -429 545
rect -383 499 -313 545
rect -267 499 -197 545
rect -151 499 -81 545
rect -35 499 35 545
rect 81 499 151 545
rect 197 499 267 545
rect 313 499 383 545
rect 429 499 499 545
rect 545 499 615 545
rect 661 499 731 545
rect 777 499 847 545
rect 893 499 963 545
rect 1009 499 1079 545
rect 1125 499 1195 545
rect 1241 499 1311 545
rect 1357 499 1427 545
rect 1473 499 1543 545
rect 1589 499 1659 545
rect 1705 499 1775 545
rect 1821 499 1891 545
rect 1937 499 2007 545
rect 2053 499 2123 545
rect 2169 499 2239 545
rect 2285 499 2355 545
rect 2401 499 2471 545
rect 2517 499 2587 545
rect 2633 499 2703 545
rect 2749 499 2819 545
rect 2865 499 2935 545
rect 2981 499 3051 545
rect 3097 499 3167 545
rect 3213 499 3283 545
rect 3329 499 3399 545
rect 3445 499 3515 545
rect 3561 499 3631 545
rect 3677 499 3747 545
rect 3793 499 3863 545
rect 3909 499 3979 545
rect 4025 499 4095 545
rect 4141 499 4211 545
rect 4257 499 4327 545
rect 4373 499 4443 545
rect 4489 499 4559 545
rect 4605 499 4675 545
rect 4721 499 4791 545
rect 4837 499 4907 545
rect 4953 499 5023 545
rect 5069 499 5139 545
rect 5185 499 5255 545
rect 5301 499 5371 545
rect 5417 499 5487 545
rect 5533 499 5603 545
rect 5649 499 5719 545
rect 5765 499 5776 545
rect -5776 429 5776 499
rect -5776 383 -5765 429
rect -5719 383 -5649 429
rect -5603 383 -5533 429
rect -5487 383 -5417 429
rect -5371 383 -5301 429
rect -5255 383 -5185 429
rect -5139 383 -5069 429
rect -5023 383 -4953 429
rect -4907 383 -4837 429
rect -4791 383 -4721 429
rect -4675 383 -4605 429
rect -4559 383 -4489 429
rect -4443 383 -4373 429
rect -4327 383 -4257 429
rect -4211 383 -4141 429
rect -4095 383 -4025 429
rect -3979 383 -3909 429
rect -3863 383 -3793 429
rect -3747 383 -3677 429
rect -3631 383 -3561 429
rect -3515 383 -3445 429
rect -3399 383 -3329 429
rect -3283 383 -3213 429
rect -3167 383 -3097 429
rect -3051 383 -2981 429
rect -2935 383 -2865 429
rect -2819 383 -2749 429
rect -2703 383 -2633 429
rect -2587 383 -2517 429
rect -2471 383 -2401 429
rect -2355 383 -2285 429
rect -2239 383 -2169 429
rect -2123 383 -2053 429
rect -2007 383 -1937 429
rect -1891 383 -1821 429
rect -1775 383 -1705 429
rect -1659 383 -1589 429
rect -1543 383 -1473 429
rect -1427 383 -1357 429
rect -1311 383 -1241 429
rect -1195 383 -1125 429
rect -1079 383 -1009 429
rect -963 383 -893 429
rect -847 383 -777 429
rect -731 383 -661 429
rect -615 383 -545 429
rect -499 383 -429 429
rect -383 383 -313 429
rect -267 383 -197 429
rect -151 383 -81 429
rect -35 383 35 429
rect 81 383 151 429
rect 197 383 267 429
rect 313 383 383 429
rect 429 383 499 429
rect 545 383 615 429
rect 661 383 731 429
rect 777 383 847 429
rect 893 383 963 429
rect 1009 383 1079 429
rect 1125 383 1195 429
rect 1241 383 1311 429
rect 1357 383 1427 429
rect 1473 383 1543 429
rect 1589 383 1659 429
rect 1705 383 1775 429
rect 1821 383 1891 429
rect 1937 383 2007 429
rect 2053 383 2123 429
rect 2169 383 2239 429
rect 2285 383 2355 429
rect 2401 383 2471 429
rect 2517 383 2587 429
rect 2633 383 2703 429
rect 2749 383 2819 429
rect 2865 383 2935 429
rect 2981 383 3051 429
rect 3097 383 3167 429
rect 3213 383 3283 429
rect 3329 383 3399 429
rect 3445 383 3515 429
rect 3561 383 3631 429
rect 3677 383 3747 429
rect 3793 383 3863 429
rect 3909 383 3979 429
rect 4025 383 4095 429
rect 4141 383 4211 429
rect 4257 383 4327 429
rect 4373 383 4443 429
rect 4489 383 4559 429
rect 4605 383 4675 429
rect 4721 383 4791 429
rect 4837 383 4907 429
rect 4953 383 5023 429
rect 5069 383 5139 429
rect 5185 383 5255 429
rect 5301 383 5371 429
rect 5417 383 5487 429
rect 5533 383 5603 429
rect 5649 383 5719 429
rect 5765 383 5776 429
rect -5776 313 5776 383
rect -5776 267 -5765 313
rect -5719 267 -5649 313
rect -5603 267 -5533 313
rect -5487 267 -5417 313
rect -5371 267 -5301 313
rect -5255 267 -5185 313
rect -5139 267 -5069 313
rect -5023 267 -4953 313
rect -4907 267 -4837 313
rect -4791 267 -4721 313
rect -4675 267 -4605 313
rect -4559 267 -4489 313
rect -4443 267 -4373 313
rect -4327 267 -4257 313
rect -4211 267 -4141 313
rect -4095 267 -4025 313
rect -3979 267 -3909 313
rect -3863 267 -3793 313
rect -3747 267 -3677 313
rect -3631 267 -3561 313
rect -3515 267 -3445 313
rect -3399 267 -3329 313
rect -3283 267 -3213 313
rect -3167 267 -3097 313
rect -3051 267 -2981 313
rect -2935 267 -2865 313
rect -2819 267 -2749 313
rect -2703 267 -2633 313
rect -2587 267 -2517 313
rect -2471 267 -2401 313
rect -2355 267 -2285 313
rect -2239 267 -2169 313
rect -2123 267 -2053 313
rect -2007 267 -1937 313
rect -1891 267 -1821 313
rect -1775 267 -1705 313
rect -1659 267 -1589 313
rect -1543 267 -1473 313
rect -1427 267 -1357 313
rect -1311 267 -1241 313
rect -1195 267 -1125 313
rect -1079 267 -1009 313
rect -963 267 -893 313
rect -847 267 -777 313
rect -731 267 -661 313
rect -615 267 -545 313
rect -499 267 -429 313
rect -383 267 -313 313
rect -267 267 -197 313
rect -151 267 -81 313
rect -35 267 35 313
rect 81 267 151 313
rect 197 267 267 313
rect 313 267 383 313
rect 429 267 499 313
rect 545 267 615 313
rect 661 267 731 313
rect 777 267 847 313
rect 893 267 963 313
rect 1009 267 1079 313
rect 1125 267 1195 313
rect 1241 267 1311 313
rect 1357 267 1427 313
rect 1473 267 1543 313
rect 1589 267 1659 313
rect 1705 267 1775 313
rect 1821 267 1891 313
rect 1937 267 2007 313
rect 2053 267 2123 313
rect 2169 267 2239 313
rect 2285 267 2355 313
rect 2401 267 2471 313
rect 2517 267 2587 313
rect 2633 267 2703 313
rect 2749 267 2819 313
rect 2865 267 2935 313
rect 2981 267 3051 313
rect 3097 267 3167 313
rect 3213 267 3283 313
rect 3329 267 3399 313
rect 3445 267 3515 313
rect 3561 267 3631 313
rect 3677 267 3747 313
rect 3793 267 3863 313
rect 3909 267 3979 313
rect 4025 267 4095 313
rect 4141 267 4211 313
rect 4257 267 4327 313
rect 4373 267 4443 313
rect 4489 267 4559 313
rect 4605 267 4675 313
rect 4721 267 4791 313
rect 4837 267 4907 313
rect 4953 267 5023 313
rect 5069 267 5139 313
rect 5185 267 5255 313
rect 5301 267 5371 313
rect 5417 267 5487 313
rect 5533 267 5603 313
rect 5649 267 5719 313
rect 5765 267 5776 313
rect -5776 197 5776 267
rect -5776 151 -5765 197
rect -5719 151 -5649 197
rect -5603 151 -5533 197
rect -5487 151 -5417 197
rect -5371 151 -5301 197
rect -5255 151 -5185 197
rect -5139 151 -5069 197
rect -5023 151 -4953 197
rect -4907 151 -4837 197
rect -4791 151 -4721 197
rect -4675 151 -4605 197
rect -4559 151 -4489 197
rect -4443 151 -4373 197
rect -4327 151 -4257 197
rect -4211 151 -4141 197
rect -4095 151 -4025 197
rect -3979 151 -3909 197
rect -3863 151 -3793 197
rect -3747 151 -3677 197
rect -3631 151 -3561 197
rect -3515 151 -3445 197
rect -3399 151 -3329 197
rect -3283 151 -3213 197
rect -3167 151 -3097 197
rect -3051 151 -2981 197
rect -2935 151 -2865 197
rect -2819 151 -2749 197
rect -2703 151 -2633 197
rect -2587 151 -2517 197
rect -2471 151 -2401 197
rect -2355 151 -2285 197
rect -2239 151 -2169 197
rect -2123 151 -2053 197
rect -2007 151 -1937 197
rect -1891 151 -1821 197
rect -1775 151 -1705 197
rect -1659 151 -1589 197
rect -1543 151 -1473 197
rect -1427 151 -1357 197
rect -1311 151 -1241 197
rect -1195 151 -1125 197
rect -1079 151 -1009 197
rect -963 151 -893 197
rect -847 151 -777 197
rect -731 151 -661 197
rect -615 151 -545 197
rect -499 151 -429 197
rect -383 151 -313 197
rect -267 151 -197 197
rect -151 151 -81 197
rect -35 151 35 197
rect 81 151 151 197
rect 197 151 267 197
rect 313 151 383 197
rect 429 151 499 197
rect 545 151 615 197
rect 661 151 731 197
rect 777 151 847 197
rect 893 151 963 197
rect 1009 151 1079 197
rect 1125 151 1195 197
rect 1241 151 1311 197
rect 1357 151 1427 197
rect 1473 151 1543 197
rect 1589 151 1659 197
rect 1705 151 1775 197
rect 1821 151 1891 197
rect 1937 151 2007 197
rect 2053 151 2123 197
rect 2169 151 2239 197
rect 2285 151 2355 197
rect 2401 151 2471 197
rect 2517 151 2587 197
rect 2633 151 2703 197
rect 2749 151 2819 197
rect 2865 151 2935 197
rect 2981 151 3051 197
rect 3097 151 3167 197
rect 3213 151 3283 197
rect 3329 151 3399 197
rect 3445 151 3515 197
rect 3561 151 3631 197
rect 3677 151 3747 197
rect 3793 151 3863 197
rect 3909 151 3979 197
rect 4025 151 4095 197
rect 4141 151 4211 197
rect 4257 151 4327 197
rect 4373 151 4443 197
rect 4489 151 4559 197
rect 4605 151 4675 197
rect 4721 151 4791 197
rect 4837 151 4907 197
rect 4953 151 5023 197
rect 5069 151 5139 197
rect 5185 151 5255 197
rect 5301 151 5371 197
rect 5417 151 5487 197
rect 5533 151 5603 197
rect 5649 151 5719 197
rect 5765 151 5776 197
rect -5776 81 5776 151
rect -5776 35 -5765 81
rect -5719 35 -5649 81
rect -5603 35 -5533 81
rect -5487 35 -5417 81
rect -5371 35 -5301 81
rect -5255 35 -5185 81
rect -5139 35 -5069 81
rect -5023 35 -4953 81
rect -4907 35 -4837 81
rect -4791 35 -4721 81
rect -4675 35 -4605 81
rect -4559 35 -4489 81
rect -4443 35 -4373 81
rect -4327 35 -4257 81
rect -4211 35 -4141 81
rect -4095 35 -4025 81
rect -3979 35 -3909 81
rect -3863 35 -3793 81
rect -3747 35 -3677 81
rect -3631 35 -3561 81
rect -3515 35 -3445 81
rect -3399 35 -3329 81
rect -3283 35 -3213 81
rect -3167 35 -3097 81
rect -3051 35 -2981 81
rect -2935 35 -2865 81
rect -2819 35 -2749 81
rect -2703 35 -2633 81
rect -2587 35 -2517 81
rect -2471 35 -2401 81
rect -2355 35 -2285 81
rect -2239 35 -2169 81
rect -2123 35 -2053 81
rect -2007 35 -1937 81
rect -1891 35 -1821 81
rect -1775 35 -1705 81
rect -1659 35 -1589 81
rect -1543 35 -1473 81
rect -1427 35 -1357 81
rect -1311 35 -1241 81
rect -1195 35 -1125 81
rect -1079 35 -1009 81
rect -963 35 -893 81
rect -847 35 -777 81
rect -731 35 -661 81
rect -615 35 -545 81
rect -499 35 -429 81
rect -383 35 -313 81
rect -267 35 -197 81
rect -151 35 -81 81
rect -35 35 35 81
rect 81 35 151 81
rect 197 35 267 81
rect 313 35 383 81
rect 429 35 499 81
rect 545 35 615 81
rect 661 35 731 81
rect 777 35 847 81
rect 893 35 963 81
rect 1009 35 1079 81
rect 1125 35 1195 81
rect 1241 35 1311 81
rect 1357 35 1427 81
rect 1473 35 1543 81
rect 1589 35 1659 81
rect 1705 35 1775 81
rect 1821 35 1891 81
rect 1937 35 2007 81
rect 2053 35 2123 81
rect 2169 35 2239 81
rect 2285 35 2355 81
rect 2401 35 2471 81
rect 2517 35 2587 81
rect 2633 35 2703 81
rect 2749 35 2819 81
rect 2865 35 2935 81
rect 2981 35 3051 81
rect 3097 35 3167 81
rect 3213 35 3283 81
rect 3329 35 3399 81
rect 3445 35 3515 81
rect 3561 35 3631 81
rect 3677 35 3747 81
rect 3793 35 3863 81
rect 3909 35 3979 81
rect 4025 35 4095 81
rect 4141 35 4211 81
rect 4257 35 4327 81
rect 4373 35 4443 81
rect 4489 35 4559 81
rect 4605 35 4675 81
rect 4721 35 4791 81
rect 4837 35 4907 81
rect 4953 35 5023 81
rect 5069 35 5139 81
rect 5185 35 5255 81
rect 5301 35 5371 81
rect 5417 35 5487 81
rect 5533 35 5603 81
rect 5649 35 5719 81
rect 5765 35 5776 81
rect -5776 -35 5776 35
rect -5776 -81 -5765 -35
rect -5719 -81 -5649 -35
rect -5603 -81 -5533 -35
rect -5487 -81 -5417 -35
rect -5371 -81 -5301 -35
rect -5255 -81 -5185 -35
rect -5139 -81 -5069 -35
rect -5023 -81 -4953 -35
rect -4907 -81 -4837 -35
rect -4791 -81 -4721 -35
rect -4675 -81 -4605 -35
rect -4559 -81 -4489 -35
rect -4443 -81 -4373 -35
rect -4327 -81 -4257 -35
rect -4211 -81 -4141 -35
rect -4095 -81 -4025 -35
rect -3979 -81 -3909 -35
rect -3863 -81 -3793 -35
rect -3747 -81 -3677 -35
rect -3631 -81 -3561 -35
rect -3515 -81 -3445 -35
rect -3399 -81 -3329 -35
rect -3283 -81 -3213 -35
rect -3167 -81 -3097 -35
rect -3051 -81 -2981 -35
rect -2935 -81 -2865 -35
rect -2819 -81 -2749 -35
rect -2703 -81 -2633 -35
rect -2587 -81 -2517 -35
rect -2471 -81 -2401 -35
rect -2355 -81 -2285 -35
rect -2239 -81 -2169 -35
rect -2123 -81 -2053 -35
rect -2007 -81 -1937 -35
rect -1891 -81 -1821 -35
rect -1775 -81 -1705 -35
rect -1659 -81 -1589 -35
rect -1543 -81 -1473 -35
rect -1427 -81 -1357 -35
rect -1311 -81 -1241 -35
rect -1195 -81 -1125 -35
rect -1079 -81 -1009 -35
rect -963 -81 -893 -35
rect -847 -81 -777 -35
rect -731 -81 -661 -35
rect -615 -81 -545 -35
rect -499 -81 -429 -35
rect -383 -81 -313 -35
rect -267 -81 -197 -35
rect -151 -81 -81 -35
rect -35 -81 35 -35
rect 81 -81 151 -35
rect 197 -81 267 -35
rect 313 -81 383 -35
rect 429 -81 499 -35
rect 545 -81 615 -35
rect 661 -81 731 -35
rect 777 -81 847 -35
rect 893 -81 963 -35
rect 1009 -81 1079 -35
rect 1125 -81 1195 -35
rect 1241 -81 1311 -35
rect 1357 -81 1427 -35
rect 1473 -81 1543 -35
rect 1589 -81 1659 -35
rect 1705 -81 1775 -35
rect 1821 -81 1891 -35
rect 1937 -81 2007 -35
rect 2053 -81 2123 -35
rect 2169 -81 2239 -35
rect 2285 -81 2355 -35
rect 2401 -81 2471 -35
rect 2517 -81 2587 -35
rect 2633 -81 2703 -35
rect 2749 -81 2819 -35
rect 2865 -81 2935 -35
rect 2981 -81 3051 -35
rect 3097 -81 3167 -35
rect 3213 -81 3283 -35
rect 3329 -81 3399 -35
rect 3445 -81 3515 -35
rect 3561 -81 3631 -35
rect 3677 -81 3747 -35
rect 3793 -81 3863 -35
rect 3909 -81 3979 -35
rect 4025 -81 4095 -35
rect 4141 -81 4211 -35
rect 4257 -81 4327 -35
rect 4373 -81 4443 -35
rect 4489 -81 4559 -35
rect 4605 -81 4675 -35
rect 4721 -81 4791 -35
rect 4837 -81 4907 -35
rect 4953 -81 5023 -35
rect 5069 -81 5139 -35
rect 5185 -81 5255 -35
rect 5301 -81 5371 -35
rect 5417 -81 5487 -35
rect 5533 -81 5603 -35
rect 5649 -81 5719 -35
rect 5765 -81 5776 -35
rect -5776 -151 5776 -81
rect -5776 -197 -5765 -151
rect -5719 -197 -5649 -151
rect -5603 -197 -5533 -151
rect -5487 -197 -5417 -151
rect -5371 -197 -5301 -151
rect -5255 -197 -5185 -151
rect -5139 -197 -5069 -151
rect -5023 -197 -4953 -151
rect -4907 -197 -4837 -151
rect -4791 -197 -4721 -151
rect -4675 -197 -4605 -151
rect -4559 -197 -4489 -151
rect -4443 -197 -4373 -151
rect -4327 -197 -4257 -151
rect -4211 -197 -4141 -151
rect -4095 -197 -4025 -151
rect -3979 -197 -3909 -151
rect -3863 -197 -3793 -151
rect -3747 -197 -3677 -151
rect -3631 -197 -3561 -151
rect -3515 -197 -3445 -151
rect -3399 -197 -3329 -151
rect -3283 -197 -3213 -151
rect -3167 -197 -3097 -151
rect -3051 -197 -2981 -151
rect -2935 -197 -2865 -151
rect -2819 -197 -2749 -151
rect -2703 -197 -2633 -151
rect -2587 -197 -2517 -151
rect -2471 -197 -2401 -151
rect -2355 -197 -2285 -151
rect -2239 -197 -2169 -151
rect -2123 -197 -2053 -151
rect -2007 -197 -1937 -151
rect -1891 -197 -1821 -151
rect -1775 -197 -1705 -151
rect -1659 -197 -1589 -151
rect -1543 -197 -1473 -151
rect -1427 -197 -1357 -151
rect -1311 -197 -1241 -151
rect -1195 -197 -1125 -151
rect -1079 -197 -1009 -151
rect -963 -197 -893 -151
rect -847 -197 -777 -151
rect -731 -197 -661 -151
rect -615 -197 -545 -151
rect -499 -197 -429 -151
rect -383 -197 -313 -151
rect -267 -197 -197 -151
rect -151 -197 -81 -151
rect -35 -197 35 -151
rect 81 -197 151 -151
rect 197 -197 267 -151
rect 313 -197 383 -151
rect 429 -197 499 -151
rect 545 -197 615 -151
rect 661 -197 731 -151
rect 777 -197 847 -151
rect 893 -197 963 -151
rect 1009 -197 1079 -151
rect 1125 -197 1195 -151
rect 1241 -197 1311 -151
rect 1357 -197 1427 -151
rect 1473 -197 1543 -151
rect 1589 -197 1659 -151
rect 1705 -197 1775 -151
rect 1821 -197 1891 -151
rect 1937 -197 2007 -151
rect 2053 -197 2123 -151
rect 2169 -197 2239 -151
rect 2285 -197 2355 -151
rect 2401 -197 2471 -151
rect 2517 -197 2587 -151
rect 2633 -197 2703 -151
rect 2749 -197 2819 -151
rect 2865 -197 2935 -151
rect 2981 -197 3051 -151
rect 3097 -197 3167 -151
rect 3213 -197 3283 -151
rect 3329 -197 3399 -151
rect 3445 -197 3515 -151
rect 3561 -197 3631 -151
rect 3677 -197 3747 -151
rect 3793 -197 3863 -151
rect 3909 -197 3979 -151
rect 4025 -197 4095 -151
rect 4141 -197 4211 -151
rect 4257 -197 4327 -151
rect 4373 -197 4443 -151
rect 4489 -197 4559 -151
rect 4605 -197 4675 -151
rect 4721 -197 4791 -151
rect 4837 -197 4907 -151
rect 4953 -197 5023 -151
rect 5069 -197 5139 -151
rect 5185 -197 5255 -151
rect 5301 -197 5371 -151
rect 5417 -197 5487 -151
rect 5533 -197 5603 -151
rect 5649 -197 5719 -151
rect 5765 -197 5776 -151
rect -5776 -267 5776 -197
rect -5776 -313 -5765 -267
rect -5719 -313 -5649 -267
rect -5603 -313 -5533 -267
rect -5487 -313 -5417 -267
rect -5371 -313 -5301 -267
rect -5255 -313 -5185 -267
rect -5139 -313 -5069 -267
rect -5023 -313 -4953 -267
rect -4907 -313 -4837 -267
rect -4791 -313 -4721 -267
rect -4675 -313 -4605 -267
rect -4559 -313 -4489 -267
rect -4443 -313 -4373 -267
rect -4327 -313 -4257 -267
rect -4211 -313 -4141 -267
rect -4095 -313 -4025 -267
rect -3979 -313 -3909 -267
rect -3863 -313 -3793 -267
rect -3747 -313 -3677 -267
rect -3631 -313 -3561 -267
rect -3515 -313 -3445 -267
rect -3399 -313 -3329 -267
rect -3283 -313 -3213 -267
rect -3167 -313 -3097 -267
rect -3051 -313 -2981 -267
rect -2935 -313 -2865 -267
rect -2819 -313 -2749 -267
rect -2703 -313 -2633 -267
rect -2587 -313 -2517 -267
rect -2471 -313 -2401 -267
rect -2355 -313 -2285 -267
rect -2239 -313 -2169 -267
rect -2123 -313 -2053 -267
rect -2007 -313 -1937 -267
rect -1891 -313 -1821 -267
rect -1775 -313 -1705 -267
rect -1659 -313 -1589 -267
rect -1543 -313 -1473 -267
rect -1427 -313 -1357 -267
rect -1311 -313 -1241 -267
rect -1195 -313 -1125 -267
rect -1079 -313 -1009 -267
rect -963 -313 -893 -267
rect -847 -313 -777 -267
rect -731 -313 -661 -267
rect -615 -313 -545 -267
rect -499 -313 -429 -267
rect -383 -313 -313 -267
rect -267 -313 -197 -267
rect -151 -313 -81 -267
rect -35 -313 35 -267
rect 81 -313 151 -267
rect 197 -313 267 -267
rect 313 -313 383 -267
rect 429 -313 499 -267
rect 545 -313 615 -267
rect 661 -313 731 -267
rect 777 -313 847 -267
rect 893 -313 963 -267
rect 1009 -313 1079 -267
rect 1125 -313 1195 -267
rect 1241 -313 1311 -267
rect 1357 -313 1427 -267
rect 1473 -313 1543 -267
rect 1589 -313 1659 -267
rect 1705 -313 1775 -267
rect 1821 -313 1891 -267
rect 1937 -313 2007 -267
rect 2053 -313 2123 -267
rect 2169 -313 2239 -267
rect 2285 -313 2355 -267
rect 2401 -313 2471 -267
rect 2517 -313 2587 -267
rect 2633 -313 2703 -267
rect 2749 -313 2819 -267
rect 2865 -313 2935 -267
rect 2981 -313 3051 -267
rect 3097 -313 3167 -267
rect 3213 -313 3283 -267
rect 3329 -313 3399 -267
rect 3445 -313 3515 -267
rect 3561 -313 3631 -267
rect 3677 -313 3747 -267
rect 3793 -313 3863 -267
rect 3909 -313 3979 -267
rect 4025 -313 4095 -267
rect 4141 -313 4211 -267
rect 4257 -313 4327 -267
rect 4373 -313 4443 -267
rect 4489 -313 4559 -267
rect 4605 -313 4675 -267
rect 4721 -313 4791 -267
rect 4837 -313 4907 -267
rect 4953 -313 5023 -267
rect 5069 -313 5139 -267
rect 5185 -313 5255 -267
rect 5301 -313 5371 -267
rect 5417 -313 5487 -267
rect 5533 -313 5603 -267
rect 5649 -313 5719 -267
rect 5765 -313 5776 -267
rect -5776 -383 5776 -313
rect -5776 -429 -5765 -383
rect -5719 -429 -5649 -383
rect -5603 -429 -5533 -383
rect -5487 -429 -5417 -383
rect -5371 -429 -5301 -383
rect -5255 -429 -5185 -383
rect -5139 -429 -5069 -383
rect -5023 -429 -4953 -383
rect -4907 -429 -4837 -383
rect -4791 -429 -4721 -383
rect -4675 -429 -4605 -383
rect -4559 -429 -4489 -383
rect -4443 -429 -4373 -383
rect -4327 -429 -4257 -383
rect -4211 -429 -4141 -383
rect -4095 -429 -4025 -383
rect -3979 -429 -3909 -383
rect -3863 -429 -3793 -383
rect -3747 -429 -3677 -383
rect -3631 -429 -3561 -383
rect -3515 -429 -3445 -383
rect -3399 -429 -3329 -383
rect -3283 -429 -3213 -383
rect -3167 -429 -3097 -383
rect -3051 -429 -2981 -383
rect -2935 -429 -2865 -383
rect -2819 -429 -2749 -383
rect -2703 -429 -2633 -383
rect -2587 -429 -2517 -383
rect -2471 -429 -2401 -383
rect -2355 -429 -2285 -383
rect -2239 -429 -2169 -383
rect -2123 -429 -2053 -383
rect -2007 -429 -1937 -383
rect -1891 -429 -1821 -383
rect -1775 -429 -1705 -383
rect -1659 -429 -1589 -383
rect -1543 -429 -1473 -383
rect -1427 -429 -1357 -383
rect -1311 -429 -1241 -383
rect -1195 -429 -1125 -383
rect -1079 -429 -1009 -383
rect -963 -429 -893 -383
rect -847 -429 -777 -383
rect -731 -429 -661 -383
rect -615 -429 -545 -383
rect -499 -429 -429 -383
rect -383 -429 -313 -383
rect -267 -429 -197 -383
rect -151 -429 -81 -383
rect -35 -429 35 -383
rect 81 -429 151 -383
rect 197 -429 267 -383
rect 313 -429 383 -383
rect 429 -429 499 -383
rect 545 -429 615 -383
rect 661 -429 731 -383
rect 777 -429 847 -383
rect 893 -429 963 -383
rect 1009 -429 1079 -383
rect 1125 -429 1195 -383
rect 1241 -429 1311 -383
rect 1357 -429 1427 -383
rect 1473 -429 1543 -383
rect 1589 -429 1659 -383
rect 1705 -429 1775 -383
rect 1821 -429 1891 -383
rect 1937 -429 2007 -383
rect 2053 -429 2123 -383
rect 2169 -429 2239 -383
rect 2285 -429 2355 -383
rect 2401 -429 2471 -383
rect 2517 -429 2587 -383
rect 2633 -429 2703 -383
rect 2749 -429 2819 -383
rect 2865 -429 2935 -383
rect 2981 -429 3051 -383
rect 3097 -429 3167 -383
rect 3213 -429 3283 -383
rect 3329 -429 3399 -383
rect 3445 -429 3515 -383
rect 3561 -429 3631 -383
rect 3677 -429 3747 -383
rect 3793 -429 3863 -383
rect 3909 -429 3979 -383
rect 4025 -429 4095 -383
rect 4141 -429 4211 -383
rect 4257 -429 4327 -383
rect 4373 -429 4443 -383
rect 4489 -429 4559 -383
rect 4605 -429 4675 -383
rect 4721 -429 4791 -383
rect 4837 -429 4907 -383
rect 4953 -429 5023 -383
rect 5069 -429 5139 -383
rect 5185 -429 5255 -383
rect 5301 -429 5371 -383
rect 5417 -429 5487 -383
rect 5533 -429 5603 -383
rect 5649 -429 5719 -383
rect 5765 -429 5776 -383
rect -5776 -499 5776 -429
rect -5776 -545 -5765 -499
rect -5719 -545 -5649 -499
rect -5603 -545 -5533 -499
rect -5487 -545 -5417 -499
rect -5371 -545 -5301 -499
rect -5255 -545 -5185 -499
rect -5139 -545 -5069 -499
rect -5023 -545 -4953 -499
rect -4907 -545 -4837 -499
rect -4791 -545 -4721 -499
rect -4675 -545 -4605 -499
rect -4559 -545 -4489 -499
rect -4443 -545 -4373 -499
rect -4327 -545 -4257 -499
rect -4211 -545 -4141 -499
rect -4095 -545 -4025 -499
rect -3979 -545 -3909 -499
rect -3863 -545 -3793 -499
rect -3747 -545 -3677 -499
rect -3631 -545 -3561 -499
rect -3515 -545 -3445 -499
rect -3399 -545 -3329 -499
rect -3283 -545 -3213 -499
rect -3167 -545 -3097 -499
rect -3051 -545 -2981 -499
rect -2935 -545 -2865 -499
rect -2819 -545 -2749 -499
rect -2703 -545 -2633 -499
rect -2587 -545 -2517 -499
rect -2471 -545 -2401 -499
rect -2355 -545 -2285 -499
rect -2239 -545 -2169 -499
rect -2123 -545 -2053 -499
rect -2007 -545 -1937 -499
rect -1891 -545 -1821 -499
rect -1775 -545 -1705 -499
rect -1659 -545 -1589 -499
rect -1543 -545 -1473 -499
rect -1427 -545 -1357 -499
rect -1311 -545 -1241 -499
rect -1195 -545 -1125 -499
rect -1079 -545 -1009 -499
rect -963 -545 -893 -499
rect -847 -545 -777 -499
rect -731 -545 -661 -499
rect -615 -545 -545 -499
rect -499 -545 -429 -499
rect -383 -545 -313 -499
rect -267 -545 -197 -499
rect -151 -545 -81 -499
rect -35 -545 35 -499
rect 81 -545 151 -499
rect 197 -545 267 -499
rect 313 -545 383 -499
rect 429 -545 499 -499
rect 545 -545 615 -499
rect 661 -545 731 -499
rect 777 -545 847 -499
rect 893 -545 963 -499
rect 1009 -545 1079 -499
rect 1125 -545 1195 -499
rect 1241 -545 1311 -499
rect 1357 -545 1427 -499
rect 1473 -545 1543 -499
rect 1589 -545 1659 -499
rect 1705 -545 1775 -499
rect 1821 -545 1891 -499
rect 1937 -545 2007 -499
rect 2053 -545 2123 -499
rect 2169 -545 2239 -499
rect 2285 -545 2355 -499
rect 2401 -545 2471 -499
rect 2517 -545 2587 -499
rect 2633 -545 2703 -499
rect 2749 -545 2819 -499
rect 2865 -545 2935 -499
rect 2981 -545 3051 -499
rect 3097 -545 3167 -499
rect 3213 -545 3283 -499
rect 3329 -545 3399 -499
rect 3445 -545 3515 -499
rect 3561 -545 3631 -499
rect 3677 -545 3747 -499
rect 3793 -545 3863 -499
rect 3909 -545 3979 -499
rect 4025 -545 4095 -499
rect 4141 -545 4211 -499
rect 4257 -545 4327 -499
rect 4373 -545 4443 -499
rect 4489 -545 4559 -499
rect 4605 -545 4675 -499
rect 4721 -545 4791 -499
rect 4837 -545 4907 -499
rect 4953 -545 5023 -499
rect 5069 -545 5139 -499
rect 5185 -545 5255 -499
rect 5301 -545 5371 -499
rect 5417 -545 5487 -499
rect 5533 -545 5603 -499
rect 5649 -545 5719 -499
rect 5765 -545 5776 -499
rect -5776 -615 5776 -545
rect -5776 -661 -5765 -615
rect -5719 -661 -5649 -615
rect -5603 -661 -5533 -615
rect -5487 -661 -5417 -615
rect -5371 -661 -5301 -615
rect -5255 -661 -5185 -615
rect -5139 -661 -5069 -615
rect -5023 -661 -4953 -615
rect -4907 -661 -4837 -615
rect -4791 -661 -4721 -615
rect -4675 -661 -4605 -615
rect -4559 -661 -4489 -615
rect -4443 -661 -4373 -615
rect -4327 -661 -4257 -615
rect -4211 -661 -4141 -615
rect -4095 -661 -4025 -615
rect -3979 -661 -3909 -615
rect -3863 -661 -3793 -615
rect -3747 -661 -3677 -615
rect -3631 -661 -3561 -615
rect -3515 -661 -3445 -615
rect -3399 -661 -3329 -615
rect -3283 -661 -3213 -615
rect -3167 -661 -3097 -615
rect -3051 -661 -2981 -615
rect -2935 -661 -2865 -615
rect -2819 -661 -2749 -615
rect -2703 -661 -2633 -615
rect -2587 -661 -2517 -615
rect -2471 -661 -2401 -615
rect -2355 -661 -2285 -615
rect -2239 -661 -2169 -615
rect -2123 -661 -2053 -615
rect -2007 -661 -1937 -615
rect -1891 -661 -1821 -615
rect -1775 -661 -1705 -615
rect -1659 -661 -1589 -615
rect -1543 -661 -1473 -615
rect -1427 -661 -1357 -615
rect -1311 -661 -1241 -615
rect -1195 -661 -1125 -615
rect -1079 -661 -1009 -615
rect -963 -661 -893 -615
rect -847 -661 -777 -615
rect -731 -661 -661 -615
rect -615 -661 -545 -615
rect -499 -661 -429 -615
rect -383 -661 -313 -615
rect -267 -661 -197 -615
rect -151 -661 -81 -615
rect -35 -661 35 -615
rect 81 -661 151 -615
rect 197 -661 267 -615
rect 313 -661 383 -615
rect 429 -661 499 -615
rect 545 -661 615 -615
rect 661 -661 731 -615
rect 777 -661 847 -615
rect 893 -661 963 -615
rect 1009 -661 1079 -615
rect 1125 -661 1195 -615
rect 1241 -661 1311 -615
rect 1357 -661 1427 -615
rect 1473 -661 1543 -615
rect 1589 -661 1659 -615
rect 1705 -661 1775 -615
rect 1821 -661 1891 -615
rect 1937 -661 2007 -615
rect 2053 -661 2123 -615
rect 2169 -661 2239 -615
rect 2285 -661 2355 -615
rect 2401 -661 2471 -615
rect 2517 -661 2587 -615
rect 2633 -661 2703 -615
rect 2749 -661 2819 -615
rect 2865 -661 2935 -615
rect 2981 -661 3051 -615
rect 3097 -661 3167 -615
rect 3213 -661 3283 -615
rect 3329 -661 3399 -615
rect 3445 -661 3515 -615
rect 3561 -661 3631 -615
rect 3677 -661 3747 -615
rect 3793 -661 3863 -615
rect 3909 -661 3979 -615
rect 4025 -661 4095 -615
rect 4141 -661 4211 -615
rect 4257 -661 4327 -615
rect 4373 -661 4443 -615
rect 4489 -661 4559 -615
rect 4605 -661 4675 -615
rect 4721 -661 4791 -615
rect 4837 -661 4907 -615
rect 4953 -661 5023 -615
rect 5069 -661 5139 -615
rect 5185 -661 5255 -615
rect 5301 -661 5371 -615
rect 5417 -661 5487 -615
rect 5533 -661 5603 -615
rect 5649 -661 5719 -615
rect 5765 -661 5776 -615
rect -5776 -731 5776 -661
rect -5776 -777 -5765 -731
rect -5719 -777 -5649 -731
rect -5603 -777 -5533 -731
rect -5487 -777 -5417 -731
rect -5371 -777 -5301 -731
rect -5255 -777 -5185 -731
rect -5139 -777 -5069 -731
rect -5023 -777 -4953 -731
rect -4907 -777 -4837 -731
rect -4791 -777 -4721 -731
rect -4675 -777 -4605 -731
rect -4559 -777 -4489 -731
rect -4443 -777 -4373 -731
rect -4327 -777 -4257 -731
rect -4211 -777 -4141 -731
rect -4095 -777 -4025 -731
rect -3979 -777 -3909 -731
rect -3863 -777 -3793 -731
rect -3747 -777 -3677 -731
rect -3631 -777 -3561 -731
rect -3515 -777 -3445 -731
rect -3399 -777 -3329 -731
rect -3283 -777 -3213 -731
rect -3167 -777 -3097 -731
rect -3051 -777 -2981 -731
rect -2935 -777 -2865 -731
rect -2819 -777 -2749 -731
rect -2703 -777 -2633 -731
rect -2587 -777 -2517 -731
rect -2471 -777 -2401 -731
rect -2355 -777 -2285 -731
rect -2239 -777 -2169 -731
rect -2123 -777 -2053 -731
rect -2007 -777 -1937 -731
rect -1891 -777 -1821 -731
rect -1775 -777 -1705 -731
rect -1659 -777 -1589 -731
rect -1543 -777 -1473 -731
rect -1427 -777 -1357 -731
rect -1311 -777 -1241 -731
rect -1195 -777 -1125 -731
rect -1079 -777 -1009 -731
rect -963 -777 -893 -731
rect -847 -777 -777 -731
rect -731 -777 -661 -731
rect -615 -777 -545 -731
rect -499 -777 -429 -731
rect -383 -777 -313 -731
rect -267 -777 -197 -731
rect -151 -777 -81 -731
rect -35 -777 35 -731
rect 81 -777 151 -731
rect 197 -777 267 -731
rect 313 -777 383 -731
rect 429 -777 499 -731
rect 545 -777 615 -731
rect 661 -777 731 -731
rect 777 -777 847 -731
rect 893 -777 963 -731
rect 1009 -777 1079 -731
rect 1125 -777 1195 -731
rect 1241 -777 1311 -731
rect 1357 -777 1427 -731
rect 1473 -777 1543 -731
rect 1589 -777 1659 -731
rect 1705 -777 1775 -731
rect 1821 -777 1891 -731
rect 1937 -777 2007 -731
rect 2053 -777 2123 -731
rect 2169 -777 2239 -731
rect 2285 -777 2355 -731
rect 2401 -777 2471 -731
rect 2517 -777 2587 -731
rect 2633 -777 2703 -731
rect 2749 -777 2819 -731
rect 2865 -777 2935 -731
rect 2981 -777 3051 -731
rect 3097 -777 3167 -731
rect 3213 -777 3283 -731
rect 3329 -777 3399 -731
rect 3445 -777 3515 -731
rect 3561 -777 3631 -731
rect 3677 -777 3747 -731
rect 3793 -777 3863 -731
rect 3909 -777 3979 -731
rect 4025 -777 4095 -731
rect 4141 -777 4211 -731
rect 4257 -777 4327 -731
rect 4373 -777 4443 -731
rect 4489 -777 4559 -731
rect 4605 -777 4675 -731
rect 4721 -777 4791 -731
rect 4837 -777 4907 -731
rect 4953 -777 5023 -731
rect 5069 -777 5139 -731
rect 5185 -777 5255 -731
rect 5301 -777 5371 -731
rect 5417 -777 5487 -731
rect 5533 -777 5603 -731
rect 5649 -777 5719 -731
rect 5765 -777 5776 -731
rect -5776 -847 5776 -777
rect -5776 -893 -5765 -847
rect -5719 -893 -5649 -847
rect -5603 -893 -5533 -847
rect -5487 -893 -5417 -847
rect -5371 -893 -5301 -847
rect -5255 -893 -5185 -847
rect -5139 -893 -5069 -847
rect -5023 -893 -4953 -847
rect -4907 -893 -4837 -847
rect -4791 -893 -4721 -847
rect -4675 -893 -4605 -847
rect -4559 -893 -4489 -847
rect -4443 -893 -4373 -847
rect -4327 -893 -4257 -847
rect -4211 -893 -4141 -847
rect -4095 -893 -4025 -847
rect -3979 -893 -3909 -847
rect -3863 -893 -3793 -847
rect -3747 -893 -3677 -847
rect -3631 -893 -3561 -847
rect -3515 -893 -3445 -847
rect -3399 -893 -3329 -847
rect -3283 -893 -3213 -847
rect -3167 -893 -3097 -847
rect -3051 -893 -2981 -847
rect -2935 -893 -2865 -847
rect -2819 -893 -2749 -847
rect -2703 -893 -2633 -847
rect -2587 -893 -2517 -847
rect -2471 -893 -2401 -847
rect -2355 -893 -2285 -847
rect -2239 -893 -2169 -847
rect -2123 -893 -2053 -847
rect -2007 -893 -1937 -847
rect -1891 -893 -1821 -847
rect -1775 -893 -1705 -847
rect -1659 -893 -1589 -847
rect -1543 -893 -1473 -847
rect -1427 -893 -1357 -847
rect -1311 -893 -1241 -847
rect -1195 -893 -1125 -847
rect -1079 -893 -1009 -847
rect -963 -893 -893 -847
rect -847 -893 -777 -847
rect -731 -893 -661 -847
rect -615 -893 -545 -847
rect -499 -893 -429 -847
rect -383 -893 -313 -847
rect -267 -893 -197 -847
rect -151 -893 -81 -847
rect -35 -893 35 -847
rect 81 -893 151 -847
rect 197 -893 267 -847
rect 313 -893 383 -847
rect 429 -893 499 -847
rect 545 -893 615 -847
rect 661 -893 731 -847
rect 777 -893 847 -847
rect 893 -893 963 -847
rect 1009 -893 1079 -847
rect 1125 -893 1195 -847
rect 1241 -893 1311 -847
rect 1357 -893 1427 -847
rect 1473 -893 1543 -847
rect 1589 -893 1659 -847
rect 1705 -893 1775 -847
rect 1821 -893 1891 -847
rect 1937 -893 2007 -847
rect 2053 -893 2123 -847
rect 2169 -893 2239 -847
rect 2285 -893 2355 -847
rect 2401 -893 2471 -847
rect 2517 -893 2587 -847
rect 2633 -893 2703 -847
rect 2749 -893 2819 -847
rect 2865 -893 2935 -847
rect 2981 -893 3051 -847
rect 3097 -893 3167 -847
rect 3213 -893 3283 -847
rect 3329 -893 3399 -847
rect 3445 -893 3515 -847
rect 3561 -893 3631 -847
rect 3677 -893 3747 -847
rect 3793 -893 3863 -847
rect 3909 -893 3979 -847
rect 4025 -893 4095 -847
rect 4141 -893 4211 -847
rect 4257 -893 4327 -847
rect 4373 -893 4443 -847
rect 4489 -893 4559 -847
rect 4605 -893 4675 -847
rect 4721 -893 4791 -847
rect 4837 -893 4907 -847
rect 4953 -893 5023 -847
rect 5069 -893 5139 -847
rect 5185 -893 5255 -847
rect 5301 -893 5371 -847
rect 5417 -893 5487 -847
rect 5533 -893 5603 -847
rect 5649 -893 5719 -847
rect 5765 -893 5776 -847
rect -5776 -963 5776 -893
rect -5776 -1009 -5765 -963
rect -5719 -1009 -5649 -963
rect -5603 -1009 -5533 -963
rect -5487 -1009 -5417 -963
rect -5371 -1009 -5301 -963
rect -5255 -1009 -5185 -963
rect -5139 -1009 -5069 -963
rect -5023 -1009 -4953 -963
rect -4907 -1009 -4837 -963
rect -4791 -1009 -4721 -963
rect -4675 -1009 -4605 -963
rect -4559 -1009 -4489 -963
rect -4443 -1009 -4373 -963
rect -4327 -1009 -4257 -963
rect -4211 -1009 -4141 -963
rect -4095 -1009 -4025 -963
rect -3979 -1009 -3909 -963
rect -3863 -1009 -3793 -963
rect -3747 -1009 -3677 -963
rect -3631 -1009 -3561 -963
rect -3515 -1009 -3445 -963
rect -3399 -1009 -3329 -963
rect -3283 -1009 -3213 -963
rect -3167 -1009 -3097 -963
rect -3051 -1009 -2981 -963
rect -2935 -1009 -2865 -963
rect -2819 -1009 -2749 -963
rect -2703 -1009 -2633 -963
rect -2587 -1009 -2517 -963
rect -2471 -1009 -2401 -963
rect -2355 -1009 -2285 -963
rect -2239 -1009 -2169 -963
rect -2123 -1009 -2053 -963
rect -2007 -1009 -1937 -963
rect -1891 -1009 -1821 -963
rect -1775 -1009 -1705 -963
rect -1659 -1009 -1589 -963
rect -1543 -1009 -1473 -963
rect -1427 -1009 -1357 -963
rect -1311 -1009 -1241 -963
rect -1195 -1009 -1125 -963
rect -1079 -1009 -1009 -963
rect -963 -1009 -893 -963
rect -847 -1009 -777 -963
rect -731 -1009 -661 -963
rect -615 -1009 -545 -963
rect -499 -1009 -429 -963
rect -383 -1009 -313 -963
rect -267 -1009 -197 -963
rect -151 -1009 -81 -963
rect -35 -1009 35 -963
rect 81 -1009 151 -963
rect 197 -1009 267 -963
rect 313 -1009 383 -963
rect 429 -1009 499 -963
rect 545 -1009 615 -963
rect 661 -1009 731 -963
rect 777 -1009 847 -963
rect 893 -1009 963 -963
rect 1009 -1009 1079 -963
rect 1125 -1009 1195 -963
rect 1241 -1009 1311 -963
rect 1357 -1009 1427 -963
rect 1473 -1009 1543 -963
rect 1589 -1009 1659 -963
rect 1705 -1009 1775 -963
rect 1821 -1009 1891 -963
rect 1937 -1009 2007 -963
rect 2053 -1009 2123 -963
rect 2169 -1009 2239 -963
rect 2285 -1009 2355 -963
rect 2401 -1009 2471 -963
rect 2517 -1009 2587 -963
rect 2633 -1009 2703 -963
rect 2749 -1009 2819 -963
rect 2865 -1009 2935 -963
rect 2981 -1009 3051 -963
rect 3097 -1009 3167 -963
rect 3213 -1009 3283 -963
rect 3329 -1009 3399 -963
rect 3445 -1009 3515 -963
rect 3561 -1009 3631 -963
rect 3677 -1009 3747 -963
rect 3793 -1009 3863 -963
rect 3909 -1009 3979 -963
rect 4025 -1009 4095 -963
rect 4141 -1009 4211 -963
rect 4257 -1009 4327 -963
rect 4373 -1009 4443 -963
rect 4489 -1009 4559 -963
rect 4605 -1009 4675 -963
rect 4721 -1009 4791 -963
rect 4837 -1009 4907 -963
rect 4953 -1009 5023 -963
rect 5069 -1009 5139 -963
rect 5185 -1009 5255 -963
rect 5301 -1009 5371 -963
rect 5417 -1009 5487 -963
rect 5533 -1009 5603 -963
rect 5649 -1009 5719 -963
rect 5765 -1009 5776 -963
rect -5776 -1079 5776 -1009
rect -5776 -1125 -5765 -1079
rect -5719 -1125 -5649 -1079
rect -5603 -1125 -5533 -1079
rect -5487 -1125 -5417 -1079
rect -5371 -1125 -5301 -1079
rect -5255 -1125 -5185 -1079
rect -5139 -1125 -5069 -1079
rect -5023 -1125 -4953 -1079
rect -4907 -1125 -4837 -1079
rect -4791 -1125 -4721 -1079
rect -4675 -1125 -4605 -1079
rect -4559 -1125 -4489 -1079
rect -4443 -1125 -4373 -1079
rect -4327 -1125 -4257 -1079
rect -4211 -1125 -4141 -1079
rect -4095 -1125 -4025 -1079
rect -3979 -1125 -3909 -1079
rect -3863 -1125 -3793 -1079
rect -3747 -1125 -3677 -1079
rect -3631 -1125 -3561 -1079
rect -3515 -1125 -3445 -1079
rect -3399 -1125 -3329 -1079
rect -3283 -1125 -3213 -1079
rect -3167 -1125 -3097 -1079
rect -3051 -1125 -2981 -1079
rect -2935 -1125 -2865 -1079
rect -2819 -1125 -2749 -1079
rect -2703 -1125 -2633 -1079
rect -2587 -1125 -2517 -1079
rect -2471 -1125 -2401 -1079
rect -2355 -1125 -2285 -1079
rect -2239 -1125 -2169 -1079
rect -2123 -1125 -2053 -1079
rect -2007 -1125 -1937 -1079
rect -1891 -1125 -1821 -1079
rect -1775 -1125 -1705 -1079
rect -1659 -1125 -1589 -1079
rect -1543 -1125 -1473 -1079
rect -1427 -1125 -1357 -1079
rect -1311 -1125 -1241 -1079
rect -1195 -1125 -1125 -1079
rect -1079 -1125 -1009 -1079
rect -963 -1125 -893 -1079
rect -847 -1125 -777 -1079
rect -731 -1125 -661 -1079
rect -615 -1125 -545 -1079
rect -499 -1125 -429 -1079
rect -383 -1125 -313 -1079
rect -267 -1125 -197 -1079
rect -151 -1125 -81 -1079
rect -35 -1125 35 -1079
rect 81 -1125 151 -1079
rect 197 -1125 267 -1079
rect 313 -1125 383 -1079
rect 429 -1125 499 -1079
rect 545 -1125 615 -1079
rect 661 -1125 731 -1079
rect 777 -1125 847 -1079
rect 893 -1125 963 -1079
rect 1009 -1125 1079 -1079
rect 1125 -1125 1195 -1079
rect 1241 -1125 1311 -1079
rect 1357 -1125 1427 -1079
rect 1473 -1125 1543 -1079
rect 1589 -1125 1659 -1079
rect 1705 -1125 1775 -1079
rect 1821 -1125 1891 -1079
rect 1937 -1125 2007 -1079
rect 2053 -1125 2123 -1079
rect 2169 -1125 2239 -1079
rect 2285 -1125 2355 -1079
rect 2401 -1125 2471 -1079
rect 2517 -1125 2587 -1079
rect 2633 -1125 2703 -1079
rect 2749 -1125 2819 -1079
rect 2865 -1125 2935 -1079
rect 2981 -1125 3051 -1079
rect 3097 -1125 3167 -1079
rect 3213 -1125 3283 -1079
rect 3329 -1125 3399 -1079
rect 3445 -1125 3515 -1079
rect 3561 -1125 3631 -1079
rect 3677 -1125 3747 -1079
rect 3793 -1125 3863 -1079
rect 3909 -1125 3979 -1079
rect 4025 -1125 4095 -1079
rect 4141 -1125 4211 -1079
rect 4257 -1125 4327 -1079
rect 4373 -1125 4443 -1079
rect 4489 -1125 4559 -1079
rect 4605 -1125 4675 -1079
rect 4721 -1125 4791 -1079
rect 4837 -1125 4907 -1079
rect 4953 -1125 5023 -1079
rect 5069 -1125 5139 -1079
rect 5185 -1125 5255 -1079
rect 5301 -1125 5371 -1079
rect 5417 -1125 5487 -1079
rect 5533 -1125 5603 -1079
rect 5649 -1125 5719 -1079
rect 5765 -1125 5776 -1079
rect -5776 -1136 5776 -1125
<< properties >>
string GDS_END 2783454
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2655258
<< end >>
