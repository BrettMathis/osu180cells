magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -2039 -309 2039 309
<< nsubdiff >>
rect -1895 105 1896 162
rect -1895 59 -1841 105
rect -1795 59 -1683 105
rect -1637 59 -1525 105
rect -1479 59 -1367 105
rect -1321 59 -1209 105
rect -1163 59 -1051 105
rect -1005 59 -893 105
rect -847 59 -735 105
rect -689 59 -577 105
rect -531 59 -418 105
rect -372 59 -260 105
rect -214 59 -102 105
rect -56 59 56 105
rect 102 59 214 105
rect 260 59 372 105
rect 418 59 531 105
rect 577 59 689 105
rect 735 59 847 105
rect 893 59 1005 105
rect 1051 59 1163 105
rect 1209 59 1321 105
rect 1367 59 1479 105
rect 1525 59 1637 105
rect 1683 59 1795 105
rect 1841 59 1896 105
rect -1895 -59 1896 59
rect -1895 -105 -1841 -59
rect -1795 -105 -1683 -59
rect -1637 -105 -1525 -59
rect -1479 -105 -1367 -59
rect -1321 -105 -1209 -59
rect -1163 -105 -1051 -59
rect -1005 -105 -893 -59
rect -847 -105 -735 -59
rect -689 -105 -577 -59
rect -531 -105 -418 -59
rect -372 -105 -260 -59
rect -214 -105 -102 -59
rect -56 -105 56 -59
rect 102 -105 214 -59
rect 260 -105 372 -59
rect 418 -105 531 -59
rect 577 -105 689 -59
rect 735 -105 847 -59
rect 893 -105 1005 -59
rect 1051 -105 1163 -59
rect 1209 -105 1321 -59
rect 1367 -105 1479 -59
rect 1525 -105 1637 -59
rect 1683 -105 1795 -59
rect 1841 -105 1896 -59
rect -1895 -162 1896 -105
<< nsubdiffcont >>
rect -1841 59 -1795 105
rect -1683 59 -1637 105
rect -1525 59 -1479 105
rect -1367 59 -1321 105
rect -1209 59 -1163 105
rect -1051 59 -1005 105
rect -893 59 -847 105
rect -735 59 -689 105
rect -577 59 -531 105
rect -418 59 -372 105
rect -260 59 -214 105
rect -102 59 -56 105
rect 56 59 102 105
rect 214 59 260 105
rect 372 59 418 105
rect 531 59 577 105
rect 689 59 735 105
rect 847 59 893 105
rect 1005 59 1051 105
rect 1163 59 1209 105
rect 1321 59 1367 105
rect 1479 59 1525 105
rect 1637 59 1683 105
rect 1795 59 1841 105
rect -1841 -105 -1795 -59
rect -1683 -105 -1637 -59
rect -1525 -105 -1479 -59
rect -1367 -105 -1321 -59
rect -1209 -105 -1163 -59
rect -1051 -105 -1005 -59
rect -893 -105 -847 -59
rect -735 -105 -689 -59
rect -577 -105 -531 -59
rect -418 -105 -372 -59
rect -260 -105 -214 -59
rect -102 -105 -56 -59
rect 56 -105 102 -59
rect 214 -105 260 -59
rect 372 -105 418 -59
rect 531 -105 577 -59
rect 689 -105 735 -59
rect 847 -105 893 -59
rect 1005 -105 1051 -59
rect 1163 -105 1209 -59
rect 1321 -105 1367 -59
rect 1479 -105 1525 -59
rect 1637 -105 1683 -59
rect 1795 -105 1841 -59
<< metal1 >>
rect -1876 105 1876 142
rect -1876 59 -1841 105
rect -1795 59 -1683 105
rect -1637 59 -1525 105
rect -1479 59 -1367 105
rect -1321 59 -1209 105
rect -1163 59 -1051 105
rect -1005 59 -893 105
rect -847 59 -735 105
rect -689 59 -577 105
rect -531 59 -418 105
rect -372 59 -260 105
rect -214 59 -102 105
rect -56 59 56 105
rect 102 59 214 105
rect 260 59 372 105
rect 418 59 531 105
rect 577 59 689 105
rect 735 59 847 105
rect 893 59 1005 105
rect 1051 59 1163 105
rect 1209 59 1321 105
rect 1367 59 1479 105
rect 1525 59 1637 105
rect 1683 59 1795 105
rect 1841 59 1876 105
rect -1876 -59 1876 59
rect -1876 -105 -1841 -59
rect -1795 -105 -1683 -59
rect -1637 -105 -1525 -59
rect -1479 -105 -1367 -59
rect -1321 -105 -1209 -59
rect -1163 -105 -1051 -59
rect -1005 -105 -893 -59
rect -847 -105 -735 -59
rect -689 -105 -577 -59
rect -531 -105 -418 -59
rect -372 -105 -260 -59
rect -214 -105 -102 -59
rect -56 -105 56 -59
rect 102 -105 214 -59
rect 260 -105 372 -59
rect 418 -105 531 -59
rect 577 -105 689 -59
rect 735 -105 847 -59
rect 893 -105 1005 -59
rect 1051 -105 1163 -59
rect 1209 -105 1321 -59
rect 1367 -105 1479 -59
rect 1525 -105 1637 -59
rect 1683 -105 1795 -59
rect 1841 -105 1876 -59
rect -1876 -142 1876 -105
<< properties >>
string GDS_END 772644
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 769312
<< end >>
