magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 918 896 1098
rect 49 710 95 918
rect 273 664 319 872
rect 477 710 523 918
rect 701 664 767 872
rect 273 618 767 664
rect 137 443 465 542
rect 366 354 418 443
rect 702 288 767 618
rect 273 242 767 288
rect 49 90 95 204
rect 273 136 319 242
rect 497 90 543 196
rect 721 136 767 242
rect 0 -90 896 90
<< labels >>
rlabel metal1 s 137 443 465 542 6 I
port 1 nsew default input
rlabel metal1 s 366 354 418 443 6 I
port 1 nsew default input
rlabel metal1 s 701 664 767 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 664 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 273 618 767 664 6 ZN
port 2 nsew default output
rlabel metal1 s 702 288 767 618 6 ZN
port 2 nsew default output
rlabel metal1 s 273 242 767 288 6 ZN
port 2 nsew default output
rlabel metal1 s 721 136 767 242 6 ZN
port 2 nsew default output
rlabel metal1 s 273 136 319 242 6 ZN
port 2 nsew default output
rlabel metal1 s 0 918 896 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 196 95 204 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 196 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 196 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 896 90 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1421662
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1418760
<< end >>
