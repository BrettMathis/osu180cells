magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4454 1094
<< pwell >>
rect -86 -86 4454 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 180 836 320
rect 940 180 1060 320
rect 1164 180 1284 320
rect 1332 180 1452 320
rect 1596 180 1716 320
rect 1864 180 1984 320
rect 2088 180 2208 320
rect 2312 180 2432 320
rect 2536 180 2656 320
rect 2760 180 2880 320
rect 3020 69 3140 333
rect 3388 69 3508 333
rect 3612 69 3732 333
rect 3836 69 3956 333
rect 4060 69 4180 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 720 593 820 793
rect 924 593 1024 793
rect 1128 593 1228 793
rect 1332 593 1432 793
rect 1536 593 1636 793
rect 1884 640 1984 840
rect 2088 640 2188 840
rect 2313 640 2413 840
rect 2532 640 2632 840
rect 2780 573 2880 939
rect 3040 573 3140 939
rect 3408 573 3508 939
rect 3612 573 3712 939
rect 3816 573 3916 939
rect 4020 573 4120 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 2940 320 3020 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 239 716 320
rect 628 193 641 239
rect 687 193 716 239
rect 628 180 716 193
rect 836 307 940 320
rect 836 261 865 307
rect 911 261 940 307
rect 836 180 940 261
rect 1060 307 1164 320
rect 1060 261 1089 307
rect 1135 261 1164 307
rect 1060 180 1164 261
rect 1284 180 1332 320
rect 1452 180 1596 320
rect 1716 239 1864 320
rect 1716 193 1745 239
rect 1791 193 1864 239
rect 1716 180 1864 193
rect 1984 307 2088 320
rect 1984 261 2013 307
rect 2059 261 2088 307
rect 1984 180 2088 261
rect 2208 307 2312 320
rect 2208 261 2237 307
rect 2283 261 2312 307
rect 2208 180 2312 261
rect 2432 307 2536 320
rect 2432 261 2461 307
rect 2507 261 2536 307
rect 2432 180 2536 261
rect 2656 239 2760 320
rect 2656 193 2685 239
rect 2731 193 2760 239
rect 2656 180 2760 193
rect 2880 180 3020 320
rect 2940 69 3020 180
rect 3140 320 3228 333
rect 3140 180 3169 320
rect 3215 180 3228 320
rect 3140 69 3228 180
rect 3300 222 3388 333
rect 3300 82 3313 222
rect 3359 82 3388 222
rect 3300 69 3388 82
rect 3508 320 3612 333
rect 3508 180 3537 320
rect 3583 180 3612 320
rect 3508 69 3612 180
rect 3732 222 3836 333
rect 3732 82 3761 222
rect 3807 82 3836 222
rect 3732 69 3836 82
rect 3956 314 4060 333
rect 3956 174 3985 314
rect 4031 174 4060 314
rect 3956 69 4060 174
rect 4180 222 4268 333
rect 4180 82 4209 222
rect 4255 82 4268 222
rect 4180 69 4268 82
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 2692 926 2780 939
rect 2692 880 2705 926
rect 2751 880 2780 926
rect 2692 840 2780 880
rect 1796 827 1884 840
rect 448 586 477 726
rect 523 586 536 726
rect 632 780 720 793
rect 632 734 645 780
rect 691 734 720 780
rect 632 593 720 734
rect 820 746 924 793
rect 820 606 849 746
rect 895 606 924 746
rect 820 593 924 606
rect 1024 746 1128 793
rect 1024 606 1053 746
rect 1099 606 1128 746
rect 1024 593 1128 606
rect 1228 780 1332 793
rect 1228 640 1257 780
rect 1303 640 1332 780
rect 1228 593 1332 640
rect 1432 780 1536 793
rect 1432 734 1461 780
rect 1507 734 1536 780
rect 1432 593 1536 734
rect 1636 780 1724 793
rect 1636 640 1665 780
rect 1711 640 1724 780
rect 1796 687 1809 827
rect 1855 687 1884 827
rect 1796 640 1884 687
rect 1984 793 2088 840
rect 1984 653 2013 793
rect 2059 653 2088 793
rect 1984 640 2088 653
rect 2188 793 2313 840
rect 2188 653 2238 793
rect 2284 653 2313 793
rect 2188 640 2313 653
rect 2413 699 2532 840
rect 2413 653 2457 699
rect 2503 653 2532 699
rect 2413 640 2532 653
rect 2632 640 2780 840
rect 1636 593 1724 640
rect 448 573 536 586
rect 2700 573 2780 640
rect 2880 632 3040 939
rect 2880 586 2911 632
rect 2957 586 3040 632
rect 2880 573 3040 586
rect 3140 926 3228 939
rect 3140 786 3169 926
rect 3215 786 3228 926
rect 3140 573 3228 786
rect 3320 926 3408 939
rect 3320 786 3333 926
rect 3379 786 3408 926
rect 3320 573 3408 786
rect 3508 726 3612 939
rect 3508 586 3537 726
rect 3583 586 3612 726
rect 3508 573 3612 586
rect 3712 926 3816 939
rect 3712 786 3741 926
rect 3787 786 3816 926
rect 3712 573 3816 786
rect 3916 726 4020 939
rect 3916 586 3945 726
rect 3991 586 4020 726
rect 3916 573 4020 586
rect 4120 926 4208 939
rect 4120 786 4149 926
rect 4195 786 4208 926
rect 4120 573 4208 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 193 687 239
rect 865 261 911 307
rect 1089 261 1135 307
rect 1745 193 1791 239
rect 2013 261 2059 307
rect 2237 261 2283 307
rect 2461 261 2507 307
rect 2685 193 2731 239
rect 3169 180 3215 320
rect 3313 82 3359 222
rect 3537 180 3583 320
rect 3761 82 3807 222
rect 3985 174 4031 314
rect 4209 82 4255 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 2705 880 2751 926
rect 477 586 523 726
rect 645 734 691 780
rect 849 606 895 746
rect 1053 606 1099 746
rect 1257 640 1303 780
rect 1461 734 1507 780
rect 1665 640 1711 780
rect 1809 687 1855 827
rect 2013 653 2059 793
rect 2238 653 2284 793
rect 2457 653 2503 699
rect 2911 586 2957 632
rect 3169 786 3215 926
rect 3333 786 3379 926
rect 3537 586 3583 726
rect 3741 786 3787 926
rect 3945 586 3991 726
rect 4149 786 4195 926
<< polysilicon >>
rect 348 909 1024 949
rect 144 849 244 893
rect 348 849 448 909
rect 720 793 820 837
rect 924 793 1024 909
rect 1128 932 2188 972
rect 2780 939 2880 983
rect 3040 939 3140 983
rect 3408 939 3508 983
rect 3612 939 3712 983
rect 3816 939 3916 983
rect 4020 939 4120 983
rect 1128 872 1228 932
rect 1128 826 1141 872
rect 1187 826 1228 872
rect 1884 840 1984 884
rect 2088 840 2188 932
rect 2313 840 2413 884
rect 2532 840 2632 884
rect 1128 793 1228 826
rect 1332 793 1432 837
rect 1536 793 1636 837
rect 144 504 244 573
rect 144 458 157 504
rect 203 458 244 504
rect 144 377 244 458
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 720 523 820 593
rect 924 549 1024 593
rect 1128 549 1228 593
rect 720 477 733 523
rect 779 477 820 523
rect 407 366 468 377
rect 348 333 468 366
rect 720 364 820 477
rect 1128 472 1168 549
rect 1020 432 1168 472
rect 1332 491 1432 593
rect 1536 549 1636 593
rect 1332 445 1373 491
rect 1419 445 1432 491
rect 1020 364 1060 432
rect 1212 399 1284 412
rect 1212 364 1225 399
rect 716 320 836 364
rect 940 320 1060 364
rect 1164 353 1225 364
rect 1271 353 1284 399
rect 1164 320 1284 353
rect 1332 364 1432 445
rect 1596 364 1636 549
rect 1884 583 1984 640
rect 1884 537 1897 583
rect 1943 537 1984 583
rect 1884 364 1984 537
rect 2088 500 2188 640
rect 2313 607 2413 640
rect 2313 561 2329 607
rect 2375 561 2413 607
rect 2313 548 2413 561
rect 2532 510 2632 640
rect 2088 460 2432 500
rect 1332 320 1452 364
rect 1596 320 1716 364
rect 1864 320 1984 364
rect 2088 399 2208 412
rect 2088 353 2105 399
rect 2151 353 2208 399
rect 2088 320 2208 353
rect 2312 320 2432 460
rect 2532 464 2573 510
rect 2619 464 2632 510
rect 2532 380 2632 464
rect 2780 399 2880 573
rect 2536 320 2656 380
rect 2780 364 2821 399
rect 2760 353 2821 364
rect 2867 353 2880 399
rect 3040 540 3140 573
rect 3040 494 3053 540
rect 3099 494 3140 540
rect 3040 377 3140 494
rect 3408 465 3508 573
rect 3612 465 3712 573
rect 3816 465 3916 573
rect 4020 465 4120 573
rect 3408 452 4120 465
rect 3408 406 3421 452
rect 3467 406 3646 452
rect 3692 406 3840 452
rect 3886 406 4120 452
rect 3408 393 4120 406
rect 3408 377 3508 393
rect 2760 320 2880 353
rect 3020 333 3140 377
rect 3388 333 3508 377
rect 3612 333 3732 393
rect 3836 333 3956 393
rect 4060 377 4120 393
rect 4060 333 4180 377
rect 124 131 244 175
rect 348 88 468 175
rect 716 136 836 180
rect 940 136 1060 180
rect 1164 88 1284 180
rect 1332 136 1452 180
rect 348 48 1284 88
rect 1596 88 1716 180
rect 1864 136 1984 180
rect 2088 136 2208 180
rect 2312 136 2432 180
rect 2536 136 2656 180
rect 2760 88 2880 180
rect 1596 48 2880 88
rect 3020 25 3140 69
rect 3388 25 3508 69
rect 3612 25 3732 69
rect 3836 25 3956 69
rect 4060 25 4180 69
<< polycontact >>
rect 1141 826 1187 872
rect 157 458 203 504
rect 361 366 407 412
rect 733 477 779 523
rect 1373 445 1419 491
rect 1225 353 1271 399
rect 1897 537 1943 583
rect 2329 561 2375 607
rect 2105 353 2151 399
rect 2573 464 2619 510
rect 2821 353 2867 399
rect 3053 494 3099 540
rect 3421 406 3467 452
rect 3646 406 3692 452
rect 3840 406 3886 452
<< metal1 >>
rect 0 926 4368 1098
rect 0 918 2705 926
rect 273 836 319 918
rect 69 739 115 750
rect 645 780 691 918
rect 273 685 319 696
rect 477 726 523 737
rect 115 599 407 634
rect 69 588 407 599
rect 142 504 315 542
rect 142 458 157 504
rect 203 458 315 504
rect 142 447 315 458
rect 361 412 407 588
rect 49 366 361 401
rect 49 355 407 366
rect 645 723 691 734
rect 737 826 1141 872
rect 1187 826 1198 872
rect 737 677 783 826
rect 1257 780 1303 791
rect 523 631 783 677
rect 849 746 911 757
rect 523 586 543 631
rect 49 320 95 355
rect 49 263 95 274
rect 477 320 543 586
rect 895 606 911 746
rect 589 523 779 542
rect 589 477 733 523
rect 589 466 779 477
rect 477 274 497 320
rect 477 263 543 274
rect 849 307 911 606
rect 849 261 865 307
rect 849 250 911 261
rect 1053 746 1099 757
rect 1461 780 1507 918
rect 1809 827 1855 918
rect 2751 918 3169 926
rect 2705 869 2751 880
rect 1461 723 1507 734
rect 1665 780 1711 791
rect 1303 640 1665 675
rect 1809 676 1855 687
rect 2013 793 2059 804
rect 1257 629 1711 640
rect 1053 583 1099 606
rect 1053 537 1897 583
rect 1943 537 1954 583
rect 1053 307 1135 537
rect 2013 491 2059 653
rect 1362 445 1373 491
rect 1419 445 2059 491
rect 1214 353 1225 399
rect 1271 353 1967 399
rect 1053 261 1089 307
rect 1053 250 1135 261
rect 273 234 319 245
rect 273 90 319 188
rect 641 239 687 250
rect 641 90 687 193
rect 1745 239 1791 250
rect 1745 90 1791 193
rect 1921 204 1967 353
rect 2013 307 2059 445
rect 2237 793 3060 804
rect 2237 653 2238 793
rect 2284 758 3060 793
rect 3215 918 3333 926
rect 3169 775 3215 786
rect 3379 918 3741 926
rect 3333 775 3379 786
rect 3787 918 4149 926
rect 3741 775 3787 786
rect 4195 918 4368 926
rect 4149 775 4195 786
rect 2237 642 2284 653
rect 2457 699 2507 710
rect 2503 653 2507 699
rect 2013 250 2059 261
rect 2105 399 2151 410
rect 2105 204 2151 353
rect 2237 307 2283 642
rect 2237 250 2283 261
rect 2329 607 2375 618
rect 2329 204 2375 561
rect 2457 307 2507 653
rect 2911 632 2968 643
rect 2957 586 2968 632
rect 2911 510 2968 586
rect 2562 464 2573 510
rect 2619 464 2968 510
rect 3014 540 3060 758
rect 3537 726 3583 737
rect 3945 726 4035 737
rect 3583 586 3945 659
rect 3991 586 4035 726
rect 3537 575 4035 586
rect 3014 494 3053 540
rect 3099 494 3110 540
rect 2922 448 2968 464
rect 3169 452 3897 455
rect 3169 448 3421 452
rect 2457 261 2461 307
rect 2457 250 2507 261
rect 2821 399 2867 410
rect 2922 406 3421 448
rect 3467 406 3646 452
rect 3692 406 3840 452
rect 3886 406 3897 452
rect 2922 403 3897 406
rect 2922 402 3215 403
rect 2821 318 2867 353
rect 3169 320 3215 402
rect 3943 331 4035 575
rect 1921 158 2375 204
rect 2685 239 2731 250
rect 2821 242 2882 318
rect 2685 90 2731 193
rect 3537 320 4035 331
rect 3169 169 3215 180
rect 3313 222 3359 233
rect 0 82 3313 90
rect 3583 314 4035 320
rect 3583 279 3985 314
rect 3537 169 3583 180
rect 3761 222 3807 233
rect 3359 82 3761 90
rect 3950 174 3985 279
rect 4031 174 4035 314
rect 3950 163 4035 174
rect 4209 222 4255 233
rect 3807 82 4209 90
rect 4255 82 4368 90
rect 0 -90 4368 82
<< labels >>
flabel metal1 s 142 447 315 542 0 FreeSans 200 0 0 0 CLKN
port 3 nsew clock input
flabel metal1 s 589 466 779 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3945 659 4035 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2821 318 2867 410 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 0 918 4368 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2685 245 2731 250 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2821 242 2882 318 1 RN
port 2 nsew default input
rlabel metal1 s 3537 659 3583 737 1 Q
port 4 nsew default output
rlabel metal1 s 3537 575 4035 659 1 Q
port 4 nsew default output
rlabel metal1 s 3943 331 4035 575 1 Q
port 4 nsew default output
rlabel metal1 s 3537 279 4035 331 1 Q
port 4 nsew default output
rlabel metal1 s 3950 169 4035 279 1 Q
port 4 nsew default output
rlabel metal1 s 3537 169 3583 279 1 Q
port 4 nsew default output
rlabel metal1 s 3950 163 4035 169 1 Q
port 4 nsew default output
rlabel metal1 s 4149 869 4195 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3741 869 3787 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3333 869 3379 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3169 869 3215 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2705 869 2751 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 869 1855 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 869 1507 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 869 691 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 869 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4149 775 4195 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3741 775 3787 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3333 775 3379 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3169 775 3215 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 775 1855 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 775 1507 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 775 691 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 723 1855 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 723 1507 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 723 691 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 723 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 685 1855 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 676 1855 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1745 245 1791 250 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 245 687 250 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2685 233 2731 245 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1745 233 1791 245 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4209 90 4255 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3761 90 3807 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3313 90 3359 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2685 90 2731 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1745 90 1791 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4368 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4368 1008
string GDS_END 1509338
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1499334
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
