magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 2900 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 570 190 630 360
rect 800 190 860 360
rect 910 190 970 360
rect 1080 190 1140 360
rect 1190 190 1250 360
rect 1420 190 1480 360
rect 1630 190 1690 360
rect 1800 190 1860 360
rect 2160 190 2220 360
rect 2480 190 2540 360
rect 2650 190 2710 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 570 700 630 1040
rect 800 700 860 1040
rect 910 700 970 1040
rect 1080 700 1140 1040
rect 1190 700 1250 1040
rect 1420 700 1480 1040
rect 1630 700 1690 1040
rect 1800 700 1860 1040
rect 2160 700 2220 1040
rect 2480 700 2540 1040
rect 2650 700 2710 1040
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 263 360 360
rect 250 217 282 263
rect 328 217 360 263
rect 250 190 360 217
rect 420 190 570 360
rect 630 263 800 360
rect 630 217 692 263
rect 738 217 800 263
rect 630 190 800 217
rect 860 190 910 360
rect 970 258 1080 360
rect 970 212 1002 258
rect 1048 212 1080 258
rect 970 190 1080 212
rect 1140 190 1190 360
rect 1250 258 1420 360
rect 1250 212 1312 258
rect 1358 212 1420 258
rect 1250 190 1420 212
rect 1480 190 1630 360
rect 1690 263 1800 360
rect 1690 217 1722 263
rect 1768 217 1800 263
rect 1690 190 1800 217
rect 1860 258 1960 360
rect 1860 212 1892 258
rect 1938 212 1960 258
rect 1860 190 1960 212
rect 2060 258 2160 360
rect 2060 212 2082 258
rect 2128 212 2160 258
rect 2060 190 2160 212
rect 2220 298 2320 360
rect 2220 252 2252 298
rect 2298 252 2320 298
rect 2220 190 2320 252
rect 2380 298 2480 360
rect 2380 252 2402 298
rect 2448 252 2480 298
rect 2380 190 2480 252
rect 2540 278 2650 360
rect 2540 232 2572 278
rect 2618 232 2650 278
rect 2540 190 2650 232
rect 2710 298 2810 360
rect 2710 252 2742 298
rect 2788 252 2810 298
rect 2710 190 2810 252
<< pdiff >>
rect 90 987 190 1040
rect 90 753 112 987
rect 158 753 190 987
rect 90 700 190 753
rect 250 1018 360 1040
rect 250 972 282 1018
rect 328 972 360 1018
rect 250 700 360 972
rect 420 700 570 1040
rect 630 1010 800 1040
rect 630 870 692 1010
rect 738 870 800 1010
rect 630 700 800 870
rect 860 700 910 1040
rect 970 1000 1080 1040
rect 970 860 1002 1000
rect 1048 860 1080 1000
rect 970 700 1080 860
rect 1140 700 1190 1040
rect 1250 1010 1420 1040
rect 1250 870 1312 1010
rect 1358 870 1420 1010
rect 1250 700 1420 870
rect 1480 700 1630 1040
rect 1690 1018 1800 1040
rect 1690 972 1722 1018
rect 1768 972 1800 1018
rect 1690 700 1800 972
rect 1860 987 1960 1040
rect 1860 753 1892 987
rect 1938 753 1960 987
rect 1860 700 1960 753
rect 2060 987 2160 1040
rect 2060 753 2082 987
rect 2128 753 2160 987
rect 2060 700 2160 753
rect 2220 987 2320 1040
rect 2220 753 2252 987
rect 2298 753 2320 987
rect 2220 700 2320 753
rect 2380 987 2480 1040
rect 2380 753 2402 987
rect 2448 753 2480 987
rect 2380 700 2480 753
rect 2540 995 2650 1040
rect 2540 855 2572 995
rect 2618 855 2650 995
rect 2540 700 2650 855
rect 2710 978 2810 1040
rect 2710 932 2742 978
rect 2788 932 2810 978
rect 2710 700 2810 932
<< ndiffc >>
rect 112 252 158 298
rect 282 217 328 263
rect 692 217 738 263
rect 1002 212 1048 258
rect 1312 212 1358 258
rect 1722 217 1768 263
rect 1892 212 1938 258
rect 2082 212 2128 258
rect 2252 252 2298 298
rect 2402 252 2448 298
rect 2572 232 2618 278
rect 2742 252 2788 298
<< pdiffc >>
rect 112 753 158 987
rect 282 972 328 1018
rect 692 870 738 1010
rect 1002 860 1048 1000
rect 1312 870 1358 1010
rect 1722 972 1768 1018
rect 1892 753 1938 987
rect 2082 753 2128 987
rect 2252 753 2298 987
rect 2402 753 2448 987
rect 2572 855 2618 995
rect 2742 932 2788 978
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
rect 1290 1178 1380 1200
rect 1290 1132 1312 1178
rect 1358 1132 1380 1178
rect 1290 1110 1380 1132
rect 1530 1178 1620 1200
rect 1530 1132 1552 1178
rect 1598 1132 1620 1178
rect 1530 1110 1620 1132
rect 1770 1178 1860 1200
rect 1770 1132 1792 1178
rect 1838 1132 1860 1178
rect 1770 1110 1860 1132
rect 2010 1178 2100 1200
rect 2010 1132 2032 1178
rect 2078 1132 2100 1178
rect 2010 1110 2100 1132
rect 2250 1178 2340 1200
rect 2250 1132 2272 1178
rect 2318 1132 2340 1178
rect 2250 1110 2340 1132
rect 2490 1178 2580 1200
rect 2490 1132 2512 1178
rect 2558 1132 2580 1178
rect 2490 1110 2580 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
rect 1312 1132 1358 1178
rect 1552 1132 1598 1178
rect 1792 1132 1838 1178
rect 2032 1132 2078 1178
rect 2272 1132 2318 1178
rect 2512 1132 2558 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 570 1040 630 1090
rect 800 1040 860 1090
rect 910 1040 970 1090
rect 1080 1040 1140 1090
rect 1190 1040 1250 1090
rect 1420 1040 1480 1090
rect 1630 1040 1690 1090
rect 1800 1040 1860 1090
rect 2160 1040 2220 1090
rect 2480 1040 2540 1090
rect 2650 1040 2710 1090
rect 190 680 250 700
rect 190 653 290 680
rect 190 607 217 653
rect 263 607 290 653
rect 360 650 420 700
rect 570 680 630 700
rect 500 658 630 680
rect 190 580 290 607
rect 340 623 450 650
rect 190 360 250 580
rect 340 577 377 623
rect 423 577 450 623
rect 500 612 532 658
rect 578 650 630 658
rect 578 612 600 650
rect 500 590 600 612
rect 340 550 450 577
rect 800 570 860 700
rect 910 680 970 700
rect 1080 680 1140 700
rect 910 610 1140 680
rect 360 360 420 550
rect 650 520 860 570
rect 650 480 710 520
rect 530 453 710 480
rect 990 470 1050 610
rect 1190 570 1250 700
rect 1420 680 1480 700
rect 1420 653 1540 680
rect 1420 650 1467 653
rect 1440 607 1467 650
rect 1513 607 1540 653
rect 1440 580 1540 607
rect 1190 520 1390 570
rect 1630 520 1690 700
rect 1800 650 1860 700
rect 1800 623 1900 650
rect 1800 577 1827 623
rect 1873 577 1900 623
rect 2160 590 2220 700
rect 2480 590 2540 700
rect 1800 550 1900 577
rect 2100 563 2220 590
rect 1340 500 1390 520
rect 530 407 567 453
rect 613 407 710 453
rect 530 400 710 407
rect 760 448 860 470
rect 760 402 787 448
rect 833 402 860 448
rect 530 380 650 400
rect 760 380 860 402
rect 570 360 630 380
rect 800 360 860 380
rect 910 460 1050 470
rect 910 448 1140 460
rect 910 402 947 448
rect 993 402 1140 448
rect 910 380 1140 402
rect 910 360 970 380
rect 1080 360 1140 380
rect 1190 448 1290 470
rect 1190 402 1217 448
rect 1263 402 1290 448
rect 1190 380 1290 402
rect 1340 453 1480 500
rect 1340 407 1397 453
rect 1443 407 1480 453
rect 1610 493 1710 520
rect 1610 447 1637 493
rect 1683 447 1710 493
rect 1610 420 1710 447
rect 1340 400 1480 407
rect 1370 380 1480 400
rect 1190 360 1250 380
rect 1420 360 1480 380
rect 1630 360 1690 420
rect 1800 360 1860 550
rect 2100 517 2127 563
rect 2173 517 2220 563
rect 2100 490 2220 517
rect 2430 563 2540 590
rect 2430 517 2457 563
rect 2503 517 2540 563
rect 2650 520 2710 700
rect 2430 490 2540 517
rect 2160 360 2220 490
rect 2480 360 2540 490
rect 2590 493 2710 520
rect 2590 447 2617 493
rect 2663 447 2710 493
rect 2590 420 2710 447
rect 2650 360 2710 420
rect 190 140 250 190
rect 360 140 420 190
rect 570 140 630 190
rect 800 140 860 190
rect 910 140 970 190
rect 1080 140 1140 190
rect 1190 140 1250 190
rect 1420 140 1480 190
rect 1630 140 1690 190
rect 1800 140 1860 190
rect 2160 140 2220 190
rect 2480 140 2540 190
rect 2650 140 2710 190
<< polycontact >>
rect 217 607 263 653
rect 377 577 423 623
rect 532 612 578 658
rect 1467 607 1513 653
rect 1827 577 1873 623
rect 567 407 613 453
rect 787 402 833 448
rect 947 402 993 448
rect 1217 402 1263 448
rect 1397 407 1443 453
rect 1637 447 1683 493
rect 2127 517 2173 563
rect 2457 517 2503 563
rect 2617 447 2663 493
<< metal1 >>
rect 0 1178 2900 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1312 1178
rect 1358 1176 1552 1178
rect 1598 1176 1792 1178
rect 1838 1176 2032 1178
rect 2078 1176 2272 1178
rect 2318 1176 2512 1178
rect 2558 1176 2900 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 1126 1132 1312 1176
rect 1366 1132 1552 1176
rect 1606 1132 1792 1176
rect 1846 1132 2032 1176
rect 2086 1132 2272 1176
rect 2326 1132 2512 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1314 1132
rect 1366 1124 1554 1132
rect 1606 1124 1794 1132
rect 1846 1124 2034 1132
rect 2086 1124 2274 1132
rect 2326 1124 2514 1132
rect 2566 1124 2900 1176
rect 0 1110 2900 1124
rect 110 987 160 1040
rect 110 753 112 987
rect 158 753 160 987
rect 280 1018 330 1110
rect 280 972 282 1018
rect 328 972 330 1018
rect 280 950 330 972
rect 660 1010 770 1040
rect 660 900 692 1010
rect 110 470 160 753
rect 100 460 160 470
rect 80 456 160 460
rect 80 404 104 456
rect 156 404 160 456
rect 80 400 160 404
rect 100 380 160 400
rect 110 298 160 380
rect 210 870 692 900
rect 738 870 770 1010
rect 210 840 770 870
rect 1000 1000 1050 1110
rect 1000 860 1002 1000
rect 1048 860 1050 1000
rect 210 660 270 840
rect 1000 820 1050 860
rect 1280 1010 1390 1040
rect 1280 896 1312 1010
rect 1280 844 1284 896
rect 1358 870 1390 1010
rect 1720 1018 1770 1110
rect 1720 972 1722 1018
rect 1768 972 1770 1018
rect 1720 950 1770 972
rect 1890 987 1940 1040
rect 1336 844 1390 870
rect 1280 840 1390 844
rect 1610 896 1710 900
rect 1610 844 1634 896
rect 1686 844 1710 896
rect 1610 840 1710 844
rect 1280 820 1340 840
rect 1630 820 1690 840
rect 1890 753 1892 987
rect 1938 753 1940 987
rect 1890 750 1940 753
rect 2080 987 2130 1110
rect 2080 753 2082 987
rect 2128 753 2130 987
rect 1890 700 2000 750
rect 2080 700 2130 753
rect 2250 987 2300 1040
rect 2250 753 2252 987
rect 2298 753 2300 987
rect 210 653 290 660
rect 210 607 217 653
rect 263 607 290 653
rect 500 658 1790 660
rect 210 600 290 607
rect 350 626 450 630
rect 210 410 270 600
rect 350 574 374 626
rect 426 574 450 626
rect 500 612 532 658
rect 578 653 1790 658
rect 578 612 1467 653
rect 500 607 1467 612
rect 1513 650 1790 653
rect 1513 630 1880 650
rect 1513 626 1900 630
rect 1513 607 1824 626
rect 500 600 1824 607
rect 350 570 450 574
rect 780 460 840 600
rect 940 460 1000 470
rect 540 456 640 460
rect 210 360 450 410
rect 540 404 564 456
rect 616 404 640 456
rect 540 400 640 404
rect 760 448 860 460
rect 760 402 787 448
rect 833 402 860 448
rect 760 400 860 402
rect 920 456 1020 460
rect 920 404 944 456
rect 996 404 1020 456
rect 1210 450 1270 600
rect 1800 574 1824 600
rect 1876 574 1900 626
rect 1800 570 1900 574
rect 1950 500 2000 700
rect 1610 496 1710 500
rect 1390 460 1450 480
rect 1380 453 1510 460
rect 920 402 947 404
rect 993 402 1020 404
rect 920 400 1020 402
rect 1190 448 1290 450
rect 1190 402 1217 448
rect 1263 402 1290 448
rect 1190 390 1290 402
rect 1380 407 1397 453
rect 1443 407 1510 453
rect 1610 444 1634 496
rect 1686 444 1710 496
rect 1610 440 1710 444
rect 1890 440 2000 500
rect 2120 563 2180 590
rect 2120 517 2127 563
rect 2173 517 2180 563
rect 1380 400 1510 407
rect 1390 380 1510 400
rect 400 330 450 360
rect 1450 366 1510 380
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 263 330 300
rect 400 280 770 330
rect 1260 326 1390 330
rect 1260 280 1284 326
rect 280 217 282 263
rect 328 217 330 263
rect 280 120 330 217
rect 660 263 770 280
rect 660 217 692 263
rect 738 217 770 263
rect 660 190 770 217
rect 1000 258 1050 280
rect 1000 212 1002 258
rect 1048 212 1050 258
rect 1000 120 1050 212
rect 1280 274 1284 280
rect 1336 274 1390 326
rect 1450 314 1454 366
rect 1506 314 1510 366
rect 1450 290 1510 314
rect 1890 366 1950 440
rect 2120 390 2180 517
rect 2250 570 2300 753
rect 2400 987 2450 1040
rect 2400 753 2402 987
rect 2448 760 2450 987
rect 2570 995 2620 1110
rect 2570 855 2572 995
rect 2618 855 2620 995
rect 2570 810 2620 855
rect 2740 978 2790 1040
rect 2740 932 2742 978
rect 2788 932 2790 978
rect 2740 900 2790 932
rect 2740 886 2850 900
rect 2740 834 2774 886
rect 2826 834 2850 886
rect 2740 830 2850 834
rect 2740 820 2840 830
rect 2448 756 2690 760
rect 2448 753 2614 756
rect 2400 704 2614 753
rect 2666 704 2690 756
rect 2400 700 2690 704
rect 2250 566 2530 570
rect 2250 514 2454 566
rect 2506 514 2530 566
rect 2250 510 2530 514
rect 1890 314 1894 366
rect 1946 314 1950 366
rect 2100 386 2200 390
rect 2100 334 2124 386
rect 2176 334 2200 386
rect 2100 330 2200 334
rect 1280 258 1390 274
rect 1280 212 1312 258
rect 1358 212 1390 258
rect 1280 190 1390 212
rect 1720 263 1770 300
rect 1720 217 1722 263
rect 1768 217 1770 263
rect 1720 120 1770 217
rect 1890 290 1950 314
rect 2250 298 2300 510
rect 2610 493 2670 700
rect 2610 447 2617 493
rect 2663 447 2670 493
rect 2610 420 2670 447
rect 1890 258 1940 290
rect 1890 212 1892 258
rect 1938 212 1940 258
rect 1890 190 1940 212
rect 2080 258 2130 280
rect 2080 212 2082 258
rect 2128 212 2130 258
rect 2080 120 2130 212
rect 2250 252 2252 298
rect 2298 252 2300 298
rect 2250 190 2300 252
rect 2400 370 2670 420
rect 2400 298 2450 370
rect 2400 252 2402 298
rect 2448 252 2450 298
rect 2400 190 2450 252
rect 2570 278 2620 320
rect 2570 232 2572 278
rect 2618 232 2620 278
rect 2570 120 2620 232
rect 2740 298 2790 820
rect 2740 252 2742 298
rect 2788 252 2790 298
rect 2740 190 2790 252
rect 0 106 2900 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2900 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2900 54
rect 0 0 2900 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 1314 1132 1358 1176
rect 1358 1132 1366 1176
rect 1554 1132 1598 1176
rect 1598 1132 1606 1176
rect 1794 1132 1838 1176
rect 1838 1132 1846 1176
rect 2034 1132 2078 1176
rect 2078 1132 2086 1176
rect 2274 1132 2318 1176
rect 2318 1132 2326 1176
rect 2514 1132 2558 1176
rect 2558 1132 2566 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 1554 1124 1606 1132
rect 1794 1124 1846 1132
rect 2034 1124 2086 1132
rect 2274 1124 2326 1132
rect 2514 1124 2566 1132
rect 104 404 156 456
rect 1284 870 1312 896
rect 1312 870 1336 896
rect 1284 844 1336 870
rect 1634 844 1686 896
rect 374 623 426 626
rect 374 577 377 623
rect 377 577 423 623
rect 423 577 426 623
rect 374 574 426 577
rect 1824 623 1876 626
rect 564 453 616 456
rect 564 407 567 453
rect 567 407 613 453
rect 613 407 616 453
rect 564 404 616 407
rect 944 448 996 456
rect 944 404 947 448
rect 947 404 993 448
rect 993 404 996 448
rect 1824 577 1827 623
rect 1827 577 1873 623
rect 1873 577 1876 623
rect 1824 574 1876 577
rect 1634 493 1686 496
rect 1634 447 1637 493
rect 1637 447 1683 493
rect 1683 447 1686 493
rect 1634 444 1686 447
rect 1284 274 1336 326
rect 1454 314 1506 366
rect 2774 834 2826 886
rect 2614 704 2666 756
rect 2454 563 2506 566
rect 2454 517 2457 563
rect 2457 517 2503 563
rect 2503 517 2506 563
rect 2454 514 2506 517
rect 1894 314 1946 366
rect 2124 334 2176 386
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 1540 1180 1620 1190
rect 1780 1180 1860 1190
rect 2020 1180 2100 1190
rect 2260 1180 2340 1190
rect 2500 1180 2580 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 1530 1176 1630 1180
rect 1530 1124 1554 1176
rect 1606 1124 1630 1176
rect 1530 1120 1630 1124
rect 1770 1176 1870 1180
rect 1770 1124 1794 1176
rect 1846 1124 1870 1176
rect 1770 1120 1870 1124
rect 2010 1176 2110 1180
rect 2010 1124 2034 1176
rect 2086 1124 2110 1176
rect 2010 1120 2110 1124
rect 2250 1176 2350 1180
rect 2250 1124 2274 1176
rect 2326 1124 2350 1176
rect 2250 1120 2350 1124
rect 2490 1176 2590 1180
rect 2490 1124 2514 1176
rect 2566 1124 2590 1176
rect 2490 1120 2590 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 1540 1110 1620 1120
rect 1780 1110 1860 1120
rect 2020 1110 2100 1120
rect 2260 1110 2340 1120
rect 2500 1110 2580 1120
rect 560 980 1510 1040
rect 350 630 450 640
rect 340 626 460 630
rect 340 574 374 626
rect 426 574 460 626
rect 340 570 460 574
rect 350 560 450 570
rect 560 470 620 980
rect 1280 910 1340 920
rect 1270 896 1350 910
rect 1270 844 1284 896
rect 1336 844 1350 896
rect 1270 830 1350 844
rect 90 460 170 470
rect 550 460 640 470
rect 930 460 1010 470
rect 80 456 180 460
rect 80 404 104 456
rect 156 404 180 456
rect 80 400 180 404
rect 540 456 640 460
rect 540 404 564 456
rect 616 404 640 456
rect 540 400 640 404
rect 920 456 1020 460
rect 920 404 944 456
rect 996 404 1020 456
rect 920 400 1020 404
rect 90 390 170 400
rect 550 390 640 400
rect 930 390 1010 400
rect 100 270 160 390
rect 940 270 1000 390
rect 1280 340 1340 830
rect 1450 380 1510 980
rect 1620 900 1700 910
rect 1610 896 2290 900
rect 1610 844 1634 896
rect 1686 844 2290 896
rect 2760 890 2840 900
rect 1610 840 2290 844
rect 1620 830 1700 840
rect 1630 510 1690 830
rect 1810 630 1890 640
rect 1800 626 1900 630
rect 1800 574 1824 626
rect 1876 574 1900 626
rect 1800 570 1900 574
rect 2230 570 2290 840
rect 2750 886 2850 890
rect 2750 834 2774 886
rect 2826 834 2850 886
rect 2750 830 2850 834
rect 2760 820 2840 830
rect 2600 760 2680 770
rect 2590 756 2690 760
rect 2590 704 2614 756
rect 2666 704 2690 756
rect 2590 700 2690 704
rect 2600 690 2680 700
rect 2440 570 2520 580
rect 1810 560 1890 570
rect 2230 566 2530 570
rect 2230 514 2454 566
rect 2506 514 2530 566
rect 2230 510 2530 514
rect 1620 500 1700 510
rect 2440 500 2520 510
rect 1610 496 1710 500
rect 1610 444 1634 496
rect 1686 444 1710 496
rect 1610 440 1710 444
rect 1620 430 1700 440
rect 2110 390 2190 400
rect 2040 386 2200 390
rect 1440 370 1520 380
rect 1880 370 1960 380
rect 1430 366 1980 370
rect 1270 330 1350 340
rect 1260 326 1350 330
rect 1260 274 1284 326
rect 1336 274 1350 326
rect 1430 314 1454 366
rect 1506 314 1894 366
rect 1946 314 1980 366
rect 1430 310 1980 314
rect 2040 334 2124 386
rect 2176 334 2200 386
rect 2040 330 2200 334
rect 2040 320 2190 330
rect 1440 300 1520 310
rect 1880 300 1960 310
rect 1260 270 1350 274
rect 100 210 1000 270
rect 1270 260 1350 270
rect 1280 240 1350 260
rect 2040 240 2100 320
rect 1280 180 2100 240
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 50 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 50 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 50 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 50 2590 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
rect 1780 40 1860 50
rect 2020 40 2100 50
rect 2260 40 2340 50
rect 2500 40 2580 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 350 560 450 640 4 D
port 1 nsew signal input
rlabel metal2 s 2760 820 2840 900 4 Q
port 2 nsew signal output
rlabel metal2 s 2600 690 2680 770 4 QN
port 3 nsew signal output
rlabel metal2 s 1810 560 1890 640 4 CLKN
port 4 nsew clock input
rlabel metal2 s 1800 570 1900 630 1 CLKN
port 4 nsew clock input
rlabel metal1 s 780 400 840 660 1 CLKN
port 4 nsew clock input
rlabel metal1 s 760 400 860 460 1 CLKN
port 4 nsew clock input
rlabel metal1 s 1210 390 1270 660 1 CLKN
port 4 nsew clock input
rlabel metal1 s 1190 390 1290 450 1 CLKN
port 4 nsew clock input
rlabel metal1 s 500 600 1790 660 1 CLKN
port 4 nsew clock input
rlabel metal1 s 500 600 1880 650 1 CLKN
port 4 nsew clock input
rlabel metal1 s 1800 570 1900 630 1 CLKN
port 4 nsew clock input
rlabel metal2 s 340 570 460 630 1 D
port 1 nsew signal input
rlabel metal1 s 350 570 450 630 1 D
port 1 nsew signal input
rlabel metal2 s 2750 830 2850 890 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 190 2790 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 820 2840 900 1 Q
port 2 nsew signal output
rlabel metal1 s 2740 830 2850 900 1 Q
port 2 nsew signal output
rlabel metal2 s 2590 700 2690 760 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 190 2450 420 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 700 2450 1040 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 370 2670 420 1 QN
port 3 nsew signal output
rlabel metal1 s 2610 370 2670 760 1 QN
port 3 nsew signal output
rlabel metal1 s 2400 700 2690 760 1 QN
port 3 nsew signal output
rlabel metal2 s 90 1120 190 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1540 1110 1620 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1530 1120 1630 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1780 1110 1860 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1770 1120 1870 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2020 1110 2100 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2010 1120 2110 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2260 1110 2340 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2250 1120 2350 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2500 1110 2580 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2490 1120 2590 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 280 950 330 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1000 820 1050 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1720 950 1770 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 2080 700 2130 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 2570 810 2620 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 1110 2900 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1780 40 1860 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1770 50 1870 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2020 40 2100 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2010 50 2110 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2260 40 2340 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2250 50 2350 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2500 40 2580 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2490 50 2590 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 280 0 330 300 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1000 0 1050 280 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1720 0 1770 300 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 2080 0 2130 280 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 2570 0 2620 320 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 0 0 2900 120 1 VSS
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2900 1230
string GDS_END 277316
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 249622
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
