magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 440 89 510
rect -31 -71 89 -1
use nmos_5p04310589983249_64x8m81  nmos_5p04310589983249_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 484
<< properties >>
string GDS_END 264518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 264268
<< end >>
