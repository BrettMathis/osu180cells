* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp9t3v3__tbuf_1 A Y EN
X0 Y a_49_56 a_44_70 VDD pmos_3p3 w=34 l=6
X1 a_49_56 EN VDD VDD pmos_3p3 w=34 l=6
X2 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X3 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X4 a_44_19 a_9_19 VSS VSS nmos_3p3 w=17 l=6
X5 a_44_70 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X6 Y EN a_44_19 VSS nmos_3p3 w=17 l=6
X7 a_49_56 EN VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
