magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 111 280 123
rect 28 94 33 111
rect 96 94 101 111
rect 130 94 135 111
rect 215 94 220 111
rect 32 73 80 79
rect 32 55 38 73
rect 43 62 69 68
rect 43 50 48 62
rect 64 53 69 62
rect 74 66 80 73
rect 117 72 199 78
rect 117 66 123 72
rect 74 60 123 66
rect 74 58 80 60
rect 117 58 123 60
rect 128 61 182 67
rect 128 53 134 61
rect 12 44 48 50
rect 53 42 59 52
rect 64 47 134 53
rect 141 42 147 55
rect 176 53 182 61
rect 193 58 199 72
rect 232 67 237 104
rect 247 94 252 111
rect 264 67 269 104
rect 232 66 238 67
rect 264 66 273 67
rect 232 60 241 66
rect 264 60 275 66
rect 232 59 238 60
rect 264 59 273 60
rect 174 47 184 53
rect 195 45 212 51
rect 195 42 201 45
rect 53 36 201 42
rect 28 12 33 28
rect 96 12 101 28
rect 130 12 135 28
rect 215 12 220 28
rect 232 19 237 59
rect 247 12 252 28
rect 264 19 269 59
rect 0 0 280 12
<< obsm1 >>
rect 11 89 16 104
rect 45 89 50 104
rect 62 94 68 104
rect 11 84 50 89
rect 113 89 118 104
rect 147 89 152 104
rect 113 84 152 89
rect 162 83 172 89
rect 156 47 166 53
rect 217 47 227 53
rect 10 19 16 29
rect 44 19 50 29
rect 62 19 68 29
rect 113 19 119 29
rect 146 19 152 29
rect 164 19 170 29
rect 249 47 259 53
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 177 112 187 118
rect 201 112 211 118
rect 225 112 235 118
rect 249 112 259 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 31 63 39 64
rect 30 57 40 63
rect 31 56 39 57
rect 12 43 22 51
rect 52 50 60 51
rect 51 44 61 50
rect 52 43 60 44
rect 232 66 240 67
rect 231 60 241 66
rect 232 59 240 60
rect 266 66 274 67
rect 265 60 275 66
rect 266 59 274 60
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< obsm2 >>
rect 62 103 68 104
rect 61 102 69 103
rect 60 96 257 102
rect 61 95 69 96
rect 75 53 81 96
rect 163 89 171 90
rect 162 83 225 89
rect 163 82 171 83
rect 157 53 165 54
rect 75 47 166 53
rect 10 28 16 29
rect 44 28 50 29
rect 62 28 68 29
rect 9 27 17 28
rect 43 27 51 28
rect 9 21 51 27
rect 9 20 17 21
rect 43 20 51 21
rect 61 27 69 28
rect 75 27 81 47
rect 157 46 165 47
rect 113 28 119 29
rect 146 28 152 29
rect 61 21 81 27
rect 112 27 120 28
rect 145 27 153 28
rect 163 27 171 28
rect 177 27 183 83
rect 219 54 225 83
rect 251 54 257 96
rect 218 46 226 54
rect 250 53 258 54
rect 249 47 259 53
rect 250 46 258 47
rect 219 45 225 46
rect 251 45 257 46
rect 112 21 153 27
rect 162 21 183 27
rect 61 20 69 21
rect 112 20 120 21
rect 145 20 153 21
rect 163 20 171 21
rect 10 19 16 20
rect 44 19 50 20
rect 62 19 68 20
rect 113 19 119 20
rect 146 19 152 20
<< labels >>
rlabel metal2 s 12 43 22 51 6 A
port 1 nsew signal input
rlabel metal1 s 12 44 48 50 6 A
port 1 nsew signal input
rlabel metal1 s 43 44 48 68 6 A
port 1 nsew signal input
rlabel metal1 s 64 47 69 68 6 A
port 1 nsew signal input
rlabel metal1 s 43 62 69 68 6 A
port 1 nsew signal input
rlabel metal1 s 64 47 134 53 6 A
port 1 nsew signal input
rlabel metal1 s 128 47 134 67 6 A
port 1 nsew signal input
rlabel metal1 s 176 47 182 67 6 A
port 1 nsew signal input
rlabel metal1 s 128 61 182 67 6 A
port 1 nsew signal input
rlabel metal1 s 174 47 184 53 6 A
port 1 nsew signal input
rlabel metal2 s 31 56 39 64 6 B
port 2 nsew signal input
rlabel metal2 s 30 57 40 63 6 B
port 2 nsew signal input
rlabel metal1 s 32 55 38 79 6 B
port 2 nsew signal input
rlabel metal1 s 74 58 80 79 6 B
port 2 nsew signal input
rlabel metal1 s 32 73 80 79 6 B
port 2 nsew signal input
rlabel metal1 s 74 60 123 66 6 B
port 2 nsew signal input
rlabel metal1 s 117 58 123 78 6 B
port 2 nsew signal input
rlabel metal1 s 193 58 199 78 6 B
port 2 nsew signal input
rlabel metal1 s 117 72 199 78 6 B
port 2 nsew signal input
rlabel metal2 s 52 43 60 51 6 CI
port 3 nsew signal input
rlabel metal2 s 51 44 61 50 6 CI
port 3 nsew signal input
rlabel metal1 s 53 36 59 52 6 CI
port 3 nsew signal input
rlabel metal1 s 141 36 147 55 6 CI
port 3 nsew signal input
rlabel metal1 s 53 36 201 42 6 CI
port 3 nsew signal input
rlabel metal1 s 195 36 201 51 6 CI
port 3 nsew signal input
rlabel metal1 s 195 45 212 51 6 CI
port 3 nsew signal input
rlabel metal2 s 266 59 274 67 6 CO
port 5 nsew signal output
rlabel metal2 s 265 60 275 66 6 CO
port 5 nsew signal output
rlabel metal1 s 264 19 269 104 6 CO
port 5 nsew signal output
rlabel metal1 s 264 59 273 67 6 CO
port 5 nsew signal output
rlabel metal1 s 264 60 275 66 6 CO
port 5 nsew signal output
rlabel metal2 s 232 59 240 67 6 S
port 4 nsew signal output
rlabel metal2 s 231 60 241 66 6 S
port 4 nsew signal output
rlabel metal1 s 232 19 237 104 6 S
port 4 nsew signal output
rlabel metal1 s 232 59 238 67 6 S
port 4 nsew signal output
rlabel metal1 s 232 60 241 66 6 S
port 4 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 178 111 186 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 177 112 187 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 202 111 210 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 201 112 211 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 226 111 234 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 225 112 235 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 250 111 258 119 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 249 112 259 118 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 28 94 33 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 96 94 101 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 130 94 135 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 215 94 220 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 247 94 252 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 0 111 280 123 6 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 28 0 33 28 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 96 0 101 28 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 130 0 135 28 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 215 0 220 28 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 247 0 252 28 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 280 12 6 VSS
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 280 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 26072
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 134
<< end >>
