magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 681 89 753
rect -31 -74 89 -1
use nmos_5p04310589983215_64x8m81  nmos_5p04310589983215_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 726
<< properties >>
string GDS_END 237692
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 237442
<< end >>
