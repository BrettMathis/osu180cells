* NGSPICE file created from gf180mcu_fd_ip_sram__sram128x8m8wm1.ext - technology: gf180mcuB

.subckt x018SRAM_cell1_cutPC_128x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_128x8m81 a_n36_52# a_444_n42# a_246_342# a_246_712# m3_n36_330#
+ a_36_n42# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt x018SRAM_cell1_dummy_128x8m81 a_n36_52# m2_90_n50# a_246_342# m2_390_n50#
+ a_246_712# m3_n36_330# w_n68_622# VSUBS
X0 a_126_298# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_246_712# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_126_298# a_36_206# a_246_712# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_126_298# a_36_206# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt new_dummyrow_unit_01_128x8m81 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# VSUBS 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50#
X018SRAM_cell1_dummy_128x8m81_10 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_11 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_12 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_13 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_14 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_15 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_0 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_1 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_3 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_2 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_4 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_5 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_6 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_7 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_8 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_9 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
.ends

.subckt new_dummyrow_unit_128x8m81 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# VSUBS 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50#
+ 018SRAM_strap1_128x8m81_1/w_n68_622#
X018SRAM_cell1_dummy_128x8m81_10 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_11 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_12 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_13 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_14 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_15 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_0 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_1 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_3 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_2 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_4 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_5 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_6 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_7 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_8 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_9 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_strap1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_128x8m81_1/a_n36_52# 018SRAM_strap1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
.ends

.subckt ldummy_128x4_128x8m81 018SRAM_cell1_dummy_128x8m81_29/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_5/a_246_342# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_5/a_246_712#
+ 018SRAM_cell1_dummy_128x8m81_17/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_18/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_19/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_13/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_6/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_1/w_n68_622# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_6/a_246_712#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_14/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_7/a_246_342# 018SRAM_cell1_dummy_128x8m81_20/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_9/w_n68_622# 018SRAM_cell1_cutPC_128x8m81_8/a_246_712#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_30/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_15/a_246_342# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_21/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_8/a_246_342#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_31/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_10/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_22/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_9/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_4/w_n68_622# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_11/m3_n36_330#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_12/m3_n36_330#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_13/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_3/w_n68_622#
+ 018SRAM_cell1_dummy_128x8m81_30/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_23/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_14/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_5/w_n68_622# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_31/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_15/m3_n36_330#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_24/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_0/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_6/w_n68_622# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_1/a_246_342# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_0/m3_n36_330# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_25/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_20/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_1/a_246_712# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_21/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_2/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_22/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_16/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_3/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_23/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_2/a_246_342# 018SRAM_cell1_dummy_128x8m81_26/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_4/m3_n36_330# 018SRAM_cell1_cutPC_128x8m81_8/w_n68_622#
+ 018SRAM_cell1_cutPC_128x8m81_9/a_246_712# 018SRAM_cell1_dummy_128x8m81_24/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_5/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_25/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_6/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_26/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_7/m3_n36_330#
+ VSS 018SRAM_cell1_dummy_128x8m81_17/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_27/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_27/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_8/m3_n36_330#
+ 018SRAM_cell1_cutPC_128x8m81_3/a_246_342# 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_28/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_3/a_246_712#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ 018SRAM_cell1_cutPC_128x8m81_9/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_29/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# 018SRAM_cell1_cutPC_128x8m81_11/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_18/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50#
+ 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_128x8m81_4/a_246_342# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_28/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_cell1_cutPC_128x8m81_4/a_246_712#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_19/m2_90_n50#
+ 018SRAM_cell1_cutPC_128x8m81_12/a_246_342# 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ VSUBS new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_16/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
X018SRAM_cell1_cutPC_128x8m81_2 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_2/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_9/a_246_712# 018SRAM_cell1_cutPC_128x8m81_2/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_9/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_128x8m81_1 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_128x8m81_1/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_128x8m81
X018SRAM_cell1_dummy_128x8m81_31 VSUBS 018SRAM_cell1_dummy_128x8m81_31/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_31/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_20 VSUBS 018SRAM_cell1_dummy_128x8m81_20/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_20/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_4 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_4/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_4/a_246_712# 018SRAM_cell1_cutPC_128x8m81_4/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_cutPC_128x8m81_3 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_3/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_3/a_246_712# 018SRAM_cell1_cutPC_128x8m81_3/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_3/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_21 VSUBS 018SRAM_cell1_dummy_128x8m81_21/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_21/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_10 VSUBS 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_5 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_5/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_5/a_246_712# 018SRAM_cell1_cutPC_128x8m81_5/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_22 VSUBS 018SRAM_cell1_dummy_128x8m81_22/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_22/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_11 VSUBS 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_6 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_6/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_6/a_246_712# 018SRAM_cell1_cutPC_128x8m81_6/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_6/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_23 VSUBS 018SRAM_cell1_dummy_128x8m81_23/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_23/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_12 VSUBS 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_7 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_7/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_8/a_246_712# 018SRAM_cell1_cutPC_128x8m81_7/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_8/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_24 VSUBS 018SRAM_cell1_dummy_128x8m81_24/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_24/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_13 VSUBS 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_8 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_8/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_8/a_246_712# 018SRAM_cell1_cutPC_128x8m81_8/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_8/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
Xnew_dummyrow_unit_01_128x8m81_0 new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ VSUBS new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# VSUBS
+ 018SRAM_cell1_128x8m81_1/w_n68_622# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# new_dummyrow_unit_01_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50#
+ new_dummyrow_unit_01_128x8m81
X018SRAM_cell1_dummy_128x8m81_25 VSUBS 018SRAM_cell1_dummy_128x8m81_25/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_25/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_14 VSUBS 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_9 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_9/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_9/a_246_712# 018SRAM_cell1_cutPC_128x8m81_9/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_9/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_26 VSUBS 018SRAM_cell1_dummy_128x8m81_26/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_26/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_15 VSUBS 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_28 VSUBS 018SRAM_cell1_dummy_128x8m81_28/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_28/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_27 VSUBS 018SRAM_cell1_dummy_128x8m81_27/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_27/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_17 VSUBS 018SRAM_cell1_dummy_128x8m81_17/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_17/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_16 VSUBS 018SRAM_cell1_dummy_128x8m81_16/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_16/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_29 VSUBS 018SRAM_cell1_dummy_128x8m81_29/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_29/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_18 VSUBS 018SRAM_cell1_dummy_128x8m81_18/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_18/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_19 VSUBS 018SRAM_cell1_dummy_128x8m81_19/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_19/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_10 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_10/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_1/a_246_712# 018SRAM_cell1_cutPC_128x8m81_10/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_cutPC_128x8m81_11 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_11/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_6/a_246_712# 018SRAM_cell1_cutPC_128x8m81_11/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_6/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_cutPC_128x8m81_12 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_12/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_3/a_246_712# 018SRAM_cell1_cutPC_128x8m81_12/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_3/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_cutPC_128x8m81_13 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_13/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_5/a_246_712# 018SRAM_cell1_cutPC_128x8m81_13/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_5/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_cutPC_128x8m81_14 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_14/a_246_342#
+ 018SRAM_cell1_128x8m81_0/w_n68_622# 018SRAM_cell1_cutPC_128x8m81_14/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_0 VSUBS 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_15 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_15/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_4/a_246_712# 018SRAM_cell1_cutPC_128x8m81_15/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_4/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_1 VSUBS 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_3 VSUBS 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_2 VSUBS 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
Xnew_dummyrow_unit_128x8m81_0 new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ VSUBS new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ VSUBS new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ new_dummyrow_unit_128x8m81
X018SRAM_cell1_dummy_128x8m81_4 VSUBS 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_5 VSUBS 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_6 VSUBS 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_7 VSUBS 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_8 VSUBS 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_0 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_0/a_246_342#
+ 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_cutPC_128x8m81_0/m3_n36_330# 018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_dummy_128x8m81_9 VSUBS 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50# VSUBS
+ 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_cutPC_128x8m81_1 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_cutPC_128x8m81_1/a_246_342#
+ 018SRAM_cell1_cutPC_128x8m81_1/a_246_712# 018SRAM_cell1_cutPC_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_cutPC_128x8m81_1/w_n68_622# VSUBS
+ x018SRAM_cell1_cutPC_128x8m81
X018SRAM_cell1_128x8m81_0 VSUBS 018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS
+ x018SRAM_cell1_128x8m81
X018SRAM_cell1_dummy_128x8m81_30 VSUBS 018SRAM_cell1_dummy_128x8m81_30/m2_90_n50#
+ VSUBS 018SRAM_cell1_dummy_128x8m81_30/m2_390_n50# 018SRAM_cell1_128x8m81_0/w_n68_622#
+ VSUBS 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_dummy_128x8m81
.ends

.subckt x018SRAM_cell1_2x_128x8m81 018SRAM_cell1_128x8m81_0/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_128x8m81_0/a_246_342#
+ 018SRAM_cell1_128x8m81_0/a_246_712# 018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_128x8m81_1/a_246_342#
+ 018SRAM_cell1_128x8m81_1/a_246_712# 018SRAM_cell1_128x8m81_0/m3_n36_330# 018SRAM_cell1_128x8m81_1/m3_n36_330#
+ VSUBS 018SRAM_cell1_128x8m81_1/a_36_n42#
X018SRAM_cell1_128x8m81_1 018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_128x8m81_1/a_246_342# 018SRAM_cell1_128x8m81_1/a_246_712# 018SRAM_cell1_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_1/w_n68_622# VSUBS x018SRAM_cell1_128x8m81
X018SRAM_cell1_128x8m81_0 018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_128x8m81_0/a_246_342# 018SRAM_cell1_128x8m81_0/a_246_712# 018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_0/w_n68_622# VSUBS x018SRAM_cell1_128x8m81
.ends

.subckt Cell_array8x8x2_128x8m81 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ VSUBS
X018SRAM_cell1_2x_128x8m81_190 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_0 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_191 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_180 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_1 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_181 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_170 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_192 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_2 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_160 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_182 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_171 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_193 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_3 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_183 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_172 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_161 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_150 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_194 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_4 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_140 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_184 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_162 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_151 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_173 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_195 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_5 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_152 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_141 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_185 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_130 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_174 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_163 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_196 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_6 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_153 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_142 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_120 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_186 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_164 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_131 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_175 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_197 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_7 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_187 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_143 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_132 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_176 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_154 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_165 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_121 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_110 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_198 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_8 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_188 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_144 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_100 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_155 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_133 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_177 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_166 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_122 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_111 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_199 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_9 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_189 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_145 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_156 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_101 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_167 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_134 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_112 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_178 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_123 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_146 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_157 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_102 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_179 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_168 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_135 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_113 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_124 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_169 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_103 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_147 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_136 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_114 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_158 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_125 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_148 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_137 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_159 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_115 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_126 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_104 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_149 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_138 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_116 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_127 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_105 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_139 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_117 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_128 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_106 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_129 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_118 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_107 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_119 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_186/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_108 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_90 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_109 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_0/a_n36_52# 018SRAM_strap1_2x_128x8m81_9/018SRAM_strap1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_91 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_80 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_70 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_92 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_81 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_60 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_71 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_93 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_82 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_250 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_50 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_61 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_72 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_94 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_83 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_251 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_240 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_51 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_62 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_73 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_40 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_95 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_84 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_252 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_230 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_241 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_96 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_30 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_52 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_63 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_74 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_41 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_85 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_231 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_220 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_253 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_242 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_97 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_31 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_20 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_53 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_75 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_64 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_42 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_86 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_221 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_254 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_232 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_210 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_243 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_98 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_32 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_54 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_76 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_65 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_21 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_10 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_43 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_87 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_200 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_233 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_222 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_255 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_211 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_244 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_99 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_88 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_55 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_77 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_66 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_22 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_11 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_33 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_44 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_201 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_223 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_234 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_212 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_245 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_56 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_78 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_67 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_23 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_45 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_34 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_89 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_12 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_202 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_235 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_224 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_213 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_246 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_57 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_79 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_68 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_46 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_35 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_13 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_24 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_203 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_225 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_236 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_214 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_247 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_58 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_69 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_25 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_14 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_47 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_36 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_204 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_237 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_248 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_226 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_215 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_26 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_59 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_15 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_37 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_48 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_205 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_227 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_216 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_249 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_238 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_27 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_16 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_49 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_38 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_206 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_239 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_217 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_228 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_28 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_17 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_39 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_207 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_229 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_218 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_29 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_18 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_8/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_219 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_255/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_208 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_19 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_209 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42# VSUBS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_0/a_n36_52# 018SRAM_cell1_2x_128x8m81_247/018SRAM_cell1_128x8m81_1/a_n36_52#
+ VSUBS 018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42# x018SRAM_cell1_2x_128x8m81
.ends

.subckt col_128a_128x8m81 WL[3] WL[2] WL[1] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+ WL[6] WL[5] WL[4] WL[15] WL[14] WL[13] WL[0] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSUBS Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
XCell_array8x8x2_128x8m81_0 Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_96/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[2] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_93/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_89/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_24/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[15] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_19/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[3] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_41/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_82/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_16/018SRAM_cell1_128x8m81_1/a_36_n42#
+ WL[4] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_43/018SRAM_cell1_128x8m81_1/a_36_n42#
+ WL[6] WL[8] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_97/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_95/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_94/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_36_n42#
+ WL[14] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_98/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_81/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[0] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_85/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_83/018SRAM_cell1_128x8m81_1/a_36_n42#
+ WL[12] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_42/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_47/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[13] WL[11] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_45/018SRAM_cell1_128x8m81_1/a_444_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[1] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_25/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_36_n42#
+ WL[9] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_12/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[10] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[5] WL[7] Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_44/018SRAM_cell1_128x8m81_1/a_36_n42#
+ Cell_array8x8x2_128x8m81_0/018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ VSUBS Cell_array8x8x2_128x8m81
.ends

.subckt nmos_5p04310590548716_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46552108_128x8m81 a_1089_n74# a_865_n74# a_641_n74# a_n31_n74# nmos_5p04310590548716_128x8m81_0/S
+ a_1537_n74# a_1313_n74# nmos_5p04310590548716_128x8m81_0/D a_417_n74# a_193_n74#
+ VSUBS
Xnmos_5p04310590548716_128x8m81_0 nmos_5p04310590548716_128x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590548716_128x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310590548716_128x8m81
.ends

.subckt pmos_5p04310590548720_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46897196_128x8m81 a_193_n74# pmos_5p04310590548720_128x8m81_0/S
+ w_n286_n142# a_n31_n74# pmos_5p04310590548720_128x8m81_0/D
Xpmos_5p04310590548720_128x8m81_0 w_n286_n142# pmos_5p04310590548720_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548720_128x8m81_0/S a_193_n74# pmos_5p04310590548720_128x8m81
.ends

.subckt nmos_5p04310590548715_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.41u l=0.6u
.ends

.subckt nmos_1p2$$46553132_128x8m81 nmos_5p04310590548715_128x8m81_0/D nmos_5p04310590548715_128x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310590548715_128x8m81_0 nmos_5p04310590548715_128x8m81_0/D a_n31_n74# nmos_5p04310590548715_128x8m81_0/S
+ VSUBS nmos_5p04310590548715_128x8m81
.ends

.subckt nmos_5p04310590548717_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
X7 S a_1568_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_1p2$$46550060_128x8m81 a_1537_n74# a_1313_n74# nmos_5p04310590548717_128x8m81_0/S
+ a_193_n74# nmos_5p04310590548717_128x8m81_0/D a_1089_n74# a_865_n74# a_n31_n74#
+ a_641_n74# a_417_n74# VSUBS
Xnmos_5p04310590548717_128x8m81_0 nmos_5p04310590548717_128x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590548717_128x8m81_0/S a_417_n74# a_193_n74# a_1537_n74#
+ a_1313_n74# a_1089_n74# VSUBS nmos_5p04310590548717_128x8m81
.ends

.subckt pmos_5p04310590548714_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46285868_128x8m81 pmos_5p04310590548714_128x8m81_0/S w_n286_n142#
+ a_n31_n73# pmos_5p04310590548714_128x8m81_0/D
Xpmos_5p04310590548714_128x8m81_0 w_n286_n142# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt pmos_5p04310590548713_128x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46286892_128x8m81 a_193_n73# a_n31_n73# a_417_n73# pmos_5p04310590548713_128x8m81_0/S
+ w_n286_n142# pmos_5p04310590548713_128x8m81_0/D
Xpmos_5p04310590548713_128x8m81_0 w_n286_n142# pmos_5p04310590548713_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548713_128x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310590548713_128x8m81
.ends

.subckt nmos_5p04310590548710_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$46551084_128x8m81 nmos_5p04310590548710_128x8m81_0/D a_n31_n73#
+ nmos_5p04310590548710_128x8m81_0/S VSUBS
Xnmos_5p04310590548710_128x8m81_0 nmos_5p04310590548710_128x8m81_0/D a_n31_n73# nmos_5p04310590548710_128x8m81_0/S
+ VSUBS nmos_5p04310590548710_128x8m81
.ends

.subckt pmos_5p04310590548719_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46898220_128x8m81 pmos_5p04310590548719_128x8m81_0/S w_n286_n142#
+ pmos_5p04310590548719_128x8m81_0/D a_n31_n74#
Xpmos_5p04310590548719_128x8m81_0 w_n286_n142# pmos_5p04310590548719_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548719_128x8m81_0/S pmos_5p04310590548719_128x8m81
.ends

.subckt pmos_5p04310590548721_128x8m81 w_n208_n120# D a_0_n44# a_672_n44# S a_448_n44#
+ a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.91u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=0.91u l=0.6u
.ends

.subckt pmos_1p2$$46896172_128x8m81 pmos_5p04310590548721_128x8m81_0/S a_668_n74#
+ a_193_n74# w_n286_n142# pmos_5p04310590548721_128x8m81_0/D a_n31_n74# a_417_n74#
Xpmos_5p04310590548721_128x8m81_0 w_n286_n142# pmos_5p04310590548721_128x8m81_0/D
+ a_n31_n74# a_668_n74# pmos_5p04310590548721_128x8m81_0/S a_417_n74# a_193_n74# pmos_5p04310590548721_128x8m81
.ends

.subckt nmos_5p04310590548712_128x8m81 D a_0_n44# a_672_n44# S a_448_n44# a_224_n44#
+ VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45107244_128x8m81 a_193_n73# nmos_5p04310590548712_128x8m81_0/S
+ a_n31_n73# a_641_n73# a_417_n73# nmos_5p04310590548712_128x8m81_0/D VSUBS
Xnmos_5p04310590548712_128x8m81_0 nmos_5p04310590548712_128x8m81_0/D a_n31_n73# a_641_n73#
+ nmos_5p04310590548712_128x8m81_0/S a_417_n73# a_193_n73# VSUBS nmos_5p04310590548712_128x8m81
.ends

.subckt pmos_5p04310590548718_128x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46549036_128x8m81 a_193_n74# pmos_5p04310590548718_128x8m81_0/S
+ w_n286_n142# a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# a_417_n74# pmos_5p04310590548718_128x8m81_0/D
Xpmos_5p04310590548718_128x8m81_0 w_n286_n142# pmos_5p04310590548718_128x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590548718_128x8m81_0/S a_417_n74# a_193_n74#
+ a_1089_n74# pmos_5p04310590548718_128x8m81
.ends

.subckt sa_128x8m81 qp wep se pcb vss d
Xnmos_1p2$$46552108_128x8m81_0 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ nmos_1p2$$46552108_128x8m81_0/nmos_5p04310590548716_128x8m81_0/D pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S vss nmos_1p2$$46552108_128x8m81
Xpmos_1p2$$46897196_128x8m81_1 se d d se pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46897196_128x8m81
Xpmos_1p2$$46897196_128x8m81_2 se d d se pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46897196_128x8m81
Xpmos_1p2$$46897196_128x8m81_3 se d d se pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46897196_128x8m81
Xnmos_1p2$$46553132_128x8m81_0 vss pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ vss vss nmos_1p2$$46553132_128x8m81
Xnmos_1p2$$46550060_128x8m81_0 se se vss se nmos_1p2$$46552108_128x8m81_0/nmos_5p04310590548716_128x8m81_0/D
+ se se se se se vss nmos_1p2$$46550060_128x8m81
Xnmos_1p2$$46553132_128x8m81_1 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ vss vss vss nmos_1p2$$46553132_128x8m81
Xpmos_1p2$$46285868_128x8m81_0 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ d pcb pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46285868_128x8m81
Xpmos_1p2$$46286892_128x8m81_0 pcb pcb pcb d d d pmos_1p2$$46286892_128x8m81
Xnmos_1p2$$46551084_128x8m81_0 vss pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ qp vss nmos_1p2$$46551084_128x8m81
Xpmos_1p2$$46898220_128x8m81_0 d d pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ d pmos_1p2$$46898220_128x8m81
Xpmos_1p2$$46898220_128x8m81_1 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ d d d pmos_1p2$$46898220_128x8m81
Xpmos_1p2$$46896172_128x8m81_0 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ d d pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46896172_128x8m81
Xnmos_1p2$$45107244_128x8m81_0 qp qp pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ qp qp vss vss nmos_1p2$$45107244_128x8m81
Xpmos_1p2$$46549036_128x8m81_0 pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ d d pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S qp qp qp pmos_1p2$$46549036_128x8m81
Xpmos_1p2$$46897196_128x8m81_0 se d d se pmos_1p2$$46898220_128x8m81_1/pmos_5p04310590548719_128x8m81_0/S
+ pmos_1p2$$46897196_128x8m81
.ends

.subckt nmos_5p0431059054875_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=11.34u l=0.6u
.ends

.subckt nmos_1p2$$46883884_128x8m81 nmos_5p0431059054875_128x8m81_0/S nmos_5p0431059054875_128x8m81_0/D
+ a_n31_n73# VSUBS
Xnmos_5p0431059054875_128x8m81_0 nmos_5p0431059054875_128x8m81_0/D a_n31_n73# nmos_5p0431059054875_128x8m81_0/S
+ VSUBS nmos_5p0431059054875_128x8m81
.ends

.subckt pmos_5p0431059054876_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt pmos_1p2$$46885932_128x8m81 a_193_n73# pmos_5p0431059054876_128x8m81_0/S a_n31_n74#
+ w_n286_n141# pmos_5p0431059054876_128x8m81_0/D
Xpmos_5p0431059054876_128x8m81_0 w_n286_n141# pmos_5p0431059054876_128x8m81_0/D a_n31_n74#
+ pmos_5p0431059054876_128x8m81_0/S a_193_n73# pmos_5p0431059054876_128x8m81
.ends

.subckt nmos_5p0431059054878_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$46563372_128x8m81 nmos_5p0431059054878_128x8m81_0/D nmos_5p0431059054878_128x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p0431059054878_128x8m81_0 nmos_5p0431059054878_128x8m81_0/D a_n31_n74# nmos_5p0431059054878_128x8m81_0/S
+ VSUBS nmos_5p0431059054878_128x8m81
.ends

.subckt pmos_5p0431059054873_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt pmos_1p2$$46273580_128x8m81 pmos_5p0431059054873_128x8m81_0/S pmos_5p0431059054873_128x8m81_0/D
+ a_193_n74# a_n31_n74# w_n286_n142#
Xpmos_5p0431059054873_128x8m81_0 w_n286_n142# pmos_5p0431059054873_128x8m81_0/D a_n31_n74#
+ pmos_5p0431059054873_128x8m81_0/S a_193_n74# pmos_5p0431059054873_128x8m81
.ends

.subckt pmos_5p0431059054874_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.61u l=0.6u
.ends

.subckt pmos_1p2$$46887980_128x8m81 pmos_5p0431059054874_128x8m81_0/D a_n31_n74# w_n286_n142#
+ pmos_5p0431059054874_128x8m81_0/S
Xpmos_5p0431059054874_128x8m81_0 w_n286_n142# pmos_5p0431059054874_128x8m81_0/D a_n31_n74#
+ pmos_5p0431059054874_128x8m81_0/S pmos_5p0431059054874_128x8m81
.ends

.subckt nmos_5p04310590548711_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.96u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_5p0431059054877_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=13.61u l=0.6u
.ends

.subckt nmos_1p2$$46884908_128x8m81 nmos_5p0431059054877_128x8m81_0/D nmos_5p0431059054877_128x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p0431059054877_128x8m81_0 nmos_5p0431059054877_128x8m81_0/D a_n31_n74# nmos_5p0431059054877_128x8m81_0/S
+ VSUBS nmos_5p0431059054877_128x8m81
.ends

.subckt pmos_5p0431059054871_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.81u l=0.6u
.ends

.subckt pmos_1p2$$46889004_128x8m81 pmos_5p0431059054871_128x8m81_0/S w_n286_n142#
+ a_n31_n74# pmos_5p0431059054871_128x8m81_0/D
Xpmos_5p0431059054871_128x8m81_0 w_n286_n142# pmos_5p0431059054871_128x8m81_0/D a_n31_n74#
+ pmos_5p0431059054871_128x8m81_0/S pmos_5p0431059054871_128x8m81
.ends

.subckt pmos_5p0431059054879_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt din_128x8m81 d db datain wep men m1_164_8068# vss pmos_5p0431059054871_128x8m81_0/D
+ vdd
Xnmos_1p2$$46883884_128x8m81_0 db pmos_5p0431059054879_128x8m81_0/S wep vss nmos_1p2$$46883884_128x8m81
Xnmos_1p2$$46883884_128x8m81_1 pmos_5p0431059054879_128x8m81_0/S vss pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ vss nmos_1p2$$46883884_128x8m81
Xnmos_1p2$$46883884_128x8m81_2 d pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ wep vss nmos_1p2$$46883884_128x8m81
Xpmos_1p2$$46885932_128x8m81_0 pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ pmos_5p0431059054876_128x8m81_0/S men vdd nmos_5p04310590548711_128x8m81_1/D pmos_1p2$$46885932_128x8m81
Xnmos_1p2$$46563372_128x8m81_0 pmos_5p0431059054876_128x8m81_0/S vss pmos_5p0431059054871_128x8m81_0/S
+ vss nmos_1p2$$46563372_128x8m81
Xnmos_1p2$$46563372_128x8m81_1 pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ vss men vss nmos_1p2$$46563372_128x8m81
Xpmos_1p2$$46273580_128x8m81_0 vdd pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ men men vdd pmos_1p2$$46273580_128x8m81
Xpmos_1p2$$46273580_128x8m81_1 vdd pmos_5p0431059054876_128x8m81_0/S pmos_5p0431059054871_128x8m81_0/S
+ pmos_5p0431059054871_128x8m81_0/S vdd pmos_1p2$$46273580_128x8m81
Xpmos_5p0431059054876_128x8m81_0 vdd vdd datain pmos_5p0431059054876_128x8m81_0/S
+ pmos_5p0431059054876_128x8m81_0/S pmos_5p0431059054876_128x8m81
Xpmos_1p2$$46887980_128x8m81_0 pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ pmos_5p0431059054871_128x8m81_0/S vdd vdd pmos_1p2$$46887980_128x8m81
Xnmos_5p04310590548711_128x8m81_0 vss datain pmos_5p0431059054876_128x8m81_0/S pmos_5p0431059054876_128x8m81_0/S
+ vss nmos_5p04310590548711_128x8m81
Xnmos_5p04310590548711_128x8m81_1 nmos_5p04310590548711_128x8m81_1/D pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ pmos_5p0431059054876_128x8m81_0/S men vss nmos_5p04310590548711_128x8m81
Xnmos_5p04310590548710_128x8m81_0 vss nmos_5p04310590548711_128x8m81_1/D pmos_5p0431059054871_128x8m81_0/S
+ vss nmos_5p04310590548710_128x8m81
Xnmos_1p2$$46884908_128x8m81_0 pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ vss pmos_5p0431059054871_128x8m81_0/S vss nmos_1p2$$46884908_128x8m81
Xpmos_1p2$$46889004_128x8m81_0 d vdd a_500_6666# pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ pmos_1p2$$46889004_128x8m81
Xpmos_5p0431059054871_128x8m81_0 vdd pmos_5p0431059054871_128x8m81_0/D nmos_5p04310590548711_128x8m81_1/D
+ pmos_5p0431059054871_128x8m81_0/S pmos_5p0431059054871_128x8m81
Xpmos_1p2$$46889004_128x8m81_1 db vdd a_500_6666# pmos_5p0431059054879_128x8m81_0/S
+ pmos_1p2$$46889004_128x8m81
Xpmos_5p0431059054879_128x8m81_0 vdd vdd pmos_1p2$$46889004_128x8m81_0/pmos_5p0431059054871_128x8m81_0/D
+ pmos_5p0431059054879_128x8m81_0/S pmos_5p0431059054879_128x8m81
X0 vdd wep a_500_6666# vdd pmos_3p3 w=1.485u l=0.6u
X1 a_500_6666# wep vss vss nmos_3p3 w=1.14u l=0.6u
X2 a_500_6666# wep vdd vdd pmos_3p3 w=1.485u l=0.6u
.ends

.subckt pmos_5p04310590548730_128x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=2.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=2.72u l=0.6u
.ends

.subckt pmos_1p2$$45095980_128x8m81 a_193_n74# pmos_5p04310590548730_128x8m81_0/D
+ a_1089_n74# a_865_n74# a_n31_n74# a_641_n74# a_1985_n74# a_1761_n74# a_417_n74#
+ w_n286_n142# a_1537_n74# a_1313_n74# pmos_5p04310590548730_128x8m81_0/S
Xpmos_5p04310590548730_128x8m81_0 w_n286_n142# pmos_5p04310590548730_128x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590548730_128x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310590548730_128x8m81
.ends

.subckt pmos_5p04310590548727_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310590548724_128x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_1p2$$46282796_128x8m81 pmos_5p04310590548724_128x8m81_0/D a_193_n74#
+ a_865_n74# a_n31_n74# a_641_n74# a_417_n74# w_n286_n142# pmos_5p04310590548724_128x8m81_0/S
Xpmos_5p04310590548724_128x8m81_0 w_n286_n142# pmos_5p04310590548724_128x8m81_0/D
+ a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590548724_128x8m81_0/S a_417_n74# a_193_n74#
+ pmos_5p04310590548724_128x8m81
.ends

.subckt nmos_5p04310590548734_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.44u l=0.6u
.ends

.subckt nmos_5p04310590548736_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_1p2$$45101100_128x8m81 nmos_5p04310590548736_128x8m81_0/S a_193_n74#
+ a_865_n74# a_n31_n74# nmos_5p04310590548736_128x8m81_0/D a_641_n74# a_417_n74# VSUBS
Xnmos_5p04310590548736_128x8m81_0 nmos_5p04310590548736_128x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590548736_128x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310590548736_128x8m81
.ends

.subckt nmos_5p04310590548733_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310590548723_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.6u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=0.6u
.ends

.subckt nmos_5p04310590548732_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_5p04310590548726_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$45102124_128x8m81 a_1313_n74# nmos_5p04310590548726_128x8m81_0/D
+ a_193_n74# a_1089_n74# nmos_5p04310590548726_128x8m81_0/S a_865_n74# a_n31_n74#
+ a_641_n74# a_417_n74# VSUBS
Xnmos_5p04310590548726_128x8m81_0 nmos_5p04310590548726_128x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590548726_128x8m81_0/S a_417_n74# a_193_n74# a_1313_n74#
+ a_1089_n74# VSUBS nmos_5p04310590548726_128x8m81
.ends

.subckt nmos_5p04310590548737_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.86u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.86u l=0.6u
.ends

.subckt nmos_1p2$$45103148_128x8m81 a_865_n73# nmos_5p04310590548737_128x8m81_0/D
+ a_193_n74# a_1089_n74# a_n31_n74# a_641_n74# a_417_n74# nmos_5p04310590548737_128x8m81_0/S
+ VSUBS
Xnmos_5p04310590548737_128x8m81_0 nmos_5p04310590548737_128x8m81_0/D a_n31_n74# a_865_n73#
+ a_641_n74# nmos_5p04310590548737_128x8m81_0/S a_417_n74# a_193_n74# a_1089_n74#
+ VSUBS nmos_5p04310590548737_128x8m81
.ends

.subckt nmos_5p04310590548729_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.61u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.61u l=0.6u
.ends

.subckt nmos_1p2$$45100076_128x8m81 nmos_5p04310590548729_128x8m81_0/S a_193_n74#
+ nmos_5p04310590548729_128x8m81_0/D a_n31_n74# VSUBS
Xnmos_5p04310590548729_128x8m81_0 nmos_5p04310590548729_128x8m81_0/D a_n31_n74# nmos_5p04310590548729_128x8m81_0/S
+ a_193_n74# VSUBS nmos_5p04310590548729_128x8m81
.ends

.subckt pmos_5p04310590548722_128x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.09u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.09u l=0.6u
.ends

.subckt pmos_1p2$$46283820_128x8m81 a_641_n74# a_1985_n74# a_1761_n74# a_417_n74#
+ pmos_5p04310590548722_128x8m81_0/S a_1537_n74# a_1313_n74# pmos_5p04310590548722_128x8m81_0/D
+ w_n286_n142# a_193_n74# a_1089_n74# a_865_n74# a_n31_n74#
Xpmos_5p04310590548722_128x8m81_0 w_n286_n142# pmos_5p04310590548722_128x8m81_0/D
+ a_1985_n74# a_n31_n74# a_865_n74# a_641_n74# pmos_5p04310590548722_128x8m81_0/S
+ a_1761_n74# a_417_n74# a_193_n74# a_1537_n74# a_1313_n74# a_1089_n74# pmos_5p04310590548722_128x8m81
.ends

.subckt nmos_5p04310590548728_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310590548731_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.41u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.41u l=0.6u
.ends

.subckt pmos_1p2$$46287916_128x8m81 pmos_5p04310590548731_128x8m81_0/D a_193_n74#
+ w_n286_n142# pmos_5p04310590548731_128x8m81_0/S a_n31_n74#
Xpmos_5p04310590548731_128x8m81_0 w_n286_n142# pmos_5p04310590548731_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548731_128x8m81_0/S a_193_n74# pmos_5p04310590548731_128x8m81
.ends

.subckt pmos_5p04310590548735_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$46284844_128x8m81 a_n31_n74# pmos_5p04310590548735_128x8m81_0/D
+ w_n286_n142# a_193_n74# pmos_5p04310590548735_128x8m81_0/S
Xpmos_5p04310590548735_128x8m81_0 w_n286_n142# pmos_5p04310590548735_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548735_128x8m81_0/S a_193_n74# pmos_5p04310590548735_128x8m81
.ends

.subckt pmos_5p04310590548738_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310590548725_128x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$46281772_128x8m81 a_n31_n73# pmos_5p04310590548725_128x8m81_0/S
+ w_n286_n142# a_193_n73# a_417_n73# pmos_5p04310590548725_128x8m81_0/D
Xpmos_5p04310590548725_128x8m81_0 w_n286_n142# pmos_5p04310590548725_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548725_128x8m81_0/S a_417_n73# a_193_n73# pmos_5p04310590548725_128x8m81
.ends

.subckt sacntl_2_128x8m81 men pcb a_4718_983# nmos_5p04310590548723_128x8m81_1/D pmos_5p04310590548727_128x8m81_2/S
+ se a_4560_1922# a_2796_670# pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_5p04310590548727_128x8m81_1/S vss vdd
Xpmos_1p2$$45095980_128x8m81_0 nmos_5p04310590548728_128x8m81_1/S se nmos_5p04310590548728_128x8m81_1/S
+ nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S
+ nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S
+ vdd nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S vdd pmos_1p2$$45095980_128x8m81
Xpmos_5p04310590548727_128x8m81_0 vdd vdd a_2796_670# pmos_5p04310590548727_128x8m81_0/S
+ pmos_5p04310590548727_128x8m81_0/S pmos_5p04310590548727_128x8m81
Xpmos_5p04310590548727_128x8m81_1 vdd vdd pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_5p04310590548727_128x8m81_1/S vss pmos_5p04310590548727_128x8m81
Xpmos_5p04310590548727_128x8m81_2 vdd vdd pmos_5p04310590548727_128x8m81_1/S pmos_5p04310590548727_128x8m81_2/S
+ pmos_5p04310590548727_128x8m81_2/S pmos_5p04310590548727_128x8m81
Xpmos_1p2$$46285868_128x8m81_0 nmos_5p04310590548728_128x8m81_1/S vdd pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ vdd pmos_1p2$$46285868_128x8m81
Xpmos_1p2$$46282796_128x8m81_0 pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ men men men men men vdd vdd pmos_1p2$$46282796_128x8m81
Xnmos_5p04310590548734_128x8m81_0 nmos_5p04310590548734_128x8m81_0/D pmos_5p04310590548727_128x8m81_1/S
+ vss vss nmos_5p04310590548734_128x8m81
Xnmos_1p2$$45101100_128x8m81_0 vss men men men pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ men men vss nmos_1p2$$45101100_128x8m81
Xpmos_1p2$$46286892_128x8m81_0 nmos_5p04310590548732_128x8m81_0/D nmos_5p04310590548732_128x8m81_0/D
+ nmos_5p04310590548732_128x8m81_0/D vdd vdd nmos_5p04310590548728_128x8m81_1/S pmos_1p2$$46286892_128x8m81
Xnmos_5p04310590548733_128x8m81_0 vss pmos_5p04310590548727_128x8m81_0/S pmos_5p04310590548738_128x8m81_0/S
+ vss nmos_5p04310590548733_128x8m81
Xnmos_5p04310590548723_128x8m81_0 vss a_2796_670# pmos_5p04310590548727_128x8m81_0/S
+ pmos_5p04310590548727_128x8m81_0/S vss nmos_5p04310590548723_128x8m81
Xnmos_5p04310590548723_128x8m81_1 nmos_5p04310590548723_128x8m81_1/D pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_5p04310590548727_128x8m81_1/S vss vss nmos_5p04310590548723_128x8m81
Xnmos_5p04310590548723_128x8m81_2 vss pmos_5p04310590548727_128x8m81_1/S pmos_5p04310590548727_128x8m81_2/S
+ pmos_5p04310590548727_128x8m81_2/S vss nmos_5p04310590548723_128x8m81
Xnmos_5p04310590548732_128x8m81_0 nmos_5p04310590548732_128x8m81_0/D nmos_5p04310590548734_128x8m81_0/D
+ vss nmos_5p04310590548734_128x8m81_0/D vss nmos_5p04310590548732_128x8m81
Xnmos_5p04310590548712_128x8m81_0 se nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S
+ vss nmos_5p04310590548728_128x8m81_1/S nmos_5p04310590548728_128x8m81_1/S vss nmos_5p04310590548712_128x8m81
Xnmos_1p2$$45102124_128x8m81_0 pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pcb pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ vss pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ vss nmos_1p2$$45102124_128x8m81
Xnmos_1p2$$45103148_128x8m81_0 nmos_5p04310590548734_128x8m81_0/D pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S
+ nmos_5p04310590548734_128x8m81_0/D pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D nmos_5p04310590548728_128x8m81_1/S
+ nmos_5p04310590548728_128x8m81_1/S vss vss nmos_1p2$$45103148_128x8m81
Xnmos_1p2$$45100076_128x8m81_0 vss pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S
+ vss nmos_1p2$$45100076_128x8m81
Xpmos_1p2$$46283820_128x8m81_0 pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S vdd pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pcb vdd pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S pmos_1p2$$46283820_128x8m81
Xnmos_5p04310590548728_128x8m81_0 nmos_5p04310590548728_128x8m81_1/D nmos_5p04310590548732_128x8m81_0/D
+ nmos_5p04310590548732_128x8m81_0/D nmos_5p04310590548732_128x8m81_0/D vss nmos_5p04310590548732_128x8m81_0/D
+ nmos_5p04310590548732_128x8m81_0/D vss nmos_5p04310590548728_128x8m81
Xnmos_5p04310590548728_128x8m81_1 nmos_5p04310590548728_128x8m81_1/D pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ nmos_5p04310590548728_128x8m81_1/S pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D vss nmos_5p04310590548728_128x8m81
Xpmos_1p2$$46287916_128x8m81_0 nmos_5p04310590548732_128x8m81_0/D nmos_5p04310590548734_128x8m81_0/D
+ vdd vdd nmos_5p04310590548734_128x8m81_0/D pmos_1p2$$46287916_128x8m81
Xpmos_1p2$$46284844_128x8m81_0 pmos_5p04310590548727_128x8m81_1/S nmos_5p04310590548734_128x8m81_0/D
+ vdd pmos_5p04310590548727_128x8m81_1/S vdd pmos_1p2$$46284844_128x8m81
Xpmos_5p04310590548738_128x8m81_0 vdd vdd pmos_5p04310590548727_128x8m81_0/S pmos_5p04310590548738_128x8m81_0/S
+ pmos_5p04310590548738_128x8m81
Xpmos_1p2$$46281772_128x8m81_0 pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_0/pmos_5p04310590548725_128x8m81_0/S vdd pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S
+ pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S vdd pmos_1p2$$46281772_128x8m81
Xpmos_1p2$$46281772_128x8m81_1 pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ pmos_1p2$$46281772_128x8m81_1/pmos_5p04310590548725_128x8m81_0/S vdd nmos_5p04310590548734_128x8m81_0/D
+ nmos_5p04310590548728_128x8m81_1/S vdd pmos_1p2$$46281772_128x8m81
.ends

.subckt nmos_5p0431059054870_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.81u l=0.6u
.ends

.subckt nmos_1p2$$47119404_128x8m81 nmos_5p0431059054870_128x8m81_0/S nmos_5p0431059054870_128x8m81_0/D
+ a_n31_n74# VSUBS
Xnmos_5p0431059054870_128x8m81_0 nmos_5p0431059054870_128x8m81_0/D a_n31_n74# nmos_5p0431059054870_128x8m81_0/S
+ VSUBS nmos_5p0431059054870_128x8m81
.ends

.subckt nmos_5p0431059054872_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.57u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=0.57u l=0.6u
.ends

.subckt ypass_gate_a_128x8m81 vss b bb db ypass d pcb a_222_11191# a_n4_11191# vdd
+ m3_n1_4331# a_447_11191# a_n80_n10# a_222_10416# m3_n1_1708# a_n4_10416# m3_n1_1160#
+ m3_n1_2030# pmos_5p0431059054871_128x8m81_1/D m3_n1_3366# a_447_10416# m3_n1_2352#
+ m3_n1_3688# m3_n1_4009# m3_n1_2674#
Xnmos_1p2$$47119404_128x8m81_0 b d ypass vss nmos_1p2$$47119404_128x8m81
Xnmos_1p2$$47119404_128x8m81_1 bb pmos_5p0431059054871_128x8m81_1/D ypass vss nmos_1p2$$47119404_128x8m81
Xpmos_1p2$$46889004_128x8m81_0 b vdd nmos_5p0431059054872_128x8m81_0/D d pmos_1p2$$46889004_128x8m81
Xpmos_5p0431059054871_128x8m81_1 vdd pmos_5p0431059054871_128x8m81_1/D nmos_5p0431059054872_128x8m81_0/D
+ bb pmos_5p0431059054871_128x8m81
Xpmos_5p0431059054871_128x8m81_0 vdd b pcb bb pmos_5p0431059054871_128x8m81
Xnmos_5p0431059054872_128x8m81_0 nmos_5p0431059054872_128x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059054872_128x8m81
X0 nmos_5p0431059054872_128x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd ypass nmos_5p0431059054872_128x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X2 a_447_11191# pcb a_222_11191# vdd pmos_3p3 w=3.41u l=0.6u
X3 a_222_11191# pcb a_n4_11191# vdd pmos_3p3 w=3.41u l=0.6u
X4 a_447_10416# pcb a_222_10416# vdd pmos_3p3 w=3.41u l=0.6u
X5 a_222_10416# pcb a_n4_10416# vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt ypass_gate_128x8m81 bb ypass d pcb db vdd m3_n1_4331# m3_n1_1708# m3_n1_1160#
+ m3_n1_2030# m3_n1_3366# m3_n1_2352# vss m3_n1_3688# m3_n1_4009# m3_n1_2674# b
Xnmos_1p2$$47119404_128x8m81_0 b d ypass vss nmos_1p2$$47119404_128x8m81
Xnmos_1p2$$47119404_128x8m81_1 bb db ypass vss nmos_1p2$$47119404_128x8m81
Xpmos_1p2$$46889004_128x8m81_0 b vdd nmos_5p0431059054872_128x8m81_0/D d pmos_1p2$$46889004_128x8m81
Xpmos_5p0431059054871_128x8m81_1 vdd db nmos_5p0431059054872_128x8m81_0/D bb pmos_5p0431059054871_128x8m81
Xpmos_5p0431059054871_128x8m81_0 vdd b pcb bb pmos_5p0431059054871_128x8m81
Xnmos_5p0431059054872_128x8m81_0 nmos_5p0431059054872_128x8m81_0/D ypass vss ypass
+ vss nmos_5p0431059054872_128x8m81
X0 nmos_5p0431059054872_128x8m81_0/D ypass vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd ypass nmos_5p0431059054872_128x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt mux821_128x8m81 a_656_7735# ypass_gate_128x8m81_0/ypass ypass_gate_128x8m81_1/ypass
+ ypass_gate_128x8m81_0/d ypass_gate_128x8m81_2/ypass ypass_gate_128x8m81_4/b ypass_gate_128x8m81_3/ypass
+ ypass_gate_a_128x8m81_0/a_222_10416# ypass_gate_128x8m81_2/d ypass_gate_128x8m81_4/ypass
+ ypass_gate_128x8m81_5/ypass ypass_gate_128x8m81_6/ypass ypass_gate_128x8m81_4/d
+ ypass_gate_128x8m81_6/db ypass_gate_a_128x8m81_0/ypass ypass_gate_128x8m81_4/db
+ ypass_gate_128x8m81_6/d ypass_gate_a_128x8m81_0/a_447_10416# ypass_gate_a_128x8m81_0/db
+ ypass_gate_128x8m81_6/m3_n1_4331# ypass_gate_a_128x8m81_0/d ypass_gate_a_128x8m81_0/b
+ ypass_gate_128x8m81_1/d ypass_gate_128x8m81_5/db ypass_gate_a_128x8m81_0/a_222_11191#
+ a_4992_424# ypass_gate_128x8m81_3/d ypass_gate_a_128x8m81_0/a_n80_n10# ypass_gate_128x8m81_6/m3_n1_1708#
+ ypass_gate_128x8m81_5/d ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vdd
+ ypass_gate_a_128x8m81_0/a_447_11191# ypass_gate_128x8m81_6/m3_n1_2674# ypass_gate_128x8m81_6/m3_n1_3688#
+ ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/vss
Xypass_gate_a_128x8m81_0 ypass_gate_128x8m81_6/vss ypass_gate_a_128x8m81_0/b ypass_gate_a_128x8m81_0/bb
+ ypass_gate_a_128x8m81_0/db ypass_gate_a_128x8m81_0/ypass ypass_gate_a_128x8m81_0/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_a_128x8m81_0/a_222_11191# ypass_gate_128x8m81_6/vdd
+ ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331# ypass_gate_a_128x8m81_0/a_447_11191#
+ ypass_gate_a_128x8m81_0/a_n80_n10# ypass_gate_a_128x8m81_0/a_222_10416# ypass_gate_128x8m81_6/m3_n1_1708#
+ ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_1/db ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_a_128x8m81_0/a_447_10416#
+ ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009#
+ ypass_gate_128x8m81_6/m3_n1_2674# ypass_gate_a_128x8m81
Xypass_gate_128x8m81_0 ypass_gate_128x8m81_0/bb ypass_gate_128x8m81_0/ypass ypass_gate_128x8m81_0/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_4/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_0/b ypass_gate_128x8m81
Xypass_gate_128x8m81_1 ypass_gate_128x8m81_1/bb ypass_gate_128x8m81_1/ypass ypass_gate_128x8m81_1/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_1/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_1/b ypass_gate_128x8m81
Xypass_gate_128x8m81_2 ypass_gate_128x8m81_2/bb ypass_gate_128x8m81_2/ypass ypass_gate_128x8m81_2/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_5/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_2/b ypass_gate_128x8m81
Xypass_gate_128x8m81_3 ypass_gate_128x8m81_3/bb ypass_gate_128x8m81_3/ypass ypass_gate_128x8m81_3/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_6/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_3/b ypass_gate_128x8m81
Xypass_gate_128x8m81_4 ypass_gate_128x8m81_4/bb ypass_gate_128x8m81_4/ypass ypass_gate_128x8m81_4/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_4/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_4/b ypass_gate_128x8m81
Xypass_gate_128x8m81_5 ypass_gate_128x8m81_5/bb ypass_gate_128x8m81_5/ypass ypass_gate_128x8m81_5/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_5/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_5/b ypass_gate_128x8m81
Xypass_gate_128x8m81_6 ypass_gate_128x8m81_6/bb ypass_gate_128x8m81_6/ypass ypass_gate_128x8m81_6/d
+ ypass_gate_128x8m81_6/pcb ypass_gate_128x8m81_6/db ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_4331#
+ ypass_gate_128x8m81_6/m3_n1_1708# ypass_gate_128x8m81_6/vdd ypass_gate_128x8m81_6/m3_n1_2030#
+ ypass_gate_128x8m81_6/m3_n1_3366# ypass_gate_128x8m81_6/m3_n1_2352# ypass_gate_128x8m81_6/vss
+ ypass_gate_128x8m81_6/m3_n1_3688# ypass_gate_128x8m81_6/m3_n1_4009# ypass_gate_128x8m81_6/m3_n1_2674#
+ ypass_gate_128x8m81_6/b ypass_gate_128x8m81
.ends

.subckt pmos_1p2$$202586156_128x8m81 pmos_5p04310590548714_128x8m81_0/S w_n286_n141#
+ pmos_5p04310590548714_128x8m81_0/D a_n31_n74#
Xpmos_5p04310590548714_128x8m81_0 w_n286_n141# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt pmos_1p2$$202583084_128x8m81 pmos_5p04310590548735_128x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310590548735_128x8m81_0/S
Xpmos_5p04310590548735_128x8m81_0 w_n286_n142# pmos_5p04310590548735_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548735_128x8m81_0/S a_193_n74# pmos_5p04310590548735_128x8m81
.ends

.subckt pmos_1p2$$202587180_128x8m81 pmos_5p04310590548714_128x8m81_0/S w_n286_n141#
+ pmos_5p04310590548714_128x8m81_0/D a_n31_n74#
Xpmos_5p04310590548714_128x8m81_0 w_n286_n141# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt pmos_5p04310590548743_128x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2u l=0.6u
.ends

.subckt nmos_5p04310590548742_128x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.8u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.8u l=0.6u
.ends

.subckt nmos_5p04310590548740_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.37u l=0.6u
.ends

.subckt nmos_1p2$$202594348_128x8m81 a_n31_n73# nmos_5p04310590548740_128x8m81_0/D
+ nmos_5p04310590548740_128x8m81_0/S VSUBS
Xnmos_5p04310590548740_128x8m81_0 nmos_5p04310590548740_128x8m81_0/D a_n31_n73# nmos_5p04310590548740_128x8m81_0/S
+ VSUBS nmos_5p04310590548740_128x8m81
.ends

.subckt nmos_1p2$$202598444_128x8m81 nmos_5p04310590548710_128x8m81_0/D nmos_5p04310590548710_128x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310590548710_128x8m81_0 nmos_5p04310590548710_128x8m81_0/D a_n31_n74# nmos_5p04310590548710_128x8m81_0/S
+ VSUBS nmos_5p04310590548710_128x8m81
.ends

.subckt pmos_5p04310590548741_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.96u l=0.6u
.ends

.subckt nmos_1p2$$202595372_128x8m81 nmos_5p0431059054878_128x8m81_0/D a_n31_n73#
+ nmos_5p0431059054878_128x8m81_0/S VSUBS
Xnmos_5p0431059054878_128x8m81_0 nmos_5p0431059054878_128x8m81_0/D a_n31_n73# nmos_5p0431059054878_128x8m81_0/S
+ VSUBS nmos_5p0431059054878_128x8m81
.ends

.subckt nmos_5p04310590548739_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt nmos_1p2$$202596396_128x8m81 nmos_5p0431059054878_128x8m81_0/D a_n31_n73#
+ nmos_5p0431059054878_128x8m81_0/S VSUBS
Xnmos_5p0431059054878_128x8m81_0 nmos_5p0431059054878_128x8m81_0/D a_n31_n73# nmos_5p0431059054878_128x8m81_0/S
+ VSUBS nmos_5p0431059054878_128x8m81
.ends

.subckt pmos_1p2$$202584108_128x8m81 pmos_5p04310590548714_128x8m81_0/S a_n31_n74#
+ w_n286_n141# pmos_5p04310590548714_128x8m81_0/D
Xpmos_5p04310590548714_128x8m81_0 w_n286_n141# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt pmos_1p2$$202585132_128x8m81 w_n256_n141# pmos_5p04310590548714_128x8m81_0/S
+ pmos_5p04310590548714_128x8m81_0/D a_n31_n74#
Xpmos_5p04310590548714_128x8m81_0 w_n256_n141# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt wen_wm1_128x8m81 GWEN vss wep wen vdd men
Xpmos_1p2$$202586156_128x8m81_0 pmos_5p04310590548741_128x8m81_0/D vdd vdd nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ pmos_1p2$$202586156_128x8m81
Xpmos_1p2$$202583084_128x8m81_0 pmos_1p2$$202583084_128x8m81_0/pmos_5p04310590548735_128x8m81_0/D
+ nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D vdd nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ vdd pmos_1p2$$202583084_128x8m81
Xpmos_5p04310590548735_128x8m81_0 vdd pmos_5p04310590548735_128x8m81_0/D pmos_5p04310590548720_128x8m81_0/S
+ vdd pmos_5p04310590548720_128x8m81_0/S pmos_5p04310590548735_128x8m81
Xpmos_1p2$$202587180_128x8m81_0 nmos_5p0431059054878_128x8m81_1/D vdd pmos_5p04310590548741_128x8m81_0/S
+ nmos_5p0431059054878_128x8m81_3/D pmos_1p2$$202587180_128x8m81
Xnmos_5p0431059054878_128x8m81_0 vss GWEN nmos_5p0431059054878_128x8m81_2/D vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_0 vdd pmos_5p04310590548714_128x8m81_2/S wen vdd pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_1 nmos_5p0431059054878_128x8m81_1/D nmos_5p0431059054878_128x8m81_2/D
+ vss vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548743_128x8m81_0 vdd wep pmos_5p04310590548735_128x8m81_0/D vdd pmos_5p04310590548735_128x8m81_0/D
+ pmos_5p04310590548735_128x8m81_0/D pmos_5p04310590548743_128x8m81
Xnmos_5p04310590548742_128x8m81_0 wep pmos_5p04310590548735_128x8m81_0/D vss pmos_5p04310590548735_128x8m81_0/D
+ pmos_5p04310590548735_128x8m81_0/D vss nmos_5p04310590548742_128x8m81
Xpmos_5p04310590548714_128x8m81_1 vdd nmos_5p0431059054878_128x8m81_1/D nmos_5p0431059054878_128x8m81_2/D
+ vdd pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_2 nmos_5p0431059054878_128x8m81_2/D wen vss vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_2 vdd nmos_5p0431059054878_128x8m81_2/D GWEN pmos_5p04310590548714_128x8m81_2/S
+ pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_3 nmos_5p0431059054878_128x8m81_3/D pmos_5p04310590548714_128x8m81_5/D
+ vss vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_3 vdd pmos_5p04310590548714_128x8m81_5/S men vdd pmos_5p04310590548714_128x8m81
Xpmos_5p04310590548714_128x8m81_4 vdd nmos_5p0431059054878_128x8m81_3/D pmos_5p04310590548714_128x8m81_5/D
+ vdd pmos_5p04310590548714_128x8m81
Xnmos_1p2$$202594348_128x8m81_0 nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ vss pmos_1p2$$202583084_128x8m81_0/pmos_5p04310590548735_128x8m81_0/D vss nmos_1p2$$202594348_128x8m81
Xpmos_5p04310590548714_128x8m81_5 vdd pmos_5p04310590548714_128x8m81_5/D vss pmos_5p04310590548714_128x8m81_5/S
+ pmos_5p04310590548714_128x8m81
Xnmos_5p04310590548740_128x8m81_0 pmos_5p04310590548735_128x8m81_0/D pmos_5p04310590548720_128x8m81_0/S
+ vss vss nmos_5p04310590548740_128x8m81
Xnmos_1p2$$202598444_128x8m81_0 pmos_5p04310590548741_128x8m81_0/S nmos_5p0431059054878_128x8m81_1/D
+ pmos_5p04310590548714_128x8m81_5/D vss nmos_1p2$$202598444_128x8m81
Xpmos_5p04310590548741_128x8m81_0 vdd pmos_5p04310590548741_128x8m81_0/D pmos_5p04310590548714_128x8m81_5/D
+ pmos_5p04310590548741_128x8m81_0/S pmos_5p04310590548741_128x8m81
Xnmos_5p04310590548740_128x8m81_1 pmos_5p04310590548714_128x8m81_5/D men vss vss nmos_5p04310590548740_128x8m81
Xnmos_1p2$$202595372_128x8m81_0 pmos_5p04310590548741_128x8m81_0/D nmos_5p0431059054878_128x8m81_3/D
+ pmos_5p04310590548741_128x8m81_0/S vss nmos_1p2$$202595372_128x8m81
Xnmos_1p2$$202595372_128x8m81_1 vss pmos_5p04310590548741_128x8m81_0/S nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ vss nmos_1p2$$202595372_128x8m81
Xnmos_5p04310590548740_128x8m81_2 vss vss pmos_5p04310590548714_128x8m81_5/D vss nmos_5p04310590548740_128x8m81
Xnmos_5p04310590548710_128x8m81_0 vss nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ pmos_5p04310590548720_128x8m81_0/S vss nmos_5p04310590548710_128x8m81
Xpmos_5p04310590548720_128x8m81_0 vdd men nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ pmos_5p04310590548720_128x8m81_0/S nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ pmos_5p04310590548720_128x8m81
Xnmos_5p04310590548739_128x8m81_0 men pmos_1p2$$202583084_128x8m81_0/pmos_5p04310590548735_128x8m81_0/D
+ pmos_5p04310590548720_128x8m81_0/S pmos_1p2$$202583084_128x8m81_0/pmos_5p04310590548735_128x8m81_0/D
+ vss nmos_5p04310590548739_128x8m81
Xnmos_1p2$$202596396_128x8m81_0 nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S vss vss nmos_1p2$$202596396_128x8m81
Xnmos_1p2$$202596396_128x8m81_1 vss nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ pmos_5p04310590548741_128x8m81_0/D vss nmos_1p2$$202596396_128x8m81
Xpmos_1p2$$202584108_128x8m81_0 nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ pmos_5p04310590548741_128x8m81_0/S vdd vdd pmos_1p2$$202584108_128x8m81
Xpmos_1p2$$202585132_128x8m81_0 vdd vdd nmos_1p2$$202596396_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ nmos_1p2$$202595372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S pmos_1p2$$202585132_128x8m81
.ends

.subckt nmos_5p04310590548746_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=2.12u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=2.12u l=0.6u
.ends

.subckt pmos_5p04310590548747_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4u l=0.6u
.ends

.subckt nmos_5p04310590548745_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310590548744_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310590548752_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.6u l=0.6u
.ends

.subckt nmos_5p04310590548750_128x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2.27u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2.27u l=0.6u
.ends

.subckt pmos_5p04310590548751_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.67u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$171625516_128x8m81 pmos_5p0431059054873_128x8m81_0/S pmos_5p0431059054873_128x8m81_0/D
+ a_193_n74# w_n286_n142# a_n31_n74# pmos_5p0431059054873_128x8m81_0/w_n208_n120#
Xpmos_5p0431059054873_128x8m81_0 pmos_5p0431059054873_128x8m81_0/w_n208_n120# pmos_5p0431059054873_128x8m81_0/D
+ a_n31_n74# pmos_5p0431059054873_128x8m81_0/S a_193_n74# pmos_5p0431059054873_128x8m81
.ends

.subckt pmos_5p04310590548749_128x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=3.78u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=3.78u l=0.6u
.ends

.subckt pmos_5p04310590548748_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.5u l=0.6u
.ends

.subckt outbuf_oe_128x8m81 qp qn se q GWE a_4913_n316# vdd vss
Xnmos_5p04310590548746_128x8m81_0 vss pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D q pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D vss nmos_5p04310590548746_128x8m81
Xpmos_5p04310590548747_128x8m81_0 vdd vdd GWE pmos_5p04310590548747_128x8m81_0/S pmos_5p04310590548747_128x8m81
Xnmos_5p04310590548745_128x8m81_0 vss pmos_5p04310590548747_128x8m81_0/S nmos_5p04310590548745_128x8m81_1/S
+ pmos_5p04310590548747_128x8m81_0/S vss nmos_5p04310590548745_128x8m81
Xnmos_5p04310590548745_128x8m81_1 pmos_5p04310590548751_128x8m81_0/D qn nmos_5p04310590548745_128x8m81_1/S
+ qn vss nmos_5p04310590548745_128x8m81
Xnmos_5p04310590548744_128x8m81_0 vss pmos_5p04310590548747_128x8m81_0/S pmos_5p04310590548748_128x8m81_0/S
+ vss nmos_5p04310590548744_128x8m81
Xnmos_5p0431059054878_128x8m81_0 nmos_5p0431059054878_128x8m81_0/D se vss vss nmos_5p0431059054878_128x8m81
Xnmos_5p04310590548733_128x8m81_0 pmos_5p04310590548738_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ vss vss nmos_5p04310590548733_128x8m81
Xnmos_5p0431059054878_128x8m81_1 vss pmos_5p04310590548738_128x8m81_0/D nmos_5p0431059054878_128x8m81_1/S
+ vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_0 vdd nmos_5p0431059054878_128x8m81_0/D se vdd pmos_5p04310590548714_128x8m81
Xnmos_5p04310590548752_128x8m81_0 vss GWE pmos_5p04310590548747_128x8m81_0/S vss nmos_5p04310590548752_128x8m81
Xpmos_5p04310590548713_128x8m81_0 vdd nmos_5p0431059054878_128x8m81_1/S se pmos_5p04310590548751_128x8m81_0/D
+ se se pmos_5p04310590548713_128x8m81
Xnmos_5p04310590548750_128x8m81_0 nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D nmos_5p0431059054878_128x8m81_0/D nmos_5p0431059054878_128x8m81_0/D
+ vss nmos_5p04310590548750_128x8m81
Xpmos_5p04310590548751_128x8m81_0 vdd pmos_5p04310590548751_128x8m81_0/D qp pmos_5p04310590548751_128x8m81_1/S
+ qp pmos_5p04310590548751_128x8m81
Xpmos_5p04310590548751_128x8m81_1 vdd vdd pmos_5p04310590548748_128x8m81_0/S pmos_5p04310590548751_128x8m81_1/S
+ pmos_5p04310590548748_128x8m81_0/S pmos_5p04310590548751_128x8m81
Xpmos_1p2$$171625516_128x8m81_0 vdd nmos_5p0431059054878_128x8m81_1/S pmos_5p04310590548738_128x8m81_0/D
+ vdd pmos_5p04310590548738_128x8m81_0/D vdd pmos_1p2$$171625516_128x8m81
Xpmos_5p04310590548749_128x8m81_0 vdd vdd pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D q pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548749_128x8m81
Xpmos_5p04310590548748_128x8m81_0 vdd vdd pmos_5p04310590548747_128x8m81_0/S pmos_5p04310590548748_128x8m81_0/S
+ pmos_5p04310590548748_128x8m81
Xpmos_5p04310590548738_128x8m81_0 vdd pmos_5p04310590548738_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D
+ vdd pmos_5p04310590548738_128x8m81
.ends

.subckt saout_m2_128x8m81 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] GWEN bb[2] bb[7] b[0] datain q pcb WEN a_5189_27176# a_5414_27176#
+ a_5189_27951# a_5414_27951# wen_wm1_128x8m81_0/GWEN sacntl_2_128x8m81_0/a_4718_983#
+ b[7] mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10# b[5] sa_128x8m81_0/wep
+ mux821_128x8m81_0/a_4992_424# b[1] b[6] bb[4] b[2] GWE bb[3] b[3] mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ bb[0] bb[1] mux821_128x8m81_0/a_656_7735# sacntl_2_128x8m81_0/a_4560_1922# outbuf_oe_128x8m81_0/a_4913_n316#
+ bb[6] mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass wen_wm1_128x8m81_0/vdd mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass
+ din_128x8m81_0/men bb[5] b[4] sa_128x8m81_0/pcb mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass vdd mux821_128x8m81_0/ypass_gate_128x8m81_6/vdd
+ mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass sacntl_2_128x8m81_0/vdd mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass
+ mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ vss
Xsa_128x8m81_0 sa_128x8m81_0/qp sa_128x8m81_0/wep sa_128x8m81_0/se sa_128x8m81_0/pcb
+ vss vdd sa_128x8m81
Xdin_128x8m81_0 vdd vdd datain sa_128x8m81_0/wep din_128x8m81_0/men sa_128x8m81_0/pcb
+ vss vdd vdd din_128x8m81
Xsacntl_2_128x8m81_0 din_128x8m81_0/men sa_128x8m81_0/pcb sacntl_2_128x8m81_0/a_4718_983#
+ vss sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_2/S sa_128x8m81_0/se sacntl_2_128x8m81_0/a_4560_1922#
+ sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_2/S sacntl_2_128x8m81_0/pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_1/S vss sacntl_2_128x8m81_0/vdd
+ sacntl_2_128x8m81
Xmux821_128x8m81_0 mux821_128x8m81_0/a_656_7735# mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass vdd mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_4/b mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass
+ a_5189_27176# vdd mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass vdd vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass
+ vdd vdd a_5414_27176# vdd mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ vdd vdd a_5189_27951# mux821_128x8m81_0/a_4992_424# vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10#
+ mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass vdd mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass sa_128x8m81_0/pcb mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/vdd a_5414_27951# mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass
+ vss mux821_128x8m81
Xwen_wm1_128x8m81_0 wen_wm1_128x8m81_0/GWEN vss sa_128x8m81_0/wep wen_wm1_128x8m81_0/wen
+ wen_wm1_128x8m81_0/vdd din_128x8m81_0/men wen_wm1_128x8m81
Xoutbuf_oe_128x8m81_0 sa_128x8m81_0/qp sa_128x8m81_0/qp sa_128x8m81_0/se q GWE outbuf_oe_128x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_128x8m81
.ends

.subckt saout_R_m2_128x8m81 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6]
+ ypass[7] men ypass[0] GWEN datain b[0] bb[5] q bb[0] pcb WEN wen_wm1_128x8m81_0/GWEN
+ sacntl_2_128x8m81_0/a_4718_983# mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass b[2]
+ sa_128x8m81_0/wep mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass b[6] mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass
+ b[1] bb[3] b[5] GWE bb[4] mux821_128x8m81_0/ypass_gate_128x8m81_4/b wen_wm1_128x8m81_0/wen
+ b[4] b[7] bb[7] bb[6] a_5189_27169# a_5414_27169# mux821_128x8m81_0/a_656_7735#
+ mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass a_5189_27944# a_5414_27944# sacntl_2_128x8m81_0/a_4560_1922#
+ outbuf_oe_128x8m81_0/a_4913_n316# bb[1] wen_wm1_128x8m81_0/vdd din_128x8m81_0/men
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass bb[2] b[3] sa_128x8m81_0/pcb mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ vdd mux821_128x8m81_0/ypass_gate_128x8m81_6/vdd mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass sacntl_2_128x8m81_0/vdd vss
Xsa_128x8m81_0 sa_128x8m81_0/qp sa_128x8m81_0/wep sa_128x8m81_0/se sa_128x8m81_0/pcb
+ vss vdd sa_128x8m81
Xdin_128x8m81_0 vdd vdd datain sa_128x8m81_0/wep din_128x8m81_0/men sa_128x8m81_0/pcb
+ vss vdd vdd din_128x8m81
Xsacntl_2_128x8m81_0 din_128x8m81_0/men sa_128x8m81_0/pcb sacntl_2_128x8m81_0/a_4718_983#
+ vss sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_2/S sa_128x8m81_0/se sacntl_2_128x8m81_0/a_4560_1922#
+ sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_2/S sacntl_2_128x8m81_0/pmos_1p2$$46282796_128x8m81_0/pmos_5p04310590548724_128x8m81_0/D
+ sacntl_2_128x8m81_0/pmos_5p04310590548727_128x8m81_1/S vss sacntl_2_128x8m81_0/vdd
+ sacntl_2_128x8m81
Xmux821_128x8m81_0 mux821_128x8m81_0/a_656_7735# mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass vdd mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_4/b mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass
+ a_5189_27169# vdd mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass vdd vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass
+ vdd vdd a_5414_27169# vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/ypass vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ vdd vdd a_5189_27944# mux821_128x8m81_0/a_4992_424# vdd mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10#
+ mux821_128x8m81_0/ypass_gate_128x8m81_3/ypass vdd mux821_128x8m81_0/ypass_gate_128x8m81_0/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/ypass sa_128x8m81_0/pcb mux821_128x8m81_0/ypass_gate_128x8m81_2/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_6/vdd a_5414_27944# mux821_128x8m81_0/ypass_gate_128x8m81_5/ypass
+ mux821_128x8m81_0/ypass_gate_128x8m81_4/ypass mux821_128x8m81_0/ypass_gate_128x8m81_1/ypass
+ vss mux821_128x8m81
Xwen_wm1_128x8m81_0 wen_wm1_128x8m81_0/GWEN vss sa_128x8m81_0/wep wen_wm1_128x8m81_0/wen
+ wen_wm1_128x8m81_0/vdd din_128x8m81_0/men wen_wm1_128x8m81
Xoutbuf_oe_128x8m81_0 sa_128x8m81_0/qp sa_128x8m81_0/qp sa_128x8m81_0/se q GWE outbuf_oe_128x8m81_0/a_4913_n316#
+ vdd vss outbuf_oe_128x8m81
.ends

.subckt saout_wm1_x4_128x8m81 ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] ypass[2]
+ b[1] b[4] b[7] b[10] b[13] b[16] b[19] b[22] b[25] b[28] b[31] din[1] din[3] din[2]
+ din[0] q[0] q[1] q[2] q[3] b[29] b[26] b[23] b[20] b[17] b[14] b[11] b[8] b[5] b[2]
+ bb[0] bb[1] bb[2] bb[3] bb[4] bb[5] bb[6] bb[7] bb[8] bb[9] bb[10] bb[11] bb[12]
+ bb[13] bb[14] bb[15] bb[16] bb[17] bb[18] bb[19] bb[20] bb[21] bb[22] bb[23] bb[24]
+ bb[25] bb[26] bb[27] bb[28] bb[29] bb[30] bb[31] b[30] b[27] b[24] b[15] b[12] b[9]
+ b[21] b[0] b[3] b[6] b[18] pcb[0] pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1] WEN[0]
+ saout_R_m2_128x8m81_1/bb[4] saout_m2_128x8m81_0/b[0] saout_R_m2_128x8m81_1/bb[1]
+ a_15501_29383# saout_m2_128x8m81_0/bb[0] saout_m2_128x8m81_0/bb[1] saout_R_m2_128x8m81_0/bb[5]
+ saout_m2_128x8m81_0/bb[6] saout_R_m2_128x8m81_1/b[4] m1_9952_31280# a_15261_28608#
+ saout_R_m2_128x8m81_0/bb[1] saout_R_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[2]
+ saout_R_m2_128x8m81_1/bb[7] saout_R_m2_128x8m81_1/bb[6] saout_R_m2_128x8m81_0/wen_wm1_128x8m81_0/wen
+ saout_m2_128x8m81_0/WEN saout_R_m2_128x8m81_0/b[2] men saout_R_m2_128x8m81_0/b[6]
+ saout_m2_128x8m81_1/bb[7] a_4701_29383# saout_R_m2_128x8m81_0/bb[3] m1_n848_31280#
+ saout_R_m2_128x8m81_0/b[5] GWE saout_R_m2_128x8m81_1/bb[0] saout_m2_128x8m81_0/bb[5]
+ saout_m2_128x8m81_0/b[4] saout_m2_128x8m81_1/b[5] saout_R_m2_128x8m81_0/bb[4] saout_m2_128x8m81_1/b[1]
+ saout_m2_128x8m81_0/bb[7] saout_m2_128x8m81_1/bb[4] a_4461_28608# saout_m2_128x8m81_1/b[2]
+ saout_R_m2_128x8m81_0/b[4] a_15501_28608# saout_R_m2_128x8m81_0/bb[0] saout_m2_128x8m81_1/bb[3]
+ saout_R_m2_128x8m81_1/bb[2] saout_R_m2_128x8m81_1/b[3] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_0/b[7] saout_m2_128x8m81_0/bb[2] saout_R_m2_128x8m81_0/bb[7]
+ saout_R_m2_128x8m81_0/bb[6] ypass[6] saout_m2_128x8m81_1/b[3] saout_R_m2_128x8m81_1/b[0]
+ saout_m2_128x8m81_1/b[6] ypass[7] saout_m2_128x8m81_1/b[0] saout_m2_128x8m81_0/b[7]
+ saout_m2_128x8m81_1/bb[0] saout_m2_128x8m81_1/bb[1] saout_R_m2_128x8m81_1/b[1] saout_R_m2_128x8m81_1/bb[5]
+ a_15261_29383# saout_m2_128x8m81_1/GWEN saout_R_m2_128x8m81_0/b[0] m1_15352_31280#
+ saout_m2_128x8m81_0/b[6] m1_4552_31280# m1_20752_31280# saout_R_m2_128x8m81_0/b[1]
+ saout_m2_128x8m81_0/b[5] saout_R_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_128x8m81_4/b
+ saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735# a_4701_28608# saout_m2_128x8m81_0/b[1]
+ saout_m2_128x8m81_0/bb[4] saout_m2_128x8m81_0/b[2] saout_m2_128x8m81_0/pcb saout_m2_128x8m81_0/bb[3]
+ saout_m2_128x8m81_1/sa_128x8m81_0/pcb saout_R_m2_128x8m81_0/bb[2] saout_R_m2_128x8m81_0/b[3]
+ saout_R_m2_128x8m81_1/b[2] saout_R_m2_128x8m81_1/sa_128x8m81_0/pcb saout_R_m2_128x8m81_1/b[6]
+ saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb saout_R_m2_128x8m81_1/bb[3] saout_m2_128x8m81_0/b[3]
+ saout_m2_128x8m81_1/bb[6] saout_R_m2_128x8m81_1/b[5] a_4461_29383# VSS saout_m2_128x8m81_1/bb[5]
+ VDD saout_m2_128x8m81_1/b[4]
Xsaout_m2_128x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] saout_m2_128x8m81_1/GWEN saout_m2_128x8m81_0/bb[2] saout_m2_128x8m81_0/bb[7]
+ saout_m2_128x8m81_0/b[0] saout_m2_128x8m81_0/datain saout_m2_128x8m81_0/q saout_m2_128x8m81_0/pcb
+ saout_m2_128x8m81_0/WEN a_4236_28608# a_4461_28608# a_4236_29383# a_4461_29383#
+ saout_m2_128x8m81_1/GWEN VSS saout_m2_128x8m81_0/b[7] saout_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10#
+ saout_m2_128x8m81_0/b[5] saout_m2_128x8m81_0/sa_128x8m81_0/wep saout_m2_128x8m81_0/mux821_128x8m81_0/a_4992_424#
+ saout_m2_128x8m81_0/b[1] saout_m2_128x8m81_0/b[6] saout_m2_128x8m81_0/bb[4] saout_m2_128x8m81_0/b[2]
+ GWE saout_m2_128x8m81_0/bb[3] saout_m2_128x8m81_0/b[3] saout_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ saout_m2_128x8m81_0/bb[0] saout_m2_128x8m81_0/bb[1] saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ VSS VSS saout_m2_128x8m81_0/bb[6] ypass[7] VDD ypass[1] men saout_m2_128x8m81_0/bb[5]
+ saout_m2_128x8m81_0/b[4] saout_m2_128x8m81_0/pcb ypass[2] ypass[4] VDD VDD ypass[5]
+ VDD ypass[6] ypass[0] ypass[3] VSS saout_m2_128x8m81
Xsaout_m2_128x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] saout_m2_128x8m81_1/GWEN saout_m2_128x8m81_1/bb[2] saout_m2_128x8m81_1/bb[7]
+ saout_m2_128x8m81_1/b[0] saout_m2_128x8m81_1/datain saout_m2_128x8m81_1/q saout_m2_128x8m81_1/pcb
+ saout_m2_128x8m81_1/WEN a_15036_28608# a_15261_28608# a_15036_29383# a_15261_29383#
+ saout_m2_128x8m81_1/GWEN VSS saout_m2_128x8m81_1/b[7] VSS saout_m2_128x8m81_1/b[5]
+ saout_m2_128x8m81_1/sa_128x8m81_0/wep VSS saout_m2_128x8m81_1/b[1] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/bb[4] saout_m2_128x8m81_1/b[2] GWE saout_m2_128x8m81_1/bb[3]
+ saout_m2_128x8m81_1/b[3] saout_m2_128x8m81_1/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ saout_m2_128x8m81_1/bb[0] saout_m2_128x8m81_1/bb[1] saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ VSS VSS saout_m2_128x8m81_1/bb[6] ypass[7] VDD ypass[1] men saout_m2_128x8m81_1/bb[5]
+ saout_m2_128x8m81_1/b[4] saout_m2_128x8m81_1/sa_128x8m81_0/pcb ypass[2] ypass[4]
+ VDD VDD ypass[5] VDD ypass[6] ypass[0] ypass[3] VSS saout_m2_128x8m81
Xsaout_R_m2_128x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] saout_m2_128x8m81_1/GWEN saout_R_m2_128x8m81_0/datain saout_R_m2_128x8m81_0/b[0]
+ saout_R_m2_128x8m81_0/bb[5] saout_R_m2_128x8m81_0/q saout_R_m2_128x8m81_0/bb[0]
+ saout_R_m2_128x8m81_0/pcb saout_R_m2_128x8m81_0/WEN saout_m2_128x8m81_1/GWEN saout_R_m2_128x8m81_0/sacntl_2_128x8m81_0/a_4718_983#
+ ypass[5] saout_R_m2_128x8m81_0/b[2] saout_R_m2_128x8m81_0/sa_128x8m81_0/wep ypass[6]
+ saout_R_m2_128x8m81_0/b[6] ypass[3] saout_R_m2_128x8m81_0/b[1] saout_R_m2_128x8m81_0/bb[3]
+ saout_R_m2_128x8m81_0/b[5] GWE saout_R_m2_128x8m81_0/bb[4] saout_R_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_128x8m81_4/b
+ saout_R_m2_128x8m81_0/wen_wm1_128x8m81_0/wen saout_R_m2_128x8m81_0/b[4] saout_R_m2_128x8m81_0/b[7]
+ saout_R_m2_128x8m81_0/bb[7] saout_R_m2_128x8m81_0/bb[6] a_15727_28608# a_15501_28608#
+ saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735# ypass[7] a_15727_29383# a_15501_29383#
+ VSS VSS saout_R_m2_128x8m81_0/bb[1] VDD men ypass[1] saout_R_m2_128x8m81_0/bb[2]
+ saout_R_m2_128x8m81_0/b[3] saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb ypass[4] VDD
+ VDD ypass[0] ypass[2] VDD VSS saout_R_m2_128x8m81
Xsaout_R_m2_128x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] saout_m2_128x8m81_1/GWEN saout_R_m2_128x8m81_1/datain saout_R_m2_128x8m81_1/b[0]
+ saout_R_m2_128x8m81_1/bb[5] saout_R_m2_128x8m81_1/q saout_R_m2_128x8m81_1/bb[0]
+ saout_R_m2_128x8m81_1/pcb saout_R_m2_128x8m81_1/WEN saout_m2_128x8m81_1/GWEN VSS
+ ypass[5] saout_R_m2_128x8m81_1/b[2] saout_R_m2_128x8m81_1/sa_128x8m81_0/wep ypass[6]
+ saout_R_m2_128x8m81_1/b[6] ypass[3] saout_R_m2_128x8m81_1/b[1] saout_R_m2_128x8m81_1/bb[3]
+ saout_R_m2_128x8m81_1/b[5] GWE saout_R_m2_128x8m81_1/bb[4] saout_R_m2_128x8m81_1/mux821_128x8m81_0/ypass_gate_128x8m81_4/b
+ saout_R_m2_128x8m81_1/wen_wm1_128x8m81_0/wen saout_R_m2_128x8m81_1/b[4] saout_R_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_1/bb[7] saout_R_m2_128x8m81_1/bb[6] a_4927_28608# a_4701_28608#
+ saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735# ypass[7] a_4927_29383# a_4701_29383#
+ VSS saout_R_m2_128x8m81_1/outbuf_oe_128x8m81_0/a_4913_n316# saout_R_m2_128x8m81_1/bb[1]
+ VDD men ypass[1] saout_R_m2_128x8m81_1/bb[2] saout_R_m2_128x8m81_1/b[3] saout_R_m2_128x8m81_1/sa_128x8m81_0/pcb
+ ypass[4] VDD VDD ypass[0] ypass[2] VDD VSS saout_R_m2_128x8m81
.ends

.subckt dcap_103_novia_128x8m81 w_n203_44# a_n67_185# a_73_103#
X0 a_n67_185# a_73_103# a_n67_185# w_n203_44# pmos_3p3 w=2.275u l=2.365u
.ends

.subckt lcol4_128_128x8m81 WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7]
+ WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] men ypass[0] ypass[1] ypass[2] ypass[3]
+ ypass[4] ypass[5] ypass[6] ypass[7] GWEN GWE din[0] din[1] din[3] din[2] q[0] q[1]
+ q[2] q[3] pcb[2] pcb[3] pcb[0] pcb[1] vdd WEN[2] WEN[1] WEN[0] col_128a_128x8m81_0/WL[0]
+ col_128a_128x8m81_0/WL[1] saout_wm1_x4_128x8m81_0/a_15501_28608# col_128a_128x8m81_0/WL[2]
+ col_128a_128x8m81_0/WL[3] col_128a_128x8m81_0/WL[4] col_128a_128x8m81_0/WL[10] col_128a_128x8m81_0/WL[5]
+ saout_wm1_x4_128x8m81_0/a_4701_29383# col_128a_128x8m81_0/WL[11] col_128a_128x8m81_0/WL[6]
+ col_128a_128x8m81_0/WL[12] col_128a_128x8m81_0/WL[7] col_128a_128x8m81_0/WL[13]
+ saout_wm1_x4_128x8m81_0/a_15261_29383# col_128a_128x8m81_0/WL[8] col_128a_128x8m81_0/WL[14]
+ saout_wm1_x4_128x8m81_0/men saout_wm1_x4_128x8m81_0/a_4461_28608# col_128a_128x8m81_0/WL[9]
+ col_128a_128x8m81_0/WL[15] saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_0/WEN saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/GWEN ldummy_128x4_128x8m81_0/VSS saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_0/wen_wm1_128x8m81_0/wen
+ saout_wm1_x4_128x8m81_0/a_15501_29383# saout_wm1_x4_128x8m81_0/a_4701_28608# saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_1/sa_128x8m81_0/pcb
+ saout_wm1_x4_128x8m81_0/a_15261_28608# saout_wm1_x4_128x8m81_0/WEN[3] saout_wm1_x4_128x8m81_0/ypass[0]
+ saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb saout_wm1_x4_128x8m81_0/a_4461_29383#
+ saout_wm1_x4_128x8m81_0/ypass[1] saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/sa_128x8m81_0/pcb
+ saout_wm1_x4_128x8m81_0/ypass[2] saout_wm1_x4_128x8m81_0/ypass[3] saout_wm1_x4_128x8m81_0/ypass[4]
+ saout_wm1_x4_128x8m81_0/GWE saout_wm1_x4_128x8m81_0/ypass[5] saout_wm1_x4_128x8m81_0/ypass[6]
+ saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_0/pcb saout_wm1_x4_128x8m81_0/ypass[7]
+ VSS VDD
Xldummy_128x4_128x8m81_0 saout_wm1_x4_128x8m81_0/b[30] saout_wm1_x4_128x8m81_0/bb[8]
+ VSS saout_wm1_x4_128x8m81_0/b[15] saout_wm1_x4_128x8m81_0/b[18] VDD saout_wm1_x4_128x8m81_0/bb[20]
+ saout_wm1_x4_128x8m81_0/bb[3] saout_wm1_x4_128x8m81_0/bb[15] saout_wm1_x4_128x8m81_0/b[9]
+ saout_wm1_x4_128x8m81_0/b[21] saout_wm1_x4_128x8m81_0/b[7] saout_wm1_x4_128x8m81_0/b[19]
+ VSS saout_wm1_x4_128x8m81_0/bb[9] VSS VDD saout_wm1_x4_128x8m81_0/bb[17] saout_wm1_x4_128x8m81_0/b[2]
+ VDD saout_wm1_x4_128x8m81_0/bb[7] saout_wm1_x4_128x8m81_0/bb[22] saout_wm1_x4_128x8m81_0/bb[20]
+ VSS saout_wm1_x4_128x8m81_0/b[10] saout_wm1_x4_128x8m81_0/b[21] VSS saout_wm1_x4_128x8m81_0/b[18]
+ saout_wm1_x4_128x8m81_0/b[16] saout_wm1_x4_128x8m81_0/b[19] VDD VDD saout_wm1_x4_128x8m81_0/bb[1]
+ saout_wm1_x4_128x8m81_0/bb[31] saout_wm1_x4_128x8m81_0/bb[18] saout_wm1_x4_128x8m81_0/b[17]
+ saout_wm1_x4_128x8m81_0/bb[11] saout_wm1_x4_128x8m81_0/bb[7] VSS saout_wm1_x4_128x8m81_0/bb[16]
+ saout_wm1_x4_128x8m81_0/bb[17] VSS saout_wm1_x4_128x8m81_0/b[24] saout_wm1_x4_128x8m81_0/bb[24]
+ saout_wm1_x4_128x8m81_0/b[0] saout_wm1_x4_128x8m81_0/b[25] saout_wm1_x4_128x8m81_0/bb[23]
+ saout_wm1_x4_128x8m81_0/bb[26] saout_wm1_x4_128x8m81_0/bb[6] saout_wm1_x4_128x8m81_0/bb[4]
+ saout_wm1_x4_128x8m81_0/bb[13] saout_wm1_x4_128x8m81_0/b[6] col_128a_128x8m81_0/WL[10]
+ saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/b[16] VSS VDD saout_wm1_x4_128x8m81_0/b[8]
+ saout_wm1_x4_128x8m81_0/bb[25] col_128a_128x8m81_0/WL[6] saout_wm1_x4_128x8m81_0/b[3]
+ col_128a_128x8m81_0/WL[8] saout_wm1_x4_128x8m81_0/bb[2] col_128a_128x8m81_0/WL[4]
+ saout_wm1_x4_128x8m81_0/b[4] saout_wm1_x4_128x8m81_0/b[1] saout_wm1_x4_128x8m81_0/b[12]
+ VDD saout_wm1_x4_128x8m81_0/b[31] saout_wm1_x4_128x8m81_0/b[24] col_128a_128x8m81_0/WL[0]
+ saout_wm1_x4_128x8m81_0/bb[0] saout_wm1_x4_128x8m81_0/b[26] saout_wm1_x4_128x8m81_0/bb[27]
+ VDD saout_wm1_x4_128x8m81_0/bb[9] saout_wm1_x4_128x8m81_0/b[23] col_128a_128x8m81_0/WL[2]
+ saout_wm1_x4_128x8m81_0/bb[8] saout_wm1_x4_128x8m81_0/b[9] saout_wm1_x4_128x8m81_0/b[14]
+ saout_wm1_x4_128x8m81_0/bb[10] saout_wm1_x4_128x8m81_0/bb[5] saout_wm1_x4_128x8m81_0/bb[25]
+ saout_wm1_x4_128x8m81_0/bb[29] VSS VDD saout_wm1_x4_128x8m81_0/b[10] saout_wm1_x4_128x8m81_0/bb[3]
+ saout_wm1_x4_128x8m81_0/bb[15] VSS saout_wm1_x4_128x8m81_0/b[28] col_128a_128x8m81_0/WL[15]
+ saout_wm1_x4_128x8m81_0/b[22] saout_wm1_x4_128x8m81_0/b[26] saout_wm1_x4_128x8m81_0/bb[18]
+ VDD saout_wm1_x4_128x8m81_0/bb[11] col_128a_128x8m81_0/WL[9] saout_wm1_x4_128x8m81_0/b[17]
+ col_128a_128x8m81_0/WL[11] saout_wm1_x4_128x8m81_0/bb[16] saout_wm1_x4_128x8m81_0/b[2]
+ saout_wm1_x4_128x8m81_0/b[22] col_128a_128x8m81_0/WL[7] saout_wm1_x4_128x8m81_0/bb[24]
+ VSS saout_wm1_x4_128x8m81_0/bb[27] saout_wm1_x4_128x8m81_0/b[20] saout_wm1_x4_128x8m81_0/b[30]
+ col_128a_128x8m81_0/WL[1] VDD VDD saout_wm1_x4_128x8m81_0/b[25] saout_wm1_x4_128x8m81_0/b[6]
+ saout_wm1_x4_128x8m81_0/bb[13] col_128a_128x8m81_0/WL[3] saout_wm1_x4_128x8m81_0/bb[26]
+ col_128a_128x8m81_0/WL[5] saout_wm1_x4_128x8m81_0/b[27] saout_wm1_x4_128x8m81_0/bb[1]
+ col_128a_128x8m81_0/WL[13] ldummy_128x4_128x8m81_0/VSS saout_wm1_x4_128x8m81_0/b[20]
+ VSS saout_wm1_x4_128x8m81_0/b[29] saout_wm1_x4_128x8m81_0/bb[31] saout_wm1_x4_128x8m81_0/bb[29]
+ col_128a_128x8m81_0/WL[14] VSS saout_wm1_x4_128x8m81_0/b[7] saout_wm1_x4_128x8m81_0/bb[21]
+ saout_wm1_x4_128x8m81_0/b[4] saout_wm1_x4_128x8m81_0/bb[28] VDD saout_wm1_x4_128x8m81_0/b[12]
+ saout_wm1_x4_128x8m81_0/bb[6] col_128a_128x8m81_0/WL[12] saout_wm1_x4_128x8m81_0/bb[30]
+ saout_wm1_x4_128x8m81_0/bb[10] saout_wm1_x4_128x8m81_0/bb[4] saout_wm1_x4_128x8m81_0/b[11]
+ saout_wm1_x4_128x8m81_0/b[27] saout_wm1_x4_128x8m81_0/b[0] VSS saout_wm1_x4_128x8m81_0/bb[21]
+ saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/b[13] saout_wm1_x4_128x8m81_0/b[29]
+ VDD VSS saout_wm1_x4_128x8m81_0/bb[19] saout_wm1_x4_128x8m81_0/b[3] saout_wm1_x4_128x8m81_0/bb[23]
+ saout_wm1_x4_128x8m81_0/b[28] saout_wm1_x4_128x8m81_0/bb[12] saout_wm1_x4_128x8m81_0/bb[5]
+ saout_wm1_x4_128x8m81_0/b[11] saout_wm1_x4_128x8m81_0/bb[28] VDD saout_wm1_x4_128x8m81_0/b[14]
+ saout_wm1_x4_128x8m81_0/bb[2] saout_wm1_x4_128x8m81_0/b[13] saout_wm1_x4_128x8m81_0/bb[30]
+ saout_wm1_x4_128x8m81_0/bb[14] saout_wm1_x4_128x8m81_0/b[1] saout_wm1_x4_128x8m81_0/bb[12]
+ saout_wm1_x4_128x8m81_0/b[31] saout_wm1_x4_128x8m81_0/b[15] saout_wm1_x4_128x8m81_0/bb[19]
+ VSS saout_wm1_x4_128x8m81_0/bb[0] saout_wm1_x4_128x8m81_0/b[8] saout_wm1_x4_128x8m81_0/bb[14]
+ VSS saout_wm1_x4_128x8m81_0/b[23] saout_wm1_x4_128x8m81_0/bb[22] VDD ldummy_128x4_128x8m81
Xcol_128a_128x8m81_0 col_128a_128x8m81_0/WL[3] col_128a_128x8m81_0/WL[2] col_128a_128x8m81_0/WL[1]
+ col_128a_128x8m81_0/WL[12] col_128a_128x8m81_0/WL[11] col_128a_128x8m81_0/WL[10]
+ col_128a_128x8m81_0/WL[9] col_128a_128x8m81_0/WL[8] col_128a_128x8m81_0/WL[7] col_128a_128x8m81_0/WL[6]
+ col_128a_128x8m81_0/WL[5] col_128a_128x8m81_0/WL[4] col_128a_128x8m81_0/WL[15] col_128a_128x8m81_0/WL[14]
+ col_128a_128x8m81_0/WL[13] col_128a_128x8m81_0/WL[0] saout_wm1_x4_128x8m81_0/b[24]
+ saout_wm1_x4_128x8m81_0/bb[11] saout_wm1_x4_128x8m81_0/bb[18] saout_wm1_x4_128x8m81_0/b[16]
+ saout_wm1_x4_128x8m81_0/bb[14] saout_wm1_x4_128x8m81_0/b[12] saout_wm1_x4_128x8m81_0/b[1]
+ saout_wm1_x4_128x8m81_0/bb[21] saout_wm1_x4_128x8m81_0/bb[4] saout_wm1_x4_128x8m81_0/bb[24]
+ saout_wm1_x4_128x8m81_0/b[10] saout_wm1_x4_128x8m81_0/bb[8] saout_wm1_x4_128x8m81_0/b[8]
+ saout_wm1_x4_128x8m81_0/bb[15] saout_wm1_x4_128x8m81_0/b[23] saout_wm1_x4_128x8m81_0/bb[1]
+ saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/bb[5] saout_wm1_x4_128x8m81_0/bb[0]
+ saout_wm1_x4_128x8m81_0/b[18] saout_wm1_x4_128x8m81_0/b[27] saout_wm1_x4_128x8m81_0/b[2]
+ saout_wm1_x4_128x8m81_0/b[21] saout_wm1_x4_128x8m81_0/bb[7] saout_wm1_x4_128x8m81_0/bb[30]
+ saout_wm1_x4_128x8m81_0/bb[27] saout_wm1_x4_128x8m81_0/bb[6] saout_wm1_x4_128x8m81_0/bb[23]
+ saout_wm1_x4_128x8m81_0/b[30] saout_wm1_x4_128x8m81_0/bb[12] saout_wm1_x4_128x8m81_0/b[3]
+ saout_wm1_x4_128x8m81_0/b[20] saout_wm1_x4_128x8m81_0/bb[31] saout_wm1_x4_128x8m81_0/bb[29]
+ saout_wm1_x4_128x8m81_0/bb[13] saout_wm1_x4_128x8m81_0/b[15] saout_wm1_x4_128x8m81_0/b[25]
+ saout_wm1_x4_128x8m81_0/b[9] saout_wm1_x4_128x8m81_0/bb[22] saout_wm1_x4_128x8m81_0/b[4]
+ saout_wm1_x4_128x8m81_0/b[26] saout_wm1_x4_128x8m81_0/b[13] saout_wm1_x4_128x8m81_0/b[7]
+ saout_wm1_x4_128x8m81_0/b[19] saout_wm1_x4_128x8m81_0/b[29] saout_wm1_x4_128x8m81_0/bb[2]
+ saout_wm1_x4_128x8m81_0/bb[9] saout_wm1_x4_128x8m81_0/b[0] saout_wm1_x4_128x8m81_0/b[11]
+ saout_wm1_x4_128x8m81_0/b[28] saout_wm1_x4_128x8m81_0/b[14] saout_wm1_x4_128x8m81_0/bb[26]
+ saout_wm1_x4_128x8m81_0/bb[17] saout_wm1_x4_128x8m81_0/bb[16] saout_wm1_x4_128x8m81_0/b[22]
+ saout_wm1_x4_128x8m81_0/bb[28] saout_wm1_x4_128x8m81_0/b[17] saout_wm1_x4_128x8m81_0/bb[10]
+ saout_wm1_x4_128x8m81_0/b[31] saout_wm1_x4_128x8m81_0/bb[25] saout_wm1_x4_128x8m81_0/bb[19]
+ saout_wm1_x4_128x8m81_0/bb[3] saout_wm1_x4_128x8m81_0/bb[20] VSS saout_wm1_x4_128x8m81_0/b[6]
+ VDD col_128a_128x8m81
Xsaout_wm1_x4_128x8m81_0 saout_wm1_x4_128x8m81_0/ypass[0] saout_wm1_x4_128x8m81_0/ypass[1]
+ saout_wm1_x4_128x8m81_0/ypass[3] saout_wm1_x4_128x8m81_0/ypass[4] saout_wm1_x4_128x8m81_0/ypass[5]
+ saout_wm1_x4_128x8m81_0/ypass[2] saout_wm1_x4_128x8m81_0/b[1] saout_wm1_x4_128x8m81_0/b[4]
+ saout_wm1_x4_128x8m81_0/b[7] saout_wm1_x4_128x8m81_0/b[10] saout_wm1_x4_128x8m81_0/b[13]
+ saout_wm1_x4_128x8m81_0/b[16] saout_wm1_x4_128x8m81_0/b[19] saout_wm1_x4_128x8m81_0/b[22]
+ saout_wm1_x4_128x8m81_0/b[25] saout_wm1_x4_128x8m81_0/b[28] saout_wm1_x4_128x8m81_0/b[31]
+ saout_wm1_x4_128x8m81_0/din[1] saout_wm1_x4_128x8m81_0/din[3] saout_wm1_x4_128x8m81_0/din[2]
+ saout_wm1_x4_128x8m81_0/din[0] saout_wm1_x4_128x8m81_0/q[0] saout_wm1_x4_128x8m81_0/q[1]
+ saout_wm1_x4_128x8m81_0/q[2] saout_wm1_x4_128x8m81_0/q[3] saout_wm1_x4_128x8m81_0/b[29]
+ saout_wm1_x4_128x8m81_0/b[26] saout_wm1_x4_128x8m81_0/b[23] saout_wm1_x4_128x8m81_0/b[20]
+ saout_wm1_x4_128x8m81_0/b[17] saout_wm1_x4_128x8m81_0/b[14] saout_wm1_x4_128x8m81_0/b[11]
+ saout_wm1_x4_128x8m81_0/b[8] saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/b[2]
+ saout_wm1_x4_128x8m81_0/bb[0] saout_wm1_x4_128x8m81_0/bb[1] saout_wm1_x4_128x8m81_0/bb[2]
+ saout_wm1_x4_128x8m81_0/bb[3] saout_wm1_x4_128x8m81_0/bb[4] saout_wm1_x4_128x8m81_0/bb[5]
+ saout_wm1_x4_128x8m81_0/bb[6] saout_wm1_x4_128x8m81_0/bb[7] saout_wm1_x4_128x8m81_0/bb[8]
+ saout_wm1_x4_128x8m81_0/bb[9] saout_wm1_x4_128x8m81_0/bb[10] saout_wm1_x4_128x8m81_0/bb[11]
+ saout_wm1_x4_128x8m81_0/bb[12] saout_wm1_x4_128x8m81_0/bb[13] saout_wm1_x4_128x8m81_0/bb[14]
+ saout_wm1_x4_128x8m81_0/bb[15] saout_wm1_x4_128x8m81_0/bb[16] saout_wm1_x4_128x8m81_0/bb[17]
+ saout_wm1_x4_128x8m81_0/bb[18] saout_wm1_x4_128x8m81_0/bb[19] saout_wm1_x4_128x8m81_0/bb[20]
+ saout_wm1_x4_128x8m81_0/bb[21] saout_wm1_x4_128x8m81_0/bb[22] saout_wm1_x4_128x8m81_0/bb[23]
+ saout_wm1_x4_128x8m81_0/bb[24] saout_wm1_x4_128x8m81_0/bb[25] saout_wm1_x4_128x8m81_0/bb[26]
+ saout_wm1_x4_128x8m81_0/bb[27] saout_wm1_x4_128x8m81_0/bb[28] saout_wm1_x4_128x8m81_0/bb[29]
+ saout_wm1_x4_128x8m81_0/bb[30] saout_wm1_x4_128x8m81_0/bb[31] saout_wm1_x4_128x8m81_0/b[30]
+ saout_wm1_x4_128x8m81_0/b[27] saout_wm1_x4_128x8m81_0/b[24] saout_wm1_x4_128x8m81_0/b[15]
+ saout_wm1_x4_128x8m81_0/b[12] saout_wm1_x4_128x8m81_0/b[9] saout_wm1_x4_128x8m81_0/b[21]
+ saout_wm1_x4_128x8m81_0/b[0] saout_wm1_x4_128x8m81_0/b[3] saout_wm1_x4_128x8m81_0/b[6]
+ saout_wm1_x4_128x8m81_0/b[18] saout_wm1_x4_128x8m81_0/pcb[0] saout_wm1_x4_128x8m81_0/pcb[1]
+ saout_wm1_x4_128x8m81_0/pcb[3] saout_wm1_x4_128x8m81_0/pcb[2] saout_wm1_x4_128x8m81_0/WEN[3]
+ saout_wm1_x4_128x8m81_0/WEN[2] saout_wm1_x4_128x8m81_0/WEN[1] saout_wm1_x4_128x8m81_0/WEN[0]
+ saout_wm1_x4_128x8m81_0/bb[20] saout_wm1_x4_128x8m81_0/b[24] saout_wm1_x4_128x8m81_0/bb[17]
+ saout_wm1_x4_128x8m81_0/a_15501_29383# saout_wm1_x4_128x8m81_0/bb[24] saout_wm1_x4_128x8m81_0/bb[25]
+ saout_wm1_x4_128x8m81_0/bb[5] saout_wm1_x4_128x8m81_0/bb[30] saout_wm1_x4_128x8m81_0/b[20]
+ VSS saout_wm1_x4_128x8m81_0/a_15261_28608# saout_wm1_x4_128x8m81_0/bb[1] saout_wm1_x4_128x8m81_0/b[23]
+ saout_wm1_x4_128x8m81_0/bb[10] saout_wm1_x4_128x8m81_0/bb[23] saout_wm1_x4_128x8m81_0/bb[22]
+ saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_0/wen_wm1_128x8m81_0/wen saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_0/WEN
+ saout_wm1_x4_128x8m81_0/b[2] saout_wm1_x4_128x8m81_0/men saout_wm1_x4_128x8m81_0/b[6]
+ saout_wm1_x4_128x8m81_0/bb[15] saout_wm1_x4_128x8m81_0/a_4701_29383# saout_wm1_x4_128x8m81_0/bb[3]
+ VSS saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/GWE saout_wm1_x4_128x8m81_0/bb[16]
+ saout_wm1_x4_128x8m81_0/bb[29] saout_wm1_x4_128x8m81_0/b[28] saout_wm1_x4_128x8m81_0/b[13]
+ saout_wm1_x4_128x8m81_0/bb[4] saout_wm1_x4_128x8m81_0/b[9] saout_wm1_x4_128x8m81_0/bb[31]
+ saout_wm1_x4_128x8m81_0/bb[12] saout_wm1_x4_128x8m81_0/a_4461_28608# saout_wm1_x4_128x8m81_0/b[10]
+ saout_wm1_x4_128x8m81_0/b[4] saout_wm1_x4_128x8m81_0/a_15501_28608# saout_wm1_x4_128x8m81_0/bb[0]
+ saout_wm1_x4_128x8m81_0/bb[11] saout_wm1_x4_128x8m81_0/bb[18] saout_wm1_x4_128x8m81_0/b[19]
+ saout_wm1_x4_128x8m81_0/b[15] saout_wm1_x4_128x8m81_0/b[7] saout_wm1_x4_128x8m81_0/bb[26]
+ saout_wm1_x4_128x8m81_0/bb[7] saout_wm1_x4_128x8m81_0/bb[6] saout_wm1_x4_128x8m81_0/ypass[6]
+ saout_wm1_x4_128x8m81_0/b[11] saout_wm1_x4_128x8m81_0/b[16] saout_wm1_x4_128x8m81_0/b[14]
+ saout_wm1_x4_128x8m81_0/ypass[7] saout_wm1_x4_128x8m81_0/b[8] saout_wm1_x4_128x8m81_0/b[31]
+ saout_wm1_x4_128x8m81_0/bb[8] saout_wm1_x4_128x8m81_0/bb[9] saout_wm1_x4_128x8m81_0/b[17]
+ saout_wm1_x4_128x8m81_0/bb[21] saout_wm1_x4_128x8m81_0/a_15261_29383# saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/GWEN
+ saout_wm1_x4_128x8m81_0/b[0] VSS saout_wm1_x4_128x8m81_0/b[30] VSS VSS saout_wm1_x4_128x8m81_0/b[1]
+ saout_wm1_x4_128x8m81_0/b[29] saout_wm1_x4_128x8m81_0/b[5] saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ saout_wm1_x4_128x8m81_0/a_4701_28608# saout_wm1_x4_128x8m81_0/b[25] saout_wm1_x4_128x8m81_0/bb[28]
+ saout_wm1_x4_128x8m81_0/b[26] saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_0/pcb saout_wm1_x4_128x8m81_0/bb[27]
+ saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/sa_128x8m81_0/pcb saout_wm1_x4_128x8m81_0/bb[2]
+ saout_wm1_x4_128x8m81_0/b[3] saout_wm1_x4_128x8m81_0/b[18] saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_1/sa_128x8m81_0/pcb
+ saout_wm1_x4_128x8m81_0/b[22] saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb
+ saout_wm1_x4_128x8m81_0/bb[19] saout_wm1_x4_128x8m81_0/b[27] saout_wm1_x4_128x8m81_0/bb[14]
+ saout_wm1_x4_128x8m81_0/b[21] saout_wm1_x4_128x8m81_0/a_4461_29383# VSS saout_wm1_x4_128x8m81_0/bb[13]
+ VDD saout_wm1_x4_128x8m81_0/b[12] saout_wm1_x4_128x8m81
Xdcap_103_novia_128x8m81_0[0] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[1] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[2] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[3] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[4] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[5] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[6] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[7] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[8] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[9] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[10] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[11] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[12] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[13] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[14] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[15] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[16] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[17] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[18] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[19] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[20] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[21] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[22] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[23] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[24] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[25] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[26] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[27] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[28] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[29] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[30] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[31] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[32] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[33] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[34] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[35] VDD VDD VSS dcap_103_novia_128x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_128x8m81 a_n36_52# a_444_n42# a_246_342# a_126_298#
+ m3_n36_330# a_36_n42# w_n68_622# VSUBS
X0 a_444_206# a_n36_52# a_444_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X1 a_36_206# a_n36_52# a_36_n42# VSUBS nmos_6p0 w=0.6u l=0.77u
X2 a_126_298# a_126_298# a_36_206# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X3 a_444_206# a_246_342# a_126_298# w_n68_622# pmos_6p0 w=0.6u l=0.6u
X4 a_246_342# a_126_298# a_36_206# VSUBS nmos_6p0 w=0.95u l=0.6u
X5 a_444_206# a_246_342# a_246_342# VSUBS nmos_6p0 w=0.95u l=0.6u
.ends

.subckt ypass_gate_128x8m81_0 vss bb db ypass pcb vdd m3_n1_4331# b m3_n1_1708# m3_n1_1160#
+ m3_n1_2030# m3_n1_3366# m3_n1_2352# m3_n1_3688# m3_n1_4009# m3_n1_2674# d a_66_539#
+ pmos_5p0431059054871_128x8m81_2/D
Xnmos_5p0431059054870_128x8m81_0 pmos_5p0431059054871_128x8m81_2/D a_66_539# bb vss
+ nmos_5p0431059054870_128x8m81
Xnmos_5p0431059054870_128x8m81_1 d a_66_539# b vss nmos_5p0431059054870_128x8m81
Xpmos_5p0431059054871_128x8m81_1 vdd b pcb bb pmos_5p0431059054871_128x8m81
Xpmos_5p0431059054871_128x8m81_0 vdd d nmos_5p0431059054872_128x8m81_0/D b pmos_5p0431059054871_128x8m81
Xpmos_5p0431059054871_128x8m81_2 vdd pmos_5p0431059054871_128x8m81_2/D nmos_5p0431059054872_128x8m81_0/D
+ bb pmos_5p0431059054871_128x8m81
Xnmos_5p0431059054872_128x8m81_0 nmos_5p0431059054872_128x8m81_0/D a_66_539# vss a_66_539#
+ vss nmos_5p0431059054872_128x8m81
X0 nmos_5p0431059054872_128x8m81_0/D a_66_539# vdd vdd pmos_3p3 w=1.485u l=0.6u
X1 vdd pcb bb vdd pmos_3p3 w=3.41u l=0.6u
X2 bb pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
X3 vdd pcb b vdd pmos_3p3 w=3.41u l=0.6u
X4 vdd a_66_539# nmos_5p0431059054872_128x8m81_0/D vdd pmos_3p3 w=1.485u l=0.6u
X5 b pcb vdd vdd pmos_3p3 w=3.41u l=0.6u
.ends

.subckt pmos_5p04310590548756_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10.64u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.64u l=0.6u
.ends

.subckt nmos_5p04310590548755_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.38u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.38u l=0.6u
.ends

.subckt nmos_5p04310590548754_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=8.5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=8.5u l=0.6u
.ends

.subckt pmos_5p04310590548753_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.51u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.51u l=0.6u
.ends

.subckt rdummy_128x4_128x8m81 tblhl pcb 018SRAM_cell1_dummy_128x8m81_29/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_1/a_126_298#
+ m3_22279_n11418# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_14/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_17/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_39/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_18/m2_390_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_15/m3_n36_330# 018SRAM_cell1_dummy_R_128x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_0/w_n68_622# 018SRAM_cell1_2x_128x8m81_4/018SRAM_cell1_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_19/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_16/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50# m3_22279_n9439#
+ m3_22426_n25051# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_128x8m81_6/a_246_342#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_20/m2_90_n50# 018SRAM_cell1_dummy_R_128x8m81_5/a_126_298#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_30/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_7/a_246_342# 018SRAM_cell1_dummy_128x8m81_40/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_40/m2_390_n50#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_R_128x8m81_1/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_41/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_21/m2_90_n50# 018SRAM_cell1_dummy_R_128x8m81_2/a_126_298#
+ 018SRAM_cell1_dummy_R_128x8m81_2/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_42/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_4/a_126_298#
+ 018SRAM_cell1_dummy_128x8m81_31/m2_90_n50# DWL 018SRAM_cell1_dummy_128x8m81_43/m2_390_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_5/w_n68_622# 018SRAM_cell1_dummy_128x8m81_41/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_8/a_246_342#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_4/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_44/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_128x8m81_5/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_45/m2_390_n50#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_0/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_22/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_46/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_6/m3_n36_330#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_32/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_47/m2_390_n50# m3_22279_n11740# 018SRAM_cell1_dummy_R_128x8m81_7/m3_n36_330#
+ 018SRAM_cell1_dummy_R_128x8m81_10/a_246_342# 018SRAM_cell1_dummy_R_128x8m81_2/w_n68_622#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_9/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_42/m2_90_n50# 018SRAM_cell1_dummy_R_128x8m81_4/w_n68_622#
+ 018SRAM_cell1_dummy_R_128x8m81_8/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_30/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_9/m3_n36_330#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_23/m2_90_n50#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/m3_n36_330# m3_22279_n9760#
+ 018SRAM_cell1_dummy_128x8m81_31/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_33/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_11/a_246_342# 018SRAM_cell1_dummy_128x8m81_32/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_43/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_33/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_34/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_24/m2_90_n50#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_0/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_35/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_34/m2_90_n50#
+ a_23341_1594# 018SRAM_cell1_dummy_R_128x8m81_12/a_246_342# 018SRAM_cell1_dummy_R_128x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_36/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_44/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_37/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_38/m2_390_n50#
+ w_22685_n22093# 018SRAM_cell1_dummy_128x8m81_25/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_20/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_39/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_9/a_126_298#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/m3_n36_330#
+ m3_22279_n11096# 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_35/m2_90_n50# 018SRAM_cell1_dummy_R_128x8m81_13/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_21/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_45/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_1/a_246_342# 018SRAM_cell1_dummy_128x8m81_22/m2_390_n50#
+ m3_22279_n10082# 018SRAM_cell1_dummy_128x8m81_16/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ vdd 018SRAM_cell1_dummy_128x8m81_23/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_26/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_24/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_36/m2_90_n50#
+ 018SRAM_cell1_2x_128x8m81_4/018SRAM_cell1_128x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_R_128x8m81_14/a_246_342#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_0/m3_n36_330# 018SRAM_cell1_dummy_128x8m81_25/m2_390_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_2/a_246_342# 018SRAM_cell1_dummy_128x8m81_46/m2_90_n50#
+ 018SRAM_cell1_dummy_R_128x8m81_9/w_n68_622# ypass_gate_128x8m81_0_0/d 018SRAM_cell1_dummy_128x8m81_26/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_17/m2_90_n50# VSS a_n257_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_27/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_27/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_6/a_126_298#
+ 018SRAM_cell1_dummy_128x8m81_28/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ m3_22279_n10774# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_37/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_29/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_15/a_246_342#
+ pmos_5p04310590548756_128x8m81_0/S 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_47/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_18/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_28/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_0/a_126_298#
+ 018SRAM_cell1_dummy_R_128x8m81_10/m3_n36_330# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ 018SRAM_cell1_dummy_128x8m81_38/m2_90_n50# 018SRAM_cell1_dummy_R_128x8m81_16/a_246_342#
+ 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50#
+ 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_6/w_n68_622#
+ 018SRAM_cell1_dummy_R_128x8m81_11/m3_n36_330# a_n257_1594# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_R_128x8m81_4/a_246_342# 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_dummy_128x8m81_19/m2_90_n50# m3_22279_n9117# 018SRAM_cell1_dummy_R_128x8m81_12/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50# 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50#
+ vss new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_cell1_dummy_R_128x8m81_13/m3_n36_330#
+ 018SRAM_cell1_dummy_128x8m81_16/m2_390_n50#
X018SRAM_cell1_128x8m81_1 a_n257_1594# 018SRAM_cell1_128x8m81_1/a_444_n42# vss 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_128x8m81
X018SRAM_cell1_dummy_128x8m81_42 a_n257_52# 018SRAM_cell1_dummy_128x8m81_42/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_42/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_20 DWL 018SRAM_cell1_dummy_128x8m81_20/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_20/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_31 DWL 018SRAM_cell1_dummy_128x8m81_31/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_31/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_10 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_10/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_0/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_10/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_0/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_2x_128x8m81_0 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_43 a_n257_52# 018SRAM_cell1_dummy_128x8m81_43/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_43/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_32 a_n257_52# 018SRAM_cell1_dummy_128x8m81_32/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_32/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_10 a_n257_52# 018SRAM_cell1_dummy_128x8m81_10/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_21 DWL 018SRAM_cell1_dummy_128x8m81_21/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_21/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_11 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_11/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_6/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_11/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_6/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
Xypass_gate_128x8m81_0_0 vss ypass_gate_128x8m81_0_0/bb ypass_gate_128x8m81_0_0/db
+ ypass_gate_128x8m81_0_0/ypass ypass_gate_128x8m81_0_0/pcb vdd m3_22279_n9117# ypass_gate_128x8m81_0_0/b
+ m3_22279_n11740# vdd m3_22279_n11418# m3_22279_n10082# m3_22279_n11096# m3_22279_n9760#
+ m3_22279_n9439# m3_22279_n10774# ypass_gate_128x8m81_0_0/d vdd ypass_gate_128x8m81_0_0/bb
+ ypass_gate_128x8m81_0
X018SRAM_cell1_dummy_128x8m81_44 a_n257_52# 018SRAM_cell1_dummy_128x8m81_44/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_44/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_33 a_n257_52# 018SRAM_cell1_dummy_128x8m81_33/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_33/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_2x_128x8m81_1 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_1/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_11 a_n257_52# 018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_22 DWL 018SRAM_cell1_dummy_128x8m81_22/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_22/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
Xpmos_5p04310590548756_128x8m81_0 w_22685_n22093# tblhl pmos_5p04310590548753_128x8m81_0/D
+ pmos_5p04310590548756_128x8m81_0/S pmos_5p04310590548753_128x8m81_0/D pmos_5p04310590548756_128x8m81
Xnmos_5p04310590548755_128x8m81_0 pmos_5p04310590548753_128x8m81_0/D ypass_gate_128x8m81_0_0/d
+ vss ypass_gate_128x8m81_0_0/d vss nmos_5p04310590548755_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_12 DWL ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_12/a_246_342#
+ 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_128x8m81_12/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_2x_128x8m81_2 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_45 a_n257_52# 018SRAM_cell1_dummy_128x8m81_45/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_45/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_34 a_n257_52# 018SRAM_cell1_dummy_128x8m81_34/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_34/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_12 a_n257_52# 018SRAM_cell1_dummy_128x8m81_12/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_12/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_23 DWL 018SRAM_cell1_dummy_128x8m81_23/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_23/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_13 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_13/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_1/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_13/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_46 a_n257_52# 018SRAM_cell1_dummy_128x8m81_46/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_46/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_35 a_n257_52# 018SRAM_cell1_dummy_128x8m81_35/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_35/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_2x_128x8m81_3 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_13 a_n257_52# 018SRAM_cell1_dummy_128x8m81_13/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_13/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_24 DWL 018SRAM_cell1_dummy_128x8m81_24/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_24/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_14 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_14/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_4/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_14/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_4/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_2x_128x8m81_4 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_4/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_4/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_47 a_n257_52# 018SRAM_cell1_dummy_128x8m81_47/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_47/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_36 a_n257_52# 018SRAM_cell1_dummy_128x8m81_36/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_36/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_14 a_n257_52# 018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_14/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_25 DWL 018SRAM_cell1_dummy_128x8m81_25/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_25/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
Xnmos_5p04310590548754_128x8m81_0 tblhl pmos_5p04310590548753_128x8m81_0/D vss pmos_5p04310590548753_128x8m81_0/D
+ vss nmos_5p04310590548754_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_15 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_15/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_15/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_37 a_n257_52# 018SRAM_cell1_dummy_128x8m81_37/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_37/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_2x_128x8m81_5 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_5/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_15 a_n257_52# 018SRAM_cell1_dummy_128x8m81_15/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_26 DWL 018SRAM_cell1_dummy_128x8m81_26/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_26/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_16 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_16/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_2/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_16/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_2/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_2x_128x8m81_6 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_6/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_38 a_n257_52# 018SRAM_cell1_dummy_128x8m81_38/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_38/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_16 DWL 018SRAM_cell1_dummy_128x8m81_16/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_16/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_27 DWL 018SRAM_cell1_dummy_128x8m81_27/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_27/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_17 a_23341_1594# ypass_gate_128x8m81_0_0/bb vss 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# ypass_gate_128x8m81_0_0/b 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_39 a_n257_52# 018SRAM_cell1_dummy_128x8m81_39/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_39/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_2x_128x8m81_7 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_1594# a_n257_1594# vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_128x8m81_1/a_444_n42#
+ vss 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_0/m3_n36_330#
+ 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/m3_n36_330# vss 018SRAM_cell1_128x8m81_1/a_36_n42#
+ x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_dummy_128x8m81_17 DWL 018SRAM_cell1_dummy_128x8m81_17/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_17/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_28 DWL 018SRAM_cell1_dummy_128x8m81_28/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_28/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_18 DWL 018SRAM_cell1_dummy_128x8m81_18/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_18/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_29 DWL 018SRAM_cell1_dummy_128x8m81_29/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_29/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_19 DWL 018SRAM_cell1_dummy_128x8m81_19/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_19/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
Xpmos_5p04310590548753_128x8m81_0 vdd pmos_5p04310590548753_128x8m81_0/D ypass_gate_128x8m81_0_0/d
+ vdd ypass_gate_128x8m81_0_0/d pmos_5p04310590548753_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_0 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_0/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_0/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_0/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_0/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_1 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_1/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_1/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_1/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_2 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_2/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_2/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_2/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_2/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_0 a_n257_52# 018SRAM_cell1_dummy_128x8m81_0/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_0/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_3 DWL ypass_gate_128x8m81_0_0/bb vss 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL ypass_gate_128x8m81_0_0/b 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_1 a_n257_52# 018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_1/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_4 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_4/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_4/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_4/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_4/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_2 a_n257_52# 018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_5 DWL ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_5/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_5/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_5/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_5/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
Xnew_dummyrow_unit_128x8m81_0 new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ DWL new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_0/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_10/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_1/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_2/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_12/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_90_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_3/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_11/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_13/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_14/m2_390_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_6/m2_390_n50#
+ vss new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_15/m2_390_n50# new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ new_dummyrow_unit_128x8m81_0/018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ new_dummyrow_unit_128x8m81
X018SRAM_cell1_dummy_128x8m81_3 a_n257_52# 018SRAM_cell1_dummy_128x8m81_3/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_3/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_6 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_6/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_6/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_6/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_6/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_4 a_n257_52# 018SRAM_cell1_dummy_128x8m81_4/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_4/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_7 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_7/a_246_342#
+ 018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_dummy_R_128x8m81_7/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_5 a_n257_52# 018SRAM_cell1_dummy_128x8m81_5/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_5/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_8 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_8/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_9/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_8/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_9/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_6 a_n257_52# 018SRAM_cell1_dummy_128x8m81_6/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_6/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_R_128x8m81_9 a_23341_1594# ypass_gate_128x8m81_0_0/bb 018SRAM_cell1_dummy_R_128x8m81_9/a_246_342#
+ 018SRAM_cell1_dummy_R_128x8m81_9/a_126_298# 018SRAM_cell1_dummy_R_128x8m81_9/m3_n36_330#
+ ypass_gate_128x8m81_0_0/b 018SRAM_cell1_dummy_R_128x8m81_9/w_n68_622# vss x018SRAM_cell1_dummy_R_128x8m81
X018SRAM_cell1_dummy_128x8m81_7 a_n257_52# 018SRAM_cell1_dummy_128x8m81_7/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_7/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_8 a_n257_52# 018SRAM_cell1_dummy_128x8m81_8/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_8/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_9 a_n257_52# 018SRAM_cell1_dummy_128x8m81_9/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_9/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_40 a_n257_52# 018SRAM_cell1_dummy_128x8m81_40/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_40/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_128x8m81_0 a_n257_52# 018SRAM_cell1_128x8m81_1/a_444_n42# vss 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/a_36_n42# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ vss x018SRAM_cell1_128x8m81
X018SRAM_cell1_dummy_128x8m81_41 a_n257_52# 018SRAM_cell1_dummy_128x8m81_41/m2_90_n50#
+ vss 018SRAM_cell1_dummy_128x8m81_41/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ a_n257_52# 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
X018SRAM_cell1_dummy_128x8m81_30 DWL 018SRAM_cell1_dummy_128x8m81_30/m2_90_n50# vss
+ 018SRAM_cell1_dummy_128x8m81_30/m2_390_n50# 018SRAM_cell1_128x8m81_1/w_n68_622#
+ DWL 018SRAM_cell1_128x8m81_1/w_n68_622# vss x018SRAM_cell1_dummy_128x8m81
.ends

.subckt rarray4_128_128x8m81 WL[9] WL[8] WL[11] WL[15] WL[0] WL[2] WL[10] WL[4] WL[3]
+ WL[14] WL[7] WL[1] WL[13] 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ b[1] 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42# bb[7] 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ b[4] 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42# b[5] 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ WL[6] 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42# b[3] 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ b[7] WL[5] WL[12] BL1B bb[4] b[6] BL VSS b[0] 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
X018SRAM_cell1_2x_128x8m81_190 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_0 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_180 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_191 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_1 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_181 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_170 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_192 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_2 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_160 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_171 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_182 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_193 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_3 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_172 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_150 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_161 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_183 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_194 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_4 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_173 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_184 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_162 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_151 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_140 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_195 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_5 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_185 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_174 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_141 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_152 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_130 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_163 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_196 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_6 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_131 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_142 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_186 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_175 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_164 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_120 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_153 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_197 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_7 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_165 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_121 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_110 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_132 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_187 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_176 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_154 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_143 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_198 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_8 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_188 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_166 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_111 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_100 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_144 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_155 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_177 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_122 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_133 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_199 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_9 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_189 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_178 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_123 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_112 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_156 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_145 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_167 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_134 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_101 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_113 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_168 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_157 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_146 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_135 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_102 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_179 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_124 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_147 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_158 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_136 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_103 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_125 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_169 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_114 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_126 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_148 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_159 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_115 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_137 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_104 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_116 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_127 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_138 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_149 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_105 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_117 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_139 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_106 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_128 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_107 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_129 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_118 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_108 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_119 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_90 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_109 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_80 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_91 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_81 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_70 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_92 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_60 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_93 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_82 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_71 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_250 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_61 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_72 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_83 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_94 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_50 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_251 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_240 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_95 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_73 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_62 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_40 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_51 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_84 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_241 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_230 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_252 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_96 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[10] WL[11] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[10] WL[11] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_74 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_63 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_41 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_30 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_52 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_85 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_231 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_253 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_220 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_242 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_97 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[12] WL[13] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_53 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_75 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_64 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_42 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_31 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_20 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_86 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_86/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_221 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_243 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_232 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_210 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_254 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_98 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[14] WL[15] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[14] WL[15] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_32 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_43 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_76 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_54 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_87 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_65 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_10 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_21 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_200 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_233 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[4] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS b[4] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_211 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_255 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_222 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_244 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_99 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[12] WL[13]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_33 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_66 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_77 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_11 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_22 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_44 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_55 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_88 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_88/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_223 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_245 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_201 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_234 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_212 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_45 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_89 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_99/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_78 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_56 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_67 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_23 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_34 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_12 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_202 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_235 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_213 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_224 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_246 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_13 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_24 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_46 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_35 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_68 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_79 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_57 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_225 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_247 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_203 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_236 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_214 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_69 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_14 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[2] WL[3] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_36 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_47 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_2/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_25 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_58 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_72/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_204 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_237 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS b[6] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_215 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_226 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_248 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_37 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_0/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_48 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_26 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_15 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_59 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_80/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_227 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_35/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS b[1] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_249 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_205 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_7/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_238 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_216 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_16 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_38 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_38/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5]
+ VSS b[3] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_49 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_67/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_27 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[0] WL[1] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_239 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_217 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_71/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_206 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_228 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_39 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_28 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS b[0] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_17 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_3/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[0] WL[1]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_207 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_229 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_218 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[6] WL[7] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_18 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_29 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[4] WL[5] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# bb[7] VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[4] WL[5] VSS b[7] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_219 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# BL1B VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ WL[8] WL[9] VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_208 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[6] WL[7]
+ VSS BL x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_19 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_33/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[2] WL[3]
+ VSS b[5] x018SRAM_cell1_2x_128x8m81
X018SRAM_cell1_2x_128x8m81_209 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622#
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9] VSS
+ 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# 018SRAM_cell1_2x_128x8m81_84/018SRAM_cell1_128x8m81_1/a_444_n42#
+ VSS 018SRAM_cell1_2x_128x8m81_9/018SRAM_cell1_128x8m81_1/w_n68_622# WL[8] WL[9]
+ VSS BL x018SRAM_cell1_2x_128x8m81
.ends

.subckt rcol4_128_128x8m81 WL[6] WL[5] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5]
+ ypass[6] DWL tblhl GWEN ypass[0] WL[11] WL[15] WL[0] WL[2] WL[12] WL[3] WL[4] WL[7]
+ WL[8] WL[9] WL[1] ypass[7] WL[10] WL[13] WL[14] din[4] din[7] q[5] q[6] q[7] din[5]
+ din[6] q[4] pcb[6] pcb[7] pcb[4] vdd WEN[4] WEN[7] pcb[5] WEN[5] WEN[6] a_17474_27175#
+ rarray4_128_128x8m81_0/WL[0] a_17474_27950# rarray4_128_128x8m81_0/WL[1] rarray4_128_128x8m81_0/WL[3]
+ rarray4_128_128x8m81_0/WL[4] rarray4_128_128x8m81_0/WL[7] rarray4_128_128x8m81_0/WL[8]
+ rdummy_128x4_128x8m81_0/VSS a_6674_27175# m3_n1_30537# a_17234_27175# a_6674_27950#
+ a_17234_27950# rarray4_128_128x8m81_0/WL[10] rdummy_128x4_128x8m81_0/pcb rarray4_128_128x8m81_0/WL[11]
+ rarray4_128_128x8m81_0/WL[14] GWE rarray4_128_128x8m81_0/WL[15] saout_R_m2_128x8m81_1/WEN
+ a_6434_27175# saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735# a_6434_27950# rdummy_128x4_128x8m81_0/DWL
+ saout_m2_128x8m81_0/pcb saout_m2_128x8m81_1/sa_128x8m81_0/pcb rdummy_128x4_128x8m81_0/a_23341_1594#
+ men saout_R_m2_128x8m81_1/pcb saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb VDD VSS
Xsaout_m2_128x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] GWEN saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_0/bb[7] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_0/datain saout_m2_128x8m81_0/q saout_m2_128x8m81_0/pcb saout_m2_128x8m81_0/WEN
+ a_17009_27175# a_17234_27175# a_17009_27950# a_17234_27950# GWEN VSS saout_m2_128x8m81_0/b[7]
+ saout_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10# saout_m2_128x8m81_0/b[5]
+ saout_m2_128x8m81_0/sa_128x8m81_0/wep saout_m2_128x8m81_0/mux821_128x8m81_0/a_4992_424#
+ saout_m2_128x8m81_0/b[1] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/bb[4] saout_m2_128x8m81_1/b[6]
+ GWE saout_m2_128x8m81_0/bb[3] saout_m2_128x8m81_0/b[3] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_0/bb[0] saout_m2_128x8m81_0/bb[1] saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ VSS VSS saout_m2_128x8m81_0/bb[6] ypass[7] VDD ypass[1] men saout_m2_128x8m81_0/bb[5]
+ saout_m2_128x8m81_0/b[4] saout_m2_128x8m81_0/pcb ypass[2] ypass[4] VDD VDD ypass[5]
+ VDD ypass[6] ypass[0] ypass[3] VSS saout_m2_128x8m81
Xsaout_m2_128x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] GWEN saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[7] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/datain saout_m2_128x8m81_1/q saout_m2_128x8m81_1/pcb saout_m2_128x8m81_1/WEN
+ a_6209_27175# a_6434_27175# a_6209_27950# a_6434_27950# GWEN saout_m2_128x8m81_1/sacntl_2_128x8m81_0/a_4718_983#
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/a_n80_n10#
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/sa_128x8m81_0/wep saout_m2_128x8m81_1/mux821_128x8m81_0/a_4992_424#
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6]
+ GWE saout_m2_128x8m81_1/bb[3] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/mux821_128x8m81_0/ypass_gate_a_128x8m81_0/b
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[1] saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ saout_m2_128x8m81_1/sacntl_2_128x8m81_0/a_4560_1922# VSS saout_m2_128x8m81_1/b[7]
+ ypass[7] VDD ypass[1] men saout_m2_128x8m81_1/bb[5] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/sa_128x8m81_0/pcb
+ ypass[2] ypass[4] VDD VDD ypass[5] VDD ypass[6] ypass[0] ypass[3] VSS saout_m2_128x8m81
Xrdummy_128x4_128x8m81_0 tblhl rdummy_128x4_128x8m81_0/pcb saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] VDD ypass[1] saout_m2_128x8m81_0/b[7] WL[9] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_0/bb[4] saout_m2_128x8m81_0/bb[7] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[6] WL[13] VSS VDD WL[9] saout_m2_128x8m81_1/b[6]
+ rarray4_128_128x8m81_0/WL[1] WL[1] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7]
+ ypass[6] VSS saout_m2_128x8m81_1/b[7] VDD VSS WL[6] saout_m2_128x8m81_1/bb[3] saout_m2_128x8m81_1/b[7]
+ VDD saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[7] VSS saout_m2_128x8m81_1/b[6]
+ rarray4_128_128x8m81_0/WL[8] saout_m2_128x8m81_0/bb[0] WL[3] saout_m2_128x8m81_1/b[7]
+ saout_m2_128x8m81_1/bb[5] WL[13] rarray4_128_128x8m81_0/WL[4] saout_m2_128x8m81_0/b[1]
+ saout_m2_128x8m81_1/b[7] VDD WL[2] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ VDD saout_m2_128x8m81_1/b[7] rdummy_128x4_128x8m81_0/DWL saout_m2_128x8m81_0/b[3]
+ VDD saout_m2_128x8m81_0/bb[1] saout_R_m2_128x8m81_1/bb[6] VSS rdummy_128x4_128x8m81_0/ypass_gate_128x8m81_0_0/d
+ rarray4_128_128x8m81_0/WL[10] saout_m2_128x8m81_0/b[5] saout_R_m2_128x8m81_1/bb[4]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] WL[4] rarray4_128_128x8m81_0/WL[14]
+ saout_m2_128x8m81_0/bb[4] WL[14] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7]
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/bb[6] WL[12] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_0/b[7] ypass[0] rarray4_128_128x8m81_0/WL[0]
+ VSS VDD saout_R_m2_128x8m81_1/bb[2] VSS saout_m2_128x8m81_1/b[6] VDD WL[6] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] WL[5]
+ saout_R_m2_128x8m81_1/bb[0] saout_m2_128x8m81_1/b[6] WL[7] ypass[5] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_0/bb[1] saout_m2_128x8m81_0/bb[0] saout_m2_128x8m81_1/b[7] VSS
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/bb[3] saout_m2_128x8m81_0/b[1] saout_R_m2_128x8m81_1/bb[6]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[7] saout_m2_128x8m81_1/b[7] saout_R_m2_128x8m81_1/bb[4]
+ saout_m2_128x8m81_1/bb[1] WL[10] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] rdummy_128x4_128x8m81_0/a_23341_1594# VSS VSS saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_0/bb[5] saout_R_m2_128x8m81_1/bb[2] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ saout_m2_128x8m81_1/b[6] VDD saout_m2_128x8m81_1/b[6] saout_R_m2_128x8m81_0/bb[2]
+ saout_R_m2_128x8m81_1/bb[0] VDD saout_m2_128x8m81_0/bb[3] WL[5] ypass[2] WL[15]
+ saout_m2_128x8m81_1/b[7] VSS saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/b[4] VSS
+ saout_R_m2_128x8m81_0/bb[0] ypass[4] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ VDD saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[3] saout_m2_128x8m81_1/b[7]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_0/bb[5] saout_m2_128x8m81_1/b[7] WL[8]
+ VSS WL[0] saout_m2_128x8m81_1/b[7] VSS saout_m2_128x8m81_1/b[6] VDD rdummy_128x4_128x8m81_0/ypass_gate_128x8m81_0_0/d
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7] rdummy_128x4_128x8m81_0/VSS m3_n1_30537#
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/bb[5] saout_R_m2_128x8m81_0/bb[6]
+ VDD saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7] ypass[3] saout_m2_128x8m81_0/b[4]
+ saout_R_m2_128x8m81_0/bb[4] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7] VSS
+ VDD WL[11] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_0/bb[7] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_R_m2_128x8m81_0/bb[2] saout_m2_128x8m81_0/b[3]
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7] VDD rarray4_128_128x8m81_0/WL[7]
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] VSS saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/b[5]
+ saout_m2_128x8m81_1/b[7] VDD rarray4_128_128x8m81_0/WL[11] VSS WL[2] VSS saout_R_m2_128x8m81_0/bb[0]
+ saout_m2_128x8m81_0/bb[4] WL[12] saout_m2_128x8m81_1/b[6] VDD saout_m2_128x8m81_1/b[7]
+ ypass[7] rarray4_128_128x8m81_0/WL[15] saout_m2_128x8m81_1/bb[1] saout_m2_128x8m81_1/b[7]
+ VSS saout_m2_128x8m81_0/bb[6] rarray4_128_128x8m81_0/WL[3] saout_R_m2_128x8m81_0/bb[6]
+ rdummy_128x4_128x8m81
Xrarray4_128_128x8m81_0 WL[9] rarray4_128_128x8m81_0/WL[8] rarray4_128_128x8m81_0/WL[11]
+ rarray4_128_128x8m81_0/WL[15] rarray4_128_128x8m81_0/WL[0] WL[2] rarray4_128_128x8m81_0/WL[10]
+ rarray4_128_128x8m81_0/WL[4] rarray4_128_128x8m81_0/WL[3] rarray4_128_128x8m81_0/WL[14]
+ rarray4_128_128x8m81_0/WL[7] rarray4_128_128x8m81_0/WL[1] WL[13] saout_m2_128x8m81_0/bb[3]
+ saout_m2_128x8m81_0/b[1] saout_R_m2_128x8m81_1/bb[6] saout_m2_128x8m81_0/bb[7] saout_R_m2_128x8m81_1/bb[0]
+ saout_m2_128x8m81_0/bb[4] saout_R_m2_128x8m81_0/bb[4] saout_m2_128x8m81_0/b[5] saout_R_m2_128x8m81_0/bb[6]
+ saout_m2_128x8m81_1/bb[5] saout_R_m2_128x8m81_0/bb[2] saout_m2_128x8m81_1/bb[3]
+ saout_m2_128x8m81_0/bb[5] saout_m2_128x8m81_1/bb[7] saout_m2_128x8m81_0/bb[1] WL[6]
+ saout_R_m2_128x8m81_1/bb[2] saout_m2_128x8m81_1/bb[1] saout_R_m2_128x8m81_0/bb[0]
+ saout_m2_128x8m81_0/b[3] saout_R_m2_128x8m81_1/bb[4] saout_m2_128x8m81_0/b[7] WL[5]
+ WL[12] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_0/b[4] saout_m2_128x8m81_0/bb[6]
+ saout_m2_128x8m81_1/b[7] VSS saout_m2_128x8m81_0/bb[0] VDD rarray4_128_128x8m81
Xdcap_103_novia_128x8m81_0[0] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[1] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[2] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[3] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[4] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[5] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[6] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[7] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[8] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[9] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[10] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[11] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[12] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[13] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[14] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[15] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[16] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[17] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[18] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[19] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[20] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[21] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[22] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[23] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[24] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[25] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[26] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[27] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[28] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[29] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[30] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[31] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[32] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[33] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[34] VDD VDD VSS dcap_103_novia_128x8m81
Xdcap_103_novia_128x8m81_0[35] VDD VDD VSS dcap_103_novia_128x8m81
Xsaout_R_m2_128x8m81_0 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] GWEN saout_R_m2_128x8m81_0/datain saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_0/q saout_R_m2_128x8m81_0/bb[0] saout_R_m2_128x8m81_0/pcb saout_R_m2_128x8m81_0/WEN
+ GWEN saout_R_m2_128x8m81_0/sacntl_2_128x8m81_0/a_4718_983# ypass[5] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_0/sa_128x8m81_0/wep ypass[6] saout_m2_128x8m81_1/b[7] ypass[3]
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] GWE saout_R_m2_128x8m81_0/bb[4]
+ saout_R_m2_128x8m81_0/mux821_128x8m81_0/ypass_gate_128x8m81_4/b saout_R_m2_128x8m81_0/wen_wm1_128x8m81_0/wen
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_R_m2_128x8m81_0/bb[6]
+ a_6900_27175# a_6674_27175# saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735# ypass[7]
+ a_6900_27950# a_6674_27950# saout_R_m2_128x8m81_0/sacntl_2_128x8m81_0/a_4560_1922#
+ saout_R_m2_128x8m81_0/outbuf_oe_128x8m81_0/a_4913_n316# saout_m2_128x8m81_1/b[7]
+ VDD men ypass[1] saout_R_m2_128x8m81_0/bb[2] saout_m2_128x8m81_1/b[6] saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb
+ ypass[4] VDD VDD ypass[0] ypass[2] VDD VSS saout_R_m2_128x8m81
Xsaout_R_m2_128x8m81_1 ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7]
+ men ypass[0] GWEN saout_R_m2_128x8m81_1/datain saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_1/q saout_R_m2_128x8m81_1/bb[0] saout_R_m2_128x8m81_1/pcb saout_R_m2_128x8m81_1/WEN
+ GWEN saout_R_m2_128x8m81_1/sacntl_2_128x8m81_0/a_4718_983# ypass[5] saout_m2_128x8m81_1/b[7]
+ saout_R_m2_128x8m81_1/sa_128x8m81_0/wep ypass[6] saout_m2_128x8m81_1/b[7] ypass[3]
+ saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] GWE saout_R_m2_128x8m81_1/bb[4]
+ saout_R_m2_128x8m81_1/mux821_128x8m81_0/ypass_gate_128x8m81_4/b saout_R_m2_128x8m81_1/wen_wm1_128x8m81_0/wen
+ saout_m2_128x8m81_1/b[7] saout_m2_128x8m81_1/b[6] saout_m2_128x8m81_1/b[7] saout_R_m2_128x8m81_1/bb[6]
+ a_17700_27175# a_17474_27175# saout_m2_128x8m81_1/mux821_128x8m81_0/a_656_7735#
+ ypass[7] a_17700_27950# a_17474_27950# saout_R_m2_128x8m81_1/sacntl_2_128x8m81_0/a_4560_1922#
+ saout_R_m2_128x8m81_1/outbuf_oe_128x8m81_0/a_4913_n316# saout_m2_128x8m81_1/b[7]
+ VDD men ypass[1] saout_R_m2_128x8m81_1/bb[2] saout_m2_128x8m81_1/b[6] saout_R_m2_128x8m81_1/pcb
+ ypass[4] VDD VDD ypass[0] ypass[2] VDD VSS saout_R_m2_128x8m81
.ends

.subckt pmos_5p04310590548796_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1u
.ends

.subckt nmos_1p2$$48629804_128x8m81 a_193_n73# a_n31_n73# nmos_5p04310590548739_128x8m81_0/S
+ nmos_5p04310590548739_128x8m81_0/D VSUBS
Xnmos_5p04310590548739_128x8m81_0 nmos_5p04310590548739_128x8m81_0/D a_n31_n73# nmos_5p04310590548739_128x8m81_0/S
+ a_193_n73# VSUBS nmos_5p04310590548739_128x8m81
.ends

.subckt pmos_5p04310590548791_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=22.68u l=0.6u
.ends

.subckt pmos_1p2$$47815724_128x8m81 pmos_5p04310590548791_128x8m81_0/D w_n286_n141#
+ a_n31_n74# pmos_5p04310590548791_128x8m81_0/S
Xpmos_5p04310590548791_128x8m81_0 w_n286_n141# pmos_5p04310590548791_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548791_128x8m81_0/S pmos_5p04310590548791_128x8m81
.ends

.subckt nmos_5p04310590548790_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=3.02u l=0.6u
.ends

.subckt nmos_1p2$$48302124_128x8m81 a_n31_n74# nmos_5p04310590548790_128x8m81_0/D
+ nmos_5p04310590548790_128x8m81_0/S VSUBS
Xnmos_5p04310590548790_128x8m81_0 nmos_5p04310590548790_128x8m81_0/D a_n31_n74# nmos_5p04310590548790_128x8m81_0/S
+ VSUBS nmos_5p04310590548790_128x8m81
.ends

.subckt nmos_5p04310590548794_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1u
.ends

.subckt nmos_5p04310590548789_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=9.98u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=9.98u l=0.6u
.ends

.subckt nmos_1p2$$48306220_128x8m81 a_417_n74# a_193_n74# nmos_5p04310590548789_128x8m81_0/S
+ nmos_5p04310590548789_128x8m81_0/D a_865_n74# a_641_n74# VSUBS a_n31_n74#
Xnmos_5p04310590548789_128x8m81_0 nmos_5p04310590548789_128x8m81_0/D a_n31_n74# a_865_n74#
+ a_641_n74# nmos_5p04310590548789_128x8m81_0/S a_417_n74# a_193_n74# VSUBS nmos_5p04310590548789_128x8m81
.ends

.subckt pmos_5p04310590548793_128x8m81 a_2464_n44# w_n208_n120# D a_2240_n44# a_3584_n44#
+ a_2016_n44# a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44#
+ a_3808_n44# a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44#
+ a_1344_n44# a_1120_n44# a_2688_n44#
X0 D a_4032_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X1 S a_4256_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X2 S a_224_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X3 D a_448_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X4 D a_0_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X5 S a_2912_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X6 D a_3136_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X7 S a_672_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X8 D a_896_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X9 S a_3360_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X10 S a_2016_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X11 D a_3584_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X12 D a_2240_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X13 S a_2464_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X14 D a_2688_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X15 S a_1120_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X16 D a_1344_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X17 S a_1568_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X18 D a_1792_n44# S w_n208_n120# pmos_6p0 w=18.37u l=0.6u
X19 S a_3808_n44# D w_n208_n120# pmos_6p0 w=18.37u l=0.6u
.ends

.subckt pmos_5p04310590548792_128x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=12.48u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=12.48u l=0.6u
.ends

.subckt pmos_5p04310590548777_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.77u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.77u l=0.6u
.ends

.subckt pmos_1p2$$48623660_128x8m81 pmos_5p04310590548777_128x8m81_0/D a_193_n74#
+ w_n286_n142# a_n31_n74# pmos_5p04310590548777_128x8m81_0/S
Xpmos_5p04310590548777_128x8m81_0 w_n286_n142# pmos_5p04310590548777_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548777_128x8m81_0/S a_193_n74# pmos_5p04310590548777_128x8m81
.ends

.subckt nmos_5p04310590548757_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.36u l=0.6u
.ends

.subckt nmos_1p2$$47342636_128x8m81 nmos_5p04310590548757_128x8m81_0/D nmos_5p04310590548757_128x8m81_0/S
+ a_n31_n73# VSUBS
Xnmos_5p04310590548757_128x8m81_0 nmos_5p04310590548757_128x8m81_0/D a_n31_n73# nmos_5p04310590548757_128x8m81_0/S
+ VSUBS nmos_5p04310590548757_128x8m81
.ends

.subckt pmos_5p04310590548795_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=19.5u l=0.6u
.ends

.subckt pmos_1p2$$48624684_128x8m81 pmos_5p04310590548795_128x8m81_0/S pmos_5p04310590548795_128x8m81_0/D
+ w_n286_n141# a_n31_n74#
Xpmos_5p04310590548795_128x8m81_0 w_n286_n141# pmos_5p04310590548795_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548795_128x8m81_0/S pmos_5p04310590548795_128x8m81
.ends

.subckt nmos_5p04310590548788_128x8m81 a_2464_n44# D a_2240_n44# a_3584_n44# a_2016_n44#
+ a_3360_n44# a_3136_n44# a_2912_n44# a_0_n44# a_4256_n44# a_4032_n44# a_3808_n44#
+ a_896_n44# a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44#
+ a_1120_n44# a_2688_n44# VSUBS
X0 S a_4256_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X1 S a_224_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X2 D a_448_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X3 D a_0_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X4 S a_2912_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X5 D a_3136_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X6 S a_672_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X7 D a_896_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X8 S a_3360_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X9 S a_2016_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X10 D a_3584_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X11 D a_2240_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X12 S a_2464_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X13 D a_2688_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X14 S a_1120_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X15 D a_1344_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X16 S a_1568_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X17 D a_1792_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
X18 S a_3808_n44# D VSUBS nmos_6p0 w=7.37u l=0.6u
X19 D a_4032_n44# S VSUBS nmos_6p0 w=7.37u l=0.6u
.ends

.subckt nmos_1p2$$48308268_128x8m81 nmos_5p04310590548788_128x8m81_0/D nmos_5p04310590548788_128x8m81_0/a_1792_n44#
+ nmos_5p04310590548788_128x8m81_0/a_1568_n44# nmos_5p04310590548788_128x8m81_0/a_0_n44#
+ nmos_5p04310590548788_128x8m81_0/a_1344_n44# nmos_5p04310590548788_128x8m81_0/a_1120_n44#
+ nmos_5p04310590548788_128x8m81_0/a_2688_n44# nmos_5p04310590548788_128x8m81_0/a_2464_n44#
+ nmos_5p04310590548788_128x8m81_0/a_2240_n44# nmos_5p04310590548788_128x8m81_0/a_2016_n44#
+ nmos_5p04310590548788_128x8m81_0/a_3584_n44# nmos_5p04310590548788_128x8m81_0/a_3360_n44#
+ nmos_5p04310590548788_128x8m81_0/S nmos_5p04310590548788_128x8m81_0/a_3136_n44#
+ nmos_5p04310590548788_128x8m81_0/a_2912_n44# nmos_5p04310590548788_128x8m81_0/a_896_n44#
+ nmos_5p04310590548788_128x8m81_0/a_672_n44# nmos_5p04310590548788_128x8m81_0/a_4256_n44#
+ nmos_5p04310590548788_128x8m81_0/a_448_n44# nmos_5p04310590548788_128x8m81_0/a_4032_n44#
+ nmos_5p04310590548788_128x8m81_0/a_224_n44# nmos_5p04310590548788_128x8m81_0/a_3808_n44#
+ VSUBS
Xnmos_5p04310590548788_128x8m81_0 nmos_5p04310590548788_128x8m81_0/a_2464_n44# nmos_5p04310590548788_128x8m81_0/D
+ nmos_5p04310590548788_128x8m81_0/a_2240_n44# nmos_5p04310590548788_128x8m81_0/a_3584_n44#
+ nmos_5p04310590548788_128x8m81_0/a_2016_n44# nmos_5p04310590548788_128x8m81_0/a_3360_n44#
+ nmos_5p04310590548788_128x8m81_0/a_3136_n44# nmos_5p04310590548788_128x8m81_0/a_2912_n44#
+ nmos_5p04310590548788_128x8m81_0/a_0_n44# nmos_5p04310590548788_128x8m81_0/a_4256_n44#
+ nmos_5p04310590548788_128x8m81_0/a_4032_n44# nmos_5p04310590548788_128x8m81_0/a_3808_n44#
+ nmos_5p04310590548788_128x8m81_0/a_896_n44# nmos_5p04310590548788_128x8m81_0/a_672_n44#
+ nmos_5p04310590548788_128x8m81_0/S nmos_5p04310590548788_128x8m81_0/a_1792_n44#
+ nmos_5p04310590548788_128x8m81_0/a_448_n44# nmos_5p04310590548788_128x8m81_0/a_224_n44#
+ nmos_5p04310590548788_128x8m81_0/a_1568_n44# nmos_5p04310590548788_128x8m81_0/a_1344_n44#
+ nmos_5p04310590548788_128x8m81_0/a_1120_n44# nmos_5p04310590548788_128x8m81_0/a_2688_n44#
+ VSUBS nmos_5p04310590548788_128x8m81
.ends

.subckt nmos_5p04310590548797_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.6u l=1.2u
.ends

.subckt pmos_5p04310590548798_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.89u l=0.6u
.ends

.subckt nmos_5p04310590548787_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.75u l=0.6u
.ends

.subckt nmos_5p04310590548785_128x8m81 D a_0_n44# a_896_n44# a_672_n44# S a_448_n44#
+ a_224_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
X5 S a_1120_n44# D VSUBS nmos_6p0 w=0.89u l=0.6u
X6 D a_1344_n44# S VSUBS nmos_6p0 w=0.89u l=0.6u
.ends

.subckt pmos_5p04310590548786_128x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.48u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.48u l=0.6u
.ends

.subckt pmos_5p04310590548784_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.84u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.84u l=0.6u
.ends

.subckt nmos_5p04310590548782_128x8m81 D a_0_n44# S a_448_n44# a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=2u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=2u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=2u l=0.6u
.ends

.subckt pmos_5p04310590548783_128x8m81 w_n208_n120# D a_0_n44# a_896_n44# a_672_n44#
+ S a_448_n44# a_224_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X5 S a_1120_n44# D w_n208_n120# pmos_6p0 w=2.2u l=0.6u
X6 D a_1344_n44# S w_n208_n120# pmos_6p0 w=2.2u l=0.6u
.ends

.subckt nmos_5p04310590548780_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.2u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.2u l=0.6u
.ends

.subckt pmos_5p04310590548781_128x8m81 w_n208_n120# D a_2016_n44# a_0_n44# a_896_n44#
+ a_672_n44# S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X3 S a_672_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X4 D a_896_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X5 S a_2016_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X6 S a_1120_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X7 D a_1344_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X8 S a_1568_n44# D w_n208_n120# pmos_6p0 w=4.72u l=0.6u
X9 D a_1792_n44# S w_n208_n120# pmos_6p0 w=4.72u l=0.6u
.ends

.subckt nmos_5p04310590548779_128x8m81 D a_2016_n44# a_0_n44# a_896_n44# a_672_n44#
+ S a_1792_n44# a_448_n44# a_224_n44# a_1568_n44# a_1344_n44# a_1120_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X1 D a_448_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X2 D a_0_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X3 S a_672_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X4 D a_896_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X5 S a_2016_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X6 S a_1120_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X7 D a_1344_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
X8 S a_1568_n44# D VSUBS nmos_6p0 w=1.92u l=0.6u
X9 D a_1792_n44# S VSUBS nmos_6p0 w=1.92u l=0.6u
.ends

.subckt wen_v2_128x8m81 clk wen GWE IGWEN vss vdd
Xnmos_5p04310590548785_128x8m81_0 pmos_5p04310590548783_128x8m81_0/D nmos_5p0431059054878_128x8m81_1/S
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S vss nmos_5p0431059054878_128x8m81_1/S
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S
+ vss nmos_5p04310590548785_128x8m81
Xpmos_5p04310590548786_128x8m81_0 vdd pmos_5p04310590548786_128x8m81_0/D wen wen wen
+ vdd wen wen wen pmos_5p04310590548786_128x8m81
Xpmos_1p2$$202586156_128x8m81_0 pmos_5p04310590548741_128x8m81_1/D vdd vdd pmos_5p04310590548714_128x8m81_2/S
+ pmos_1p2$$202586156_128x8m81
Xpmos_5p04310590548784_128x8m81_0 vdd pmos_5p04310590548784_128x8m81_0/D pmos_5p04310590548714_128x8m81_2/S
+ vdd pmos_5p04310590548714_128x8m81_2/S pmos_5p04310590548784_128x8m81
Xnmos_5p04310590548782_128x8m81_0 pmos_5p04310590548786_128x8m81_0/D wen vss wen wen
+ vss nmos_5p04310590548782_128x8m81
Xpmos_1p2$$202587180_128x8m81_0 nmos_5p0431059054878_128x8m81_2/S vdd pmos_5p04310590548741_128x8m81_1/S
+ nmos_5p0431059054878_128x8m81_4/D pmos_1p2$$202587180_128x8m81
Xpmos_5p04310590548783_128x8m81_0 vdd pmos_5p04310590548783_128x8m81_0/D nmos_5p0431059054878_128x8m81_1/S
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S vdd nmos_5p0431059054878_128x8m81_1/S
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/S
+ pmos_5p04310590548783_128x8m81
Xnmos_5p0431059054878_128x8m81_0 vss pmos_5p04310590548783_128x8m81_0/D nmos_5p0431059054878_128x8m81_1/D
+ vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_0 vdd vdd pmos_5p04310590548783_128x8m81_0/D nmos_5p0431059054878_128x8m81_1/D
+ pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_1 nmos_5p0431059054878_128x8m81_1/D nmos_5p0431059054878_128x8m81_3/D
+ nmos_5p0431059054878_128x8m81_1/S vss nmos_5p0431059054878_128x8m81
Xnmos_5p0431059054878_128x8m81_2 vss wen nmos_5p0431059054878_128x8m81_2/S vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_1 vdd nmos_5p0431059054878_128x8m81_3/D clk vdd pmos_5p04310590548714_128x8m81
Xpmos_5p04310590548714_128x8m81_2 vdd vdd pmos_5p04310590548741_128x8m81_1/S pmos_5p04310590548714_128x8m81_2/S
+ pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_3 nmos_5p0431059054878_128x8m81_3/D clk vss vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_3 vdd vdd wen nmos_5p0431059054878_128x8m81_2/S pmos_5p04310590548714_128x8m81
Xnmos_5p0431059054878_128x8m81_4 nmos_5p0431059054878_128x8m81_4/D nmos_5p0431059054878_128x8m81_3/D
+ vss vss nmos_5p0431059054878_128x8m81
Xpmos_5p04310590548714_128x8m81_4 vdd nmos_5p0431059054878_128x8m81_4/D nmos_5p0431059054878_128x8m81_3/D
+ vdd pmos_5p04310590548714_128x8m81
Xnmos_5p04310590548780_128x8m81_0 pmos_5p04310590548784_128x8m81_0/D pmos_5p04310590548714_128x8m81_2/S
+ vss pmos_5p04310590548714_128x8m81_2/S vss nmos_5p04310590548780_128x8m81
Xpmos_5p04310590548781_128x8m81_0 vdd GWE pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D vdd pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548781_128x8m81
Xpmos_5p04310590548781_128x8m81_1 vdd IGWEN pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D vdd pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548781_128x8m81
Xpmos_5p04310590548741_128x8m81_0 vdd nmos_5p0431059054878_128x8m81_1/D nmos_5p0431059054878_128x8m81_4/D
+ nmos_5p0431059054878_128x8m81_1/S pmos_5p04310590548741_128x8m81
Xpmos_5p04310590548741_128x8m81_1 vdd pmos_5p04310590548741_128x8m81_1/D nmos_5p0431059054878_128x8m81_3/D
+ pmos_5p04310590548741_128x8m81_1/S pmos_5p04310590548741_128x8m81
Xnmos_1p2$$202595372_128x8m81_0 vss pmos_5p04310590548741_128x8m81_1/S pmos_5p04310590548714_128x8m81_2/S
+ vss nmos_1p2$$202595372_128x8m81
Xnmos_1p2$$202595372_128x8m81_1 pmos_5p04310590548741_128x8m81_1/D nmos_5p0431059054878_128x8m81_4/D
+ pmos_5p04310590548741_128x8m81_1/S vss nmos_1p2$$202595372_128x8m81
Xnmos_5p04310590548710_128x8m81_0 pmos_5p04310590548741_128x8m81_1/S nmos_5p0431059054878_128x8m81_3/D
+ nmos_5p0431059054878_128x8m81_2/S vss nmos_5p04310590548710_128x8m81
Xnmos_5p04310590548779_128x8m81_0 GWE pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D vss pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D
+ pmos_5p04310590548783_128x8m81_0/D pmos_5p04310590548783_128x8m81_0/D vss nmos_5p04310590548779_128x8m81
Xnmos_5p04310590548779_128x8m81_1 IGWEN pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D vss pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D
+ pmos_5p04310590548786_128x8m81_0/D pmos_5p04310590548786_128x8m81_0/D vss nmos_5p04310590548779_128x8m81
Xpmos_5p04310590548720_128x8m81_0 vdd pmos_5p04310590548784_128x8m81_0/D nmos_5p0431059054878_128x8m81_3/D
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_3/D pmos_5p04310590548720_128x8m81
Xnmos_5p04310590548739_128x8m81_0 pmos_5p04310590548784_128x8m81_0/D nmos_5p0431059054878_128x8m81_4/D
+ nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_4/D vss nmos_5p04310590548739_128x8m81
Xnmos_1p2$$202596396_128x8m81_0 vss pmos_5p04310590548714_128x8m81_2/S pmos_5p04310590548741_128x8m81_1/D
+ vss nmos_1p2$$202596396_128x8m81
.ends

.subckt pmos_5p04310590548778_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=0.9u l=1.2u
.ends

.subckt pmos_1p2$$47330348_128x8m81 pmos_5p04310590548741_128x8m81_0/S pmos_5p04310590548741_128x8m81_0/D
+ a_n31_n73# w_n286_n141#
Xpmos_5p04310590548741_128x8m81_0 w_n286_n141# pmos_5p04310590548741_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548741_128x8m81_0/S pmos_5p04310590548741_128x8m81
.ends

.subckt gen_512x8_128x8m81 tblhl cen clk WEN GWE pmos_5p04310590548792_128x8m81_0/D
+ wen_v2_128x8m81_0/wen wen_v2_128x8m81_0/IGWEN VSS men VDD
Xpmos_5p04310590548796_128x8m81_0 VDD pmos_5p04310590548796_128x8m81_0/D pmos_5p04310590548778_128x8m81_1/D
+ VDD pmos_5p04310590548796_128x8m81
Xnmos_1p2$$48629804_128x8m81_0 nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S VSS pmos_5p04310590548751_128x8m81_0/D
+ VSS nmos_1p2$$48629804_128x8m81
Xpmos_1p2$$47815724_128x8m81_7 VDD VDD pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81
Xnmos_1p2$$48302124_128x8m81_0 pmos_5p04310590548798_128x8m81_0/D pmos_1p2$$48623660_128x8m81_0/pmos_5p04310590548777_128x8m81_0/D
+ VSS VSS nmos_1p2$$48302124_128x8m81
Xnmos_5p04310590548794_128x8m81_0 pmos_5p04310590548796_128x8m81_0/D pmos_5p04310590548778_128x8m81_1/D
+ VSS VSS nmos_5p04310590548794_128x8m81
Xpmos_1p2$$46285868_128x8m81_0 VDD VDD nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S
+ nmos_1p2$$46563372_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D pmos_1p2$$46285868_128x8m81
Xnmos_1p2$$48306220_128x8m81_0 pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S VSS pmos_5p04310590548792_128x8m81_0/D
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ VSS pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S nmos_1p2$$48306220_128x8m81
Xnmos_1p2$$46563372_128x8m81_0 nmos_1p2$$46563372_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ VSS nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S VSS nmos_1p2$$46563372_128x8m81
Xpmos_1p2$$46285868_128x8m81_1 nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ VDD nmos_1p2$$46563372_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D cen pmos_1p2$$46285868_128x8m81
Xnmos_1p2$$46563372_128x8m81_1 pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S nmos_1p2$$46563372_128x8m81_0/nmos_5p0431059054878_128x8m81_0/D
+ VSS nmos_1p2$$46563372_128x8m81
Xnmos_1p2$$46563372_128x8m81_2 VSS pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D VSS nmos_1p2$$46563372_128x8m81
Xpmos_1p2$$46273580_128x8m81_0 VDD pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D
+ pmos_5p04310590548751_128x8m81_0/D pmos_5p04310590548751_128x8m81_0/D VDD pmos_1p2$$46273580_128x8m81
Xpmos_5p04310590548793_128x8m81_0 pmos_5p04310590548792_128x8m81_0/D VDD men pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D VDD pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548793_128x8m81
Xnmos_1p2$$46551084_128x8m81_0 cen nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S
+ nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S VSS nmos_1p2$$46551084_128x8m81
Xpmos_5p04310590548792_128x8m81_0 VDD pmos_5p04310590548792_128x8m81_0/D pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S VDD pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_5p04310590548792_128x8m81
Xpmos_1p2$$48623660_128x8m81_0 pmos_1p2$$48623660_128x8m81_0/pmos_5p04310590548777_128x8m81_0/D
+ pmos_5p04310590548798_128x8m81_0/D VDD pmos_5p04310590548798_128x8m81_0/D VDD pmos_1p2$$48623660_128x8m81
Xnmos_1p2$$47342636_128x8m81_0 nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S
+ VSS clk VSS nmos_1p2$$47342636_128x8m81
Xnmos_1p2$$47342636_128x8m81_1 VSS nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S
+ men VSS nmos_1p2$$47342636_128x8m81
Xpmos_5p04310590548751_128x8m81_0 VDD pmos_5p04310590548751_128x8m81_0/D nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ VDD nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S pmos_5p04310590548751_128x8m81
Xpmos_1p2$$48624684_128x8m81_0 VDD pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S
+ VDD pmos_5p04310590548751_128x8m81_0/D pmos_1p2$$48624684_128x8m81
Xnmos_1p2$$48308268_128x8m81_0 men pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ VSS pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D pmos_5p04310590548792_128x8m81_0/D
+ VSS nmos_1p2$$48308268_128x8m81
Xpmos_1p2$$48624684_128x8m81_1 VDD pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S
+ VDD pmos_1p2$$48623660_128x8m81_0/pmos_5p04310590548777_128x8m81_0/D pmos_1p2$$48624684_128x8m81
Xpmos_1p2$$48624684_128x8m81_2 pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S
+ VDD VDD clk pmos_1p2$$48624684_128x8m81
Xnmos_5p04310590548797_128x8m81_0 pmos_5p04310590548778_128x8m81_0/D clk VSS VSS nmos_5p04310590548797_128x8m81
Xpmos_5p04310590548798_128x8m81_0 VDD pmos_5p04310590548798_128x8m81_0/D pmos_5p04310590548796_128x8m81_0/D
+ VDD pmos_5p04310590548798_128x8m81
Xpmos_1p2$$47815724_128x8m81_0 VDD VDD tblhl pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81
Xnmos_5p04310590548787_128x8m81_0 pmos_5p04310590548798_128x8m81_0/D pmos_5p04310590548796_128x8m81_0/D
+ VSS VSS nmos_5p04310590548787_128x8m81
Xwen_v2_128x8m81_0 clk wen_v2_128x8m81_0/wen wen_v2_128x8m81_0/GWE wen_v2_128x8m81_0/IGWEN
+ VSS VDD wen_v2_128x8m81
Xnmos_5p04310590548797_128x8m81_1 pmos_5p04310590548778_128x8m81_1/D pmos_5p04310590548778_128x8m81_0/D
+ VSS VSS nmos_5p04310590548797_128x8m81
Xpmos_1p2$$47815724_128x8m81_1 pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S
+ VDD pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S VDD pmos_1p2$$47815724_128x8m81
Xpmos_5p04310590548778_128x8m81_0 VDD pmos_5p04310590548778_128x8m81_0/D clk VDD pmos_5p04310590548778_128x8m81
Xpmos_1p2$$47815724_128x8m81_2 pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S
+ VDD tblhl VDD pmos_1p2$$47815724_128x8m81
Xpmos_5p04310590548778_128x8m81_1 VDD pmos_5p04310590548778_128x8m81_1/D pmos_5p04310590548778_128x8m81_0/D
+ VDD pmos_5p04310590548778_128x8m81
Xpmos_1p2$$47815724_128x8m81_3 VDD VDD pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81
Xpmos_1p2$$47815724_128x8m81_4 pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ VDD pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S VDD pmos_1p2$$47815724_128x8m81
Xpmos_1p2$$47815724_128x8m81_5 pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S
+ VDD pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S VDD pmos_1p2$$47815724_128x8m81
Xpmos_1p2$$47330348_128x8m81_0 nmos_1p2$$46563372_128x8m81_1/nmos_5p0431059054878_128x8m81_0/S
+ pmos_1p2$$46273580_128x8m81_0/pmos_5p0431059054873_128x8m81_0/D nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S
+ VDD pmos_1p2$$47330348_128x8m81
Xpmos_1p2$$47815724_128x8m81_6 VDD VDD pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S
+ pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$47815724_128x8m81
X0 VSS pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S a_11293_484# VSS nmos_6p0 w=18.145u l=0.6u
X1 a_9646_262# pmos_1p2$$48623660_128x8m81_0/pmos_5p04310590548777_128x8m81_0/D VSS VSS nmos_6p0 w=22.68u l=0.6u
X2 pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S a_10845_484# VSS nmos_6p0 w=18.145u l=0.6u
X3 a_12578_3205# tblhl pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S VSS nmos_6p0 w=4.54u l=0.6u
X4 pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S pmos_5p04310590548751_128x8m81_0/D a_9870_262# VSS nmos_6p0 w=22.68u l=0.6u
X5 a_11293_484# pmos_1p2$$48624684_128x8m81_2/pmos_5p04310590548795_128x8m81_0/S pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S VSS nmos_6p0 w=18.145u l=0.6u
X6 a_12130_3205# pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S VSS VSS nmos_6p0 w=4.54u l=0.6u
X7 a_10845_484# pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S VSS VSS nmos_6p0 w=18.145u l=0.6u
X8 pmos_1p2$$47815724_128x8m81_3/pmos_5p04310590548791_128x8m81_0/S tblhl a_12130_3205# VSS nmos_6p0 w=4.54u l=0.6u
X9 nmos_1p2$$47342636_128x8m81_1/nmos_5p04310590548757_128x8m81_0/S clk a_5174_6131# VDD pmos_6p0 w=2.28u l=0.595u
X10 VSS pmos_1p2$$47815724_128x8m81_7/pmos_5p04310590548791_128x8m81_0/S a_12578_3205# VSS nmos_6p0 w=4.54u l=0.6u
X11 a_9870_262# clk a_9646_262# VSS nmos_6p0 w=22.68u l=0.6u
X12 a_5174_6131# men VDD VDD pmos_6p0 w=2.28u l=0.595u
.ends

.subckt nmos_1p2$$46551084_157_128x8m81 nmos_5p04310590548710_128x8m81_0/D a_n31_n74#
+ nmos_5p04310590548710_128x8m81_0/S VSUBS
Xnmos_5p04310590548710_128x8m81_0 nmos_5p04310590548710_128x8m81_0/D a_n31_n74# nmos_5p04310590548710_128x8m81_0/S
+ VSUBS nmos_5p04310590548710_128x8m81
.ends

.subckt pmos_5p04310590548762_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=4.54u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=4.54u l=0.6u
.ends

.subckt pmos_1p2$$47331372_128x8m81 pmos_5p04310590548762_128x8m81_0/D a_n30_n74#
+ pmos_5p04310590548762_128x8m81_0/S w_n286_n142# a_194_n74#
Xpmos_5p04310590548762_128x8m81_0 w_n286_n142# pmos_5p04310590548762_128x8m81_0/D
+ a_n30_n74# pmos_5p04310590548762_128x8m81_0/S a_194_n74# pmos_5p04310590548762_128x8m81
.ends

.subckt pmos_1p2$$46285868_160_128x8m81 pmos_5p04310590548714_128x8m81_0/S a_n31_n74#
+ w_n286_n142# pmos_5p04310590548714_128x8m81_0/D
Xpmos_5p04310590548714_128x8m81_0 w_n286_n142# pmos_5p04310590548714_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548714_128x8m81_0/S pmos_5p04310590548714_128x8m81
.ends

.subckt pmos_1p2$$47330348_161_128x8m81 pmos_5p04310590548741_128x8m81_0/S pmos_5p04310590548741_128x8m81_0/D
+ a_n31_191# w_n286_n141#
Xpmos_5p04310590548741_128x8m81_0 w_n286_n141# pmos_5p04310590548741_128x8m81_0/D
+ a_n31_191# pmos_5p04310590548741_128x8m81_0/S pmos_5p04310590548741_128x8m81
.ends

.subckt nmos_5p04310590548763_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=1.82u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=1.82u l=0.6u
.ends

.subckt nmos_1p2$$47329324_128x8m81 a_194_n74# nmos_5p04310590548763_128x8m81_0/D
+ nmos_5p04310590548763_128x8m81_0/S a_n30_n74# VSUBS
Xnmos_5p04310590548763_128x8m81_0 nmos_5p04310590548763_128x8m81_0/D a_n30_n74# nmos_5p04310590548763_128x8m81_0/S
+ a_194_n74# VSUBS nmos_5p04310590548763_128x8m81
.ends

.subckt alatch_128x8m81 enb en ab a vdd vss
Xnmos_1p2$$46551084_157_128x8m81_0 a en nmos_5p0431059054878_128x8m81_1/S vss nmos_1p2$$46551084_157_128x8m81
Xpmos_1p2$$47331372_128x8m81_0 ab nmos_5p0431059054878_128x8m81_1/S vdd vdd nmos_5p0431059054878_128x8m81_1/S
+ pmos_1p2$$47331372_128x8m81
Xnmos_5p0431059054878_128x8m81_0 vss ab nmos_5p0431059054878_128x8m81_1/D vss nmos_5p0431059054878_128x8m81
Xnmos_5p0431059054878_128x8m81_1 nmos_5p0431059054878_128x8m81_1/D enb nmos_5p0431059054878_128x8m81_1/S
+ vss nmos_5p0431059054878_128x8m81
Xpmos_1p2$$46285868_160_128x8m81_0 nmos_5p0431059054878_128x8m81_1/S enb vdd a pmos_1p2$$46285868_160_128x8m81
Xpmos_1p2$$47330348_161_128x8m81_0 nmos_5p0431059054878_128x8m81_1/S nmos_5p0431059054878_128x8m81_1/D
+ en vdd pmos_1p2$$47330348_161_128x8m81
Xpmos_1p2$$47330348_161_128x8m81_1 nmos_5p0431059054878_128x8m81_1/D vdd ab vdd pmos_1p2$$47330348_161_128x8m81
Xnmos_1p2$$47329324_128x8m81_0 nmos_5p0431059054878_128x8m81_1/S ab vss nmos_5p0431059054878_128x8m81_1/S
+ vss nmos_1p2$$47329324_128x8m81
.ends

.subckt nmos_5p04310590548761_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=4.54u l=0.6u
.ends

.subckt nmos_1p2$$47514668_128x8m81 nmos_5p04310590548761_128x8m81_0/S nmos_5p04310590548761_128x8m81_0/D
+ a_n30_n73# VSUBS
Xnmos_5p04310590548761_128x8m81_0 nmos_5p04310590548761_128x8m81_0/D a_n30_n73# nmos_5p04310590548761_128x8m81_0/S
+ VSUBS nmos_5p04310590548761_128x8m81
.ends

.subckt ypredec1_bot_128x8m81 m1_n14_3279# alatch_128x8m81_0/a alatch_128x8m81_0/en
+ m1_n14_2674# alatch_128x8m81_0/enb m1_n14_2876# m1_n14_3078# m1_n14_3481# pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ m1_n14_2472# pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D alatch_128x8m81_0/vdd
+ alatch_128x8m81_0/vss pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
Xalatch_128x8m81_0 alatch_128x8m81_0/enb alatch_128x8m81_0/en alatch_128x8m81_0/ab
+ alatch_128x8m81_0/a alatch_128x8m81_0/vdd alatch_128x8m81_0/vss alatch_128x8m81
Xpmos_1p2$$46887980_128x8m81_0 pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S pmos_1p2$$46887980_128x8m81
Xpmos_1p2$$46887980_128x8m81_1 pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ alatch_128x8m81_0/ab pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S pmos_1p2$$46887980_128x8m81
Xnmos_1p2$$47514668_128x8m81_0 alatch_128x8m81_0/vss pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D alatch_128x8m81_0/vss
+ nmos_1p2$$47514668_128x8m81
Xnmos_1p2$$47514668_128x8m81_1 alatch_128x8m81_0/vss pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ alatch_128x8m81_0/ab alatch_128x8m81_0/vss nmos_1p2$$47514668_128x8m81
.ends

.subckt nmos_5p04310590548758_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=9.08u l=0.6u
.ends

.subckt pmos_5p04310590548759_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=20u l=0.6u
.ends

.subckt ypredec1_ys_128x8m81 a_254_2184# pmos_5p04310590548759_128x8m81_1/S nmos_5p04310590548758_128x8m81_1/D
+ nmos_5p04310590548758_128x8m81_3/D nmos_5p04310590548758_128x8m81_2/S pmos_5p04310590548759_128x8m81_3/S
+ pmos_5p04310590548759_128x8m81_3/D VSUBS
Xnmos_5p04310590548758_128x8m81_1 nmos_5p04310590548758_128x8m81_1/D pmos_5p04310590548759_128x8m81_0/D
+ pmos_5p04310590548759_128x8m81_1/S VSUBS nmos_5p04310590548758_128x8m81
Xnmos_5p04310590548758_128x8m81_0 pmos_5p04310590548759_128x8m81_3/S pmos_5p04310590548759_128x8m81_0/D
+ nmos_5p04310590548758_128x8m81_1/D VSUBS nmos_5p04310590548758_128x8m81
Xpmos_5p04310590548759_128x8m81_0 pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81_0/D
+ a_254_2184# pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81
Xnmos_5p04310590548758_128x8m81_2 pmos_5p04310590548759_128x8m81_0/D a_254_2184# nmos_5p04310590548758_128x8m81_2/S
+ VSUBS nmos_5p04310590548758_128x8m81
Xpmos_5p04310590548759_128x8m81_1 pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81_3/D
+ pmos_5p04310590548759_128x8m81_0/D pmos_5p04310590548759_128x8m81_1/S pmos_5p04310590548759_128x8m81
Xnmos_5p04310590548758_128x8m81_3 nmos_5p04310590548758_128x8m81_3/D pmos_5p04310590548759_128x8m81_0/D
+ pmos_5p04310590548759_128x8m81_3/S VSUBS nmos_5p04310590548758_128x8m81
Xpmos_5p04310590548759_128x8m81_3 pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81_3/D
+ pmos_5p04310590548759_128x8m81_0/D pmos_5p04310590548759_128x8m81_3/S pmos_5p04310590548759_128x8m81
Xpmos_5p04310590548759_128x8m81_2 pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81_3/S
+ pmos_5p04310590548759_128x8m81_0/D pmos_5p04310590548759_128x8m81_3/D pmos_5p04310590548759_128x8m81
.ends

.subckt nmos_5p04310590548760_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=1.91u l=0.6u
.ends

.subckt pmos_5p04310590548765_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.77u l=0.6u
.ends

.subckt pmos_1p2$$47820844_128x8m81 pmos_5p04310590548765_128x8m81_0/S pmos_5p04310590548765_128x8m81_0/D
+ w_n286_n141# a_n30_n74#
Xpmos_5p04310590548765_128x8m81_0 w_n286_n141# pmos_5p04310590548765_128x8m81_0/D
+ a_n30_n74# pmos_5p04310590548765_128x8m81_0/S pmos_5p04310590548765_128x8m81
.ends

.subckt pmos_5p04310590548764_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.67u l=0.6u
.ends

.subckt pmos_1p2$$47821868_128x8m81 pmos_5p04310590548764_128x8m81_0/S pmos_5p04310590548764_128x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310590548764_128x8m81_0 w_n286_n142# pmos_5p04310590548764_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548764_128x8m81_0/S pmos_5p04310590548764_128x8m81
.ends

.subckt ypredec1_xa_128x8m81 m1_n58_n4290# m1_n58_n4895# pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ m1_n58_n5097# m3_n1_n7124# a_644_n6680# m1_n58_n4492# m1_n58_n4088# a_421_n4311#
+ a_n1_81# a_197_n5120# m1_n58_n4694# pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ M3_M2$$47819820_128x8m81_0/VSUBS
Xnmos_1p2$$46551084_128x8m81_0 pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D M3_M2$$47819820_128x8m81_0/VSUBS
+ M3_M2$$47819820_128x8m81_0/VSUBS nmos_1p2$$46551084_128x8m81
Xnmos_1p2$$46551084_128x8m81_1 M3_M2$$47819820_128x8m81_0/VSUBS pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D
+ pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S M3_M2$$47819820_128x8m81_0/VSUBS
+ nmos_1p2$$46551084_128x8m81
Xnmos_1p2$$46551084_128x8m81_2 pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D M3_M2$$47819820_128x8m81_0/VSUBS
+ M3_M2$$47819820_128x8m81_0/VSUBS nmos_1p2$$46551084_128x8m81
Xpmos_1p2$$47820844_128x8m81_1 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D pmos_1p2$$47820844_128x8m81
Xpmos_1p2$$47820844_128x8m81_0 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D pmos_1p2$$47820844_128x8m81
Xpmos_1p2$$47820844_128x8m81_2 pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D pmos_1p2$$47820844_128x8m81
Xpmos_1p2$$47821868_128x8m81_0 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ a_197_n5120# pmos_1p2$$47821868_128x8m81
Xpmos_1p2$$47821868_128x8m81_2 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ a_644_n6680# pmos_1p2$$47821868_128x8m81
Xpmos_1p2$$47821868_128x8m81_1 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D
+ pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ a_421_n4311# pmos_1p2$$47821868_128x8m81
X0 pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/D a_644_n6680# a_542_n6607# M3_M2$$47819820_128x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X1 a_318_n6607# a_197_n5120# M3_M2$$47819820_128x8m81_0/VSUBS M3_M2$$47819820_128x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
X2 a_542_n6607# a_421_n4311# a_318_n6607# M3_M2$$47819820_128x8m81_0/VSUBS nmos_3p3 w=6.81u l=0.6u
.ends

.subckt ypredec1_xax8_128x8m81 ypredec1_xa_128x8m81_7/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_6/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_2/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_5/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_1/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_0/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xa_128x8m81_6/a_n1_81# a_527_2758# ypredec1_xa_128x8m81_3/a_n1_81# ypredec1_xa_128x8m81_4/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_6100_2150# ypredec1_xa_128x8m81_0/a_n1_81# a_975_1949# a_6324_2352# ypredec1_xa_128x8m81_7/a_n1_81#
+ ypredec1_xa_128x8m81_3/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_751_2554# a_303_2957# VSUBS ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
Xypredec1_xa_128x8m81_1 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_1/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_6324_2352# a_751_2554# a_303_2957# a_6100_2150# VSUBS a_751_2554#
+ a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_0 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_0/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_6324_2352# a_751_2554# a_303_2957# a_527_2758# ypredec1_xa_128x8m81_0/a_n1_81#
+ a_751_2554# a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_2 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_2/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_303_2957# a_751_2554# a_303_2957# a_6100_2150# VSUBS a_751_2554#
+ a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_3 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_3/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_303_2957# a_751_2554# a_303_2957# a_527_2758# ypredec1_xa_128x8m81_3/a_n1_81#
+ a_751_2554# a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_4 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_4/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_6324_2352# a_751_2554# a_303_2957# a_527_2758# ypredec1_xa_128x8m81_4/a_n1_81#
+ a_975_1949# a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_5 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_5/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_6324_2352# a_751_2554# a_303_2957# a_6100_2150# VSUBS a_975_1949#
+ a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_6 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_6/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_303_2957# a_751_2554# a_303_2957# a_6100_2150# ypredec1_xa_128x8m81_6/a_n1_81#
+ a_975_1949# a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
Xypredec1_xa_128x8m81_7 a_527_2758# a_6100_2150# ypredec1_xa_128x8m81_7/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ a_975_1949# VSUBS a_303_2957# a_751_2554# a_303_2957# a_527_2758# ypredec1_xa_128x8m81_7/a_n1_81#
+ a_975_1949# a_6324_2352# ypredec1_xa_128x8m81_7/pmos_1p2$$47821868_128x8m81_2/pmos_5p04310590548764_128x8m81_0/S
+ VSUBS ypredec1_xa_128x8m81
.ends

.subckt pmos_5p04310590548766_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.71u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.71u l=0.6u
.ends

.subckt pmos_1p2$$47109164_128x8m81 a_n31_341# pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ pmos_5p04310590548766_128x8m81_0/D pmos_5p04310590548766_128x8m81_0/S a_193_341#
Xpmos_5p04310590548766_128x8m81_0 pmos_5p04310590548766_128x8m81_0/w_n208_n120# pmos_5p04310590548766_128x8m81_0/D
+ a_n31_341# pmos_5p04310590548766_128x8m81_0/S a_193_341# pmos_5p04310590548766_128x8m81
.ends

.subckt ypredec1_128x8m81 ly[5] ly[4] ly[7] ly[3] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd
+ pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120# ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D
+ pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S
Xypredec1_bot_128x8m81_2 ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ A[1] nmos_5p04310590548760_128x8m81_1/D ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/enb ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ ypredec1_bot_128x8m81
Xypredec1_ys_128x8m81_4 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_6/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[4] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[4] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_5 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_2/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[5] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[5] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_6 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_7/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[6] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[6] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_7 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_1/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[1] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[1] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_8 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_4/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[2] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[2] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_9 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_0/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[3] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[3] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_10 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_6/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[4] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[4] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_11 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_2/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[5] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[5] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_12 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_7/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[6] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[6] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_13 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_3/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[7] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[7] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_14 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_5/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ry[0] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ry[0] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_15 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_3/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[7] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[7] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xnmos_1p2$$47342636_128x8m81_0 ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/alatch_128x8m81_0/enb
+ nmos_5p04310590548760_128x8m81_1/D ypredec1_ys_128x8m81_9/VSUBS nmos_1p2$$47342636_128x8m81
Xnmos_5p04310590548760_128x8m81_0 ypredec1_ys_128x8m81_9/VSUBS clk nmos_5p04310590548760_128x8m81_1/D
+ ypredec1_ys_128x8m81_9/VSUBS nmos_5p04310590548760_128x8m81
Xnmos_5p04310590548760_128x8m81_1 nmos_5p04310590548760_128x8m81_1/D men ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81_9/VSUBS nmos_5p04310590548760_128x8m81
Xypredec1_xax8_128x8m81_0 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_7/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_6/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_2/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_5/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_1/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_0/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_4/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_3/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ ypredec1_xax8_128x8m81
Xypredec1_ys_128x8m81_0 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_5/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[0] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[0] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_1 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_1/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[1] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[1] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_ys_128x8m81_2 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_4/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[2] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[2] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
Xypredec1_bot_128x8m81_0 ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ A[0] nmos_5p04310590548760_128x8m81_1/D ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/enb ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ ypredec1_bot_128x8m81
Xpmos_1p2$$47109164_128x8m81_0 nmos_5p04310590548760_128x8m81_1/D pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/enb pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S
+ nmos_5p04310590548760_128x8m81_1/D pmos_1p2$$47109164_128x8m81
Xypredec1_bot_128x8m81_1 ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ A[2] nmos_5p04310590548760_128x8m81_1/D ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/enb ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_0/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_1/pmos_1p2$$46887980_128x8m81_0/pmos_5p0431059054874_128x8m81_0/D
+ ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd ypredec1_ys_128x8m81_9/VSUBS ypredec1_bot_128x8m81_2/pmos_1p2$$46887980_128x8m81_1/pmos_5p0431059054874_128x8m81_0/S
+ ypredec1_bot_128x8m81
Xypredec1_ys_128x8m81_3 ypredec1_xax8_128x8m81_0/ypredec1_xa_128x8m81_0/pmos_1p2$$47820844_128x8m81_2/pmos_5p04310590548765_128x8m81_0/S
+ ly[3] ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS ypredec1_ys_128x8m81_9/VSUBS
+ ly[3] ypredec1_ys_128x8m81_9/pmos_5p04310590548759_128x8m81_3/D ypredec1_ys_128x8m81_9/VSUBS
+ ypredec1_ys_128x8m81
X0 a_7843_267# clk nmos_5p04310590548760_128x8m81_1/D pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X1 nmos_5p04310590548760_128x8m81_1/D clk a_7395_267# pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X2 a_7395_267# men pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S pmos_3p3 w=2.275u l=0.6u
X3 pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S men a_7843_267# pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/S pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310590548776_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=10.43u l=0.6u
.ends

.subckt pmos_1p2$$47512620_128x8m81 pmos_5p04310590548776_128x8m81_0/S a_n30_n74#
+ pmos_5p04310590548776_128x8m81_0/D w_n286_n142#
Xpmos_5p04310590548776_128x8m81_0 w_n286_n142# pmos_5p04310590548776_128x8m81_0/D
+ a_n30_n74# pmos_5p04310590548776_128x8m81_0/S pmos_5p04310590548776_128x8m81
.ends

.subckt pmos_5p04310590548772_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=11.34u l=0.6u
.ends

.subckt pmos_1p2$$47513644_128x8m81 pmos_5p04310590548772_128x8m81_0/D a_n30_n74#
+ w_n286_n141# pmos_5p04310590548772_128x8m81_0/S
Xpmos_5p04310590548772_128x8m81_0 w_n286_n141# pmos_5p04310590548772_128x8m81_0/D
+ a_n30_n74# pmos_5p04310590548772_128x8m81_0/S pmos_5p04310590548772_128x8m81
.ends

.subckt xpredec1_xa_128x8m81 a_197_n10255# m1_n58_n7539# a_421_n10255# m1_n58_n6933#
+ a_645_n10255# m1_n58_n7135# m1_n58_n6530# m1_n58_n7337# a_n1_81# pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ m1_n58_n6732# pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S M3_M2$$47333420_128x8m81_1/VSUBS
Xpmos_1p2$$47512620_128x8m81_0 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ a_645_n10255# pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47512620_128x8m81
Xpmos_1p2$$47512620_128x8m81_1 pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D
+ a_421_n10255# pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47512620_128x8m81
Xpmos_1p2$$47512620_128x8m81_2 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ a_197_n10255# pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47512620_128x8m81
Xnmos_1p2$$47514668_128x8m81_0 M3_M2$$47333420_128x8m81_1/VSUBS pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D M3_M2$$47333420_128x8m81_1/VSUBS
+ nmos_1p2$$47514668_128x8m81
Xnmos_1p2$$47514668_128x8m81_1 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ M3_M2$$47333420_128x8m81_1/VSUBS pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D
+ M3_M2$$47333420_128x8m81_1/VSUBS nmos_1p2$$47514668_128x8m81
Xnmos_1p2$$47514668_128x8m81_2 M3_M2$$47333420_128x8m81_1/VSUBS pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D M3_M2$$47333420_128x8m81_1/VSUBS
+ nmos_1p2$$47514668_128x8m81
Xpmos_1p2$$47513644_128x8m81_0 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D pmos_1p2$$47513644_128x8m81
Xpmos_1p2$$47513644_128x8m81_1 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S pmos_1p2$$47513644_128x8m81
Xpmos_1p2$$47513644_128x8m81_2 pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47513644_128x8m81_2/pmos_5p04310590548772_128x8m81_0/S pmos_1p2$$47513644_128x8m81
X0 pmos_1p2$$47512620_128x8m81_2/pmos_5p04310590548776_128x8m81_0/D a_645_n10255# a_541_n10182# M3_M2$$47333420_128x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X1 a_317_n10182# a_197_n10255# M3_M2$$47333420_128x8m81_1/VSUBS M3_M2$$47333420_128x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
X2 a_541_n10182# a_421_n10255# a_317_n10182# M3_M2$$47333420_128x8m81_1/VSUBS nmos_3p3 w=12.475u l=0.6u
.ends

.subckt nmos_5p04310590548775_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.58u l=0.6u
.ends

.subckt nmos_1p2$$47336492_128x8m81 nmos_5p04310590548775_128x8m81_0/D a_n31_n74#
+ nmos_5p04310590548775_128x8m81_0/S VSUBS
Xnmos_5p04310590548775_128x8m81_0 nmos_5p04310590548775_128x8m81_0/D a_n31_n74# nmos_5p04310590548775_128x8m81_0/S
+ VSUBS nmos_5p04310590548775_128x8m81
.ends

.subckt pmos_5p04310590548774_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=16.33u l=0.6u
.ends

.subckt pmos_1p2$$47337516_128x8m81 pmos_5p04310590548774_128x8m81_0/D pmos_5p04310590548774_128x8m81_0/S
+ a_n31_n73# w_n286_n141#
Xpmos_5p04310590548774_128x8m81_0 w_n286_n141# pmos_5p04310590548774_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548774_128x8m81_0/S pmos_5p04310590548774_128x8m81
.ends

.subckt xpredec1_bot_128x8m81 pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ alatch_128x8m81_0/a alatch_128x8m81_0/en m1_n106_2472# m1_n106_3279# alatch_128x8m81_0/enb
+ pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D m1_n106_2674# alatch_128x8m81_0/vdd
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/S m1_n106_2876# m1_n106_3078#
+ m1_n106_3481# VSUBS
Xnmos_1p2$$47336492_128x8m81_0 pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D VSUBS VSUBS nmos_1p2$$47336492_128x8m81
Xpmos_1p2$$47337516_128x8m81_0 pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/S pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/S pmos_1p2$$47337516_128x8m81
Xnmos_1p2$$47336492_128x8m81_1 pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ alatch_128x8m81_0/ab VSUBS VSUBS nmos_1p2$$47336492_128x8m81
Xpmos_1p2$$47337516_128x8m81_1 pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/S alatch_128x8m81_0/ab
+ pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/S pmos_1p2$$47337516_128x8m81
Xalatch_128x8m81_0 alatch_128x8m81_0/enb alatch_128x8m81_0/en alatch_128x8m81_0/ab
+ alatch_128x8m81_0/a alatch_128x8m81_0/vdd VSUBS alatch_128x8m81
.ends

.subckt xpredec1_128x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1] A[0]
+ clk pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ w_7178_9364# vss vdd
Xxpredec1_xa_128x8m81_1 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_xa_128x8m81_1/a_n1_81# x[1] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_xa_128x8m81_0 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vss x[3] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_xa_128x8m81_2 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vss x[5] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_bot_128x8m81_0 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ A[0] nmos_5p04310590548760_128x8m81_1/D xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/alatch_128x8m81_0/enb xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vdd vdd xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vss xpredec1_bot_128x8m81
Xxpredec1_xa_128x8m81_3 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_xa_128x8m81_3/a_n1_81# x[7] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_bot_128x8m81_1 xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ A[2] nmos_5p04310590548760_128x8m81_1/D xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/alatch_128x8m81_0/enb xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vdd vdd xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vss xpredec1_bot_128x8m81
Xxpredec1_xa_128x8m81_4 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vss x[2] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_bot_128x8m81_2 xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ A[1] nmos_5p04310590548760_128x8m81_1/D xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/alatch_128x8m81_0/enb xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vdd vdd xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vss xpredec1_bot_128x8m81
Xxpredec1_xa_128x8m81_5 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vss x[0] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_xa_128x8m81_6 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ vss x[4] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xxpredec1_xa_128x8m81_7 xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_0/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_1/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_0/pmos_5p04310590548774_128x8m81_0/D
+ xpredec1_xa_128x8m81_7/a_n1_81# x[6] xpredec1_bot_128x8m81_2/pmos_1p2$$47337516_128x8m81_1/pmos_5p04310590548774_128x8m81_0/D
+ vdd vss xpredec1_xa_128x8m81
Xnmos_1p2$$47342636_128x8m81_0 vss xpredec1_bot_128x8m81_2/alatch_128x8m81_0/enb nmos_5p04310590548760_128x8m81_1/D
+ vss nmos_1p2$$47342636_128x8m81
Xnmos_5p04310590548760_128x8m81_0 vss clk nmos_5p04310590548760_128x8m81_1/D vss nmos_5p04310590548760_128x8m81
Xnmos_5p04310590548760_128x8m81_1 nmos_5p04310590548760_128x8m81_1/D men vss vss nmos_5p04310590548760_128x8m81
Xpmos_1p2$$47109164_128x8m81_0 nmos_5p04310590548760_128x8m81_1/D pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ xpredec1_bot_128x8m81_2/alatch_128x8m81_0/enb vdd nmos_5p04310590548760_128x8m81_1/D
+ pmos_1p2$$47109164_128x8m81
X0 nmos_5p04310590548760_128x8m81_1/D clk a_7553_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X1 a_7553_9505# men vdd w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X2 a_8001_9505# clk nmos_5p04310590548760_128x8m81_1/D w_7178_9364# pmos_3p3 w=2.275u l=0.6u
X3 vdd men a_8001_9505# w_7178_9364# pmos_3p3 w=2.275u l=0.6u
.ends

.subckt pmos_5p04310590548773_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=1.14u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.14u l=0.6u
.ends

.subckt nmos_5p04310590548770_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=7.04u l=0.6u
.ends

.subckt nmos_5p04310590548769_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=5.22u l=0.6u
.ends

.subckt nmos_1p2$$47502380_128x8m81 nmos_5p04310590548769_128x8m81_0/D nmos_5p04310590548769_128x8m81_0/S
+ a_n31_n74# VSUBS
Xnmos_5p04310590548769_128x8m81_0 nmos_5p04310590548769_128x8m81_0/D a_n31_n74# nmos_5p04310590548769_128x8m81_0/S
+ VSUBS nmos_5p04310590548769_128x8m81
.ends

.subckt pmos_5p04310590548768_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=17.69u l=0.6u
.ends

.subckt pmos_1p2$$47503404_128x8m81 a_n31_n73# pmos_5p04310590548768_128x8m81_0/S
+ w_n286_n141# pmos_5p04310590548768_128x8m81_0/D
Xpmos_5p04310590548768_128x8m81_0 w_n286_n141# pmos_5p04310590548768_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548768_128x8m81_0/S pmos_5p04310590548768_128x8m81
.ends

.subckt pmos_5p04310590548767_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=13.16u l=0.6u
.ends

.subckt pmos_1p2$$47504428_128x8m81 pmos_5p04310590548767_128x8m81_0/D a_n31_n73#
+ pmos_5p04310590548767_128x8m81_0/w_n208_n120# pmos_5p04310590548767_128x8m81_0/S
+ w_n286_n142#
Xpmos_5p04310590548767_128x8m81_0 pmos_5p04310590548767_128x8m81_0/w_n208_n120# pmos_5p04310590548767_128x8m81_0/D
+ a_n31_n73# pmos_5p04310590548767_128x8m81_0/S pmos_5p04310590548767_128x8m81
.ends

.subckt xpredec0_bot_128x8m81 alatch_128x8m81_0/a alatch_128x8m81_0/en pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ m1_n106_2472# nmos_5p04310590548770_128x8m81_0/D alatch_128x8m81_0/enb m1_n106_2674#
+ alatch_128x8m81_0/vdd m1_n106_2876# pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S
+ m1_n106_3078# VSUBS
Xalatch_128x8m81_0 alatch_128x8m81_0/enb alatch_128x8m81_0/en alatch_128x8m81_0/ab
+ alatch_128x8m81_0/a alatch_128x8m81_0/vdd VSUBS alatch_128x8m81
Xnmos_5p04310590548770_128x8m81_0 nmos_5p04310590548770_128x8m81_0/D alatch_128x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310590548770_128x8m81
Xnmos_1p2$$47502380_128x8m81_0 pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ VSUBS nmos_5p04310590548770_128x8m81_0/D VSUBS nmos_1p2$$47502380_128x8m81
Xpmos_1p2$$47503404_128x8m81_0 alatch_128x8m81_0/ab pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S
+ pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S nmos_5p04310590548770_128x8m81_0/D
+ pmos_1p2$$47503404_128x8m81
Xpmos_1p2$$47504428_128x8m81_0 pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ nmos_5p04310590548770_128x8m81_0/D pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S
+ pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/S
+ pmos_1p2$$47504428_128x8m81
.ends

.subckt pmos_5p04310590548771_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=15.2u l=0.6u
.ends

.subckt pmos_1p2$$47642668_128x8m81 w_n546_n142# pmos_5p04310590548771_128x8m81_0/S
+ pmos_5p04310590548771_128x8m81_0/D a_n31_n74#
Xpmos_5p04310590548771_128x8m81_0 w_n546_n142# pmos_5p04310590548771_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548771_128x8m81_0/S pmos_5p04310590548771_128x8m81
.ends

.subckt pmos_1p2$$47643692_128x8m81 pmos_5p04310590548771_128x8m81_0/S pmos_5p04310590548771_128x8m81_0/D
+ w_n286_n142# a_n31_n74#
Xpmos_5p04310590548771_128x8m81_0 w_n286_n142# pmos_5p04310590548771_128x8m81_0/D
+ a_n31_n74# pmos_5p04310590548771_128x8m81_0/S pmos_5p04310590548771_128x8m81
.ends

.subckt nmos_1p2$$47641644_128x8m81 a_n31_n73# nmos_5p04310590548761_128x8m81_0/S
+ nmos_5p04310590548761_128x8m81_0/D VSUBS
Xnmos_5p04310590548761_128x8m81_0 nmos_5p04310590548761_128x8m81_0/D a_n31_n73# nmos_5p04310590548761_128x8m81_0/S
+ VSUBS nmos_5p04310590548761_128x8m81
.ends

.subckt xpredec0_xa_128x8m81 nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ m1_342_3273# a_875_414# m3_855_1044# a_651_414# m1_342_3474# pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/S
+ m3_153_8117# nmos_1p2$$47641644_128x8m81_3/nmos_5p04310590548761_128x8m81_0/D m1_342_3071#
+ m1_342_3676# pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ M3_M2$$47644716_128x8m81_2/VSUBS
Xpmos_1p2$$47642668_128x8m81_0 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ a_875_414# pmos_1p2$$47642668_128x8m81
Xpmos_1p2$$47643692_128x8m81_0 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ a_651_414# pmos_1p2$$47643692_128x8m81
Xnmos_1p2$$47641644_128x8m81_0 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D
+ M3_M2$$47644716_128x8m81_2/VSUBS nmos_1p2$$47641644_128x8m81
Xnmos_1p2$$47641644_128x8m81_1 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ nmos_1p2$$47641644_128x8m81_3/nmos_5p04310590548761_128x8m81_0/D pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D
+ M3_M2$$47644716_128x8m81_2/VSUBS nmos_1p2$$47641644_128x8m81
Xnmos_1p2$$47641644_128x8m81_2 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D nmos_1p2$$47641644_128x8m81_3/nmos_5p04310590548761_128x8m81_0/D
+ M3_M2$$47644716_128x8m81_2/VSUBS nmos_1p2$$47641644_128x8m81
Xnmos_1p2$$47641644_128x8m81_3 pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D nmos_1p2$$47641644_128x8m81_3/nmos_5p04310590548761_128x8m81_0/D
+ M3_M2$$47644716_128x8m81_2/VSUBS nmos_1p2$$47641644_128x8m81
Xpmos_1p2$$47513644_128x8m81_0 pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D pmos_1p2$$47513644_128x8m81
Xpmos_1p2$$47513644_128x8m81_1 pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/S pmos_1p2$$47513644_128x8m81
Xpmos_1p2$$47513644_128x8m81_2 pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/S
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D pmos_1p2$$47513644_128x8m81
Xpmos_1p2$$47513644_128x8m81_3 pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/D
+ pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/D
+ pmos_1p2$$47513644_128x8m81_3/pmos_5p04310590548772_128x8m81_0/S pmos_1p2$$47513644_128x8m81
X0 a_771_486# a_651_414# pmos_1p2$$47643692_128x8m81_0/pmos_5p04310590548771_128x8m81_0/S M3_M2$$47644716_128x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
X1 M3_M2$$47644716_128x8m81_2/VSUBS a_875_414# a_771_486# M3_M2$$47644716_128x8m81_2/VSUBS nmos_3p3 w=12.25u l=0.6u
.ends

.subckt xpredec0_128x8m81 A[0] men x[1] x[2] x[3] A[1] clk xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ x[0] vdd vss
Xnmos_1p2$$46563372_128x8m81_0 vss pmos_5p04310590548773_128x8m81_0/D nmos_5p04310590548740_128x8m81_1/S
+ vss nmos_1p2$$46563372_128x8m81
Xpmos_5p04310590548773_128x8m81_0 vdd pmos_5p04310590548773_128x8m81_0/D nmos_5p04310590548740_128x8m81_1/S
+ vdd nmos_5p04310590548740_128x8m81_1/S pmos_5p04310590548773_128x8m81
Xxpredec0_bot_128x8m81_0 A[0] nmos_5p04310590548740_128x8m81_1/S xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D pmos_5p04310590548773_128x8m81_0/D
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D vdd xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D vss xpredec0_bot_128x8m81
Xxpredec0_xa_128x8m81_0 xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd vss vss xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D x[0] vdd vss xpredec0_xa_128x8m81
Xxpredec0_bot_128x8m81_1 A[1] nmos_5p04310590548740_128x8m81_1/S xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D pmos_5p04310590548773_128x8m81_0/D
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D vdd xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D vss xpredec0_bot_128x8m81
Xxpredec0_xa_128x8m81_1 xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd vss vss xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D x[2] vdd vss xpredec0_xa_128x8m81
Xxpredec0_xa_128x8m81_2 xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd vss vss xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D x[1] vdd vss xpredec0_xa_128x8m81
Xxpredec0_xa_128x8m81_3 xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_0/nmos_5p04310590548770_128x8m81_0/D
+ vdd xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D xpredec0_bot_128x8m81_1/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ vdd vss vss xpredec0_bot_128x8m81_0/pmos_1p2$$47504428_128x8m81_0/pmos_5p04310590548767_128x8m81_0/D
+ xpredec0_bot_128x8m81_1/nmos_5p04310590548770_128x8m81_0/D x[3] vdd vss xpredec0_xa_128x8m81
Xnmos_5p04310590548740_128x8m81_1 vss clk nmos_5p04310590548740_128x8m81_1/S vss nmos_5p04310590548740_128x8m81
Xnmos_5p04310590548740_128x8m81_0 nmos_5p04310590548740_128x8m81_1/S men vss vss nmos_5p04310590548740_128x8m81
X0 vdd men a_4894_9505# vdd pmos_3p3 w=1.705u l=0.6u
X1 a_4446_9505# men vdd vdd pmos_3p3 w=1.705u l=0.6u
X2 a_4894_9505# clk nmos_5p04310590548740_128x8m81_1/S vdd pmos_3p3 w=1.705u l=0.6u
X3 nmos_5p04310590548740_128x8m81_1/S clk a_4446_9505# vdd pmos_3p3 w=1.705u l=0.6u
.ends

.subckt prexdec_top_128x8m81 clk A[2] A[6] A[4] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1]
+ xb[2] xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1] xpredec1_128x8m81_0/pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ xpredec0_128x8m81_0/xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_128x8m81_0/xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_128x8m81_1/xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_128x8m81_1/xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xc[0] xpredec1_128x8m81_0/w_7178_9364# men VSUBS xpredec1_128x8m81_0/vdd
Xxpredec1_128x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] clk xpredec1_128x8m81_0/pmos_1p2$$47109164_128x8m81_0/pmos_5p04310590548766_128x8m81_0/w_n208_n120#
+ xpredec1_128x8m81_0/w_7178_9364# VSUBS xpredec1_128x8m81_0/vdd xpredec1_128x8m81
Xxpredec0_128x8m81_1 A[5] men xc[1] xc[2] xc[3] A[6] clk xpredec0_128x8m81_1/xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_128x8m81_1/xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xc[0] xpredec1_128x8m81_0/vdd VSUBS xpredec0_128x8m81
Xxpredec0_128x8m81_0 A[3] men xb[1] xb[2] xb[3] A[4] clk xpredec0_128x8m81_0/xpredec0_xa_128x8m81_3/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xpredec0_128x8m81_0/xpredec0_xa_128x8m81_2/nmos_1p2$$47641644_128x8m81_0/nmos_5p04310590548761_128x8m81_0/S
+ xb[0] xpredec1_128x8m81_0/vdd VSUBS xpredec0_128x8m81
.ends

.subckt control_512x8_128x8m81 VSS VDD RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[5] xa[4] xa[3] xa[2] A[0] CEN xb[1] xc[3] xc[1] xc[2] xc[0]
+ xa[0] xa[1] A[9] A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWE gen_512x8_128x8m81_0/tblhl
+ gen_512x8_128x8m81_0/wen_v2_128x8m81_0/wen gen_512x8_128x8m81_0/WEN xa[6] ypredec1_128x8m81_0/ly[2]
+ ypredec1_128x8m81_0/ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd men prexdec_top_128x8m81_0/xpredec1_128x8m81_0/vdd
+ VSUBS gen_512x8_128x8m81_0/VDD
Xgen_512x8_128x8m81_0 gen_512x8_128x8m81_0/tblhl CEN CLK gen_512x8_128x8m81_0/WEN
+ GWE gen_512x8_128x8m81_0/pmos_5p04310590548792_128x8m81_0/D gen_512x8_128x8m81_0/wen_v2_128x8m81_0/wen
+ IGWEN VSUBS men gen_512x8_128x8m81_0/VDD gen_512x8_128x8m81
Xypredec1_128x8m81_0 ypredec1_128x8m81_0/ly[5] ypredec1_128x8m81_0/ly[4] ypredec1_128x8m81_0/ly[7]
+ ypredec1_128x8m81_0/ly[3] ypredec1_128x8m81_0/ly[2] ypredec1_128x8m81_0/ly[1] ypredec1_128x8m81_0/ly[0]
+ RYS[0] RYS[1] RYS[2] RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_128x8m81_0/ly[6]
+ men A[0] A[1] A[2] CLK ypredec1_128x8m81_0/ypredec1_bot_128x8m81_2/alatch_128x8m81_0/vdd
+ gen_512x8_128x8m81_0/VDD gen_512x8_128x8m81_0/VDD VSUBS gen_512x8_128x8m81_0/VDD
+ gen_512x8_128x8m81_0/VDD ypredec1_128x8m81
Xprexdec_top_128x8m81_0 CLK A[5] A[9] A[7] xb[3] xa[0] xc[1] xc[2] xc[3] xb[1] xb[2]
+ xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] prexdec_top_128x8m81_0/xpredec1_128x8m81_0/vdd
+ VSUBS VSUBS VSUBS VSUBS xc[0] prexdec_top_128x8m81_0/xpredec1_128x8m81_0/vdd men
+ VSUBS prexdec_top_128x8m81_0/xpredec1_128x8m81_0/vdd prexdec_top_128x8m81
.ends

.subckt pmoscap_W2_5_R270_128x8m81 w_n60_n407# a_81_507# m3_509_n1#
X0 a_81_507# M1_POLY2$$204395564_128x8m81_0/VSUBS a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt pmoscap_W2_5_477_R270_128x8m81 m3_489_n1# m3_1409_n1# w_n60_n407# a_81_507#
X0 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
X1 a_81_507# a_49_1969# a_81_507# w_n60_n407# pmos_3p3 w=5.495u l=3.94u
.ends

.subckt nmos_5p043105905487111_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=2.64u l=0.6u
.ends

.subckt nmos_5p043105905487101_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=6.59u l=0.6u
.ends

.subckt nmos_1p2$$204215340_128x8m81 nmos_5p043105905487101_128x8m81_0/S a_n31_n71#
+ nmos_5p043105905487101_128x8m81_0/D VSUBS
Xnmos_5p043105905487101_128x8m81_0 nmos_5p043105905487101_128x8m81_0/D a_n31_n71#
+ nmos_5p043105905487101_128x8m81_0/S VSUBS nmos_5p043105905487101_128x8m81
.ends

.subckt pmos_5p043105905487106_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=3.3u l=0.6u
.ends

.subckt pmos_1p2$$49271852_R270_128x8m81 w_n296_n137# pmos_5p043105905487106_128x8m81_0/S
+ pmos_5p043105905487106_128x8m81_0/D a_193_n71# a_n31_n71#
Xpmos_5p043105905487106_128x8m81_0 w_n296_n137# pmos_5p043105905487106_128x8m81_0/D
+ a_n31_n71# pmos_5p043105905487106_128x8m81_0/S a_193_n71# pmos_5p043105905487106_128x8m81
.ends

.subckt pmos_5p043105905487103_128x8m81 w_n208_n120# D a_0_n44# S a_448_n44# a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=10u l=0.6u
X1 D a_448_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
X2 D a_0_n44# S w_n208_n120# pmos_6p0 w=10u l=0.6u
.ends

.subckt pmos_1p2$$49270828_R270_128x8m81 w_n296_n137# pmos_5p043105905487103_128x8m81_0/D
+ a_193_n71# a_n31_n71# pmos_5p043105905487103_128x8m81_0/S a_417_n71#
Xpmos_5p043105905487103_128x8m81_0 w_n296_n137# pmos_5p043105905487103_128x8m81_0/D
+ a_n31_n71# pmos_5p043105905487103_128x8m81_0/S a_417_n71# a_193_n71# pmos_5p043105905487103_128x8m81
.ends

.subckt pmos_5p043105905487105_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=2.62u l=0.6u
.ends

.subckt pmos_5p043105905487104_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=5.5u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=5.5u l=0.6u
.ends

.subckt pmos_1p2$$49272876_R270_128x8m81 w_n296_n137# pmos_5p043105905487104_128x8m81_0/S
+ a_n31_n71# a_193_n71# pmos_5p043105905487104_128x8m81_0/D
Xpmos_5p043105905487104_128x8m81_0 w_n296_n137# pmos_5p043105905487104_128x8m81_0/D
+ a_n31_n71# pmos_5p043105905487104_128x8m81_0/S a_193_n71# pmos_5p043105905487104_128x8m81
.ends

.subckt nmos_5p043105905487109_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=3.3u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=3.3u l=0.6u
.ends

.subckt nmos_1p2$$49277996_R270_128x8m81 nmos_5p04310590548744_128x8m81_0/D a_n31_n71#
+ nmos_5p04310590548744_128x8m81_0/S VSUBS
Xnmos_5p04310590548744_128x8m81_0 nmos_5p04310590548744_128x8m81_0/D a_n31_n71# nmos_5p04310590548744_128x8m81_0/S
+ VSUBS nmos_5p04310590548744_128x8m81
.ends

.subckt nmos_5p043105905487108_128x8m81 D a_0_n44# S a_224_n44# VSUBS
X0 S a_224_n44# D VSUBS nmos_6p0 w=5u l=0.6u
X1 D a_0_n44# S VSUBS nmos_6p0 w=5u l=0.6u
.ends

.subckt nmos_5p043105905487107_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=0.66u l=0.6u
.ends

.subckt pmos_5p043105905487110_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=1.59u l=0.6u
.ends

.subckt xdec_128x8m81 LWL xc xb xa m2_16621_n223# m2_17754_n223# m2_11825_n223# m2_12202_n223#
+ m2_12958_n223# m2_15487_n223# m2_12580_n223# m2_15110_n223# m2_11069_n223# m2_15865_n223#
+ m2_16243_n223# m2_10314_n223# m2_16998_n223# m2_17376_n223# vdd m2_11447_n223# RWL
+ vss m2_10691_n223# men
Xpmos_1p2$$49271852_R270_128x8m81_0 vdd nmos_5p043105905487109_128x8m81_0/S men pmos_5p043105905487105_128x8m81_2/S
+ pmos_5p043105905487105_128x8m81_2/S pmos_1p2$$49271852_R270_128x8m81
Xpmos_1p2$$49270828_R270_128x8m81_0 vdd vdd pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D
+ pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D LWL pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D
+ pmos_1p2$$49270828_R270_128x8m81
Xpmos_5p043105905487105_128x8m81_0 vdd pmos_5p043105905487105_128x8m81_2/S xb vdd
+ pmos_5p043105905487105_128x8m81
Xpmos_5p043105905487105_128x8m81_1 vdd vdd xc pmos_5p043105905487105_128x8m81_2/S
+ pmos_5p043105905487105_128x8m81
Xpmos_5p043105905487105_128x8m81_2 vdd vdd xa pmos_5p043105905487105_128x8m81_2/S
+ pmos_5p043105905487105_128x8m81
Xpmos_1p2$$49272876_R270_128x8m81_0 vdd vdd nmos_5p043105905487109_128x8m81_0/S nmos_5p043105905487109_128x8m81_0/S
+ pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D pmos_1p2$$49272876_R270_128x8m81
Xnmos_5p043105905487109_128x8m81_0 men pmos_5p043105905487110_128x8m81_0/S nmos_5p043105905487109_128x8m81_0/S
+ pmos_5p043105905487110_128x8m81_0/S vss nmos_5p043105905487109_128x8m81
Xnmos_1p2$$49277996_R270_128x8m81_0 vss pmos_5p043105905487105_128x8m81_2/S nmos_5p043105905487109_128x8m81_0/S
+ vss nmos_1p2$$49277996_R270_128x8m81
Xpmos_1p2$$49272876_R270_128x8m81_1 vdd vdd nmos_5p043105905487109_128x8m81_0/S nmos_5p043105905487109_128x8m81_0/S
+ pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D pmos_1p2$$49272876_R270_128x8m81
Xpmos_5p043105905487103_128x8m81_0 vdd vdd pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D
+ RWL pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D
+ pmos_5p043105905487103_128x8m81
Xnmos_5p043105905487108_128x8m81_0 LWL pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D
+ vss pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D vss nmos_5p043105905487108_128x8m81
Xnmos_5p043105905487108_128x8m81_1 RWL pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D
+ vss pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D vss nmos_5p043105905487108_128x8m81
Xnmos_5p043105905487107_128x8m81_0 vss pmos_5p043105905487105_128x8m81_2/S pmos_5p043105905487110_128x8m81_0/S
+ vss nmos_5p043105905487107_128x8m81
Xpmos_5p043105905487110_128x8m81_0 vdd vdd pmos_5p043105905487105_128x8m81_2/S pmos_5p043105905487110_128x8m81_0/S
+ pmos_5p043105905487110_128x8m81
X0 a_13291_624# xb a_13291_400# vss nmos_3p3 w=3.15u l=0.6u
X1 vss xc a_13291_624# vss nmos_3p3 w=3.15u l=0.6u
X2 a_13291_400# xa pmos_5p043105905487105_128x8m81_2/S vss nmos_3p3 w=3.15u l=0.6u
X3 vss nmos_5p043105905487109_128x8m81_0/S pmos_1p2$$49272876_R270_128x8m81_0/pmos_5p043105905487104_128x8m81_0/D vss nmos_3p3 w=5u l=0.6u
X4 vss nmos_5p043105905487109_128x8m81_0/S pmos_1p2$$49272876_R270_128x8m81_1/pmos_5p043105905487104_128x8m81_0/D vss nmos_3p3 w=5u l=0.6u
.ends

.subckt xdec8_128x8m81 RWL[0] LWL[5] LWL[2] RWL[5] RWL[4] RWL[2] RWL[1] RWL[7] LWL[6]
+ LWL[0] LWL[3] xa[5] xa[2] xa[1] xa[7] xa[4] xdec_128x8m81_7/m2_17376_n223# RWL[3]
+ xdec_128x8m81_7/m2_11447_n223# LWL[1] xdec_128x8m81_7/m2_17754_n223# xdec_128x8m81_7/m2_11825_n223#
+ xdec_128x8m81_3/RWL xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_15865_n223#
+ LWL[7] xc xdec_128x8m81_7/m2_10691_n223# xdec_128x8m81_7/m2_16243_n223# xa[3] xdec_128x8m81_7/m2_12580_n223#
+ xb RWL[6] xa[0] xdec_128x8m81_7/m2_10314_n223# xa[6] xdec_128x8m81_7/m2_16621_n223#
+ LWL[4] xdec_128x8m81_7/m2_12958_n223# men xdec_128x8m81_7/m2_15110_n223# xdec_128x8m81_7/m2_16998_n223#
+ vdd xdec_128x8m81_7/m2_15487_n223# vss xdec_128x8m81_7/m2_11069_n223#
Xxdec_128x8m81_0 LWL[6] xc xb xa[6] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[6] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_1 LWL[4] xc xb xa[4] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[4] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_2 LWL[2] xc xb xa[2] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[2] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_3 LWL[0] xc xb xa[0] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# xdec_128x8m81_3/RWL vss xdec_128x8m81_7/m2_10691_n223#
+ men xdec_128x8m81
Xxdec_128x8m81_4 LWL[7] xc xb xa[7] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[7] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_5 LWL[5] xc xb xa[5] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[5] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_6 LWL[3] xc xb xa[3] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[3] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
Xxdec_128x8m81_7 LWL[1] xc xb xa[1] xdec_128x8m81_7/m2_16621_n223# xdec_128x8m81_7/m2_17754_n223#
+ xdec_128x8m81_7/m2_11825_n223# xdec_128x8m81_7/m2_12202_n223# xdec_128x8m81_7/m2_12958_n223#
+ xdec_128x8m81_7/m2_15487_n223# xdec_128x8m81_7/m2_12580_n223# xdec_128x8m81_7/m2_15110_n223#
+ xdec_128x8m81_7/m2_11069_n223# xdec_128x8m81_7/m2_15865_n223# xdec_128x8m81_7/m2_16243_n223#
+ xdec_128x8m81_7/m2_10314_n223# xdec_128x8m81_7/m2_16998_n223# xdec_128x8m81_7/m2_17376_n223#
+ vdd xdec_128x8m81_7/m2_11447_n223# RWL[1] vss xdec_128x8m81_7/m2_10691_n223# men
+ xdec_128x8m81
.ends

.subckt xdec16_128x8_128x8m81 LWL[7] RWL[15] RWL[14] RWL[12] LWL[9] LWL[2] LWL[3]
+ LWL[4] LWL[5] RWL[11] RWL[9] RWL[8] RWL[7] RWL[5] RWL[1] RWL[0] LWL[15] LWL[12]
+ RWL[4] RWL[6] xa[2] xa[0] xa[3] xa[4] xa[5] xa[6] xa[7] xb[3] xb[2] xb[1] xb[0]
+ xc xdec8_128x8m81_1/xdec_128x8m81_7/m2_10314_n223# xdec8_128x8m81_0/xdec_128x8m81_3/RWL
+ xdec8_128x8m81_1/xdec_128x8m81_7/m2_10691_n223# LWL[10] xdec8_128x8m81_1/xdec_128x8m81_7/m2_11069_n223#
+ RWL[2] LWL[0] men RWL[13] LWL[6] LWL[11] RWL[10] LWL[8] xa[1] RWL[3] LWL[13] LWL[1]
+ LWL[14] xdec8_128x8m81_1/xdec_128x8m81_3/RWL VSUBS xdec8_128x8m81_1/vdd
Xxdec8_128x8m81_0 RWL[8] LWL[13] LWL[10] RWL[13] RWL[12] RWL[10] RWL[9] RWL[15] LWL[14]
+ LWL[8] LWL[11] xa[5] xa[2] xa[1] xa[7] xa[4] xa[1] RWL[11] xc LWL[9] xa[0] xb[3]
+ xdec8_128x8m81_0/xdec_128x8m81_3/RWL xb[2] xa[5] LWL[15] xc xdec8_128x8m81_1/xdec_128x8m81_7/m2_10691_n223#
+ xa[4] xa[3] xb[1] xb[1] RWL[14] xa[0] xdec8_128x8m81_1/xdec_128x8m81_7/m2_10314_n223#
+ xa[6] xa[3] LWL[12] xb[0] men xa[7] xa[2] xdec8_128x8m81_1/vdd xa[6] VSUBS xdec8_128x8m81_1/xdec_128x8m81_7/m2_11069_n223#
+ xdec8_128x8m81
Xxdec8_128x8m81_1 xdec8_128x8m81_1/RWL[0] LWL[5] LWL[2] RWL[5] RWL[4] RWL[2] RWL[1]
+ RWL[7] LWL[6] LWL[0] LWL[3] xa[5] xa[2] xa[1] xa[7] xa[4] xa[1] RWL[3] xc LWL[1]
+ xa[0] xb[3] xdec8_128x8m81_1/xdec_128x8m81_3/RWL xb[2] xa[5] LWL[7] xc xdec8_128x8m81_1/xdec_128x8m81_7/m2_10691_n223#
+ xa[4] xa[3] xb[1] xb[0] RWL[6] xa[0] xdec8_128x8m81_1/xdec_128x8m81_7/m2_10314_n223#
+ xa[6] xa[3] LWL[4] xb[0] men xa[7] xa[2] xdec8_128x8m81_1/vdd xa[6] VSUBS xdec8_128x8m81_1/xdec_128x8m81_7/m2_11069_n223#
+ xdec8_128x8m81
.ends

.subckt nmos_5p04310590548799_128x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nmos_6p0 w=10.11u l=0.6u
.ends

.subckt nmos_1p2$$204213292_R90_128x8m81 nmos_5p04310590548799_128x8m81_0/D a_n31_n71#
+ nmos_5p04310590548799_128x8m81_0/S VSUBS
Xnmos_5p04310590548799_128x8m81_0 nmos_5p04310590548799_128x8m81_0/D a_n31_n71# nmos_5p04310590548799_128x8m81_0/S
+ VSUBS nmos_5p04310590548799_128x8m81
.ends

.subckt pmos_5p043105905487100_128x8m81 w_n208_n120# D a_0_n44# S
X0 D a_0_n44# S w_n208_n120# pmos_6p0 w=6.59u l=0.6u
.ends

.subckt pmos_5p043105905487102_128x8m81 w_n208_n120# D a_0_n44# S a_224_n44#
X0 S a_224_n44# D w_n208_n120# pmos_6p0 w=12.63u l=0.6u
X1 D a_0_n44# S w_n208_n120# pmos_6p0 w=12.63u l=0.6u
.ends

.subckt pmos_1p2$$204216364_128x8m81 pmos_5p043105905487102_128x8m81_0/D a_193_n71#
+ a_n31_n71# w_n296_n137# pmos_5p043105905487102_128x8m81_0/S
Xpmos_5p043105905487102_128x8m81_0 w_n296_n137# pmos_5p043105905487102_128x8m81_0/D
+ a_n31_n71# pmos_5p043105905487102_128x8m81_0/S a_193_n71# pmos_5p043105905487102_128x8m81
.ends

.subckt pmos_1p2$$204217388_R90_128x8m81 w_n295_n137# pmos_5p043105905487100_128x8m81_0/S
+ a_n31_n71# pmos_5p043105905487100_128x8m81_0/D
Xpmos_5p043105905487100_128x8m81_0 w_n295_n137# pmos_5p043105905487100_128x8m81_0/D
+ a_n31_n71# pmos_5p043105905487100_128x8m81_0/S pmos_5p043105905487100_128x8m81
.ends

.subckt xdec16_128_128x8m81 DRWL RWL[3] RWL[5] RWL[7] RWL[8] RWL[9] RWL[10] RWL[11]
+ RWL[13] RWL[15] LWL[13] LWL[15] LWL[5] LWL[8] LWL[9] LWL[6] LWL[7] DLWL xb[0] xb[1]
+ xb[2] xb[3] xa[7] xa[6] xa[5] xa[4] xa[0] xa[3] xa[2] xc[1] LWL[11] RWL[1] RWL[6]
+ RWL[4] LWL[14] RWL[2] LWL[12] RWL[0] LWL[10] men LWL[4] LWL[2] LWL[0] LWL[3] RWL[14]
+ RWL[12] LWL[1] vdd xa[1] xc[0] vss
Xpmoscap_W2_5_R270_128x8m81_0 vdd vdd DLWL pmoscap_W2_5_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_10 RWL[11] RWL[10] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_R270_128x8m81_1 vdd vdd DRWL pmoscap_W2_5_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_0 LWL[15] LWL[14] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_11 RWL[9] RWL[8] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_1 LWL[13] LWL[12] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_12 RWL[7] RWL[6] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_2 LWL[11] LWL[10] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_14 RWL[3] RWL[2] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_13 RWL[5] RWL[4] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_3 LWL[9] LWL[8] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_15 RWL[1] RWL[0] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xnmos_5p043105905487111_128x8m81_0 vss pmos_5p043105905487100_128x8m81_0/D pmos_5p043105905487100_128x8m81_1/S
+ vss nmos_5p043105905487111_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_4 LWL[7] LWL[6] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_5 LWL[5] LWL[4] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xnmos_1p2$$204215340_128x8m81_0 pmos_5p043105905487100_128x8m81_0/D vdd men vss nmos_1p2$$204215340_128x8m81
Xnmos_5p043105905487111_128x8m81_1 vss pmos_5p043105905487100_128x8m81_0/D nmos_5p043105905487111_128x8m81_1/S
+ vss nmos_5p043105905487111_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_6 LWL[3] LWL[2] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_7 LWL[1] LWL[0] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xxdec16_128x8_128x8m81_0 LWL[7] RWL[15] RWL[14] RWL[12] LWL[9] LWL[2] LWL[3] LWL[4]
+ LWL[5] RWL[11] RWL[9] RWL[8] RWL[7] RWL[5] RWL[1] RWL[0] LWL[15] LWL[12] RWL[4]
+ RWL[6] xa[2] xa[0] xa[3] xa[4] xa[5] xa[6] xa[7] xb[3] xb[2] xb[1] xb[0] xc[0] vdd
+ RWL[8] vdd LWL[10] xc[1] RWL[2] LWL[0] men RWL[13] LWL[6] LWL[11] RWL[10] LWL[8]
+ xa[1] RWL[3] LWL[13] LWL[1] LWL[14] RWL[0] vss vdd xdec16_128x8_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_8 RWL[15] RWL[14] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xnmos_1p2$$204213292_R90_128x8m81_0 vss nmos_5p043105905487111_128x8m81_1/S DLWL vss
+ nmos_1p2$$204213292_R90_128x8m81
Xpmoscap_W2_5_477_R270_128x8m81_9 RWL[13] RWL[12] vdd vdd pmoscap_W2_5_477_R270_128x8m81
Xnmos_5p04310590548799_128x8m81_0 vss pmos_5p043105905487100_128x8m81_1/S DRWL vss
+ nmos_5p04310590548799_128x8m81
Xpmos_5p043105905487100_128x8m81_0 vdd pmos_5p043105905487100_128x8m81_0/D vss men
+ pmos_5p043105905487100_128x8m81
Xpmos_1p2$$204216364_128x8m81_0 DRWL pmos_5p043105905487100_128x8m81_1/S pmos_5p043105905487100_128x8m81_1/S
+ vdd vdd pmos_1p2$$204216364_128x8m81
Xpmos_5p043105905487100_128x8m81_1 vdd vdd pmos_5p043105905487100_128x8m81_0/D pmos_5p043105905487100_128x8m81_1/S
+ pmos_5p043105905487100_128x8m81
Xpmos_1p2$$204216364_128x8m81_1 DLWL nmos_5p043105905487111_128x8m81_1/S nmos_5p043105905487111_128x8m81_1/S
+ vdd vdd pmos_1p2$$204216364_128x8m81
Xpmos_1p2$$204217388_R90_128x8m81_0 vdd nmos_5p043105905487111_128x8m81_1/S pmos_5p043105905487100_128x8m81_0/D
+ vdd pmos_1p2$$204217388_R90_128x8m81
.ends

.subckt gf180mcu_fd_ip_sram__sram128x8m8wm1 VSS CLK D[0] A[2] A[1] A[0] Q[2] Q[3]
+ CEN A[5] A[6] A[4] WEN[3] D[7] Q[7] D[3] D[1] D[2] A[3] Q[1] Q[6] D[5] Q[4] WEN[5]
+ WEN[2] WEN[1] WEN[4] WEN[7] WEN[6] D[4] D[6] Q[5] Q[0] GWEN WEN[0]
Xlcol4_128_128x8m81_0 lcol4_128_128x8m81_0/WL[15] lcol4_128_128x8m81_0/WL[14] lcol4_128_128x8m81_0/WL[13]
+ lcol4_128_128x8m81_0/WL[12] lcol4_128_128x8m81_0/WL[11] lcol4_128_128x8m81_0/WL[10]
+ lcol4_128_128x8m81_0/WL[9] lcol4_128_128x8m81_0/WL[8] lcol4_128_128x8m81_0/WL[7]
+ lcol4_128_128x8m81_0/WL[6] lcol4_128_128x8m81_0/WL[5] lcol4_128_128x8m81_0/WL[4]
+ lcol4_128_128x8m81_0/WL[3] lcol4_128_128x8m81_0/WL[2] lcol4_128_128x8m81_0/WL[1]
+ lcol4_128_128x8m81_0/WL[0] lcol4_128_128x8m81_0/men lcol4_128_128x8m81_0/ypass[0]
+ lcol4_128_128x8m81_0/ypass[1] lcol4_128_128x8m81_0/ypass[2] lcol4_128_128x8m81_0/ypass[3]
+ lcol4_128_128x8m81_0/ypass[4] lcol4_128_128x8m81_0/ypass[5] lcol4_128_128x8m81_0/ypass[6]
+ lcol4_128_128x8m81_0/ypass[7] lcol4_128_128x8m81_0/GWEN lcol4_128_128x8m81_0/GWE
+ D[0] D[1] D[3] D[2] Q[0] Q[1] Q[2] Q[3] lcol4_128_128x8m81_0/pcb[2] lcol4_128_128x8m81_0/pcb[3]
+ lcol4_128_128x8m81_0/pcb[0] lcol4_128_128x8m81_0/pcb[1] VSS WEN[1] WEN[2] WEN[3]
+ xdec16_128_128x8m81_0/LWL[0] xdec16_128_128x8m81_0/LWL[1] VSS xdec16_128_128x8m81_0/LWL[2]
+ xdec16_128_128x8m81_0/LWL[3] xdec16_128_128x8m81_0/LWL[4] xdec16_128_128x8m81_0/LWL[10]
+ xdec16_128_128x8m81_0/LWL[5] VSS xdec16_128_128x8m81_0/LWL[11] xdec16_128_128x8m81_0/LWL[6]
+ xdec16_128_128x8m81_0/LWL[12] xdec16_128_128x8m81_0/LWL[7] xdec16_128_128x8m81_0/LWL[13]
+ VSS xdec16_128_128x8m81_0/LWL[8] xdec16_128_128x8m81_0/LWL[14] rcol4_128_128x8m81_0/men
+ VSS xdec16_128_128x8m81_0/LWL[9] xdec16_128_128x8m81_0/LWL[15] WEN[0] VSS rcol4_128_128x8m81_0/GWEN
+ VSS WEN[3] VSS VSS lcol4_128_128x8m81_0/saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_1/sa_128x8m81_0/pcb
+ VSS WEN[0] control_512x8_128x8m81_0/LYS[0] lcol4_128_128x8m81_0/saout_wm1_x4_128x8m81_0/saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb
+ VSS control_512x8_128x8m81_0/LYS[1] lcol4_128_128x8m81_0/saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_1/sa_128x8m81_0/pcb
+ control_512x8_128x8m81_0/LYS[2] control_512x8_128x8m81_0/LYS[3] control_512x8_128x8m81_0/LYS[4]
+ rcol4_128_128x8m81_0/GWE control_512x8_128x8m81_0/LYS[5] control_512x8_128x8m81_0/LYS[6]
+ lcol4_128_128x8m81_0/saout_wm1_x4_128x8m81_0/saout_m2_128x8m81_0/pcb control_512x8_128x8m81_0/LYS[7]
+ VSS VSS lcol4_128_128x8m81
Xrcol4_128_128x8m81_0 rcol4_128_128x8m81_0/WL[6] rcol4_128_128x8m81_0/WL[5] rcol4_128_128x8m81_0/ypass[1]
+ rcol4_128_128x8m81_0/ypass[2] rcol4_128_128x8m81_0/ypass[3] rcol4_128_128x8m81_0/ypass[4]
+ rcol4_128_128x8m81_0/ypass[5] rcol4_128_128x8m81_0/ypass[6] rcol4_128_128x8m81_0/DWL
+ rcol4_128_128x8m81_0/tblhl rcol4_128_128x8m81_0/GWEN rcol4_128_128x8m81_0/ypass[0]
+ rcol4_128_128x8m81_0/WL[11] rcol4_128_128x8m81_0/WL[15] rcol4_128_128x8m81_0/WL[0]
+ rcol4_128_128x8m81_0/WL[2] rcol4_128_128x8m81_0/WL[12] rcol4_128_128x8m81_0/WL[3]
+ rcol4_128_128x8m81_0/WL[4] rcol4_128_128x8m81_0/WL[7] rcol4_128_128x8m81_0/WL[8]
+ rcol4_128_128x8m81_0/WL[9] rcol4_128_128x8m81_0/WL[1] rcol4_128_128x8m81_0/ypass[7]
+ rcol4_128_128x8m81_0/WL[10] rcol4_128_128x8m81_0/WL[13] rcol4_128_128x8m81_0/WL[14]
+ D[4] D[7] Q[5] Q[6] Q[7] D[5] D[6] Q[4] rcol4_128_128x8m81_0/pcb[6] rcol4_128_128x8m81_0/pcb[7]
+ rcol4_128_128x8m81_0/pcb[4] rcol4_128_128x8m81_0/vdd WEN[7] WEN[4] rcol4_128_128x8m81_0/pcb[5]
+ WEN[6] WEN[5] VSS rcol4_128_128x8m81_0/WL[0] VSS rcol4_128_128x8m81_0/WL[1] rcol4_128_128x8m81_0/WL[3]
+ rcol4_128_128x8m81_0/WL[4] rcol4_128_128x8m81_0/WL[7] rcol4_128_128x8m81_0/WL[8]
+ VSS VSS VSS VSS VSS VSS rcol4_128_128x8m81_0/WL[10] rcol4_128_128x8m81_0/saout_R_m2_128x8m81_1/pcb
+ rcol4_128_128x8m81_0/WL[11] rcol4_128_128x8m81_0/WL[14] rcol4_128_128x8m81_0/GWE
+ rcol4_128_128x8m81_0/WL[15] WEN[7] VSS VSS VSS rcol4_128_128x8m81_0/DWL rcol4_128_128x8m81_0/saout_m2_128x8m81_0/pcb
+ rcol4_128_128x8m81_0/saout_m2_128x8m81_1/sa_128x8m81_0/pcb VSS rcol4_128_128x8m81_0/men
+ rcol4_128_128x8m81_0/saout_R_m2_128x8m81_1/pcb rcol4_128_128x8m81_0/saout_R_m2_128x8m81_0/sa_128x8m81_0/pcb
+ VSS VSS rcol4_128_128x8m81
Xcontrol_512x8_128x8m81_0 VSS VSS rcol4_128_128x8m81_0/ypass[7] rcol4_128_128x8m81_0/ypass[6]
+ rcol4_128_128x8m81_0/ypass[5] rcol4_128_128x8m81_0/ypass[4] rcol4_128_128x8m81_0/ypass[3]
+ rcol4_128_128x8m81_0/ypass[2] rcol4_128_128x8m81_0/ypass[1] rcol4_128_128x8m81_0/ypass[0]
+ control_512x8_128x8m81_0/LYS[0] control_512x8_128x8m81_0/LYS[1] control_512x8_128x8m81_0/LYS[2]
+ control_512x8_128x8m81_0/LYS[3] control_512x8_128x8m81_0/LYS[6] control_512x8_128x8m81_0/LYS[5]
+ control_512x8_128x8m81_0/LYS[4] control_512x8_128x8m81_0/LYS[7] rcol4_128_128x8m81_0/tblhl
+ rcol4_128_128x8m81_0/GWEN xdec16_128_128x8m81_0/xb[3] xdec16_128_128x8m81_0/xb[2]
+ xdec16_128_128x8m81_0/xb[0] xdec16_128_128x8m81_0/xa[7] xdec16_128_128x8m81_0/xa[5]
+ xdec16_128_128x8m81_0/xa[4] xdec16_128_128x8m81_0/xa[3] xdec16_128_128x8m81_0/xa[2]
+ A[0] CEN xdec16_128_128x8m81_0/xb[1] control_512x8_128x8m81_0/xc[3] xdec16_128_128x8m81_0/xc[1]
+ control_512x8_128x8m81_0/xc[2] control_512x8_128x8m81_0/xc[0] xdec16_128_128x8m81_0/xa[0]
+ xdec16_128_128x8m81_0/xa[1] VSS VSS CLK A[2] A[1] A[6] A[3] A[4] A[5] VSS rcol4_128_128x8m81_0/GWE
+ rcol4_128_128x8m81_0/tblhl GWEN GWEN xdec16_128_128x8m81_0/xa[6] control_512x8_128x8m81_0/LYS[2]
+ VSS rcol4_128_128x8m81_0/men VSS VSS VSS control_512x8_128x8m81
Xxdec16_128_128x8m81_0 rcol4_128_128x8m81_0/DWL rcol4_128_128x8m81_0/WL[3] rcol4_128_128x8m81_0/WL[5]
+ rcol4_128_128x8m81_0/WL[7] rcol4_128_128x8m81_0/WL[8] rcol4_128_128x8m81_0/WL[9]
+ rcol4_128_128x8m81_0/WL[10] rcol4_128_128x8m81_0/WL[11] rcol4_128_128x8m81_0/WL[13]
+ rcol4_128_128x8m81_0/WL[15] xdec16_128_128x8m81_0/LWL[13] xdec16_128_128x8m81_0/LWL[15]
+ xdec16_128_128x8m81_0/LWL[5] xdec16_128_128x8m81_0/LWL[8] xdec16_128_128x8m81_0/LWL[9]
+ xdec16_128_128x8m81_0/LWL[6] xdec16_128_128x8m81_0/LWL[7] xdec16_128_128x8m81_0/DLWL
+ xdec16_128_128x8m81_0/xb[0] xdec16_128_128x8m81_0/xb[1] xdec16_128_128x8m81_0/xb[2]
+ xdec16_128_128x8m81_0/xb[3] xdec16_128_128x8m81_0/xa[7] xdec16_128_128x8m81_0/xa[6]
+ xdec16_128_128x8m81_0/xa[5] xdec16_128_128x8m81_0/xa[4] xdec16_128_128x8m81_0/xa[0]
+ xdec16_128_128x8m81_0/xa[3] xdec16_128_128x8m81_0/xa[2] xdec16_128_128x8m81_0/xc[1]
+ xdec16_128_128x8m81_0/LWL[11] rcol4_128_128x8m81_0/WL[1] rcol4_128_128x8m81_0/WL[6]
+ rcol4_128_128x8m81_0/WL[4] xdec16_128_128x8m81_0/LWL[14] rcol4_128_128x8m81_0/WL[2]
+ xdec16_128_128x8m81_0/LWL[12] rcol4_128_128x8m81_0/WL[0] xdec16_128_128x8m81_0/LWL[10]
+ rcol4_128_128x8m81_0/men xdec16_128_128x8m81_0/LWL[4] xdec16_128_128x8m81_0/LWL[2]
+ xdec16_128_128x8m81_0/LWL[0] xdec16_128_128x8m81_0/LWL[3] rcol4_128_128x8m81_0/WL[14]
+ rcol4_128_128x8m81_0/WL[12] xdec16_128_128x8m81_0/LWL[1] VSS xdec16_128_128x8m81_0/xa[1]
+ VSS VSS xdec16_128_128x8m81
.ends

