magic
tech gf180mcuB
timestamp 1669390400
<< properties >>
string GDS_END 1409468
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1403704
<< end >>
