magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect 272 69800 2172 70000
rect 2752 69800 4802 70000
rect 5122 69800 7172 70000
rect 7828 69800 9878 70000
rect 10198 69800 12248 70000
rect 12828 69800 14728 70000
<< metal3 >>
rect 0 68400 200 69678
rect 14800 68400 15000 69678
rect 0 66800 200 68200
rect 14800 66800 15000 68200
rect 0 65200 200 66600
rect 14800 65200 15000 66600
rect 0 63600 200 65000
rect 14800 63600 15000 65000
rect 0 62000 200 63400
rect 14800 62000 15000 63400
rect 0 60400 200 61800
rect 14800 60400 15000 61800
rect 0 58800 200 60200
rect 14800 58800 15000 60200
rect 0 57200 200 58600
rect 14800 57200 15000 58600
rect 0 55600 200 57000
rect 14800 55600 15000 57000
rect 0 54000 200 55400
rect 14800 54000 15000 55400
rect 0 52400 200 53800
rect 14800 52400 15000 53800
rect 0 50800 200 52200
rect 14800 50800 15000 52200
rect 0 49200 200 50600
rect 14800 49200 15000 50600
rect 0 46000 200 49000
rect 14800 46000 15000 49000
rect 0 42800 200 45800
rect 14800 42800 15000 45800
rect 0 41200 200 42600
rect 14800 41200 15000 42600
rect 0 39600 200 41000
rect 14800 39600 15000 41000
rect 0 36400 200 39400
rect 14800 36400 15000 39400
rect 0 33200 200 36200
rect 14800 33200 15000 36200
rect 0 30000 200 33000
rect 14800 30000 15000 33000
rect 0 26800 200 29800
rect 14800 26800 15000 29800
rect 0 25200 200 26600
rect 14800 25200 15000 26600
rect 0 23600 200 25000
rect 14800 23600 15000 25000
rect 0 20400 200 23400
rect 14800 20400 15000 23400
rect 0 17200 200 20200
rect 14800 17200 15000 20200
rect 0 14000 200 17000
rect 14800 14000 15000 17000
<< metal4 >>
rect 0 68400 200 69678
rect 14800 68400 15000 69678
rect 0 66800 200 68200
rect 14800 66800 15000 68200
rect 0 65200 200 66600
rect 14800 65200 15000 66600
rect 0 63600 200 65000
rect 14800 63600 15000 65000
rect 0 62000 200 63400
rect 14800 62000 15000 63400
rect 0 60400 200 61800
rect 14800 60400 15000 61800
rect 0 58800 200 60200
rect 14800 58800 15000 60200
rect 0 57200 200 58600
rect 14800 57200 15000 58600
rect 0 55600 200 57000
rect 14800 55600 15000 57000
rect 0 54000 200 55400
rect 14800 54000 15000 55400
rect 0 52400 200 53800
rect 14800 52400 15000 53800
rect 0 50800 200 52200
rect 14800 50800 15000 52200
rect 0 49200 200 50600
rect 14800 49200 15000 50600
rect 0 46000 200 49000
rect 14800 46000 15000 49000
rect 0 42800 200 45800
rect 14800 42800 15000 45800
rect 0 41200 200 42600
rect 14800 41200 15000 42600
rect 0 39600 200 41000
rect 14800 39600 15000 41000
rect 0 36400 200 39400
rect 14800 36400 15000 39400
rect 0 33200 200 36200
rect 14800 33200 15000 36200
rect 0 30000 200 33000
rect 14800 30000 15000 33000
rect 0 26800 200 29800
rect 14800 26800 15000 29800
rect 0 25200 200 26600
rect 14800 25200 15000 26600
rect 0 23600 200 25000
rect 14800 23600 15000 25000
rect 0 20400 200 23400
rect 14800 20400 15000 23400
rect 0 17200 200 20200
rect 14800 17200 15000 20200
rect 0 14000 200 17000
rect 14800 14000 15000 17000
<< metal5 >>
rect 0 68400 200 69678
rect 14800 68400 15000 69678
rect 0 66800 200 68200
rect 14800 66800 15000 68200
rect 0 65200 200 66600
rect 14800 65200 15000 66600
rect 0 63600 200 65000
rect 14800 63600 15000 65000
rect 0 62000 200 63400
rect 14800 62000 15000 63400
rect 0 60400 200 61800
rect 14800 60400 15000 61800
rect 0 58800 200 60200
rect 14800 58800 15000 60200
rect 0 57200 200 58600
rect 14800 57200 15000 58600
rect 0 55600 200 57000
rect 14800 55600 15000 57000
rect 0 54000 200 55400
rect 14800 54000 15000 55400
rect 0 52400 200 53800
rect 14800 52400 15000 53800
rect 0 50800 200 52200
rect 14800 50800 15000 52200
rect 0 49200 200 50600
rect 14800 49200 15000 50600
rect 0 46000 200 49000
rect 14800 46000 15000 49000
rect 0 42800 200 45800
rect 14800 42800 15000 45800
rect 0 41200 200 42600
rect 14800 41200 15000 42600
rect 0 39600 200 41000
rect 14800 39600 15000 41000
rect 0 36400 200 39400
rect 14800 36400 15000 39400
rect 0 33200 200 36200
rect 14800 33200 15000 36200
rect 0 30000 200 33000
rect 14800 30000 15000 33000
rect 0 26800 200 29800
rect 14800 26800 15000 29800
rect 0 25200 200 26600
rect 14800 25200 15000 26600
rect 0 23600 200 25000
rect 14800 23600 15000 25000
rect 0 20400 200 23400
rect 14800 20400 15000 23400
rect 0 17200 200 20200
rect 14800 17200 15000 20200
rect 0 14000 200 17000
rect 14800 14000 15000 17000
use 5LM_METAL_RAIL_PAD_60  5LM_METAL_RAIL_PAD_60_0
timestamp 1669390400
transform 1 0 0 0 1 0
box -32 0 15032 69968
use GF_NI_DVSS_BASE  GF_NI_DVSS_BASE_0
timestamp 1669390400
transform 1 0 11 0 1 12400
box -11 0 14989 57600
<< labels >>
rlabel metal5 s 14800 20400 15000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 17200 15000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 14000 15000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 25200 15000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 39600 15000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 46000 15000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 49200 15000 50600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 57200 15000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 60400 15000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 63600 15000 65000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 65200 15000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 68400 15000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14800 23600 15000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 36400 15000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 33200 15000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 30000 15000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 26800 15000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 42800 15000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 41200 15000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 55600 15000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 54000 15000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 52400 15000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 58800 15000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 66800 15000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 14800 50800 15000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal5 s 14800 62000 15000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 14800 20400 15000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 17200 15000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 14000 15000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 25200 15000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 39600 15000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 46000 15000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 49200 15000 50600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 57200 15000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 60400 15000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 63600 15000 65000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 65200 15000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 68400 15000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14800 23600 15000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 36400 15000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 33200 15000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 30000 15000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 26800 15000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 42800 15000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 41200 15000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 55600 15000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 54000 15000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 52400 15000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 58800 15000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 66800 15000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14800 50800 15000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 14800 62000 15000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 14800 20400 15000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 17200 15000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 14000 15000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 25200 15000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 39600 15000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 46000 15000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 49200 15000 50600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 57200 15000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 60400 15000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 63600 15000 65000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 65200 15000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 68400 15000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14800 23600 15000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 36400 15000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 33200 15000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 30000 15000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 26800 15000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 42800 15000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 41200 15000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 55600 15000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 54000 15000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 52400 15000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 58800 15000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 66800 15000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 14800 50800 15000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 14800 62000 15000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal2 s 272 69800 2172 70000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 2752 69800 4802 70000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 5122 69800 7172 70000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 7828 69800 9878 70000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 10198 69800 12248 70000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 68400 200 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 200 69678 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 65200 200 66600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 63600 200 65000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 49200 200 50600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 68400 200 69678 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 65200 200 66600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 63600 200 65000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 49200 200 50600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal2 s 12828 69800 14728 70000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string GDS_END 4985370
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4981582
string LEFclass PAD POWER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
