magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -2594 355 2594 393
rect -2594 299 -2558 355
rect -2502 299 -2347 355
rect -2291 299 -2136 355
rect -2080 299 -1926 355
rect -1870 299 -1715 355
rect -1659 299 -1504 355
rect -1448 299 -1293 355
rect -1237 299 -1082 355
rect -1026 299 -872 355
rect -816 299 -661 355
rect -605 299 -450 355
rect -394 299 -239 355
rect -183 299 -28 355
rect 28 299 183 355
rect 239 299 394 355
rect 450 299 605 355
rect 661 299 816 355
rect 872 299 1026 355
rect 1082 299 1237 355
rect 1293 299 1448 355
rect 1504 299 1659 355
rect 1715 299 1870 355
rect 1926 299 2080 355
rect 2136 299 2291 355
rect 2347 299 2502 355
rect 2558 299 2594 355
rect -2594 137 2594 299
rect -2594 81 -2558 137
rect -2502 81 -2347 137
rect -2291 81 -2136 137
rect -2080 81 -1926 137
rect -1870 81 -1715 137
rect -1659 81 -1504 137
rect -1448 81 -1293 137
rect -1237 81 -1082 137
rect -1026 81 -872 137
rect -816 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 816 137
rect 872 81 1026 137
rect 1082 81 1237 137
rect 1293 81 1448 137
rect 1504 81 1659 137
rect 1715 81 1870 137
rect 1926 81 2080 137
rect 2136 81 2291 137
rect 2347 81 2502 137
rect 2558 81 2594 137
rect -2594 -81 2594 81
rect -2594 -137 -2558 -81
rect -2502 -137 -2347 -81
rect -2291 -137 -2136 -81
rect -2080 -137 -1926 -81
rect -1870 -137 -1715 -81
rect -1659 -137 -1504 -81
rect -1448 -137 -1293 -81
rect -1237 -137 -1082 -81
rect -1026 -137 -872 -81
rect -816 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 816 -81
rect 872 -137 1026 -81
rect 1082 -137 1237 -81
rect 1293 -137 1448 -81
rect 1504 -137 1659 -81
rect 1715 -137 1870 -81
rect 1926 -137 2080 -81
rect 2136 -137 2291 -81
rect 2347 -137 2502 -81
rect 2558 -137 2594 -81
rect -2594 -299 2594 -137
rect -2594 -355 -2558 -299
rect -2502 -355 -2347 -299
rect -2291 -355 -2136 -299
rect -2080 -355 -1926 -299
rect -1870 -355 -1715 -299
rect -1659 -355 -1504 -299
rect -1448 -355 -1293 -299
rect -1237 -355 -1082 -299
rect -1026 -355 -872 -299
rect -816 -355 -661 -299
rect -605 -355 -450 -299
rect -394 -355 -239 -299
rect -183 -355 -28 -299
rect 28 -355 183 -299
rect 239 -355 394 -299
rect 450 -355 605 -299
rect 661 -355 816 -299
rect 872 -355 1026 -299
rect 1082 -355 1237 -299
rect 1293 -355 1448 -299
rect 1504 -355 1659 -299
rect 1715 -355 1870 -299
rect 1926 -355 2080 -299
rect 2136 -355 2291 -299
rect 2347 -355 2502 -299
rect 2558 -355 2594 -299
rect -2594 -393 2594 -355
<< via2 >>
rect -2558 299 -2502 355
rect -2347 299 -2291 355
rect -2136 299 -2080 355
rect -1926 299 -1870 355
rect -1715 299 -1659 355
rect -1504 299 -1448 355
rect -1293 299 -1237 355
rect -1082 299 -1026 355
rect -872 299 -816 355
rect -661 299 -605 355
rect -450 299 -394 355
rect -239 299 -183 355
rect -28 299 28 355
rect 183 299 239 355
rect 394 299 450 355
rect 605 299 661 355
rect 816 299 872 355
rect 1026 299 1082 355
rect 1237 299 1293 355
rect 1448 299 1504 355
rect 1659 299 1715 355
rect 1870 299 1926 355
rect 2080 299 2136 355
rect 2291 299 2347 355
rect 2502 299 2558 355
rect -2558 81 -2502 137
rect -2347 81 -2291 137
rect -2136 81 -2080 137
rect -1926 81 -1870 137
rect -1715 81 -1659 137
rect -1504 81 -1448 137
rect -1293 81 -1237 137
rect -1082 81 -1026 137
rect -872 81 -816 137
rect -661 81 -605 137
rect -450 81 -394 137
rect -239 81 -183 137
rect -28 81 28 137
rect 183 81 239 137
rect 394 81 450 137
rect 605 81 661 137
rect 816 81 872 137
rect 1026 81 1082 137
rect 1237 81 1293 137
rect 1448 81 1504 137
rect 1659 81 1715 137
rect 1870 81 1926 137
rect 2080 81 2136 137
rect 2291 81 2347 137
rect 2502 81 2558 137
rect -2558 -137 -2502 -81
rect -2347 -137 -2291 -81
rect -2136 -137 -2080 -81
rect -1926 -137 -1870 -81
rect -1715 -137 -1659 -81
rect -1504 -137 -1448 -81
rect -1293 -137 -1237 -81
rect -1082 -137 -1026 -81
rect -872 -137 -816 -81
rect -661 -137 -605 -81
rect -450 -137 -394 -81
rect -239 -137 -183 -81
rect -28 -137 28 -81
rect 183 -137 239 -81
rect 394 -137 450 -81
rect 605 -137 661 -81
rect 816 -137 872 -81
rect 1026 -137 1082 -81
rect 1237 -137 1293 -81
rect 1448 -137 1504 -81
rect 1659 -137 1715 -81
rect 1870 -137 1926 -81
rect 2080 -137 2136 -81
rect 2291 -137 2347 -81
rect 2502 -137 2558 -81
rect -2558 -355 -2502 -299
rect -2347 -355 -2291 -299
rect -2136 -355 -2080 -299
rect -1926 -355 -1870 -299
rect -1715 -355 -1659 -299
rect -1504 -355 -1448 -299
rect -1293 -355 -1237 -299
rect -1082 -355 -1026 -299
rect -872 -355 -816 -299
rect -661 -355 -605 -299
rect -450 -355 -394 -299
rect -239 -355 -183 -299
rect -28 -355 28 -299
rect 183 -355 239 -299
rect 394 -355 450 -299
rect 605 -355 661 -299
rect 816 -355 872 -299
rect 1026 -355 1082 -299
rect 1237 -355 1293 -299
rect 1448 -355 1504 -299
rect 1659 -355 1715 -299
rect 1870 -355 1926 -299
rect 2080 -355 2136 -299
rect 2291 -355 2347 -299
rect 2502 -355 2558 -299
<< metal3 >>
rect -2594 355 2594 393
rect -2594 299 -2558 355
rect -2502 299 -2347 355
rect -2291 299 -2136 355
rect -2080 299 -1926 355
rect -1870 299 -1715 355
rect -1659 299 -1504 355
rect -1448 299 -1293 355
rect -1237 299 -1082 355
rect -1026 299 -872 355
rect -816 299 -661 355
rect -605 299 -450 355
rect -394 299 -239 355
rect -183 299 -28 355
rect 28 299 183 355
rect 239 299 394 355
rect 450 299 605 355
rect 661 299 816 355
rect 872 299 1026 355
rect 1082 299 1237 355
rect 1293 299 1448 355
rect 1504 299 1659 355
rect 1715 299 1870 355
rect 1926 299 2080 355
rect 2136 299 2291 355
rect 2347 299 2502 355
rect 2558 299 2594 355
rect -2594 137 2594 299
rect -2594 81 -2558 137
rect -2502 81 -2347 137
rect -2291 81 -2136 137
rect -2080 81 -1926 137
rect -1870 81 -1715 137
rect -1659 81 -1504 137
rect -1448 81 -1293 137
rect -1237 81 -1082 137
rect -1026 81 -872 137
rect -816 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 816 137
rect 872 81 1026 137
rect 1082 81 1237 137
rect 1293 81 1448 137
rect 1504 81 1659 137
rect 1715 81 1870 137
rect 1926 81 2080 137
rect 2136 81 2291 137
rect 2347 81 2502 137
rect 2558 81 2594 137
rect -2594 -81 2594 81
rect -2594 -137 -2558 -81
rect -2502 -137 -2347 -81
rect -2291 -137 -2136 -81
rect -2080 -137 -1926 -81
rect -1870 -137 -1715 -81
rect -1659 -137 -1504 -81
rect -1448 -137 -1293 -81
rect -1237 -137 -1082 -81
rect -1026 -137 -872 -81
rect -816 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 816 -81
rect 872 -137 1026 -81
rect 1082 -137 1237 -81
rect 1293 -137 1448 -81
rect 1504 -137 1659 -81
rect 1715 -137 1870 -81
rect 1926 -137 2080 -81
rect 2136 -137 2291 -81
rect 2347 -137 2502 -81
rect 2558 -137 2594 -81
rect -2594 -299 2594 -137
rect -2594 -355 -2558 -299
rect -2502 -355 -2347 -299
rect -2291 -355 -2136 -299
rect -2080 -355 -1926 -299
rect -1870 -355 -1715 -299
rect -1659 -355 -1504 -299
rect -1448 -355 -1293 -299
rect -1237 -355 -1082 -299
rect -1026 -355 -872 -299
rect -816 -355 -661 -299
rect -605 -355 -450 -299
rect -394 -355 -239 -299
rect -183 -355 -28 -299
rect 28 -355 183 -299
rect 239 -355 394 -299
rect 450 -355 605 -299
rect 661 -355 816 -299
rect 872 -355 1026 -299
rect 1082 -355 1237 -299
rect 1293 -355 1448 -299
rect 1504 -355 1659 -299
rect 1715 -355 1870 -299
rect 1926 -355 2080 -299
rect 2136 -355 2291 -299
rect 2347 -355 2502 -299
rect 2558 -355 2594 -299
rect -2594 -393 2594 -355
<< properties >>
string GDS_END 645080
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 638548
<< end >>
