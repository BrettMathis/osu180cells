magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 2438 1094
<< pwell >>
rect -86 -86 2438 453
<< mvnmos >>
rect 124 149 244 307
rect 384 167 504 307
rect 552 167 672 307
rect 776 167 896 307
rect 944 167 1064 307
rect 1204 149 1324 307
rect 1372 149 1492 307
rect 1746 175 1866 333
rect 2015 69 2135 333
<< mvpmos >>
rect 144 597 244 873
rect 384 673 484 873
rect 532 673 632 873
rect 736 673 836 873
rect 916 673 1016 873
rect 1204 597 1304 873
rect 1408 597 1508 873
rect 1775 573 1875 849
rect 2015 573 2115 939
<< mvndiff >>
rect 36 226 124 307
rect 36 180 49 226
rect 95 180 124 226
rect 36 149 124 180
rect 244 226 384 307
rect 244 180 273 226
rect 319 180 384 226
rect 244 167 384 180
rect 504 167 552 307
rect 672 226 776 307
rect 672 180 701 226
rect 747 180 776 226
rect 672 167 776 180
rect 896 167 944 307
rect 1064 226 1204 307
rect 1064 180 1093 226
rect 1139 180 1204 226
rect 1064 167 1204 180
rect 244 149 324 167
rect 1124 149 1204 167
rect 1324 149 1372 307
rect 1492 226 1580 307
rect 1492 180 1521 226
rect 1567 180 1580 226
rect 1492 149 1580 180
rect 1658 234 1746 333
rect 1658 188 1671 234
rect 1717 188 1746 234
rect 1658 175 1746 188
rect 1866 233 2015 333
rect 1866 187 1940 233
rect 1986 187 2015 233
rect 1866 175 2015 187
rect 1935 69 2015 175
rect 2135 320 2223 333
rect 2135 180 2164 320
rect 2210 180 2223 320
rect 2135 69 2223 180
<< mvpdiff >>
rect 56 835 144 873
rect 56 695 69 835
rect 115 695 144 835
rect 56 597 144 695
rect 244 835 384 873
rect 244 695 273 835
rect 319 695 384 835
rect 244 673 384 695
rect 484 673 532 873
rect 632 835 736 873
rect 632 695 661 835
rect 707 695 736 835
rect 632 673 736 695
rect 836 673 916 873
rect 1016 835 1204 873
rect 1016 695 1045 835
rect 1091 695 1204 835
rect 1016 673 1204 695
rect 244 597 324 673
rect 1124 597 1204 673
rect 1304 835 1408 873
rect 1304 695 1333 835
rect 1379 695 1408 835
rect 1304 597 1408 695
rect 1508 835 1596 873
rect 1935 849 2015 939
rect 1508 695 1537 835
rect 1583 695 1596 835
rect 1508 597 1596 695
rect 1687 835 1775 849
rect 1687 695 1700 835
rect 1746 695 1775 835
rect 1687 573 1775 695
rect 1875 835 2015 849
rect 1875 695 1914 835
rect 1960 695 2015 835
rect 1875 573 2015 695
rect 2115 835 2203 939
rect 2115 695 2144 835
rect 2190 695 2203 835
rect 2115 573 2203 695
<< mvndiffc >>
rect 49 180 95 226
rect 273 180 319 226
rect 701 180 747 226
rect 1093 180 1139 226
rect 1521 180 1567 226
rect 1671 188 1717 234
rect 1940 187 1986 233
rect 2164 180 2210 320
<< mvpdiffc >>
rect 69 695 115 835
rect 273 695 319 835
rect 661 695 707 835
rect 1045 695 1091 835
rect 1333 695 1379 835
rect 1537 695 1583 835
rect 1700 695 1746 835
rect 1914 695 1960 835
rect 2144 695 2190 835
<< polysilicon >>
rect 2015 939 2115 983
rect 144 873 244 917
rect 384 873 484 917
rect 532 873 632 917
rect 736 873 836 917
rect 916 873 1016 917
rect 1204 873 1304 917
rect 1408 873 1508 917
rect 144 432 244 597
rect 144 386 157 432
rect 203 386 244 432
rect 144 351 244 386
rect 124 307 244 351
rect 384 432 484 673
rect 532 627 632 673
rect 532 581 545 627
rect 591 581 632 627
rect 736 640 836 673
rect 736 594 749 640
rect 795 594 836 640
rect 916 629 1016 673
rect 736 581 836 594
rect 532 533 632 581
rect 532 493 896 533
rect 384 386 397 432
rect 443 386 484 432
rect 384 351 484 386
rect 552 432 672 445
rect 552 386 613 432
rect 659 386 672 432
rect 384 307 504 351
rect 552 307 672 386
rect 776 307 896 493
rect 944 432 1016 629
rect 1775 849 1875 893
rect 944 386 957 432
rect 1003 386 1016 432
rect 944 351 1016 386
rect 1204 432 1304 597
rect 1408 553 1508 597
rect 1408 445 1492 553
rect 1775 529 1875 573
rect 1775 445 1865 529
rect 1204 386 1217 432
rect 1263 386 1304 432
rect 1204 351 1304 386
rect 1372 432 1492 445
rect 1372 386 1385 432
rect 1431 386 1492 432
rect 944 307 1064 351
rect 1204 307 1324 351
rect 1372 307 1492 386
rect 1746 432 1865 445
rect 1746 386 1759 432
rect 1805 386 1865 432
rect 1746 377 1865 386
rect 2015 432 2115 573
rect 2015 386 2028 432
rect 2074 386 2115 432
rect 2015 377 2115 386
rect 1746 333 1866 377
rect 2015 333 2135 377
rect 124 105 244 149
rect 384 123 504 167
rect 552 123 672 167
rect 776 123 896 167
rect 944 123 1064 167
rect 1204 105 1324 149
rect 1372 105 1492 149
rect 1746 131 1866 175
rect 2015 25 2135 69
<< polycontact >>
rect 157 386 203 432
rect 545 581 591 627
rect 749 594 795 640
rect 397 386 443 432
rect 613 386 659 432
rect 957 386 1003 432
rect 1217 386 1263 432
rect 1385 386 1431 432
rect 1759 386 1805 432
rect 2028 386 2074 432
<< metal1 >>
rect 0 918 2352 1098
rect 49 835 115 846
rect 49 695 69 835
rect 49 638 115 695
rect 273 835 319 918
rect 273 684 319 695
rect 661 835 898 846
rect 707 800 898 835
rect 661 684 707 695
rect 49 627 591 638
rect 49 581 545 627
rect 49 570 591 581
rect 738 594 749 640
rect 795 594 806 640
rect 49 226 95 570
rect 142 478 659 524
rect 142 432 203 478
rect 613 432 659 478
rect 142 386 157 432
rect 142 354 203 386
rect 366 386 397 432
rect 443 386 454 432
rect 366 242 454 386
rect 738 418 806 594
rect 659 386 806 418
rect 613 366 806 386
rect 852 237 898 800
rect 1045 835 1091 918
rect 1045 684 1091 695
rect 1333 835 1379 846
rect 1333 535 1379 695
rect 1537 835 1583 918
rect 1537 684 1583 695
rect 1700 835 1746 846
rect 1700 641 1746 695
rect 1914 835 1960 918
rect 1914 684 1960 695
rect 2144 835 2210 846
rect 2190 695 2210 835
rect 1700 595 1897 641
rect 1125 524 1379 535
rect 1125 489 1567 524
rect 1125 443 1171 489
rect 1349 478 1567 489
rect 1521 443 1567 478
rect 957 432 1171 443
rect 1003 386 1171 432
rect 957 375 1171 386
rect 1217 432 1263 443
rect 1521 432 1805 443
rect 1217 329 1263 386
rect 49 169 95 180
rect 273 226 319 237
rect 273 90 319 180
rect 701 226 898 237
rect 747 215 898 226
rect 1001 283 1263 329
rect 1374 386 1385 432
rect 1431 386 1442 432
rect 1001 215 1047 283
rect 1374 242 1442 386
rect 1521 386 1759 432
rect 1521 375 1805 386
rect 1851 387 1897 595
rect 2028 432 2074 443
rect 1851 386 2028 387
rect 747 180 1047 215
rect 701 169 1047 180
rect 1093 226 1139 237
rect 1093 90 1139 180
rect 1521 226 1567 375
rect 1851 358 2074 386
rect 1848 341 2074 358
rect 1848 245 1894 341
rect 1521 169 1567 180
rect 1671 234 1894 245
rect 2144 320 2210 695
rect 1717 188 1894 234
rect 1671 177 1894 188
rect 1940 233 1986 244
rect 1940 90 1986 187
rect 2144 180 2164 320
rect 2144 169 2210 180
rect 0 -90 2352 90
<< labels >>
flabel metal1 s 366 242 454 432 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 738 524 806 640 0 FreeSans 200 0 0 0 E
port 2 nsew clock input
flabel metal1 s 2144 169 2210 846 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 1374 242 1442 432 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 2352 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1940 237 1986 244 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 738 478 806 524 1 E
port 2 nsew clock input
rlabel metal1 s 142 478 659 524 1 E
port 2 nsew clock input
rlabel metal1 s 738 418 806 478 1 E
port 2 nsew clock input
rlabel metal1 s 613 418 659 478 1 E
port 2 nsew clock input
rlabel metal1 s 142 418 203 478 1 E
port 2 nsew clock input
rlabel metal1 s 613 366 806 418 1 E
port 2 nsew clock input
rlabel metal1 s 142 366 203 418 1 E
port 2 nsew clock input
rlabel metal1 s 142 354 203 366 1 E
port 2 nsew clock input
rlabel metal1 s 1914 684 1960 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1537 684 1583 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1045 684 1091 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 684 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1940 90 1986 237 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1093 90 1139 237 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 237 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2352 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2352 1008
string GDS_END 1034528
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1028492
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
