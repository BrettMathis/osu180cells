magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -81 106 81 112
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -112 81 -106
<< via1 >>
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
<< metal2 >>
rect -81 106 81 112
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -112 81 -106
<< properties >>
string GDS_END 2001788
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2000888
<< end >>
