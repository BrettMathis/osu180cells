magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -156 2270 4862 3006
rect -156 0 4862 694
<< mvpdiff >>
rect 1782 2411 1839 2603
rect 2083 2411 2140 2603
<< mvpsubdiff >>
rect -39 2021 45 2040
rect -39 1881 -20 2021
rect 26 1881 45 2021
rect -39 1862 45 1881
rect 4842 2021 4926 2040
rect 4842 1881 4861 2021
rect 4907 1881 4926 2021
rect 4842 1862 4926 1881
rect -39 1094 45 1113
rect -39 954 -20 1094
rect 26 954 45 1094
rect -39 935 45 954
rect 1422 1094 1506 1113
rect 1422 954 1441 1094
rect 1487 954 1506 1094
rect 1422 935 1506 954
rect 2144 1094 2228 1113
rect 2144 954 2163 1094
rect 2209 954 2228 1094
rect 3359 1094 3443 1113
rect 2144 935 2228 954
rect 3359 954 3378 1094
rect 3424 954 3443 1094
rect 3359 935 3443 954
<< mvnsubdiff >>
rect -77 2754 77 2811
rect -77 2708 -23 2754
rect 23 2708 77 2754
rect -77 2590 77 2708
rect -77 2544 -23 2590
rect 23 2544 77 2590
rect -77 2488 77 2544
rect 4629 2754 4783 2811
rect 4629 2708 4683 2754
rect 4729 2708 4783 2754
rect 4629 2590 4783 2708
rect 4629 2544 4683 2590
rect 4729 2544 4783 2590
rect 4629 2488 4783 2544
rect -77 471 77 528
rect -77 425 -23 471
rect 23 425 77 471
rect -77 307 77 425
rect -77 261 -23 307
rect 23 261 77 307
rect -77 205 77 261
rect 1389 471 1543 528
rect 1389 425 1443 471
rect 1489 425 1543 471
rect 1389 307 1543 425
rect 1389 261 1443 307
rect 1489 261 1543 307
rect 1389 205 1543 261
rect 3324 471 3478 528
rect 3324 425 3378 471
rect 3424 425 3478 471
rect 3324 307 3478 425
rect 3324 261 3378 307
rect 3424 261 3478 307
rect 3665 461 3749 480
rect 3665 321 3684 461
rect 3730 321 3749 461
rect 3665 302 3749 321
rect 3324 205 3478 261
<< mvpsubdiffcont >>
rect -20 1881 26 2021
rect 4861 1881 4907 2021
rect -20 954 26 1094
rect 1441 954 1487 1094
rect 2163 954 2209 1094
rect 3378 954 3424 1094
<< mvnsubdiffcont >>
rect -23 2708 23 2754
rect -23 2544 23 2590
rect 4683 2708 4729 2754
rect 4683 2544 4729 2590
rect -23 425 23 471
rect -23 261 23 307
rect 1443 425 1489 471
rect 1443 261 1489 307
rect 3378 425 3424 471
rect 3378 261 3424 307
rect 3684 321 3730 461
<< polysilicon >>
rect 1025 3027 1999 3088
rect 295 2998 473 3017
rect 295 2952 314 2998
rect 454 2952 473 2998
rect 295 2933 473 2952
rect 353 2865 473 2933
rect 577 2865 697 2938
rect 1025 2892 1145 3027
rect 1879 2604 1999 3027
rect 353 2079 473 2411
rect 353 2054 472 2079
rect 353 1708 473 1781
rect 577 1647 697 2411
rect 1025 2323 1145 2387
rect 774 2304 1145 2323
rect 774 2258 793 2304
rect 933 2258 1145 2304
rect 774 2239 1145 2258
rect 1025 2072 1145 2239
rect 1239 2332 1819 2351
rect 1239 2192 1258 2332
rect 1304 2290 1819 2332
rect 1304 2192 1323 2290
rect 1756 2253 1819 2290
rect 2218 2323 2338 2387
rect 2218 2304 2562 2323
rect 2218 2258 2403 2304
rect 2543 2258 2562 2304
rect 1756 2192 2114 2253
rect 2218 2239 2562 2258
rect 1239 2173 1323 2192
rect 2218 2151 2338 2239
rect 1025 2054 1144 2072
rect 1025 1856 1144 1862
rect 577 1628 755 1647
rect 577 1582 596 1628
rect 736 1582 755 1628
rect 577 1563 755 1582
rect 1025 1617 1145 1856
rect 2666 1733 2785 2947
rect 2665 1711 2785 1733
rect 2271 1692 2785 1711
rect 2271 1646 2290 1692
rect 2430 1646 2785 1692
rect 2271 1627 2785 1646
rect 2890 1711 3010 2384
rect 3338 2323 3458 2511
rect 3562 2351 3682 2511
rect 4010 2351 4130 2411
rect 4234 2351 4354 2411
rect 3562 2323 4578 2351
rect 3338 2321 4578 2323
rect 3199 2302 4578 2321
rect 3199 2256 3218 2302
rect 3358 2290 4578 2302
rect 3358 2256 3682 2290
rect 3199 2237 3682 2256
rect 3562 2129 3682 2237
rect 4458 2129 4578 2290
rect 2890 1692 3068 1711
rect 2890 1646 2909 1692
rect 3049 1646 3068 1692
rect 2890 1627 3068 1646
rect 3483 1617 3661 1635
rect 4010 1617 4130 1660
rect 4234 1617 4354 1654
rect 1025 1556 1652 1617
rect 3483 1616 4354 1617
rect 3483 1570 3502 1616
rect 3642 1570 4354 1616
rect 3483 1551 4354 1570
rect 1784 1435 1904 1454
rect 577 1397 755 1416
rect 577 1351 596 1397
rect 736 1351 755 1397
rect 577 1332 755 1351
rect 353 590 473 1014
rect 577 590 697 1332
rect 1784 1295 1822 1435
rect 1868 1295 1904 1435
rect 1784 1161 1904 1295
rect 1025 790 1145 904
rect 847 771 1145 790
rect 847 725 866 771
rect 1006 725 1145 771
rect 847 706 1145 725
rect 1025 589 1145 706
rect 1784 765 1904 904
rect 2544 790 2664 960
rect 2407 771 2664 790
rect 1784 660 2128 765
rect 2407 725 2426 771
rect 2566 765 2664 771
rect 2768 765 2888 960
rect 2992 765 3112 960
rect 2566 725 3112 765
rect 2407 706 3112 725
rect 1784 589 1904 660
rect 2008 593 2128 660
rect 2544 660 3112 706
rect 2544 589 2664 660
rect 2768 589 2888 660
rect 2992 589 3112 660
rect 353 60 473 120
rect 295 41 473 60
rect 295 -5 314 41
rect 454 -5 473 41
rect 295 -24 473 -5
<< polycontact >>
rect 314 2952 454 2998
rect 793 2258 933 2304
rect 1258 2192 1304 2332
rect 2403 2258 2543 2304
rect 596 1582 736 1628
rect 2290 1646 2430 1692
rect 3218 2256 3358 2302
rect 2909 1646 3049 1692
rect 3502 1570 3642 1616
rect 596 1351 736 1397
rect 1822 1295 1868 1435
rect 866 725 1006 771
rect 2426 725 2566 771
rect 314 -5 454 41
<< metal1 >>
rect 303 3154 4245 3287
rect 303 2998 465 3154
rect 303 2952 314 2998
rect 454 2952 465 2998
rect 303 2941 465 2952
rect -65 2784 65 2825
rect -65 2732 -26 2784
rect 26 2732 65 2784
rect -65 2708 -23 2732
rect 23 2708 65 2732
rect -65 2590 65 2708
rect -65 2566 -23 2590
rect 23 2566 65 2590
rect -65 2514 -26 2566
rect 26 2514 65 2566
rect -65 2474 65 2514
rect 236 2773 366 2865
rect 236 2721 275 2773
rect 327 2721 366 2773
rect 236 2555 366 2721
rect 236 2503 275 2555
rect 327 2503 366 2555
rect 236 2420 366 2503
rect 691 2331 806 2865
rect 908 2814 1037 2865
rect 908 2773 1038 2814
rect 908 2721 947 2773
rect 999 2721 1038 2773
rect 908 2555 1038 2721
rect 908 2503 947 2555
rect 999 2503 1038 2555
rect 908 2463 1038 2503
rect 908 2420 1037 2463
rect 467 2315 806 2331
rect 1132 2343 1261 2865
rect 1416 2732 1544 2865
rect 1416 2680 1454 2732
rect 1506 2680 1544 2732
rect 1416 2515 1544 2680
rect 1416 2463 1454 2515
rect 1506 2463 1544 2515
rect 1132 2332 1315 2343
rect 467 2304 944 2315
rect 467 2258 793 2304
rect 933 2258 944 2304
rect 467 2247 944 2258
rect -65 2082 65 2123
rect -65 2030 -26 2082
rect 26 2030 65 2082
rect -65 2021 65 2030
rect -65 1881 -20 2021
rect 26 1881 65 2021
rect -65 1864 65 1881
rect -65 1812 -26 1864
rect 26 1812 65 1864
rect -65 1772 65 1812
rect 236 2082 366 2123
rect 236 2030 275 2082
rect 327 2030 366 2082
rect 236 1864 366 2030
rect 236 1812 275 1864
rect 327 1812 366 1864
rect 236 1772 366 1812
rect 467 1781 582 2247
rect 1132 2192 1258 2332
rect 1304 2192 1315 2332
rect 1132 2181 1315 2192
rect 1416 2297 1544 2463
rect 1416 2245 1454 2297
rect 1506 2245 1544 2297
rect 685 2081 813 2122
rect 685 2029 723 2081
rect 775 2029 813 2081
rect 685 1895 813 2029
rect 685 1843 723 1895
rect 775 1843 813 1895
rect 685 1642 813 1843
rect 909 2081 1037 2122
rect 909 2029 947 2081
rect 999 2029 1037 2081
rect 909 1895 1037 2029
rect 909 1843 947 1895
rect 999 1843 1037 1895
rect 1132 1863 1261 2181
rect 1416 2079 1544 2245
rect 1416 2027 1454 2079
rect 1506 2027 1544 2079
rect 909 1803 1037 1843
rect 1416 1862 1544 2027
rect 1416 1810 1454 1862
rect 1506 1810 1544 1862
rect 582 1630 813 1642
rect 582 1578 594 1630
rect 646 1628 726 1630
rect 646 1578 726 1582
rect 778 1578 813 1630
rect 1416 1579 1544 1810
rect 1640 2603 1768 2865
rect 2143 2603 2189 2865
rect 1640 2411 1849 2603
rect 2028 2411 2189 2603
rect 2324 2773 2454 2865
rect 2324 2721 2363 2773
rect 2415 2721 2454 2773
rect 2324 2555 2454 2721
rect 2324 2503 2363 2555
rect 2415 2503 2454 2555
rect 2324 2420 2454 2503
rect 1640 2132 1768 2411
rect 1640 1940 1999 2132
rect 2143 1940 2189 2411
rect 2549 2315 2677 2865
rect 2772 2773 2902 2865
rect 2772 2721 2811 2773
rect 2863 2721 2902 2773
rect 2772 2555 2902 2721
rect 2772 2503 2811 2555
rect 2863 2503 2902 2555
rect 2772 2420 2902 2503
rect 2392 2304 2677 2315
rect 2392 2258 2403 2304
rect 2543 2258 2677 2304
rect 2392 2247 2677 2258
rect 2325 2081 2453 2122
rect 2325 2029 2363 2081
rect 2415 2029 2453 2081
rect 1640 1703 1768 1940
rect 2325 1895 2453 2029
rect 2325 1843 2363 1895
rect 2415 1843 2453 1895
rect 2325 1803 2453 1843
rect 2549 1703 2677 2247
rect 2997 2313 3125 2865
rect 3220 2816 3350 2857
rect 3220 2764 3259 2816
rect 3311 2764 3350 2816
rect 3220 2598 3350 2764
rect 3220 2546 3259 2598
rect 3311 2546 3350 2598
rect 3220 2506 3350 2546
rect 2997 2302 3369 2313
rect 2997 2256 3218 2302
rect 3358 2256 3369 2302
rect 2997 2245 3369 2256
rect 2773 2081 2901 2122
rect 2773 2029 2811 2081
rect 2863 2029 2901 2081
rect 2773 1895 2901 2029
rect 2997 1940 3125 2245
rect 2773 1843 2811 1895
rect 2863 1843 2901 1895
rect 2773 1803 2901 1843
rect 1640 1692 2453 1703
rect 1640 1646 2290 1692
rect 2430 1646 2453 1692
rect 1640 1635 2453 1646
rect 2549 1692 3068 1703
rect 2549 1646 2909 1692
rect 3049 1646 3068 1692
rect 2549 1635 3068 1646
rect 582 1566 813 1578
rect 1174 1533 1544 1579
rect 3445 1627 3573 2867
rect 3668 2816 3798 2857
rect 3668 2764 3707 2816
rect 3759 2764 3798 2816
rect 3668 2598 3798 2764
rect 3668 2546 3707 2598
rect 3759 2546 3798 2598
rect 3668 2506 3798 2546
rect 3893 2331 4021 2865
rect 4117 2814 4245 3154
rect 4116 2773 4246 2814
rect 4116 2721 4155 2773
rect 4207 2721 4246 2773
rect 4116 2555 4246 2721
rect 4116 2503 4155 2555
rect 4207 2503 4246 2555
rect 4116 2463 4246 2503
rect 4117 2420 4245 2463
rect 4341 2331 4469 2865
rect 4641 2784 4771 2825
rect 4641 2732 4680 2784
rect 4732 2732 4771 2784
rect 4641 2708 4683 2732
rect 4729 2708 4771 2732
rect 4641 2590 4771 2708
rect 4641 2566 4683 2590
rect 4729 2566 4771 2590
rect 4641 2514 4680 2566
rect 4732 2514 4771 2566
rect 4641 2474 4771 2514
rect 3893 2211 4469 2331
rect 3669 2081 3797 2122
rect 3669 2029 3707 2081
rect 3759 2029 3797 2081
rect 3669 1895 3797 2029
rect 3669 1843 3707 1895
rect 3759 1843 3797 1895
rect 3669 1803 3797 1843
rect 3445 1616 3653 1627
rect 3445 1570 3502 1616
rect 3642 1570 3653 1616
rect 3445 1559 3653 1570
rect 582 1399 790 1411
rect 582 1347 594 1399
rect 646 1397 726 1399
rect 646 1347 726 1351
rect 778 1347 790 1399
rect 582 1335 790 1347
rect -65 1164 65 1205
rect -65 1112 -26 1164
rect 26 1112 65 1164
rect -65 1094 65 1112
rect -65 954 -20 1094
rect 26 954 65 1094
rect -65 946 65 954
rect -65 894 -26 946
rect 26 894 65 946
rect -65 854 65 894
rect 236 1163 366 1204
rect 236 1111 275 1163
rect 327 1111 366 1163
rect 236 945 366 1111
rect 685 1163 813 1204
rect 685 1111 723 1163
rect 775 1111 813 1163
rect 236 893 275 945
rect 327 893 366 945
rect 236 853 366 893
rect 502 771 548 1097
rect 685 977 813 1111
rect 685 925 723 977
rect 775 925 813 977
rect 685 885 813 925
rect 908 1163 1036 1204
rect 908 1111 946 1163
rect 998 1111 1036 1163
rect 908 977 1036 1111
rect 908 925 946 977
rect 998 925 1036 977
rect 908 885 1036 925
rect 855 771 1017 782
rect 502 725 866 771
rect 1006 725 1017 771
rect -65 501 65 542
rect -65 449 -26 501
rect 26 449 65 501
rect -65 425 -23 449
rect 23 425 65 449
rect -65 307 65 425
rect -65 283 -23 307
rect 23 283 65 307
rect -65 231 -26 283
rect 26 231 65 283
rect -65 191 65 231
rect 236 490 366 574
rect 726 538 772 725
rect 855 714 1017 725
rect 236 438 275 490
rect 327 438 366 490
rect 236 272 366 438
rect 236 220 275 272
rect 327 220 366 272
rect 236 120 366 220
rect 907 486 1037 574
rect 907 434 946 486
rect 998 434 1037 486
rect 1174 463 1220 1533
rect 3893 1446 4021 2211
rect 4116 2039 4246 2122
rect 4116 1987 4155 2039
rect 4207 1987 4246 2039
rect 4116 1821 4246 1987
rect 4116 1769 4155 1821
rect 4207 1769 4246 1821
rect 4116 1677 4246 1769
rect 4341 1446 4469 2211
rect 4564 2082 4694 2131
rect 4564 2030 4603 2082
rect 4655 2030 4694 2082
rect 4564 1864 4694 2030
rect 4564 1812 4603 1864
rect 4655 1812 4694 1864
rect 4564 1677 4694 1812
rect 4816 2082 4946 2123
rect 4816 2030 4855 2082
rect 4907 2030 4946 2082
rect 4816 2021 4946 2030
rect 4816 1881 4861 2021
rect 4907 1881 4946 2021
rect 4816 1864 4946 1881
rect 4816 1812 4855 1864
rect 4907 1812 4946 1864
rect 4816 1772 4946 1812
rect 1811 1435 4469 1446
rect 1811 1295 1822 1435
rect 1868 1400 4469 1435
rect 1868 1295 1879 1400
rect 1811 1284 1879 1295
rect 1401 1164 1531 1205
rect 1401 1112 1440 1164
rect 1492 1112 1531 1164
rect 1401 1094 1531 1112
rect 1401 954 1441 1094
rect 1487 954 1531 1094
rect 1401 946 1531 954
rect 1401 894 1440 946
rect 1492 894 1531 946
rect 1401 854 1531 894
rect 1668 1163 1796 1204
rect 1668 1111 1706 1163
rect 1758 1111 1796 1163
rect 1668 977 1796 1111
rect 2119 1164 2249 1205
rect 2119 1112 2158 1164
rect 2210 1112 2249 1164
rect 2119 1094 2249 1112
rect 1668 925 1706 977
rect 1758 925 1796 977
rect 1668 885 1796 925
rect 1933 771 1979 999
rect 2119 954 2163 1094
rect 2209 954 2249 1094
rect 2119 946 2249 954
rect 2119 894 2158 946
rect 2210 894 2249 946
rect 2119 854 2249 894
rect 2428 1163 2556 1204
rect 2428 1111 2466 1163
rect 2518 1111 2556 1163
rect 2428 977 2556 1111
rect 2876 1163 3004 1204
rect 2876 1111 2914 1163
rect 2966 1111 3004 1163
rect 2428 925 2466 977
rect 2518 925 2556 977
rect 2428 885 2556 925
rect 2693 785 2739 999
rect 2876 977 3004 1111
rect 3336 1164 3466 1205
rect 3336 1112 3375 1164
rect 3427 1112 3466 1164
rect 3336 1094 3466 1112
rect 2876 925 2914 977
rect 2966 925 3004 977
rect 2876 885 3004 925
rect 3141 785 3187 999
rect 3336 954 3378 1094
rect 3424 954 3466 1094
rect 3336 946 3466 954
rect 3336 894 3375 946
rect 3427 894 3466 946
rect 3336 854 3466 894
rect 2415 771 2577 782
rect 1933 725 2426 771
rect 2566 725 2577 771
rect 1401 501 1531 542
rect 907 300 1037 434
rect 907 248 946 300
rect 998 248 1037 300
rect 907 120 1037 248
rect 1401 449 1440 501
rect 1492 449 1531 501
rect 1401 425 1443 449
rect 1489 425 1531 449
rect 1401 307 1531 425
rect 1401 283 1443 307
rect 1489 283 1531 307
rect 1401 231 1440 283
rect 1492 231 1531 283
rect 1401 191 1531 231
rect 1667 486 1797 574
rect 1933 538 1979 725
rect 2415 714 2577 725
rect 2693 665 3617 785
rect 1667 434 1706 486
rect 1758 434 1797 486
rect 1667 300 1797 434
rect 1667 248 1706 300
rect 1758 248 1797 300
rect 1667 120 1797 248
rect 2115 486 2245 574
rect 2115 434 2154 486
rect 2206 434 2245 486
rect 2115 300 2245 434
rect 2115 248 2154 300
rect 2206 248 2245 300
rect 2115 120 2245 248
rect 2427 486 2557 574
rect 2693 538 2739 665
rect 2427 434 2466 486
rect 2518 434 2557 486
rect 2427 300 2557 434
rect 2427 248 2466 300
rect 2518 248 2557 300
rect 2427 120 2557 248
rect 2875 486 3005 574
rect 3141 538 3187 665
rect 2875 434 2914 486
rect 2966 434 3005 486
rect 2875 300 3005 434
rect 2875 248 2914 300
rect 2966 248 3005 300
rect 2875 120 3005 248
rect 3336 501 3466 542
rect 3336 449 3375 501
rect 3427 449 3466 501
rect 3336 425 3378 449
rect 3424 425 3466 449
rect 3336 307 3466 425
rect 3336 283 3378 307
rect 3424 283 3466 307
rect 3336 231 3375 283
rect 3427 231 3466 283
rect 3336 191 3466 231
rect 3646 501 3776 542
rect 3646 461 3685 501
rect 3646 321 3684 461
rect 3737 449 3776 501
rect 3730 321 3776 449
rect 3646 283 3776 321
rect 3646 231 3685 283
rect 3737 231 3776 283
rect 3646 191 3776 231
rect 0 41 465 52
rect 0 -5 314 41
rect 454 -5 465 41
rect 0 -24 465 -5
<< via1 >>
rect -26 2754 26 2784
rect -26 2732 -23 2754
rect -23 2732 23 2754
rect 23 2732 26 2754
rect -26 2544 -23 2566
rect -23 2544 23 2566
rect 23 2544 26 2566
rect -26 2514 26 2544
rect 275 2721 327 2773
rect 275 2503 327 2555
rect 947 2721 999 2773
rect 947 2503 999 2555
rect 1454 2680 1506 2732
rect 1454 2463 1506 2515
rect -26 2030 26 2082
rect -26 1812 26 1864
rect 275 2030 327 2082
rect 275 1812 327 1864
rect 1454 2245 1506 2297
rect 723 2029 775 2081
rect 723 1843 775 1895
rect 947 2029 999 2081
rect 947 1843 999 1895
rect 1454 2027 1506 2079
rect 1454 1810 1506 1862
rect 594 1628 646 1630
rect 726 1628 778 1630
rect 594 1582 596 1628
rect 596 1582 646 1628
rect 726 1582 736 1628
rect 736 1582 778 1628
rect 594 1578 646 1582
rect 726 1578 778 1582
rect 2363 2721 2415 2773
rect 2363 2503 2415 2555
rect 2811 2721 2863 2773
rect 2811 2503 2863 2555
rect 2363 2029 2415 2081
rect 2363 1843 2415 1895
rect 3259 2764 3311 2816
rect 3259 2546 3311 2598
rect 2811 2029 2863 2081
rect 2811 1843 2863 1895
rect 3707 2764 3759 2816
rect 3707 2546 3759 2598
rect 4155 2721 4207 2773
rect 4155 2503 4207 2555
rect 4680 2754 4732 2784
rect 4680 2732 4683 2754
rect 4683 2732 4729 2754
rect 4729 2732 4732 2754
rect 4680 2544 4683 2566
rect 4683 2544 4729 2566
rect 4729 2544 4732 2566
rect 4680 2514 4732 2544
rect 3707 2029 3759 2081
rect 3707 1843 3759 1895
rect 594 1397 646 1399
rect 726 1397 778 1399
rect 594 1351 596 1397
rect 596 1351 646 1397
rect 726 1351 736 1397
rect 736 1351 778 1397
rect 594 1347 646 1351
rect 726 1347 778 1351
rect -26 1112 26 1164
rect -26 894 26 946
rect 275 1111 327 1163
rect 723 1111 775 1163
rect 275 893 327 945
rect 723 925 775 977
rect 946 1111 998 1163
rect 946 925 998 977
rect -26 471 26 501
rect -26 449 -23 471
rect -23 449 23 471
rect 23 449 26 471
rect -26 261 -23 283
rect -23 261 23 283
rect 23 261 26 283
rect -26 231 26 261
rect 275 438 327 490
rect 275 220 327 272
rect 946 434 998 486
rect 4155 1987 4207 2039
rect 4155 1769 4207 1821
rect 4603 2030 4655 2082
rect 4603 1812 4655 1864
rect 4855 2030 4907 2082
rect 4855 1812 4907 1864
rect 1440 1112 1492 1164
rect 1440 894 1492 946
rect 1706 1111 1758 1163
rect 2158 1112 2210 1164
rect 1706 925 1758 977
rect 2158 894 2210 946
rect 2466 1111 2518 1163
rect 2914 1111 2966 1163
rect 2466 925 2518 977
rect 3375 1112 3427 1164
rect 2914 925 2966 977
rect 3375 894 3427 946
rect 946 248 998 300
rect 1440 471 1492 501
rect 1440 449 1443 471
rect 1443 449 1489 471
rect 1489 449 1492 471
rect 1440 261 1443 283
rect 1443 261 1489 283
rect 1489 261 1492 283
rect 1440 231 1492 261
rect 1706 434 1758 486
rect 1706 248 1758 300
rect 2154 434 2206 486
rect 2154 248 2206 300
rect 2466 434 2518 486
rect 2466 248 2518 300
rect 2914 434 2966 486
rect 2914 248 2966 300
rect 3375 471 3427 501
rect 3375 449 3378 471
rect 3378 449 3424 471
rect 3424 449 3427 471
rect 3375 261 3378 283
rect 3378 261 3424 283
rect 3424 261 3427 283
rect 3375 231 3427 261
rect 3685 461 3737 501
rect 3685 449 3730 461
rect 3730 449 3737 461
rect 3685 231 3737 283
<< metal2 >>
rect -65 2786 65 2825
rect -65 2730 -28 2786
rect 28 2730 65 2786
rect -65 2568 65 2730
rect -65 2512 -28 2568
rect 28 2512 65 2568
rect -65 2474 65 2512
rect 236 2775 366 2814
rect 236 2719 273 2775
rect 329 2719 366 2775
rect 236 2557 366 2719
rect 236 2501 273 2557
rect 329 2501 366 2557
rect 236 2463 366 2501
rect 908 2775 1038 2814
rect 908 2719 945 2775
rect 1001 2719 1038 2775
rect 908 2557 1038 2719
rect 908 2501 945 2557
rect 1001 2501 1038 2557
rect 908 2463 1038 2501
rect 1416 2732 1544 2865
rect 3220 2818 3350 2857
rect 1416 2680 1454 2732
rect 1506 2680 1544 2732
rect 1416 2515 1544 2680
rect 1416 2463 1454 2515
rect 1506 2463 1544 2515
rect 2324 2775 2454 2814
rect 2324 2719 2361 2775
rect 2417 2719 2454 2775
rect 2324 2557 2454 2719
rect 2324 2501 2361 2557
rect 2417 2501 2454 2557
rect 2324 2463 2454 2501
rect 2772 2775 2902 2814
rect 2772 2719 2809 2775
rect 2865 2719 2902 2775
rect 2772 2557 2902 2719
rect 2772 2501 2809 2557
rect 2865 2501 2902 2557
rect 3220 2762 3257 2818
rect 3313 2762 3350 2818
rect 3220 2600 3350 2762
rect 3220 2544 3257 2600
rect 3313 2544 3350 2600
rect 3220 2506 3350 2544
rect 3668 2818 3798 2857
rect 3668 2762 3705 2818
rect 3761 2762 3798 2818
rect 3668 2600 3798 2762
rect 3668 2544 3705 2600
rect 3761 2544 3798 2600
rect 3668 2506 3798 2544
rect 4116 2773 4246 2863
rect 4116 2721 4155 2773
rect 4207 2721 4246 2773
rect 4116 2555 4246 2721
rect 2772 2463 2902 2501
rect 4116 2503 4155 2555
rect 4207 2503 4246 2555
rect 1416 2297 1544 2463
rect 1416 2245 1454 2297
rect 1506 2245 1544 2297
rect -65 2084 65 2123
rect -65 2028 -28 2084
rect 28 2028 65 2084
rect -65 1866 65 2028
rect -65 1810 -28 1866
rect 28 1810 65 1866
rect -65 1772 65 1810
rect 236 2084 366 2123
rect 236 2028 273 2084
rect 329 2028 366 2084
rect 236 1866 366 2028
rect 236 1810 273 1866
rect 329 1810 366 1866
rect 236 1772 366 1810
rect 685 2083 813 2122
rect 685 2027 721 2083
rect 777 2027 813 2083
rect 685 1897 813 2027
rect 685 1841 721 1897
rect 777 1841 813 1897
rect 685 1803 813 1841
rect 909 2083 1037 2122
rect 909 2027 945 2083
rect 1001 2027 1037 2083
rect 909 1897 1037 2027
rect 909 1841 945 1897
rect 1001 1841 1037 1897
rect 909 1803 1037 1841
rect 1416 2079 1544 2245
rect 1416 2027 1454 2079
rect 1506 2027 1544 2079
rect 1416 1862 1544 2027
rect 1416 1810 1454 1862
rect 1506 1810 1544 1862
rect 1416 1685 1544 1810
rect 2325 2083 2453 2122
rect 2325 2027 2361 2083
rect 2417 2027 2453 2083
rect 2325 1897 2453 2027
rect 2325 1841 2361 1897
rect 2417 1841 2453 1897
rect 2325 1803 2453 1841
rect 2773 2083 2901 2122
rect 2773 2027 2809 2083
rect 2865 2027 2901 2083
rect 2773 1897 2901 2027
rect 2773 1841 2809 1897
rect 2865 1841 2901 1897
rect 2773 1803 2901 1841
rect 3669 2083 3797 2122
rect 3669 2027 3705 2083
rect 3761 2027 3797 2083
rect 3669 1897 3797 2027
rect 3669 1841 3705 1897
rect 3761 1841 3797 1897
rect 3669 1803 3797 1841
rect 4116 2039 4246 2503
rect 4641 2786 4771 2825
rect 4641 2730 4678 2786
rect 4734 2730 4771 2786
rect 4641 2568 4771 2730
rect 4641 2512 4678 2568
rect 4734 2512 4771 2568
rect 4641 2474 4771 2512
rect 4116 1987 4155 2039
rect 4207 1987 4246 2039
rect 4116 1821 4246 1987
rect 4116 1769 4155 1821
rect 4207 1769 4246 1821
rect 4564 2084 4694 2123
rect 4564 2028 4601 2084
rect 4657 2028 4694 2084
rect 4564 1866 4694 2028
rect 4564 1810 4601 1866
rect 4657 1810 4694 1866
rect 4564 1772 4694 1810
rect 4816 2084 4946 2123
rect 4816 2028 4853 2084
rect 4909 2028 4946 2084
rect 4816 1866 4946 2028
rect 4816 1810 4853 1866
rect 4909 1810 4946 1866
rect 4816 1772 4946 1810
rect 4116 1685 4246 1769
rect 582 1632 790 1642
rect 582 1576 592 1632
rect 648 1576 724 1632
rect 780 1576 790 1632
rect 582 1566 790 1576
rect 582 1401 790 1411
rect 582 1345 592 1401
rect 648 1345 724 1401
rect 780 1345 790 1401
rect 582 1335 790 1345
rect -65 1166 65 1205
rect -65 1110 -28 1166
rect 28 1110 65 1166
rect -65 948 65 1110
rect -65 892 -28 948
rect 28 892 65 948
rect -65 854 65 892
rect 236 1165 366 1204
rect 236 1109 273 1165
rect 329 1109 366 1165
rect 236 947 366 1109
rect 236 891 273 947
rect 329 891 366 947
rect 236 853 366 891
rect 684 1165 814 1204
rect 684 1109 721 1165
rect 777 1109 814 1165
rect 684 977 814 1109
rect 684 947 723 977
rect 775 947 814 977
rect 684 891 721 947
rect 777 891 814 947
rect 684 853 814 891
rect 907 1165 1037 1204
rect 907 1109 944 1165
rect 1000 1109 1037 1165
rect 907 977 1037 1109
rect 907 947 946 977
rect 998 947 1037 977
rect 907 891 944 947
rect 1000 891 1037 947
rect 907 853 1037 891
rect 1401 1166 1531 1205
rect 1401 1110 1438 1166
rect 1494 1110 1531 1166
rect 1401 948 1531 1110
rect 1401 892 1438 948
rect 1494 892 1531 948
rect 1401 854 1531 892
rect 1667 1165 1797 1204
rect 1667 1109 1704 1165
rect 1760 1109 1797 1165
rect 1667 977 1797 1109
rect 1667 947 1706 977
rect 1758 947 1797 977
rect 1667 891 1704 947
rect 1760 891 1797 947
rect 1667 853 1797 891
rect 2119 1166 2249 1205
rect 2119 1110 2156 1166
rect 2212 1110 2249 1166
rect 2119 948 2249 1110
rect 2119 892 2156 948
rect 2212 892 2249 948
rect 2119 854 2249 892
rect 2427 1165 2557 1204
rect 2427 1109 2464 1165
rect 2520 1109 2557 1165
rect 2427 977 2557 1109
rect 2427 947 2466 977
rect 2518 947 2557 977
rect 2427 891 2464 947
rect 2520 891 2557 947
rect 2427 853 2557 891
rect 2875 1165 3005 1204
rect 2875 1109 2912 1165
rect 2968 1109 3005 1165
rect 2875 977 3005 1109
rect 2875 947 2914 977
rect 2966 947 3005 977
rect 2875 891 2912 947
rect 2968 891 3005 947
rect 2875 853 3005 891
rect 3336 1166 3466 1205
rect 3336 1110 3373 1166
rect 3429 1110 3466 1166
rect 3336 948 3466 1110
rect 3336 892 3373 948
rect 3429 892 3466 948
rect 3336 854 3466 892
rect -65 503 65 542
rect -65 447 -28 503
rect 28 447 65 503
rect -65 285 65 447
rect -65 229 -28 285
rect 28 229 65 285
rect -65 191 65 229
rect 236 492 366 531
rect 236 436 273 492
rect 329 436 366 492
rect 236 274 366 436
rect 236 218 273 274
rect 329 218 366 274
rect 236 180 366 218
rect 907 488 1037 527
rect 907 432 944 488
rect 1000 432 1037 488
rect 907 300 1037 432
rect 907 270 946 300
rect 998 270 1037 300
rect 907 214 944 270
rect 1000 214 1037 270
rect 907 176 1037 214
rect 1401 503 1531 542
rect 1401 447 1438 503
rect 1494 447 1531 503
rect 1401 285 1531 447
rect 1401 229 1438 285
rect 1494 229 1531 285
rect 1401 191 1531 229
rect 1667 488 1797 527
rect 1667 432 1704 488
rect 1760 432 1797 488
rect 1667 300 1797 432
rect 1667 270 1706 300
rect 1758 270 1797 300
rect 1667 214 1704 270
rect 1760 214 1797 270
rect 1667 176 1797 214
rect 2115 488 2245 527
rect 2115 432 2152 488
rect 2208 432 2245 488
rect 2115 300 2245 432
rect 2115 270 2154 300
rect 2206 270 2245 300
rect 2115 214 2152 270
rect 2208 214 2245 270
rect 2115 176 2245 214
rect 2427 488 2557 527
rect 2427 432 2464 488
rect 2520 432 2557 488
rect 2427 300 2557 432
rect 2427 270 2466 300
rect 2518 270 2557 300
rect 2427 214 2464 270
rect 2520 214 2557 270
rect 2427 176 2557 214
rect 2875 488 3005 527
rect 2875 432 2912 488
rect 2968 432 3005 488
rect 2875 300 3005 432
rect 2875 270 2914 300
rect 2966 270 3005 300
rect 2875 214 2912 270
rect 2968 214 3005 270
rect 2875 176 3005 214
rect 3336 503 3466 542
rect 3336 447 3373 503
rect 3429 447 3466 503
rect 3336 285 3466 447
rect 3336 229 3373 285
rect 3429 229 3466 285
rect 3336 191 3466 229
rect 3646 503 3776 542
rect 3646 447 3683 503
rect 3739 447 3776 503
rect 3646 285 3776 447
rect 3646 229 3683 285
rect 3739 229 3776 285
rect 3646 191 3776 229
<< via2 >>
rect -28 2784 28 2786
rect -28 2732 -26 2784
rect -26 2732 26 2784
rect 26 2732 28 2784
rect -28 2730 28 2732
rect -28 2566 28 2568
rect -28 2514 -26 2566
rect -26 2514 26 2566
rect 26 2514 28 2566
rect -28 2512 28 2514
rect 273 2773 329 2775
rect 273 2721 275 2773
rect 275 2721 327 2773
rect 327 2721 329 2773
rect 273 2719 329 2721
rect 273 2555 329 2557
rect 273 2503 275 2555
rect 275 2503 327 2555
rect 327 2503 329 2555
rect 273 2501 329 2503
rect 945 2773 1001 2775
rect 945 2721 947 2773
rect 947 2721 999 2773
rect 999 2721 1001 2773
rect 945 2719 1001 2721
rect 945 2555 1001 2557
rect 945 2503 947 2555
rect 947 2503 999 2555
rect 999 2503 1001 2555
rect 945 2501 1001 2503
rect 2361 2773 2417 2775
rect 2361 2721 2363 2773
rect 2363 2721 2415 2773
rect 2415 2721 2417 2773
rect 2361 2719 2417 2721
rect 2361 2555 2417 2557
rect 2361 2503 2363 2555
rect 2363 2503 2415 2555
rect 2415 2503 2417 2555
rect 2361 2501 2417 2503
rect 2809 2773 2865 2775
rect 2809 2721 2811 2773
rect 2811 2721 2863 2773
rect 2863 2721 2865 2773
rect 2809 2719 2865 2721
rect 2809 2555 2865 2557
rect 2809 2503 2811 2555
rect 2811 2503 2863 2555
rect 2863 2503 2865 2555
rect 2809 2501 2865 2503
rect 3257 2816 3313 2818
rect 3257 2764 3259 2816
rect 3259 2764 3311 2816
rect 3311 2764 3313 2816
rect 3257 2762 3313 2764
rect 3257 2598 3313 2600
rect 3257 2546 3259 2598
rect 3259 2546 3311 2598
rect 3311 2546 3313 2598
rect 3257 2544 3313 2546
rect 3705 2816 3761 2818
rect 3705 2764 3707 2816
rect 3707 2764 3759 2816
rect 3759 2764 3761 2816
rect 3705 2762 3761 2764
rect 3705 2598 3761 2600
rect 3705 2546 3707 2598
rect 3707 2546 3759 2598
rect 3759 2546 3761 2598
rect 3705 2544 3761 2546
rect -28 2082 28 2084
rect -28 2030 -26 2082
rect -26 2030 26 2082
rect 26 2030 28 2082
rect -28 2028 28 2030
rect -28 1864 28 1866
rect -28 1812 -26 1864
rect -26 1812 26 1864
rect 26 1812 28 1864
rect -28 1810 28 1812
rect 273 2082 329 2084
rect 273 2030 275 2082
rect 275 2030 327 2082
rect 327 2030 329 2082
rect 273 2028 329 2030
rect 273 1864 329 1866
rect 273 1812 275 1864
rect 275 1812 327 1864
rect 327 1812 329 1864
rect 273 1810 329 1812
rect 721 2081 777 2083
rect 721 2029 723 2081
rect 723 2029 775 2081
rect 775 2029 777 2081
rect 721 2027 777 2029
rect 721 1895 777 1897
rect 721 1843 723 1895
rect 723 1843 775 1895
rect 775 1843 777 1895
rect 721 1841 777 1843
rect 945 2081 1001 2083
rect 945 2029 947 2081
rect 947 2029 999 2081
rect 999 2029 1001 2081
rect 945 2027 1001 2029
rect 945 1895 1001 1897
rect 945 1843 947 1895
rect 947 1843 999 1895
rect 999 1843 1001 1895
rect 945 1841 1001 1843
rect 2361 2081 2417 2083
rect 2361 2029 2363 2081
rect 2363 2029 2415 2081
rect 2415 2029 2417 2081
rect 2361 2027 2417 2029
rect 2361 1895 2417 1897
rect 2361 1843 2363 1895
rect 2363 1843 2415 1895
rect 2415 1843 2417 1895
rect 2361 1841 2417 1843
rect 2809 2081 2865 2083
rect 2809 2029 2811 2081
rect 2811 2029 2863 2081
rect 2863 2029 2865 2081
rect 2809 2027 2865 2029
rect 2809 1895 2865 1897
rect 2809 1843 2811 1895
rect 2811 1843 2863 1895
rect 2863 1843 2865 1895
rect 2809 1841 2865 1843
rect 3705 2081 3761 2083
rect 3705 2029 3707 2081
rect 3707 2029 3759 2081
rect 3759 2029 3761 2081
rect 3705 2027 3761 2029
rect 3705 1895 3761 1897
rect 3705 1843 3707 1895
rect 3707 1843 3759 1895
rect 3759 1843 3761 1895
rect 3705 1841 3761 1843
rect 4678 2784 4734 2786
rect 4678 2732 4680 2784
rect 4680 2732 4732 2784
rect 4732 2732 4734 2784
rect 4678 2730 4734 2732
rect 4678 2566 4734 2568
rect 4678 2514 4680 2566
rect 4680 2514 4732 2566
rect 4732 2514 4734 2566
rect 4678 2512 4734 2514
rect 4601 2082 4657 2084
rect 4601 2030 4603 2082
rect 4603 2030 4655 2082
rect 4655 2030 4657 2082
rect 4601 2028 4657 2030
rect 4601 1864 4657 1866
rect 4601 1812 4603 1864
rect 4603 1812 4655 1864
rect 4655 1812 4657 1864
rect 4601 1810 4657 1812
rect 4853 2082 4909 2084
rect 4853 2030 4855 2082
rect 4855 2030 4907 2082
rect 4907 2030 4909 2082
rect 4853 2028 4909 2030
rect 4853 1864 4909 1866
rect 4853 1812 4855 1864
rect 4855 1812 4907 1864
rect 4907 1812 4909 1864
rect 4853 1810 4909 1812
rect 592 1630 648 1632
rect 592 1578 594 1630
rect 594 1578 646 1630
rect 646 1578 648 1630
rect 592 1576 648 1578
rect 724 1630 780 1632
rect 724 1578 726 1630
rect 726 1578 778 1630
rect 778 1578 780 1630
rect 724 1576 780 1578
rect 592 1399 648 1401
rect 592 1347 594 1399
rect 594 1347 646 1399
rect 646 1347 648 1399
rect 592 1345 648 1347
rect 724 1399 780 1401
rect 724 1347 726 1399
rect 726 1347 778 1399
rect 778 1347 780 1399
rect 724 1345 780 1347
rect -28 1164 28 1166
rect -28 1112 -26 1164
rect -26 1112 26 1164
rect 26 1112 28 1164
rect -28 1110 28 1112
rect -28 946 28 948
rect -28 894 -26 946
rect -26 894 26 946
rect 26 894 28 946
rect -28 892 28 894
rect 273 1163 329 1165
rect 273 1111 275 1163
rect 275 1111 327 1163
rect 327 1111 329 1163
rect 273 1109 329 1111
rect 273 945 329 947
rect 273 893 275 945
rect 275 893 327 945
rect 327 893 329 945
rect 273 891 329 893
rect 721 1163 777 1165
rect 721 1111 723 1163
rect 723 1111 775 1163
rect 775 1111 777 1163
rect 721 1109 777 1111
rect 721 925 723 947
rect 723 925 775 947
rect 775 925 777 947
rect 721 891 777 925
rect 944 1163 1000 1165
rect 944 1111 946 1163
rect 946 1111 998 1163
rect 998 1111 1000 1163
rect 944 1109 1000 1111
rect 944 925 946 947
rect 946 925 998 947
rect 998 925 1000 947
rect 944 891 1000 925
rect 1438 1164 1494 1166
rect 1438 1112 1440 1164
rect 1440 1112 1492 1164
rect 1492 1112 1494 1164
rect 1438 1110 1494 1112
rect 1438 946 1494 948
rect 1438 894 1440 946
rect 1440 894 1492 946
rect 1492 894 1494 946
rect 1438 892 1494 894
rect 1704 1163 1760 1165
rect 1704 1111 1706 1163
rect 1706 1111 1758 1163
rect 1758 1111 1760 1163
rect 1704 1109 1760 1111
rect 1704 925 1706 947
rect 1706 925 1758 947
rect 1758 925 1760 947
rect 1704 891 1760 925
rect 2156 1164 2212 1166
rect 2156 1112 2158 1164
rect 2158 1112 2210 1164
rect 2210 1112 2212 1164
rect 2156 1110 2212 1112
rect 2156 946 2212 948
rect 2156 894 2158 946
rect 2158 894 2210 946
rect 2210 894 2212 946
rect 2156 892 2212 894
rect 2464 1163 2520 1165
rect 2464 1111 2466 1163
rect 2466 1111 2518 1163
rect 2518 1111 2520 1163
rect 2464 1109 2520 1111
rect 2464 925 2466 947
rect 2466 925 2518 947
rect 2518 925 2520 947
rect 2464 891 2520 925
rect 2912 1163 2968 1165
rect 2912 1111 2914 1163
rect 2914 1111 2966 1163
rect 2966 1111 2968 1163
rect 2912 1109 2968 1111
rect 2912 925 2914 947
rect 2914 925 2966 947
rect 2966 925 2968 947
rect 2912 891 2968 925
rect 3373 1164 3429 1166
rect 3373 1112 3375 1164
rect 3375 1112 3427 1164
rect 3427 1112 3429 1164
rect 3373 1110 3429 1112
rect 3373 946 3429 948
rect 3373 894 3375 946
rect 3375 894 3427 946
rect 3427 894 3429 946
rect 3373 892 3429 894
rect -28 501 28 503
rect -28 449 -26 501
rect -26 449 26 501
rect 26 449 28 501
rect -28 447 28 449
rect -28 283 28 285
rect -28 231 -26 283
rect -26 231 26 283
rect 26 231 28 283
rect -28 229 28 231
rect 273 490 329 492
rect 273 438 275 490
rect 275 438 327 490
rect 327 438 329 490
rect 273 436 329 438
rect 273 272 329 274
rect 273 220 275 272
rect 275 220 327 272
rect 327 220 329 272
rect 273 218 329 220
rect 944 486 1000 488
rect 944 434 946 486
rect 946 434 998 486
rect 998 434 1000 486
rect 944 432 1000 434
rect 944 248 946 270
rect 946 248 998 270
rect 998 248 1000 270
rect 944 214 1000 248
rect 1438 501 1494 503
rect 1438 449 1440 501
rect 1440 449 1492 501
rect 1492 449 1494 501
rect 1438 447 1494 449
rect 1438 283 1494 285
rect 1438 231 1440 283
rect 1440 231 1492 283
rect 1492 231 1494 283
rect 1438 229 1494 231
rect 1704 486 1760 488
rect 1704 434 1706 486
rect 1706 434 1758 486
rect 1758 434 1760 486
rect 1704 432 1760 434
rect 1704 248 1706 270
rect 1706 248 1758 270
rect 1758 248 1760 270
rect 1704 214 1760 248
rect 2152 486 2208 488
rect 2152 434 2154 486
rect 2154 434 2206 486
rect 2206 434 2208 486
rect 2152 432 2208 434
rect 2152 248 2154 270
rect 2154 248 2206 270
rect 2206 248 2208 270
rect 2152 214 2208 248
rect 2464 486 2520 488
rect 2464 434 2466 486
rect 2466 434 2518 486
rect 2518 434 2520 486
rect 2464 432 2520 434
rect 2464 248 2466 270
rect 2466 248 2518 270
rect 2518 248 2520 270
rect 2464 214 2520 248
rect 2912 486 2968 488
rect 2912 434 2914 486
rect 2914 434 2966 486
rect 2966 434 2968 486
rect 2912 432 2968 434
rect 2912 248 2914 270
rect 2914 248 2966 270
rect 2966 248 2968 270
rect 2912 214 2968 248
rect 3373 501 3429 503
rect 3373 449 3375 501
rect 3375 449 3427 501
rect 3427 449 3429 501
rect 3373 447 3429 449
rect 3373 283 3429 285
rect 3373 231 3375 283
rect 3375 231 3427 283
rect 3427 231 3429 283
rect 3373 229 3429 231
rect 3683 501 3739 503
rect 3683 449 3685 501
rect 3685 449 3737 501
rect 3737 449 3739 501
rect 3683 447 3739 449
rect 3683 283 3739 285
rect 3683 231 3685 283
rect 3685 231 3737 283
rect 3737 231 3739 283
rect 3683 229 3739 231
<< metal3 >>
rect -65 2818 4862 2866
rect -65 2786 3257 2818
rect -65 2730 -28 2786
rect 28 2775 3257 2786
rect 28 2730 273 2775
rect -65 2719 273 2730
rect 329 2719 945 2775
rect 1001 2719 2361 2775
rect 2417 2719 2809 2775
rect 2865 2762 3257 2775
rect 3313 2762 3705 2818
rect 3761 2786 4862 2818
rect 3761 2762 4678 2786
rect 2865 2730 4678 2762
rect 4734 2730 4862 2786
rect 2865 2719 4862 2730
rect -65 2600 4862 2719
rect -65 2568 3257 2600
rect -65 2512 -28 2568
rect 28 2557 3257 2568
rect 28 2512 273 2557
rect -65 2501 273 2512
rect 329 2501 945 2557
rect 1001 2501 2361 2557
rect 2417 2501 2809 2557
rect 2865 2544 3257 2557
rect 3313 2544 3705 2600
rect 3761 2568 4862 2600
rect 3761 2544 4678 2568
rect 2865 2512 4678 2544
rect 4734 2512 4862 2568
rect 2865 2501 4862 2512
rect -65 2411 4862 2501
rect -65 2084 4946 2123
rect -65 2028 -28 2084
rect 28 2028 273 2084
rect 329 2083 4601 2084
rect 329 2028 721 2083
rect -65 2027 721 2028
rect 777 2027 945 2083
rect 1001 2027 2361 2083
rect 2417 2027 2809 2083
rect 2865 2027 3705 2083
rect 3761 2028 4601 2083
rect 4657 2028 4853 2084
rect 4909 2028 4946 2084
rect 3761 2027 4946 2028
rect -65 1897 4946 2027
rect -65 1866 721 1897
rect -65 1810 -28 1866
rect 28 1810 273 1866
rect 329 1841 721 1866
rect 777 1841 945 1897
rect 1001 1841 2361 1897
rect 2417 1841 2809 1897
rect 2865 1841 3705 1897
rect 3761 1866 4946 1897
rect 3761 1841 4601 1866
rect 329 1810 4601 1841
rect 4657 1810 4853 1866
rect 4909 1810 4946 1866
rect -65 1772 4946 1810
rect -65 1632 4862 1648
rect -65 1576 592 1632
rect 648 1576 724 1632
rect 780 1576 4862 1632
rect -65 1560 4862 1576
rect -65 1401 4862 1411
rect -65 1345 592 1401
rect 648 1345 724 1401
rect 780 1345 4862 1401
rect -65 1335 4862 1345
rect -65 1204 65 1205
rect 1401 1204 1531 1205
rect 2119 1204 2249 1205
rect 3336 1204 3466 1205
rect -65 1166 4862 1204
rect -65 1110 -28 1166
rect 28 1165 1438 1166
rect 28 1110 273 1165
rect -65 1109 273 1110
rect 329 1109 721 1165
rect 777 1109 944 1165
rect 1000 1110 1438 1165
rect 1494 1165 2156 1166
rect 1494 1110 1704 1165
rect 1000 1109 1704 1110
rect 1760 1110 2156 1165
rect 2212 1165 3373 1166
rect 2212 1110 2464 1165
rect 1760 1109 2464 1110
rect 2520 1109 2912 1165
rect 2968 1110 3373 1165
rect 3429 1110 4862 1166
rect 2968 1109 4862 1110
rect -65 948 4862 1109
rect -65 892 -28 948
rect 28 947 1438 948
rect 28 892 273 947
rect -65 891 273 892
rect 329 891 721 947
rect 777 891 944 947
rect 1000 892 1438 947
rect 1494 947 2156 948
rect 1494 892 1704 947
rect 1000 891 1704 892
rect 1760 892 2156 947
rect 2212 947 3373 948
rect 2212 892 2464 947
rect 1760 891 2464 892
rect 2520 891 2912 947
rect 2968 892 3373 947
rect 3429 892 4862 948
rect 2968 891 4862 892
rect -65 853 4862 891
rect -65 503 4862 583
rect -65 447 -28 503
rect 28 492 1438 503
rect 28 447 273 492
rect -65 436 273 447
rect 329 488 1438 492
rect 329 436 944 488
rect -65 432 944 436
rect 1000 447 1438 488
rect 1494 488 3373 503
rect 1494 447 1704 488
rect 1000 432 1704 447
rect 1760 432 2152 488
rect 2208 432 2464 488
rect 2520 432 2912 488
rect 2968 447 3373 488
rect 3429 447 3683 503
rect 3739 447 4862 503
rect 2968 432 4862 447
rect -65 285 4862 432
rect -65 229 -28 285
rect 28 274 1438 285
rect 28 229 273 274
rect -65 218 273 229
rect 329 270 1438 274
rect 329 218 944 270
rect -65 214 944 218
rect 1000 229 1438 270
rect 1494 270 3373 285
rect 1494 229 1704 270
rect 1000 214 1704 229
rect 1760 214 2152 270
rect 2208 214 2464 270
rect 2520 214 2912 270
rect 2968 229 3373 270
rect 3429 229 3683 285
rect 3739 229 4862 285
rect 2968 214 4862 229
rect -65 128 4862 214
use M1_NACTIVE$$202392620_128x8m81  M1_NACTIVE$$202392620_128x8m81_0
timestamp 1669390400
transform 1 0 3401 0 1 366
box 0 0 1 1
use M1_NACTIVE$$202392620_128x8m81  M1_NACTIVE$$202392620_128x8m81_1
timestamp 1669390400
transform 1 0 1466 0 1 366
box 0 0 1 1
use M1_NACTIVE$$202392620_128x8m81  M1_NACTIVE$$202392620_128x8m81_2
timestamp 1669390400
transform 1 0 0 0 1 366
box 0 0 1 1
use M1_NACTIVE$$202392620_128x8m81  M1_NACTIVE$$202392620_128x8m81_3
timestamp 1669390400
transform 1 0 0 0 1 2649
box 0 0 1 1
use M1_NACTIVE$$202392620_128x8m81  M1_NACTIVE$$202392620_128x8m81_4
timestamp 1669390400
transform 1 0 4706 0 1 2649
box 0 0 1 1
use M1_NACTIVE4310590548738_128x8m81  M1_NACTIVE4310590548738_128x8m81_0
timestamp 1669390400
transform 1 0 3707 0 1 391
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_0
timestamp 1669390400
transform 1 0 3401 0 1 1024
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_1
timestamp 1669390400
transform 1 0 3 0 1 1024
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_2
timestamp 1669390400
transform 1 0 1464 0 1 1024
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_3
timestamp 1669390400
transform 1 0 2186 0 1 1024
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_4
timestamp 1669390400
transform 1 0 3 0 1 1951
box 0 0 1 1
use M1_PACTIVE4310590548728_128x8m81  M1_PACTIVE4310590548728_128x8m81_5
timestamp 1669390400
transform 1 0 4884 0 1 1951
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_0
timestamp 1669390400
transform 1 0 2496 0 1 748
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_1
timestamp 1669390400
transform 0 -1 1845 1 0 1365
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_2
timestamp 1669390400
transform 1 0 384 0 1 18
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_3
timestamp 1669390400
transform 1 0 666 0 1 1374
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_4
timestamp 1669390400
transform 1 0 936 0 1 748
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_5
timestamp 1669390400
transform 1 0 666 0 1 1605
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_6
timestamp 1669390400
transform 1 0 384 0 1 2975
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1669390400
transform 0 -1 863 1 0 2281
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1669390400
transform 1 0 1281 0 1 2262
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1669390400
transform 0 -1 3288 1 0 2279
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_3
timestamp 1669390400
transform 0 -1 2979 1 0 1669
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_4
timestamp 1669390400
transform 0 -1 3572 1 0 1593
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_5
timestamp 1669390400
transform 0 -1 2473 1 0 2281
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_6
timestamp 1669390400
transform 0 -1 2360 1 0 1669
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_0
timestamp 1669390400
transform 1 0 2940 0 1 367
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_1
timestamp 1669390400
transform 1 0 2492 0 1 1044
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_2
timestamp 1669390400
transform 1 0 2492 0 1 367
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_3
timestamp 1669390400
transform 1 0 2940 0 1 1044
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_4
timestamp 1669390400
transform 1 0 749 0 1 1044
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_5
timestamp 1669390400
transform 1 0 972 0 1 1044
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_6
timestamp 1669390400
transform 1 0 972 0 1 367
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_7
timestamp 1669390400
transform 1 0 1732 0 1 367
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_8
timestamp 1669390400
transform 1 0 1732 0 1 1044
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_9
timestamp 1669390400
transform 1 0 2180 0 1 367
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_10
timestamp 1669390400
transform 1 0 749 0 1 1962
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_11
timestamp 1669390400
transform 1 0 973 0 1 1962
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_12
timestamp 1669390400
transform 1 0 2837 0 1 1962
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_13
timestamp 1669390400
transform 1 0 3733 0 1 1962
box 0 0 1 1
use M2_M1$$202395692_128x8m81  M2_M1$$202395692_128x8m81_14
timestamp 1669390400
transform 1 0 2389 0 1 1962
box 0 0 1 1
use M2_M1$$202396716_128x8m81  M2_M1$$202396716_128x8m81_0
timestamp 1669390400
transform 1 0 1480 0 1 2271
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_0
timestamp 1669390400
transform 1 0 3401 0 1 1029
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_1
timestamp 1669390400
transform 1 0 3401 0 1 366
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_2
timestamp 1669390400
transform 1 0 3711 0 1 366
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_3
timestamp 1669390400
transform 1 0 1466 0 1 1029
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_4
timestamp 1669390400
transform 1 0 2184 0 1 1029
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_5
timestamp 1669390400
transform 1 0 1466 0 1 366
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_6
timestamp 1669390400
transform 1 0 0 0 1 366
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_7
timestamp 1669390400
transform 1 0 301 0 1 355
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_8
timestamp 1669390400
transform 1 0 0 0 1 1029
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_9
timestamp 1669390400
transform 1 0 301 0 1 1028
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_10
timestamp 1669390400
transform 1 0 0 0 1 2649
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_11
timestamp 1669390400
transform 1 0 301 0 1 2638
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_12
timestamp 1669390400
transform 1 0 301 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_13
timestamp 1669390400
transform 1 0 973 0 1 2638
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_14
timestamp 1669390400
transform 1 0 0 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_15
timestamp 1669390400
transform 1 0 0 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_16
timestamp 1669390400
transform 1 0 3733 0 1 2681
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_17
timestamp 1669390400
transform 1 0 3285 0 1 2681
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_18
timestamp 1669390400
transform 1 0 2837 0 1 2638
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_19
timestamp 1669390400
transform 1 0 4181 0 1 2638
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_20
timestamp 1669390400
transform 1 0 4629 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_21
timestamp 1669390400
transform 1 0 4706 0 1 2649
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_22
timestamp 1669390400
transform 1 0 4881 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_23
timestamp 1669390400
transform 1 0 4881 0 1 1947
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_24
timestamp 1669390400
transform 1 0 4181 0 1 1904
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_25
timestamp 1669390400
transform 1 0 2389 0 1 2638
box 0 0 1 1
use M2_M14310590548736_128x8m81  M2_M14310590548736_128x8m81_0
timestamp 1669390400
transform 1 0 686 0 1 1373
box 0 0 1 1
use M2_M14310590548736_128x8m81  M2_M14310590548736_128x8m81_1
timestamp 1669390400
transform 1 0 686 0 1 1604
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_0
timestamp 1669390400
transform 1 0 2940 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_1
timestamp 1669390400
transform 1 0 2940 0 1 351
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_2
timestamp 1669390400
transform 1 0 3711 0 1 366
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_3
timestamp 1669390400
transform 1 0 3401 0 1 366
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_4
timestamp 1669390400
transform 1 0 2492 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_5
timestamp 1669390400
transform 1 0 2492 0 1 351
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_6
timestamp 1669390400
transform 1 0 3401 0 1 1029
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_7
timestamp 1669390400
transform 1 0 1466 0 1 366
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_8
timestamp 1669390400
transform 1 0 2184 0 1 1029
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_9
timestamp 1669390400
transform 1 0 1466 0 1 1029
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_10
timestamp 1669390400
transform 1 0 0 0 1 366
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_11
timestamp 1669390400
transform 1 0 301 0 1 355
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_12
timestamp 1669390400
transform 1 0 0 0 1 1029
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_13
timestamp 1669390400
transform 1 0 972 0 1 351
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_14
timestamp 1669390400
transform 1 0 1732 0 1 351
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_15
timestamp 1669390400
transform 1 0 1732 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_16
timestamp 1669390400
transform 1 0 2180 0 1 351
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_17
timestamp 1669390400
transform 1 0 749 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_18
timestamp 1669390400
transform 1 0 972 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_19
timestamp 1669390400
transform 1 0 301 0 1 1028
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_20
timestamp 1669390400
transform 1 0 973 0 1 2638
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_21
timestamp 1669390400
transform 1 0 0 0 1 2649
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_22
timestamp 1669390400
transform 1 0 0 0 1 1947
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_23
timestamp 1669390400
transform 1 0 301 0 1 2638
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_24
timestamp 1669390400
transform 1 0 301 0 1 1947
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_25
timestamp 1669390400
transform 1 0 4881 0 1 1947
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_26
timestamp 1669390400
transform 1 0 3733 0 1 2681
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_27
timestamp 1669390400
transform 1 0 3285 0 1 2681
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_28
timestamp 1669390400
transform 1 0 2837 0 1 2638
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_29
timestamp 1669390400
transform 1 0 4629 0 1 1947
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_30
timestamp 1669390400
transform 1 0 4706 0 1 2649
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_31
timestamp 1669390400
transform 1 0 2389 0 1 2638
box 0 0 1 1
use M3_M2$$202397740_128x8m81  M3_M2$$202397740_128x8m81_0
timestamp 1669390400
transform 1 0 749 0 1 1962
box 0 0 1 1
use M3_M2$$202397740_128x8m81  M3_M2$$202397740_128x8m81_1
timestamp 1669390400
transform 1 0 973 0 1 1962
box 0 0 1 1
use M3_M2$$202397740_128x8m81  M3_M2$$202397740_128x8m81_2
timestamp 1669390400
transform 1 0 3733 0 1 1962
box 0 0 1 1
use M3_M2$$202397740_128x8m81  M3_M2$$202397740_128x8m81_3
timestamp 1669390400
transform 1 0 2837 0 1 1962
box 0 0 1 1
use M3_M2$$202397740_128x8m81  M3_M2$$202397740_128x8m81_4
timestamp 1669390400
transform 1 0 2389 0 1 1962
box 0 0 1 1
use M3_M24310590548737_128x8m81  M3_M24310590548737_128x8m81_0
timestamp 1669390400
transform 1 0 686 0 1 1373
box 0 0 1 1
use M3_M24310590548737_128x8m81  M3_M24310590548737_128x8m81_1
timestamp 1669390400
transform 1 0 686 0 1 1604
box 0 0 1 1
use nmos_1p2$$202594348_128x8m81  nmos_1p2$$202594348_128x8m81_0
timestamp 1669390400
transform 1 0 3593 0 1 1858
box -119 -73 177 346
use nmos_1p2$$202595372_128x8m81  nmos_1p2$$202595372_128x8m81_0
timestamp 1669390400
transform 1 0 2025 0 1 1940
box -119 -73 177 264
use nmos_1p2$$202595372_128x8m81  nmos_1p2$$202595372_128x8m81_1
timestamp 1669390400
transform 1 0 2697 0 1 1940
box -119 -73 177 264
use nmos_1p2$$202596396_128x8m81  nmos_1p2$$202596396_128x8m81_0
timestamp 1669390400
transform 1 0 2921 0 1 1940
box -119 -73 177 264
use nmos_1p2$$202596396_128x8m81  nmos_1p2$$202596396_128x8m81_1
timestamp 1669390400
transform 1 0 2249 0 1 1940
box -119 -73 177 264
use nmos_1p2$$202598444_128x8m81  nmos_1p2$$202598444_128x8m81_0
timestamp 1669390400
transform 1 0 1563 0 1 1677
box -119 -74 177 527
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_0
timestamp 1669390400
transform 1 0 577 0 -1 1204
box -88 -44 208 236
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_1
timestamp 1669390400
transform 1 0 1025 0 -1 1122
box -88 -44 208 236
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_2
timestamp 1669390400
transform 1 0 353 0 -1 1204
box -88 -44 208 236
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_3
timestamp 1669390400
transform 1 0 1025 0 1 1863
box -88 -44 208 236
use nmos_5p04310590548710_128x8m81  nmos_5p04310590548710_128x8m81_0
timestamp 1669390400
transform 1 0 4458 0 1 1677
box -88 -44 208 498
use nmos_5p04310590548739_128x8m81  nmos_5p04310590548739_128x8m81_0
timestamp 1669390400
transform 1 0 4010 0 1 1677
box -88 -44 432 498
use nmos_5p04310590548740_128x8m81  nmos_5p04310590548740_128x8m81_0
timestamp 1669390400
transform 1 0 1784 0 -1 1122
box -88 -44 208 318
use nmos_5p04310590548740_128x8m81  nmos_5p04310590548740_128x8m81_1
timestamp 1669390400
transform 1 0 353 0 1 1781
box -88 -44 208 318
use nmos_5p04310590548740_128x8m81  nmos_5p04310590548740_128x8m81_2
timestamp 1669390400
transform 1 0 577 0 1 1781
box -88 -44 208 318
use nmos_5p04310590548742_128x8m81  nmos_5p04310590548742_128x8m81_0
timestamp 1669390400
transform 1 0 2544 0 -1 1122
box -88 -44 656 204
use pmos_1p2$$202583084_128x8m81  pmos_1p2$$202583084_128x8m81_0
timestamp 1669390400
transform 1 0 3369 0 1 2525
box -286 -142 568 482
use pmos_1p2$$202584108_128x8m81  pmos_1p2$$202584108_128x8m81_0
timestamp 1669390400
transform 1 0 2697 0 1 2411
box -286 -141 297 595
use pmos_1p2$$202585132_128x8m81  pmos_1p2$$202585132_128x8m81_0
timestamp 1669390400
transform 1 0 2921 0 1 2411
box -256 -141 344 595
use pmos_1p2$$202586156_128x8m81  pmos_1p2$$202586156_128x8m81_0
timestamp 1669390400
transform 1 0 2249 0 1 2411
box -286 -141 344 595
use pmos_1p2$$202587180_128x8m81  pmos_1p2$$202587180_128x8m81_0
timestamp 1669390400
transform 1 0 1563 0 1 2411
box -286 -141 344 595
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_0
timestamp 1669390400
transform 1 0 353 0 -1 574
box -208 -120 328 574
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_1
timestamp 1669390400
transform 1 0 1025 0 -1 574
box -208 -120 328 574
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_2
timestamp 1669390400
transform 1 0 577 0 -1 574
box -208 -120 328 574
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_3
timestamp 1669390400
transform 1 0 353 0 1 2411
box -208 -120 328 574
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_4
timestamp 1669390400
transform 1 0 1025 0 1 2411
box -208 -120 328 574
use pmos_5p04310590548714_128x8m81  pmos_5p04310590548714_128x8m81_5
timestamp 1669390400
transform 1 0 577 0 1 2411
box -208 -120 328 574
use pmos_5p04310590548720_128x8m81  pmos_5p04310590548720_128x8m81_0
timestamp 1669390400
transform 1 0 4010 0 1 2411
box -208 -120 552 574
use pmos_5p04310590548735_128x8m81  pmos_5p04310590548735_128x8m81_0
timestamp 1669390400
transform 1 0 1784 0 -1 574
box -208 -120 552 462
use pmos_5p04310590548741_128x8m81  pmos_5p04310590548741_128x8m81_0
timestamp 1669390400
transform 1 0 1879 0 1 2411
box -208 -120 328 312
use pmos_5p04310590548743_128x8m81  pmos_5p04310590548743_128x8m81_0
timestamp 1669390400
transform 1 0 2544 0 -1 574
box -208 -120 776 520
<< labels >>
rlabel metal3 s 136 1062 136 1062 4 vss
port 1 nsew
rlabel metal3 s 649 1366 649 1366 4 GWEN
port 2 nsew
rlabel metal3 s 136 1947 136 1947 4 vss
port 1 nsew
rlabel metal3 s 136 2638 136 2638 4 vdd
port 3 nsew
rlabel metal3 s 649 1597 649 1597 4 VSS
port 4 nsew
rlabel metal3 s 136 430 136 430 4 vdd
port 3 nsew
rlabel metal1 s 356 3089 356 3089 4 men
port 5 nsew
rlabel metal1 s 3165 800 3165 800 4 wep
port 6 nsew
rlabel metal1 s 356 30 356 30 4 wen
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 4862 3287
string GDS_END 427552
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 412762
string path 15.820 2.690 15.820 4.995 
<< end >>
