magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 1141 7525 1771 7858
rect 311 6743 1771 7525
rect 1141 5102 1771 6743
rect 1978 1577 2607 1593
rect 298 1370 2607 1577
rect -223 580 2607 1370
rect 297 579 1152 580
rect 1977 579 2607 580
rect 298 498 1152 579
rect 1978 -51 2607 579
<< nmos >>
rect 720 7664 840 7892
<< pmos >>
rect 605 7088 725 7385
rect 878 7088 998 7385
<< ndiff >>
rect 581 7779 720 7892
rect 581 7733 625 7779
rect 671 7733 720 7779
rect 581 7664 720 7733
rect 840 7779 978 7892
rect 840 7733 888 7779
rect 934 7733 978 7779
rect 840 7664 978 7733
<< pdiff >>
rect 487 7260 605 7385
rect 487 7214 530 7260
rect 576 7214 605 7260
rect 487 7088 605 7214
rect 725 7260 878 7385
rect 725 7214 794 7260
rect 840 7214 878 7260
rect 725 7088 878 7214
rect 998 7260 1116 7385
rect 998 7214 1027 7260
rect 1073 7214 1116 7260
rect 998 7088 1116 7214
<< ndiffc >>
rect 625 7733 671 7779
rect 888 7733 934 7779
<< pdiffc >>
rect 530 7214 576 7260
rect 794 7214 840 7260
rect 1027 7214 1073 7260
<< psubdiff >>
rect -80 1714 80 1774
rect -80 1668 -23 1714
rect 23 1668 80 1714
rect -80 1608 80 1668
rect -9 319 75 338
rect -9 179 10 319
rect 56 179 75 319
rect -9 160 75 179
<< nsubdiff >>
rect 1323 7750 1595 7769
rect 1323 7704 1342 7750
rect 1576 7704 1595 7750
rect 1323 7685 1595 7704
rect -78 1166 78 1223
rect -78 1120 -23 1166
rect 23 1120 78 1166
rect -78 1002 78 1120
rect -78 956 -23 1002
rect 23 956 78 1002
rect -78 899 78 956
<< psubdiffcont >>
rect -23 1668 23 1714
rect 10 179 56 319
<< nsubdiffcont >>
rect 1342 7704 1576 7750
rect -23 1120 23 1166
rect -23 956 23 1002
<< polysilicon >>
rect 720 7892 840 7965
rect 720 7602 840 7664
rect 593 7595 840 7602
rect 593 7556 998 7595
rect 593 7510 667 7556
rect 713 7510 998 7556
rect 593 7465 998 7510
rect 605 7455 998 7465
rect 605 7385 725 7455
rect 878 7385 998 7455
rect 605 7016 725 7088
rect 878 7016 998 7088
rect 711 6890 905 6936
rect 711 6844 785 6890
rect 831 6844 905 6890
rect 711 6726 905 6844
rect 500 6666 1068 6726
rect 52 4735 172 5340
rect 1396 5093 1516 5340
rect 1251 5092 1516 5093
rect 1120 5047 1516 5092
rect 1120 5001 1193 5047
rect 1239 5001 1516 5047
rect 1120 4956 1516 5001
rect 1251 4955 1516 4956
rect 1396 4735 1516 4955
rect 500 2453 1068 2479
rect 500 2407 653 2453
rect 699 2407 1068 2453
rect 500 2388 1068 2407
rect 1381 2240 1501 2259
rect 1381 2194 1418 2240
rect 1464 2194 1501 2240
rect 1381 2099 1501 2194
rect 16 1968 208 2013
rect 16 1922 89 1968
rect 135 1922 208 1968
rect 16 1877 208 1922
rect 1381 1824 1501 1983
rect 663 1549 783 1807
rect 1381 1764 1725 1824
rect 1381 1658 1501 1764
rect 1605 1658 1725 1764
rect 553 1495 897 1549
rect 553 1488 673 1495
rect 777 1488 897 1495
rect 2233 1452 2353 1731
rect 1048 1215 1240 1260
rect 1048 1169 1121 1215
rect 1167 1184 1240 1215
rect 1167 1169 1725 1184
rect 553 1120 673 1169
rect 1048 1124 1725 1169
rect 1604 1123 1725 1124
rect 479 1075 673 1120
rect 479 1029 552 1075
rect 598 1044 673 1075
rect 598 1029 1501 1044
rect 479 984 1501 1029
rect 553 983 1501 984
rect 1605 942 1725 1123
rect 276 529 470 568
rect 553 529 673 639
rect 777 567 897 639
rect 1381 568 1501 683
rect 276 522 673 529
rect 276 476 350 522
rect 396 476 673 522
rect 276 469 673 476
rect 276 431 470 469
rect 288 430 470 431
rect 553 362 673 469
rect 721 522 913 567
rect 721 476 794 522
rect 840 476 913 522
rect 1381 507 1725 568
rect 721 431 913 476
rect 1102 457 1186 466
rect 1102 447 1501 457
rect 777 360 897 431
rect 1102 401 1121 447
rect 1167 401 1501 447
rect 1102 397 1501 401
rect 1102 382 1186 397
rect 1381 366 1501 397
rect 1605 336 1725 507
rect 2233 8 2353 90
rect 2233 -38 2270 8
rect 2316 -38 2353 8
rect 2233 -57 2353 -38
<< polycontact >>
rect 667 7510 713 7556
rect 785 6844 831 6890
rect 1193 5001 1239 5047
rect 653 2407 699 2453
rect 1418 2194 1464 2240
rect 89 1922 135 1968
rect 1121 1169 1167 1215
rect 552 1029 598 1075
rect 350 476 396 522
rect 794 476 840 522
rect 1121 401 1167 447
rect 2270 -38 2316 8
<< metal1 >>
rect 355 8811 2067 8836
rect 355 8759 405 8811
rect 457 8759 591 8811
rect 643 8759 1422 8811
rect 1474 8759 1608 8811
rect 1660 8759 2067 8811
rect 355 8739 2067 8759
rect 355 8623 2067 8627
rect 355 8603 2301 8623
rect 355 8551 785 8603
rect 837 8551 971 8603
rect 1023 8551 2023 8603
rect 2075 8551 2209 8603
rect 2261 8551 2301 8603
rect 355 8531 2301 8551
rect 355 8530 2067 8531
rect 606 8418 735 8419
rect 45 8378 2067 8418
rect 45 8326 644 8378
rect 696 8326 2067 8378
rect 45 8281 2067 8326
rect 164 8068 1580 8164
rect 590 7969 1090 7970
rect 590 7929 1168 7969
rect 590 7895 1096 7929
rect 590 7779 686 7895
rect 1076 7877 1096 7895
rect 1148 7877 1168 7929
rect 590 7733 625 7779
rect 671 7733 686 7779
rect 590 7673 686 7733
rect 803 7779 969 7815
rect 803 7733 888 7779
rect 934 7733 969 7779
rect 803 7696 969 7733
rect 1076 7743 1168 7877
rect 467 7556 725 7593
rect 467 7553 667 7556
rect 467 7501 644 7553
rect 713 7510 725 7556
rect 696 7501 725 7510
rect 467 7460 725 7501
rect 803 7376 875 7696
rect 1076 7691 1096 7743
rect 1148 7691 1168 7743
rect 1331 7750 1587 7761
rect 1331 7704 1342 7750
rect 1576 7729 1587 7750
rect 1576 7704 1591 7729
rect 1331 7693 1591 7704
rect 1076 7650 1168 7691
rect 1545 7468 1591 7693
rect 495 7260 592 7364
rect 495 7214 530 7260
rect 576 7214 592 7260
rect 495 7097 592 7214
rect 759 7260 875 7376
rect 759 7214 794 7260
rect 840 7214 875 7260
rect 759 7097 875 7214
rect 519 6750 592 7097
rect 803 6904 875 7097
rect 751 6890 875 6904
rect 751 6844 785 6890
rect 831 6844 875 6890
rect 751 6830 875 6844
rect 992 7260 1108 7376
rect 992 7214 1027 7260
rect 1073 7214 1108 7260
rect 992 7097 1108 7214
rect 992 6750 1064 7097
rect 519 6676 1064 6750
rect 397 6546 489 6586
rect 397 6494 417 6546
rect 469 6494 489 6546
rect 397 6360 489 6494
rect 397 6308 417 6360
rect 469 6308 489 6360
rect 397 6267 489 6308
rect 850 6546 942 6586
rect 850 6494 870 6546
rect 922 6494 942 6546
rect 850 6360 942 6494
rect 850 6308 870 6360
rect 922 6308 942 6360
rect 850 6267 942 6308
rect 166 5084 282 5519
rect 614 5084 730 5519
rect 1330 5372 1402 5519
rect 1062 5252 1402 5372
rect 166 5047 1253 5084
rect 166 5001 1193 5047
rect 1239 5001 1253 5047
rect 166 4964 1253 5001
rect 166 4708 282 4964
rect 400 4755 492 4795
rect 400 4703 420 4755
rect 472 4703 492 4755
rect 614 4708 730 4964
rect 1330 4798 1402 5252
rect 1995 4809 2155 7747
rect 850 4755 942 4795
rect 400 4569 492 4703
rect 400 4517 420 4569
rect 472 4517 492 4569
rect 400 4476 492 4517
rect 850 4703 870 4755
rect 922 4703 942 4755
rect 850 4569 942 4703
rect 1062 4678 1402 4798
rect 850 4517 870 4569
rect 922 4517 942 4569
rect 850 4476 942 4517
rect 1510 2597 2155 4809
rect 618 2453 906 2467
rect 618 2407 653 2453
rect 699 2443 906 2453
rect 618 2391 655 2407
rect 707 2391 906 2443
rect 618 2371 906 2391
rect 359 2240 2204 2291
rect 359 2194 1418 2240
rect 1464 2194 2204 2240
rect 359 2171 2204 2194
rect 359 1985 475 2171
rect 54 1968 475 1985
rect 54 1922 89 1968
rect 135 1922 475 1968
rect 54 1865 475 1922
rect -71 1754 71 1765
rect -71 1714 275 1754
rect -71 1713 -23 1714
rect 23 1713 275 1714
rect -71 1661 -27 1713
rect 25 1661 185 1713
rect 237 1661 275 1713
rect -71 1620 275 1661
rect -71 1617 71 1620
rect 825 1608 897 1991
rect 695 1534 1180 1608
rect 695 1217 767 1534
rect 1108 1215 1180 1534
rect -58 1166 58 1203
rect -58 1120 -23 1166
rect 23 1120 58 1166
rect -58 1002 58 1120
rect 1108 1169 1121 1215
rect 1167 1169 1180 1215
rect 1270 1183 1386 1427
rect 1286 1182 1380 1183
rect -58 956 -23 1002
rect 23 956 58 1002
rect 227 1075 633 1094
rect 227 1029 552 1075
rect 598 1029 633 1075
rect 227 985 633 1029
rect -58 920 58 956
rect -47 919 47 920
rect 194 522 409 559
rect 194 476 350 522
rect 396 476 409 522
rect 194 439 409 476
rect 487 536 559 715
rect 487 522 874 536
rect 487 476 794 522
rect 840 476 874 522
rect 487 462 874 476
rect -1 319 67 330
rect -1 179 10 319
rect 56 179 67 319
rect 487 246 559 462
rect 694 291 787 331
rect 694 239 714 291
rect 766 239 787 291
rect 694 199 787 239
rect 694 198 783 199
rect -1 89 67 179
rect 700 89 772 198
rect -1 15 772 89
rect 952 89 1024 831
rect 1108 447 1180 1169
rect 1494 1103 1610 1944
rect 1720 1461 1812 1502
rect 1720 1427 1740 1461
rect 1718 1409 1740 1427
rect 1792 1427 1812 1461
rect 1792 1409 1834 1427
rect 1718 1275 1834 1409
rect 1718 1223 1740 1275
rect 1792 1223 1834 1275
rect 2158 1248 2204 2171
rect 2409 1849 2465 2158
rect 1718 1183 1834 1223
rect 1494 983 1834 1103
rect 1108 401 1121 447
rect 1167 401 1180 447
rect 1108 390 1180 401
rect 1306 89 1352 808
rect 952 15 1352 89
rect 1530 19 1576 794
rect 1718 145 1834 983
rect 1530 8 2327 19
rect 1530 -38 2270 8
rect 2316 -38 2327 8
rect 1530 -55 2327 -38
<< via1 >>
rect 405 8759 457 8811
rect 591 8759 643 8811
rect 1422 8759 1474 8811
rect 1608 8759 1660 8811
rect 785 8551 837 8603
rect 971 8551 1023 8603
rect 2023 8551 2075 8603
rect 2209 8551 2261 8603
rect 644 8326 696 8378
rect 1096 7877 1148 7929
rect 644 7510 667 7553
rect 667 7510 696 7553
rect 644 7501 696 7510
rect 1096 7691 1148 7743
rect 417 6494 469 6546
rect 417 6308 469 6360
rect 870 6494 922 6546
rect 870 6308 922 6360
rect 420 4703 472 4755
rect 420 4517 472 4569
rect 870 4703 922 4755
rect 870 4517 922 4569
rect 655 2407 699 2443
rect 699 2407 707 2443
rect 655 2391 707 2407
rect -27 1668 -23 1713
rect -23 1668 23 1713
rect 23 1668 25 1713
rect -27 1661 25 1668
rect 185 1661 237 1713
rect 714 239 766 291
rect 1740 1409 1792 1461
rect 1740 1223 1792 1275
<< metal2 >>
rect 1191 8997 1286 8999
rect 396 8831 491 8836
rect 375 8811 683 8831
rect 375 8759 405 8811
rect 457 8759 591 8811
rect 643 8759 683 8811
rect 375 8739 683 8759
rect 396 6546 491 8739
rect 884 8627 974 8949
rect 849 8623 974 8627
rect 755 8603 1063 8623
rect 755 8551 785 8603
rect 837 8551 971 8603
rect 1023 8551 1063 8603
rect 755 8531 1063 8551
rect 849 8530 974 8531
rect 605 8380 735 8419
rect 605 8324 642 8380
rect 698 8324 735 8380
rect 605 8285 735 8324
rect 396 6494 417 6546
rect 469 6494 491 6546
rect 396 6360 491 6494
rect 396 6308 417 6360
rect 469 6308 491 6360
rect 396 4795 491 6308
rect 623 7553 717 8285
rect 623 7501 644 7553
rect 696 7501 717 7553
rect 396 4755 492 4795
rect 396 4703 420 4755
rect 472 4703 492 4755
rect 396 4569 492 4703
rect 396 4517 420 4569
rect 472 4517 492 4569
rect 396 4477 492 4517
rect 623 2464 717 7501
rect 849 6546 943 8530
rect 1191 7970 1285 8997
rect 1503 8831 1593 8949
rect 1392 8811 1700 8831
rect 1392 8759 1422 8811
rect 1474 8759 1608 8811
rect 1660 8759 1700 8811
rect 1392 8739 1700 8759
rect 2123 8623 2212 8949
rect 1993 8603 2301 8623
rect 1993 8551 2023 8603
rect 2075 8551 2209 8603
rect 2261 8551 2301 8603
rect 1993 8531 2301 8551
rect 2123 8530 2212 8531
rect 1075 7929 1285 7970
rect 1075 7877 1096 7929
rect 1148 7877 1285 7929
rect 1075 7873 1285 7877
rect 1075 7743 1169 7873
rect 1075 7691 1096 7743
rect 1148 7691 1169 7743
rect 1075 7650 1169 7691
rect 849 6494 870 6546
rect 922 6494 943 6546
rect 849 6360 943 6494
rect 849 6308 870 6360
rect 922 6308 943 6360
rect 849 4755 943 6308
rect 849 4703 870 4755
rect 922 4703 943 4755
rect 849 4569 943 4703
rect 849 4517 870 4569
rect 922 4517 943 4569
rect 849 4477 943 4517
rect 620 2443 747 2464
rect 620 2391 655 2443
rect 707 2391 747 2443
rect 620 2371 747 2391
rect 1097 1890 1191 1928
rect 1097 1834 1116 1890
rect 1172 1834 1191 1890
rect -65 1715 275 1754
rect -65 1659 -29 1715
rect 27 1659 183 1715
rect 239 1659 275 1715
rect -65 1620 275 1659
rect 1097 1704 1191 1834
rect 1097 1648 1116 1704
rect 1172 1648 1191 1704
rect 694 316 787 331
rect 1097 316 1191 1648
rect 1720 1461 1812 1501
rect 1720 1409 1740 1461
rect 1792 1409 1812 1461
rect 1720 1316 1812 1409
rect 1719 1277 1812 1316
rect 1719 1221 1738 1277
rect 1794 1221 1812 1277
rect 1719 1091 1812 1221
rect 1719 1035 1738 1091
rect 1794 1035 1812 1091
rect 1719 997 1812 1035
rect 693 291 1191 316
rect 693 239 714 291
rect 766 239 1191 291
rect 693 219 1191 239
rect 694 199 787 219
<< via2 >>
rect 642 8378 698 8380
rect 642 8326 644 8378
rect 644 8326 696 8378
rect 696 8326 698 8378
rect 642 8324 698 8326
rect 1116 1834 1172 1890
rect -29 1713 27 1715
rect -29 1661 -27 1713
rect -27 1661 25 1713
rect 25 1661 27 1713
rect -29 1659 27 1661
rect 183 1713 239 1715
rect 183 1661 185 1713
rect 185 1661 237 1713
rect 237 1661 239 1713
rect 183 1659 239 1661
rect 1116 1648 1172 1704
rect 1738 1275 1794 1277
rect 1738 1223 1740 1275
rect 1740 1223 1792 1275
rect 1792 1223 1794 1275
rect 1738 1221 1794 1223
rect 1738 1035 1794 1091
<< metal3 >>
rect 605 8380 735 8419
rect 605 8324 642 8380
rect 698 8324 735 8380
rect 605 8285 735 8324
rect -47 5186 2456 7908
rect -47 1890 2456 4900
rect -47 1834 1116 1890
rect 1172 1834 2456 1890
rect -47 1754 2456 1834
rect -65 1715 2456 1754
rect -65 1659 -29 1715
rect 27 1659 183 1715
rect 239 1704 2456 1715
rect 239 1659 1116 1704
rect -65 1648 1116 1659
rect 1172 1648 2456 1704
rect -65 1620 2456 1648
rect -47 1498 2456 1620
rect -47 1277 2456 1348
rect -47 1221 1738 1277
rect 1794 1221 2456 1277
rect -47 1091 2456 1221
rect -47 1035 1738 1091
rect 1794 1035 2456 1091
rect -47 631 2456 1035
use M1_NWELL08_512x8m81  M1_NWELL08_512x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 1061
box 0 0 1 1
use M1_NWELL4310591302032_512x8m81  M1_NWELL4310591302032_512x8m81_0
timestamp 1669390400
transform 1 0 1459 0 1 7727
box 0 0 1 1
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_0
timestamp 1669390400
transform 1 0 33 0 1 249
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1669390400
transform 1 0 676 0 1 2430
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1669390400
transform 1 0 1144 0 1 424
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1669390400
transform 1 0 2293 0 1 -15
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1669390400
transform 1 0 1441 0 1 2217
box 0 0 1 1
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 1691
box 0 0 1 1
use M1_PSUB$$46892076_512x8m81  M1_PSUB$$46892076_512x8m81_0
timestamp 1669390400
transform 1 0 2066 0 1 5225
box -80 -2530 80 2531
use M1_PSUB$$46893100_512x8m81  M1_PSUB$$46893100_512x8m81_0
timestamp 1669390400
transform 1 0 1908 0 1 3756
box -80 -1061 80 1062
use M2_M1$$43375660_R90_512x8m81  M2_M1$$43375660_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 105 1 0 1687
box 0 0 1 1
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1669390400
transform 1 0 670 0 1 8352
box 0 0 1 1
use M3_M2$$43368492_R90_512x8m81  M3_M2$$43368492_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 105 1 0 1687
box 0 0 1 1
use M3_M2$$46895148_512x8m81  M3_M2$$46895148_512x8m81_0
timestamp 1669390400
transform 1 0 670 0 1 8352
box 0 0 1 1
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_0
timestamp 1669390400
transform 1 0 1412 0 -1 2099
box -119 -74 177 264
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_1
timestamp 1669390400
transform 1 0 694 0 1 1807
box -119 -74 177 264
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_0
timestamp 1669390400
transform 1 0 979 0 1 2539
box -119 -73 177 2341
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_1
timestamp 1669390400
transform 1 0 1427 0 1 2539
box -119 -73 177 2341
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_2
timestamp 1669390400
transform 1 0 531 0 1 2539
box -119 -73 177 2341
use nmos_1p2$$46884908_512x8m81  nmos_1p2$$46884908_512x8m81_0
timestamp 1669390400
transform 1 0 83 0 1 2086
box -119 -74 177 2794
use nmos_5p04310591302010_512x8m81  nmos_5p04310591302010_512x8m81_0
timestamp 1669390400
transform 1 0 2233 0 -1 2185
box -88 -44 208 498
use nmos_5p04310591302011_512x8m81  nmos_5p04310591302011_512x8m81_0
timestamp 1669390400
transform 1 0 553 0 -1 358
box -88 -44 432 236
use nmos_5p04310591302011_512x8m81  nmos_5p04310591302011_512x8m81_1
timestamp 1669390400
transform 1 0 1381 0 1 145
box -88 -44 432 236
use pmos_1p2$$46273580_512x8m81  pmos_1p2$$46273580_512x8m81_0
timestamp 1669390400
transform 1 0 584 0 -1 1435
box -286 -142 568 348
use pmos_1p2$$46273580_512x8m81  pmos_1p2$$46273580_512x8m81_1
timestamp 1669390400
transform 1 0 1412 0 -1 1628
box -286 -142 568 348
use pmos_1p2$$46885932_512x8m81  pmos_1p2$$46885932_512x8m81_0
timestamp 1669390400
transform 1 0 1412 0 1 721
box -286 -141 568 332
use pmos_1p2$$46887980_512x8m81  pmos_1p2$$46887980_512x8m81_0
timestamp 1669390400
transform 1 0 83 0 1 5244
box -286 -142 344 2862
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_0
timestamp 1669390400
transform 1 0 531 0 1 5244
box -286 -142 343 1502
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_1
timestamp 1669390400
transform 1 0 979 0 1 5244
box -286 -142 343 1502
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1669390400
transform 1 0 2233 0 1 91
box -208 -120 328 1482
use pmos_5p0431059130206_512x8m81  pmos_5p0431059130206_512x8m81_0
timestamp 1669390400
transform 1 0 553 0 1 639
box -208 -120 552 312
use pmos_5p0431059130209_512x8m81  pmos_5p0431059130209_512x8m81_0
timestamp 1669390400
transform 1 0 1396 0 1 5244
box -208 -120 328 2388
use po_m1_512x8m81  po_m1_512x8m81_0
timestamp 1669390400
transform -1 0 883 0 -1 567
box 0 0 1 1
use po_m1_512x8m81  po_m1_512x8m81_1
timestamp 1669390400
transform 1 0 742 0 -1 6935
box 0 0 1 1
use po_m1_512x8m81  po_m1_512x8m81_2
timestamp 1669390400
transform 1 0 509 0 1 984
box 0 0 1 1
use po_m1_512x8m81  po_m1_512x8m81_3
timestamp 1669390400
transform 1 0 46 0 1 1877
box 0 0 1 1
use po_m1_R90_512x8m81  po_m1_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 1282 1 0 4956
box 0 0 1 1
use po_m1_R90_512x8m81  po_m1_R90_512x8m81_1
timestamp 1669390400
transform 0 -1 1210 1 0 1124
box 0 0 1 1
use po_m1_R270_512x8m81  po_m1_R270_512x8m81_0
timestamp 1669390400
transform 0 1 307 -1 0 567
box 0 0 1 1
use po_m1_R270_512x8m81  po_m1_R270_512x8m81_1
timestamp 1669390400
transform 0 1 624 -1 0 7601
box 0 0 1 1
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1669390400
transform -1 0 808 0 -1 966
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1669390400
transform -1 0 990 0 -1 1315
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1669390400
transform -1 0 1379 0 -1 1315
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1669390400
transform 1 0 -46 0 1 3523
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1669390400
transform 1 0 1511 0 1 2607
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1669390400
transform 1 0 -46 0 1 4471
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1669390400
transform 1 0 1511 0 1 4471
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1669390400
transform 1 0 1511 0 1 3523
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1669390400
transform 1 0 -46 0 1 898
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1669390400
transform 1 0 575 0 1 1755
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1669390400
transform 1 0 2449 0 1 927
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1669390400
transform 1 0 1524 0 1 5466
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1669390400
transform 1 0 -46 0 1 5466
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1669390400
transform 1 0 1524 0 1 6957
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1669390400
transform 1 0 -46 0 1 7522
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1669390400
transform 1 0 -46 0 1 6923
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1669390400
transform 1 0 2449 0 1 1850
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1669390400
transform 1 0 1293 0 1 1755
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1669390400
transform 1 0 -46 0 1 2607
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1669390400
transform 1 0 1034 0 1 7057
box 0 -1 93 308
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 558 1 0 1220
box 0 -1 93 308
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_1
timestamp 1669390400
transform 0 -1 1612 1 0 7681
box 0 -1 93 308
use via1_512x8m81  via1_512x8m81_0
timestamp 1669390400
transform 1 0 694 0 1 199
box 0 0 1 1
use via1_512x8m81  via1_512x8m81_1
timestamp 1669390400
transform 1 0 624 0 1 7461
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 747 1 0 2371
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1669390400
transform -1 0 1812 0 -1 1501
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1669390400
transform 1 0 850 0 1 6268
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1669390400
transform 1 0 397 0 1 6268
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1669390400
transform 1 0 1076 0 1 7651
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1669390400
transform 1 0 400 0 1 4477
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1669390400
transform 1 0 850 0 1 4477
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 2301 1 0 8531
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1669390400
transform 0 -1 1700 1 0 8739
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1669390400
transform 0 -1 1063 1 0 8531
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1669390400
transform 0 -1 683 1 0 8739
box 0 0 1 1
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1669390400
transform -1 0 1812 0 -1 1315
box 0 0 1 1
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1669390400
transform 1 0 1098 0 1 1610
box 0 0 1 1
<< labels >>
rlabel metal3 s 1557 3224 1557 3224 4 vss
port 1 nsew
rlabel metal3 s 1487 5955 1487 5955 4 vdd
port 2 nsew
rlabel metal3 s 1337 918 1337 918 4 vdd
port 2 nsew
rlabel metal2 s 435 7996 435 7996 4 d
port 3 nsew
rlabel metal2 s 887 7996 887 7996 4 db
port 4 nsew
rlabel metal2 s 1228 8197 1228 8197 4 vss
port 1 nsew
rlabel metal1 s 376 508 376 508 4 datain
port 5 nsew
rlabel metal1 s 1050 8363 1050 8363 4 wep
port 6 nsew
rlabel metal1 s 571 1056 571 1056 4 men
port 7 nsew
rlabel metal1 s 1254 8798 1254 8798 4 d
port 3 nsew
rlabel metal1 s 1394 8594 1394 8594 4 db
port 4 nsew
<< properties >>
string GDS_END 435698
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 425536
<< end >>
