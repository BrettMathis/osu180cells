magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4342 1094
<< pwell >>
rect -86 -86 4342 453
<< mvnmos >>
rect 134 69 254 333
rect 358 69 478 333
rect 582 69 702 333
rect 806 69 926 333
rect 1030 69 1150 333
rect 1254 69 1374 333
rect 1478 69 1598 333
rect 1702 69 1822 333
rect 1926 69 2046 333
rect 2150 69 2270 333
rect 2374 69 2494 333
rect 2598 69 2718 333
rect 2822 69 2942 333
rect 3046 69 3166 333
rect 3270 69 3390 333
rect 3494 69 3614 333
rect 3718 69 3838 333
rect 3942 69 4062 333
<< mvpmos >>
rect 134 573 234 939
rect 358 573 458 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1254 573 1354 939
rect 1478 573 1578 939
rect 1702 573 1802 939
rect 1926 573 2026 939
rect 2150 573 2250 939
rect 2374 573 2474 939
rect 2598 573 2698 939
rect 2822 573 2922 939
rect 3046 573 3146 939
rect 3270 573 3370 939
rect 3494 573 3594 939
rect 3718 573 3818 939
rect 3942 573 4042 939
<< mvndiff >>
rect 46 287 134 333
rect 46 147 59 287
rect 105 147 134 287
rect 46 69 134 147
rect 254 287 358 333
rect 254 147 283 287
rect 329 147 358 287
rect 254 69 358 147
rect 478 287 582 333
rect 478 147 507 287
rect 553 147 582 287
rect 478 69 582 147
rect 702 287 806 333
rect 702 147 731 287
rect 777 147 806 287
rect 702 69 806 147
rect 926 287 1030 333
rect 926 147 955 287
rect 1001 147 1030 287
rect 926 69 1030 147
rect 1150 287 1254 333
rect 1150 147 1179 287
rect 1225 147 1254 287
rect 1150 69 1254 147
rect 1374 287 1478 333
rect 1374 147 1403 287
rect 1449 147 1478 287
rect 1374 69 1478 147
rect 1598 287 1702 333
rect 1598 147 1627 287
rect 1673 147 1702 287
rect 1598 69 1702 147
rect 1822 287 1926 333
rect 1822 147 1851 287
rect 1897 147 1926 287
rect 1822 69 1926 147
rect 2046 287 2150 333
rect 2046 147 2075 287
rect 2121 147 2150 287
rect 2046 69 2150 147
rect 2270 287 2374 333
rect 2270 147 2299 287
rect 2345 147 2374 287
rect 2270 69 2374 147
rect 2494 287 2598 333
rect 2494 147 2523 287
rect 2569 147 2598 287
rect 2494 69 2598 147
rect 2718 287 2822 333
rect 2718 147 2747 287
rect 2793 147 2822 287
rect 2718 69 2822 147
rect 2942 287 3046 333
rect 2942 147 2971 287
rect 3017 147 3046 287
rect 2942 69 3046 147
rect 3166 287 3270 333
rect 3166 147 3195 287
rect 3241 147 3270 287
rect 3166 69 3270 147
rect 3390 287 3494 333
rect 3390 147 3419 287
rect 3465 147 3494 287
rect 3390 69 3494 147
rect 3614 287 3718 333
rect 3614 147 3643 287
rect 3689 147 3718 287
rect 3614 69 3718 147
rect 3838 287 3942 333
rect 3838 147 3867 287
rect 3913 147 3942 287
rect 3838 69 3942 147
rect 4062 287 4150 333
rect 4062 147 4091 287
rect 4137 147 4150 287
rect 4062 69 4150 147
<< mvpdiff >>
rect 46 861 134 939
rect 46 721 59 861
rect 105 721 134 861
rect 46 573 134 721
rect 234 861 358 939
rect 234 721 283 861
rect 329 721 358 861
rect 234 573 358 721
rect 458 861 582 939
rect 458 721 487 861
rect 533 721 582 861
rect 458 573 582 721
rect 682 861 806 939
rect 682 721 711 861
rect 757 721 806 861
rect 682 573 806 721
rect 906 861 1030 939
rect 906 721 935 861
rect 981 721 1030 861
rect 906 573 1030 721
rect 1130 861 1254 939
rect 1130 721 1164 861
rect 1210 721 1254 861
rect 1130 573 1254 721
rect 1354 861 1478 939
rect 1354 721 1383 861
rect 1429 721 1478 861
rect 1354 573 1478 721
rect 1578 861 1702 939
rect 1578 721 1627 861
rect 1673 721 1702 861
rect 1578 573 1702 721
rect 1802 926 1926 939
rect 1802 786 1831 926
rect 1877 786 1926 926
rect 1802 573 1926 786
rect 2026 861 2150 939
rect 2026 721 2055 861
rect 2101 721 2150 861
rect 2026 573 2150 721
rect 2250 861 2374 939
rect 2250 721 2279 861
rect 2325 721 2374 861
rect 2250 573 2374 721
rect 2474 861 2598 939
rect 2474 721 2503 861
rect 2549 721 2598 861
rect 2474 573 2598 721
rect 2698 861 2822 939
rect 2698 721 2727 861
rect 2773 721 2822 861
rect 2698 573 2822 721
rect 2922 861 3046 939
rect 2922 721 2951 861
rect 2997 721 3046 861
rect 2922 573 3046 721
rect 3146 861 3270 939
rect 3146 721 3175 861
rect 3221 721 3270 861
rect 3146 573 3270 721
rect 3370 861 3494 939
rect 3370 721 3399 861
rect 3445 721 3494 861
rect 3370 573 3494 721
rect 3594 861 3718 939
rect 3594 721 3623 861
rect 3669 721 3718 861
rect 3594 573 3718 721
rect 3818 861 3942 939
rect 3818 721 3847 861
rect 3893 721 3942 861
rect 3818 573 3942 721
rect 4042 861 4130 939
rect 4042 721 4071 861
rect 4117 721 4130 861
rect 4042 573 4130 721
<< mvndiffc >>
rect 59 147 105 287
rect 283 147 329 287
rect 507 147 553 287
rect 731 147 777 287
rect 955 147 1001 287
rect 1179 147 1225 287
rect 1403 147 1449 287
rect 1627 147 1673 287
rect 1851 147 1897 287
rect 2075 147 2121 287
rect 2299 147 2345 287
rect 2523 147 2569 287
rect 2747 147 2793 287
rect 2971 147 3017 287
rect 3195 147 3241 287
rect 3419 147 3465 287
rect 3643 147 3689 287
rect 3867 147 3913 287
rect 4091 147 4137 287
<< mvpdiffc >>
rect 59 721 105 861
rect 283 721 329 861
rect 487 721 533 861
rect 711 721 757 861
rect 935 721 981 861
rect 1164 721 1210 861
rect 1383 721 1429 861
rect 1627 721 1673 861
rect 1831 786 1877 926
rect 2055 721 2101 861
rect 2279 721 2325 861
rect 2503 721 2549 861
rect 2727 721 2773 861
rect 2951 721 2997 861
rect 3175 721 3221 861
rect 3399 721 3445 861
rect 3623 721 3669 861
rect 3847 721 3893 861
rect 4071 721 4117 861
<< polysilicon >>
rect 134 939 234 983
rect 358 939 458 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1254 939 1354 983
rect 1478 939 1578 983
rect 1702 939 1802 983
rect 1926 939 2026 983
rect 2150 939 2250 983
rect 2374 939 2474 983
rect 2598 939 2698 983
rect 2822 939 2922 983
rect 3046 939 3146 983
rect 3270 939 3370 983
rect 3494 939 3594 983
rect 3718 939 3818 983
rect 3942 939 4042 983
rect 134 513 234 573
rect 358 513 458 573
rect 582 513 682 573
rect 806 513 906 573
rect 1030 513 1130 573
rect 1254 513 1354 573
rect 24 500 1354 513
rect 24 454 37 500
rect 1117 454 1354 500
rect 24 441 1354 454
rect 134 333 254 441
rect 358 333 478 441
rect 582 333 702 441
rect 806 333 926 441
rect 1030 439 1354 441
rect 1030 333 1150 439
rect 1254 377 1354 439
rect 1478 513 1578 573
rect 1702 513 1802 573
rect 1926 513 2026 573
rect 2150 513 2250 573
rect 2374 513 2474 573
rect 2598 513 2698 573
rect 1478 511 2698 513
rect 2822 513 2922 573
rect 3046 513 3146 573
rect 3270 513 3370 573
rect 3494 513 3594 573
rect 3718 513 3818 573
rect 3942 513 4042 573
rect 2822 511 4042 513
rect 1478 500 4042 511
rect 1478 454 1491 500
rect 2571 454 2846 500
rect 3926 454 4042 500
rect 1478 441 4042 454
rect 1254 333 1374 377
rect 1478 333 1598 441
rect 1702 333 1822 441
rect 1926 333 2046 441
rect 2150 333 2270 441
rect 2374 333 2494 441
rect 2598 333 2718 441
rect 2822 333 2942 441
rect 3046 333 3166 441
rect 3270 333 3390 441
rect 3494 333 3614 441
rect 3718 333 3838 441
rect 3942 377 4042 441
rect 3942 333 4062 377
rect 134 25 254 69
rect 358 25 478 69
rect 582 25 702 69
rect 806 25 926 69
rect 1030 25 1150 69
rect 1254 25 1374 69
rect 1478 25 1598 69
rect 1702 25 1822 69
rect 1926 25 2046 69
rect 2150 25 2270 69
rect 2374 25 2494 69
rect 2598 25 2718 69
rect 2822 25 2942 69
rect 3046 25 3166 69
rect 3270 25 3390 69
rect 3494 25 3614 69
rect 3718 25 3838 69
rect 3942 25 4062 69
<< polycontact >>
rect 37 454 1117 500
rect 1491 454 2571 500
rect 2846 454 3926 500
<< metal1 >>
rect 0 926 4256 1098
rect 0 918 1831 926
rect 59 861 105 918
rect 59 710 105 721
rect 283 861 329 872
rect 283 664 329 721
rect 487 861 533 918
rect 487 710 533 721
rect 711 861 757 872
rect 711 664 757 721
rect 935 861 981 918
rect 935 710 981 721
rect 1164 861 1245 872
rect 1210 721 1245 861
rect 1164 664 1245 721
rect 1383 861 1429 918
rect 1383 710 1429 721
rect 1627 861 1673 872
rect 1877 918 4256 926
rect 1831 775 1877 786
rect 2055 861 2101 872
rect 283 576 1245 664
rect 26 500 1128 530
rect 26 454 37 500
rect 1117 454 1128 500
rect 1179 500 1245 576
rect 1627 664 1673 721
rect 2055 664 2101 721
rect 2279 861 2325 918
rect 2279 710 2325 721
rect 2503 861 2549 872
rect 2503 664 2549 721
rect 2727 861 2773 918
rect 2727 710 2773 721
rect 2951 861 2997 872
rect 2951 664 2997 721
rect 3175 861 3221 918
rect 3175 710 3221 721
rect 3399 861 3445 872
rect 3399 664 3445 721
rect 3623 861 3669 918
rect 3623 710 3669 721
rect 3847 861 3893 872
rect 3847 664 3893 721
rect 4071 861 4117 918
rect 4071 710 4117 721
rect 1627 568 3893 664
rect 1179 454 1491 500
rect 2571 454 2582 500
rect 1179 408 1245 454
rect 2700 408 2800 568
rect 2846 500 3926 511
rect 2846 443 3926 454
rect 283 344 1245 408
rect 59 287 105 298
rect 59 90 105 147
rect 283 287 329 344
rect 283 136 329 147
rect 507 287 553 298
rect 507 90 553 147
rect 731 287 777 344
rect 731 136 777 147
rect 955 287 1001 298
rect 955 90 1001 147
rect 1179 287 1245 344
rect 1627 397 2800 408
rect 1627 351 3913 397
rect 1225 147 1245 287
rect 1179 136 1245 147
rect 1403 287 1449 298
rect 1403 90 1449 147
rect 1627 287 1673 351
rect 1627 136 1673 147
rect 1851 287 1897 298
rect 1851 90 1897 147
rect 2075 287 2121 351
rect 2075 136 2121 147
rect 2299 287 2345 298
rect 2299 90 2345 147
rect 2477 287 2569 351
rect 2477 147 2523 287
rect 2477 136 2569 147
rect 2747 287 2793 298
rect 2747 90 2793 147
rect 2971 287 3017 351
rect 2971 136 3017 147
rect 3195 287 3241 298
rect 3195 90 3241 147
rect 3419 287 3465 351
rect 3419 136 3465 147
rect 3643 287 3689 298
rect 3643 90 3689 147
rect 3867 287 3913 351
rect 3867 136 3913 147
rect 4091 287 4137 298
rect 4091 90 4137 147
rect 0 -90 4256 90
<< labels >>
flabel metal1 s 26 454 1128 530 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 4256 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 4091 90 4137 298 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3847 664 3893 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
rlabel metal1 s 3399 664 3445 872 1 Z
port 2 nsew default output
rlabel metal1 s 2951 664 2997 872 1 Z
port 2 nsew default output
rlabel metal1 s 2503 664 2549 872 1 Z
port 2 nsew default output
rlabel metal1 s 2055 664 2101 872 1 Z
port 2 nsew default output
rlabel metal1 s 1627 664 1673 872 1 Z
port 2 nsew default output
rlabel metal1 s 1627 568 3893 664 1 Z
port 2 nsew default output
rlabel metal1 s 2700 408 2800 568 1 Z
port 2 nsew default output
rlabel metal1 s 1627 397 2800 408 1 Z
port 2 nsew default output
rlabel metal1 s 1627 351 3913 397 1 Z
port 2 nsew default output
rlabel metal1 s 3867 136 3913 351 1 Z
port 2 nsew default output
rlabel metal1 s 3419 136 3465 351 1 Z
port 2 nsew default output
rlabel metal1 s 2971 136 3017 351 1 Z
port 2 nsew default output
rlabel metal1 s 2477 136 2569 351 1 Z
port 2 nsew default output
rlabel metal1 s 2075 136 2121 351 1 Z
port 2 nsew default output
rlabel metal1 s 1627 136 1673 351 1 Z
port 2 nsew default output
rlabel metal1 s 4071 775 4117 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3623 775 3669 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3175 775 3221 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2727 775 2773 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2279 775 2325 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1831 775 1877 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1383 775 1429 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 935 775 981 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 487 775 533 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 59 775 105 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4071 710 4117 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3623 710 3669 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3175 710 3221 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2727 710 2773 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2279 710 2325 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1383 710 1429 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 935 710 981 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 487 710 533 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 59 710 105 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3643 90 3689 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3195 90 3241 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2747 90 2793 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2299 90 2345 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1851 90 1897 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1403 90 1449 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 955 90 1001 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 507 90 553 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 59 90 105 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4256 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 1008
string GDS_END 1268398
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1257256
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
