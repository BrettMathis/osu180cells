magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 150
<< mvndiff >>
rect -88 98 0 150
rect -88 52 -75 98
rect -29 52 0 98
rect -88 0 0 52
rect 120 98 208 150
rect 120 52 149 98
rect 195 52 208 98
rect 120 0 208 52
<< mvndiffc >>
rect -75 52 -29 98
rect 149 52 195 98
<< polysilicon >>
rect 0 150 120 194
rect 0 -44 120 0
<< metal1 >>
rect -75 98 -29 150
rect -75 0 -29 52
rect 149 98 195 150
rect 149 0 195 52
<< labels >>
flabel metal1 s -52 75 -52 75 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 75 172 75 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 921886
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 920862
<< end >>
