magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 147 8 159
rect 0 -3 8 9
<< labels >>
rlabel metal1 s 0 147 8 159 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -3 8 9 6 VSS
port 2 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 -3 8 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 342076
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 341800
<< end >>
