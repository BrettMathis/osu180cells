magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 2600 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 520 190 580 360
rect 690 190 750 360
rect 800 190 860 360
rect 970 190 1030 360
rect 1080 190 1140 360
rect 1250 190 1310 360
rect 1360 190 1420 360
rect 1530 190 1590 360
rect 1850 190 1910 360
rect 2170 190 2230 360
rect 2340 190 2400 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 520 1090 580 1430
rect 690 1090 750 1430
rect 800 1090 860 1430
rect 970 1090 1030 1430
rect 1080 1090 1140 1430
rect 1250 1090 1310 1430
rect 1360 1090 1420 1430
rect 1530 1090 1590 1430
rect 1850 1090 1910 1430
rect 2170 1090 2230 1430
rect 2340 1090 2400 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 520 360
rect 580 298 690 360
rect 580 252 612 298
rect 658 252 690 298
rect 580 190 690 252
rect 750 190 800 360
rect 860 258 970 360
rect 860 212 892 258
rect 938 212 970 258
rect 860 190 970 212
rect 1030 190 1080 360
rect 1140 298 1250 360
rect 1140 252 1172 298
rect 1218 252 1250 298
rect 1140 190 1250 252
rect 1310 190 1360 360
rect 1420 298 1530 360
rect 1420 252 1452 298
rect 1498 252 1530 298
rect 1420 190 1530 252
rect 1590 298 1690 360
rect 1590 252 1622 298
rect 1668 252 1690 298
rect 1590 190 1690 252
rect 1750 263 1850 360
rect 1750 217 1772 263
rect 1818 217 1850 263
rect 1750 190 1850 217
rect 1910 298 2010 360
rect 1910 252 1942 298
rect 1988 252 2010 298
rect 1910 190 2010 252
rect 2070 298 2170 360
rect 2070 252 2092 298
rect 2138 252 2170 298
rect 2070 190 2170 252
rect 2230 298 2340 360
rect 2230 252 2262 298
rect 2308 252 2340 298
rect 2230 190 2340 252
rect 2400 298 2500 360
rect 2400 252 2432 298
rect 2478 252 2500 298
rect 2400 190 2500 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1090 520 1430
rect 580 1377 690 1430
rect 580 1143 612 1377
rect 658 1143 690 1377
rect 580 1090 690 1143
rect 750 1090 800 1430
rect 860 1377 970 1430
rect 860 1143 892 1377
rect 938 1143 970 1377
rect 860 1090 970 1143
rect 1030 1090 1080 1430
rect 1140 1405 1250 1430
rect 1140 1265 1172 1405
rect 1218 1265 1250 1405
rect 1140 1090 1250 1265
rect 1310 1090 1360 1430
rect 1420 1405 1530 1430
rect 1420 1265 1452 1405
rect 1498 1265 1530 1405
rect 1420 1090 1530 1265
rect 1590 1377 1690 1430
rect 1590 1143 1622 1377
rect 1668 1143 1690 1377
rect 1590 1090 1690 1143
rect 1750 1377 1850 1430
rect 1750 1143 1772 1377
rect 1818 1143 1850 1377
rect 1750 1090 1850 1143
rect 1910 1377 2010 1430
rect 1910 1143 1942 1377
rect 1988 1143 2010 1377
rect 1910 1090 2010 1143
rect 2070 1377 2170 1430
rect 2070 1143 2092 1377
rect 2138 1143 2170 1377
rect 2070 1090 2170 1143
rect 2230 1377 2340 1430
rect 2230 1143 2262 1377
rect 2308 1143 2340 1377
rect 2230 1090 2340 1143
rect 2400 1377 2500 1430
rect 2400 1143 2432 1377
rect 2478 1143 2500 1377
rect 2400 1090 2500 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 612 252 658 298
rect 892 212 938 258
rect 1172 252 1218 298
rect 1452 252 1498 298
rect 1622 252 1668 298
rect 1772 217 1818 263
rect 1942 252 1988 298
rect 2092 252 2138 298
rect 2262 252 2308 298
rect 2432 252 2478 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 612 1143 658 1377
rect 892 1143 938 1377
rect 1172 1265 1218 1405
rect 1452 1265 1498 1405
rect 1622 1143 1668 1377
rect 1772 1143 1818 1377
rect 1942 1143 1988 1377
rect 2092 1143 2138 1377
rect 2262 1143 2308 1377
rect 2432 1143 2478 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
rect 1290 1568 1380 1590
rect 1290 1522 1312 1568
rect 1358 1522 1380 1568
rect 1290 1500 1380 1522
rect 1530 1568 1620 1590
rect 1530 1522 1552 1568
rect 1598 1522 1620 1568
rect 1530 1500 1620 1522
rect 1770 1568 1860 1590
rect 1770 1522 1792 1568
rect 1838 1522 1860 1568
rect 1770 1500 1860 1522
rect 2010 1568 2100 1590
rect 2010 1522 2032 1568
rect 2078 1522 2100 1568
rect 2010 1500 2100 1522
rect 2250 1568 2340 1590
rect 2250 1522 2272 1568
rect 2318 1522 2340 1568
rect 2250 1500 2340 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
rect 1552 1522 1598 1568
rect 1792 1522 1838 1568
rect 2032 1522 2078 1568
rect 2272 1522 2318 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 520 1430 580 1480
rect 690 1430 750 1480
rect 800 1430 860 1480
rect 970 1430 1030 1480
rect 1080 1430 1140 1480
rect 1250 1430 1310 1480
rect 1360 1430 1420 1480
rect 1530 1430 1590 1480
rect 1850 1430 1910 1480
rect 2170 1430 2230 1480
rect 2340 1430 2400 1480
rect 190 910 250 1090
rect 190 883 310 910
rect 190 837 237 883
rect 283 837 310 883
rect 190 810 310 837
rect 190 360 250 810
rect 360 780 420 1090
rect 520 910 580 1090
rect 520 883 620 910
rect 520 837 547 883
rect 593 837 620 883
rect 520 810 620 837
rect 360 753 480 780
rect 360 707 407 753
rect 453 707 480 753
rect 360 680 480 707
rect 360 360 420 680
rect 690 640 750 1090
rect 800 1040 860 1090
rect 970 1040 1030 1090
rect 800 1013 1030 1040
rect 800 970 837 1013
rect 810 967 837 970
rect 883 970 1030 1013
rect 883 967 910 970
rect 810 920 910 967
rect 1080 640 1140 1090
rect 1250 910 1310 1090
rect 1210 883 1310 910
rect 1210 837 1237 883
rect 1283 837 1310 883
rect 1210 810 1310 837
rect 1360 780 1420 1090
rect 1530 910 1590 1090
rect 1530 883 1630 910
rect 1530 837 1557 883
rect 1603 837 1630 883
rect 1530 810 1630 837
rect 1350 753 1460 780
rect 1350 707 1377 753
rect 1423 707 1460 753
rect 1350 680 1460 707
rect 1210 640 1310 650
rect 520 623 1310 640
rect 520 580 1237 623
rect 520 360 580 580
rect 1210 577 1237 580
rect 1283 577 1310 623
rect 1210 550 1310 577
rect 650 493 750 520
rect 810 500 910 520
rect 650 447 677 493
rect 723 447 750 493
rect 650 420 750 447
rect 690 360 750 420
rect 800 493 1030 500
rect 800 447 837 493
rect 883 447 1030 493
rect 800 420 1030 447
rect 800 360 860 420
rect 970 360 1030 420
rect 1080 483 1180 510
rect 1080 437 1107 483
rect 1153 437 1180 483
rect 1080 410 1180 437
rect 1080 360 1140 410
rect 1250 360 1310 550
rect 1360 360 1420 680
rect 1530 360 1590 810
rect 1850 650 1910 1090
rect 2170 650 2230 1090
rect 2340 910 2400 1090
rect 2280 883 2400 910
rect 2280 837 2307 883
rect 2353 837 2400 883
rect 2280 810 2400 837
rect 1790 623 1910 650
rect 1790 577 1817 623
rect 1863 577 1910 623
rect 1790 550 1910 577
rect 2110 623 2230 650
rect 2110 577 2157 623
rect 2203 577 2230 623
rect 2110 550 2230 577
rect 1850 360 1910 550
rect 2170 360 2230 550
rect 2340 360 2400 810
rect 190 140 250 190
rect 360 140 420 190
rect 520 140 580 190
rect 690 140 750 190
rect 800 140 860 190
rect 970 140 1030 190
rect 1080 140 1140 190
rect 1250 140 1310 190
rect 1360 140 1420 190
rect 1530 140 1590 190
rect 1850 140 1910 190
rect 2170 140 2230 190
rect 2340 140 2400 190
<< polycontact >>
rect 237 837 283 883
rect 547 837 593 883
rect 407 707 453 753
rect 837 967 883 1013
rect 1237 837 1283 883
rect 1557 837 1603 883
rect 1377 707 1423 753
rect 1237 577 1283 623
rect 677 447 723 493
rect 837 447 883 493
rect 1107 437 1153 483
rect 2307 837 2353 883
rect 1817 577 1863 623
rect 2157 577 2203 623
<< metal1 >>
rect 0 1568 2600 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1552 1568
rect 1598 1566 1792 1568
rect 1838 1566 2032 1568
rect 2078 1566 2272 1568
rect 2318 1566 2600 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 1366 1522 1552 1566
rect 1606 1522 1792 1566
rect 1846 1522 2032 1566
rect 2086 1522 2272 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1794 1522
rect 1846 1514 2034 1522
rect 2086 1514 2274 1522
rect 2326 1514 2600 1566
rect 0 1470 2600 1514
rect 110 1377 160 1430
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 520 160 1143
rect 280 1377 330 1470
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 1060 330 1143
rect 610 1377 660 1430
rect 610 1143 612 1377
rect 658 1143 660 1377
rect 610 1040 660 1143
rect 890 1377 940 1470
rect 890 1143 892 1377
rect 938 1143 940 1377
rect 1170 1405 1220 1430
rect 1170 1265 1172 1405
rect 1218 1265 1220 1405
rect 1170 1240 1220 1265
rect 890 1060 940 1143
rect 990 1190 1220 1240
rect 1450 1405 1500 1470
rect 1450 1265 1452 1405
rect 1498 1265 1500 1405
rect 1450 1210 1500 1265
rect 1620 1377 1670 1430
rect 280 990 660 1040
rect 810 1013 910 1020
rect 280 890 330 990
rect 810 967 837 1013
rect 883 967 910 1013
rect 810 960 910 967
rect 210 883 330 890
rect 210 837 237 883
rect 283 837 330 883
rect 210 830 330 837
rect 100 496 160 520
rect 100 444 104 496
rect 156 444 160 496
rect 280 500 330 830
rect 520 886 750 890
rect 520 883 674 886
rect 520 837 547 883
rect 593 837 674 883
rect 520 834 674 837
rect 726 834 750 886
rect 520 800 750 834
rect 380 756 480 760
rect 380 704 404 756
rect 456 704 480 756
rect 380 670 480 704
rect 670 500 730 800
rect 830 500 890 960
rect 990 740 1040 1190
rect 1620 1143 1622 1377
rect 1668 1143 1670 1377
rect 1340 1016 1440 1020
rect 1340 964 1364 1016
rect 1416 964 1440 1016
rect 1340 960 1440 964
rect 1620 1000 1670 1143
rect 1770 1377 1820 1470
rect 1770 1143 1772 1377
rect 1818 1143 1820 1377
rect 1770 1060 1820 1143
rect 1940 1377 1990 1430
rect 1940 1143 1942 1377
rect 1988 1143 1990 1377
rect 980 690 1040 740
rect 1100 886 1310 890
rect 1100 834 1234 886
rect 1286 834 1310 886
rect 1100 800 1310 834
rect 280 450 480 500
rect 100 420 160 444
rect 110 298 160 420
rect 400 360 480 450
rect 650 493 750 500
rect 650 447 677 493
rect 723 447 750 493
rect 650 410 750 447
rect 810 496 910 500
rect 810 444 834 496
rect 886 444 910 496
rect 810 440 910 444
rect 980 370 1030 690
rect 1100 490 1160 800
rect 1360 760 1420 960
rect 1620 950 1780 1000
rect 1530 886 1630 890
rect 1530 834 1554 886
rect 1606 834 1630 886
rect 1530 800 1630 834
rect 1720 760 1780 950
rect 1350 756 1460 760
rect 1350 704 1374 756
rect 1426 704 1460 756
rect 1350 700 1460 704
rect 1620 710 1780 760
rect 1360 690 1440 700
rect 1210 626 1310 630
rect 1210 574 1234 626
rect 1286 574 1310 626
rect 1210 570 1310 574
rect 1620 626 1680 710
rect 1810 630 1870 650
rect 1940 630 1990 1143
rect 2090 1377 2140 1430
rect 2090 1143 2092 1377
rect 2138 1143 2140 1377
rect 2090 890 2140 1143
rect 2260 1377 2310 1470
rect 2260 1143 2262 1377
rect 2308 1143 2310 1377
rect 2260 1060 2310 1143
rect 2430 1377 2480 1430
rect 2430 1143 2432 1377
rect 2478 1143 2480 1377
rect 2430 1030 2480 1143
rect 2430 1016 2530 1030
rect 2430 964 2454 1016
rect 2506 964 2530 1016
rect 2430 930 2530 964
rect 2430 920 2520 930
rect 2090 886 2380 890
rect 2090 834 2304 886
rect 2356 834 2380 886
rect 2090 800 2380 834
rect 1620 574 1624 626
rect 1676 574 1680 626
rect 1620 550 1680 574
rect 1790 623 1890 630
rect 1790 577 1817 623
rect 1863 577 1890 623
rect 1790 570 1890 577
rect 1940 626 2230 630
rect 1940 574 2154 626
rect 2206 574 2230 626
rect 1940 570 2230 574
rect 1080 483 1180 490
rect 1080 437 1107 483
rect 1153 437 1180 483
rect 1080 400 1180 437
rect 980 366 1250 370
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 400 310 660 360
rect 980 320 1174 366
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 610 298 660 310
rect 610 252 612 298
rect 658 252 660 298
rect 1170 314 1174 320
rect 1226 314 1250 366
rect 1170 310 1250 314
rect 1170 298 1220 310
rect 610 190 660 252
rect 890 258 940 280
rect 890 212 892 258
rect 938 212 940 258
rect 890 120 940 212
rect 1170 252 1172 298
rect 1218 252 1220 298
rect 1170 190 1220 252
rect 1450 298 1500 360
rect 1450 252 1452 298
rect 1498 252 1500 298
rect 1450 120 1500 252
rect 1620 298 1670 550
rect 1810 400 1870 570
rect 1790 396 1890 400
rect 1790 344 1814 396
rect 1866 344 1890 396
rect 1790 340 1890 344
rect 1620 252 1622 298
rect 1668 252 1670 298
rect 1940 298 1990 570
rect 2310 460 2360 800
rect 1620 190 1670 252
rect 1770 263 1820 290
rect 1770 217 1772 263
rect 1818 217 1820 263
rect 1770 120 1820 217
rect 1940 252 1942 298
rect 1988 252 1990 298
rect 1940 190 1990 252
rect 2090 380 2360 460
rect 2090 298 2140 380
rect 2090 252 2092 298
rect 2138 252 2140 298
rect 2090 160 2140 252
rect 2260 298 2310 360
rect 2260 252 2262 298
rect 2308 252 2310 298
rect 2260 120 2310 252
rect 2430 298 2480 920
rect 2430 252 2432 298
rect 2478 252 2480 298
rect 2430 160 2480 252
rect 0 106 2600 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2600 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2600 54
rect 0 -30 2600 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 1554 1522 1598 1566
rect 1598 1522 1606 1566
rect 1794 1522 1838 1566
rect 1838 1522 1846 1566
rect 2034 1522 2078 1566
rect 2078 1522 2086 1566
rect 2274 1522 2318 1566
rect 2318 1522 2326 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 1794 1514 1846 1522
rect 2034 1514 2086 1522
rect 2274 1514 2326 1522
rect 104 444 156 496
rect 674 834 726 886
rect 404 753 456 756
rect 404 707 407 753
rect 407 707 453 753
rect 453 707 456 753
rect 404 704 456 707
rect 1364 964 1416 1016
rect 1234 883 1286 886
rect 1234 837 1237 883
rect 1237 837 1283 883
rect 1283 837 1286 883
rect 1234 834 1286 837
rect 834 493 886 496
rect 834 447 837 493
rect 837 447 883 493
rect 883 447 886 493
rect 834 444 886 447
rect 1554 883 1606 886
rect 1554 837 1557 883
rect 1557 837 1603 883
rect 1603 837 1606 883
rect 1554 834 1606 837
rect 1374 753 1426 756
rect 1374 707 1377 753
rect 1377 707 1423 753
rect 1423 707 1426 753
rect 1374 704 1426 707
rect 1234 623 1286 626
rect 1234 577 1237 623
rect 1237 577 1283 623
rect 1283 577 1286 623
rect 1234 574 1286 577
rect 2454 964 2506 1016
rect 2304 883 2356 886
rect 2304 837 2307 883
rect 2307 837 2353 883
rect 2353 837 2356 883
rect 2304 834 2356 837
rect 1624 574 1676 626
rect 2154 623 2206 626
rect 2154 577 2157 623
rect 2157 577 2203 623
rect 2203 577 2206 623
rect 2154 574 2206 577
rect 1174 314 1226 366
rect 1814 344 1866 396
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect 1780 1570 1860 1580
rect 2020 1570 2100 1580
rect 2260 1570 2340 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1480 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1480 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1480 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1480 1390 1514
rect 1530 1566 1630 1570
rect 1530 1514 1554 1566
rect 1606 1514 1630 1566
rect 1530 1480 1630 1514
rect 1770 1566 1870 1570
rect 1770 1514 1794 1566
rect 1846 1514 1870 1566
rect 1770 1480 1870 1514
rect 2010 1566 2110 1570
rect 2010 1514 2034 1566
rect 2086 1514 2110 1566
rect 2010 1480 2110 1514
rect 2250 1566 2350 1570
rect 2250 1514 2274 1566
rect 2326 1514 2350 1566
rect 2250 1480 2350 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 580 1470 660 1480
rect 820 1470 900 1480
rect 1060 1470 1140 1480
rect 1300 1470 1380 1480
rect 1540 1470 1620 1480
rect 1780 1470 1860 1480
rect 2020 1470 2100 1480
rect 2260 1470 2340 1480
rect 1350 1020 1430 1030
rect 2440 1020 2520 1030
rect 1340 1016 1980 1020
rect 1340 964 1364 1016
rect 1416 964 1980 1016
rect 1340 960 1980 964
rect 1350 950 1430 960
rect 650 890 740 900
rect 1210 890 1310 900
rect 1540 890 1620 900
rect 650 886 1630 890
rect 650 834 674 886
rect 726 834 1234 886
rect 1286 834 1554 886
rect 1606 834 1630 886
rect 650 800 1630 834
rect 650 790 740 800
rect 1210 790 1310 800
rect 1540 790 1620 800
rect 380 760 480 770
rect 1360 760 1440 770
rect 350 756 510 760
rect 350 704 404 756
rect 456 704 510 756
rect 350 670 510 704
rect 1350 756 1450 760
rect 1350 704 1374 756
rect 1426 704 1450 756
rect 1350 700 1450 704
rect 1360 690 1440 700
rect 380 660 480 670
rect 1220 630 1300 640
rect 1610 630 1690 640
rect 1920 630 1980 960
rect 2430 1016 2530 1020
rect 2430 964 2454 1016
rect 2506 964 2530 1016
rect 2430 930 2530 964
rect 2440 920 2520 930
rect 2290 890 2370 900
rect 2280 886 2380 890
rect 2280 834 2304 886
rect 2356 834 2380 886
rect 2280 800 2380 834
rect 2290 790 2370 800
rect 2140 630 2220 640
rect 1210 626 1710 630
rect 1210 574 1234 626
rect 1286 574 1624 626
rect 1676 574 1710 626
rect 1210 570 1710 574
rect 1920 626 2230 630
rect 1920 574 2154 626
rect 2206 574 2230 626
rect 1920 570 2230 574
rect 1220 560 1300 570
rect 1610 560 1690 570
rect 2140 560 2220 570
rect 90 500 170 510
rect 820 500 900 510
rect 80 496 910 500
rect 80 444 104 496
rect 156 444 834 496
rect 886 444 910 496
rect 80 440 910 444
rect 90 430 170 440
rect 820 430 900 440
rect 1800 400 1880 410
rect 1700 396 1890 400
rect 1160 370 1240 380
rect 1700 370 1814 396
rect 1150 366 1814 370
rect 1150 314 1174 366
rect 1226 344 1814 366
rect 1866 344 1890 396
rect 1226 340 1890 344
rect 1226 330 1880 340
rect 1226 314 1760 330
rect 1150 310 1760 314
rect 1160 300 1240 310
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 20 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 20 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 20 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 20 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 20 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 20 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 20 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 20 2350 54
rect 100 10 180 20
rect 340 10 420 20
rect 580 10 660 20
rect 820 10 900 20
rect 1060 10 1140 20
rect 1300 10 1380 20
rect 1540 10 1620 20
rect 1780 10 1860 20
rect 2020 10 2100 20
rect 2260 10 2340 20
<< labels >>
rlabel metal2 s 100 10 180 90 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 100 1470 180 1550 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 380 660 480 740 4 D
port 1 nsew signal input
rlabel metal2 s 2440 920 2520 1000 4 Q
port 2 nsew signal output
rlabel metal2 s 2290 790 2370 870 4 QN
port 3 nsew signal output
rlabel metal2 s 650 790 740 870 4 CLK
port 4 nsew clock input
rlabel metal2 s 1210 790 1310 870 1 CLK
port 4 nsew clock input
rlabel metal2 s 1540 790 1620 870 1 CLK
port 4 nsew clock input
rlabel metal2 s 650 800 1630 860 1 CLK
port 4 nsew clock input
rlabel metal1 s 670 410 730 860 1 CLK
port 4 nsew clock input
rlabel metal1 s 650 410 750 470 1 CLK
port 4 nsew clock input
rlabel metal1 s 520 800 750 860 1 CLK
port 4 nsew clock input
rlabel metal1 s 1100 400 1160 860 1 CLK
port 4 nsew clock input
rlabel metal1 s 1080 400 1180 460 1 CLK
port 4 nsew clock input
rlabel metal1 s 1100 800 1310 860 1 CLK
port 4 nsew clock input
rlabel metal1 s 1530 800 1630 860 1 CLK
port 4 nsew clock input
rlabel metal2 s 350 670 510 730 1 D
port 1 nsew signal input
rlabel metal1 s 380 670 480 730 1 D
port 1 nsew signal input
rlabel metal2 s 2430 930 2530 990 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 160 2480 1400 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 920 2520 1000 1 Q
port 2 nsew signal output
rlabel metal1 s 2430 930 2530 1000 1 Q
port 2 nsew signal output
rlabel metal2 s 2280 800 2380 860 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 160 2140 430 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 800 2140 1400 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 380 2360 430 1 QN
port 3 nsew signal output
rlabel metal1 s 2310 380 2360 860 1 QN
port 3 nsew signal output
rlabel metal1 s 2090 800 2380 860 1 QN
port 3 nsew signal output
rlabel metal2 s 90 1480 190 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 1470 660 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 570 1480 670 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 820 1470 900 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 810 1480 910 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1060 1470 1140 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1050 1480 1150 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1300 1470 1380 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1290 1480 1390 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1540 1470 1620 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1530 1480 1630 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1780 1470 1860 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1770 1480 1870 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2020 1470 2100 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2010 1480 2110 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2260 1470 2340 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 2250 1480 2350 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 280 1060 330 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 890 1060 940 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1450 1210 1500 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1770 1060 1820 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 2260 1060 2310 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 1470 2600 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 580 10 660 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 570 20 670 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 820 10 900 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 810 20 910 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1060 10 1140 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1050 20 1150 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1300 10 1380 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1290 20 1390 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1540 10 1620 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1530 20 1630 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1780 10 1860 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1770 20 1870 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2020 10 2100 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2010 20 2110 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2260 10 2340 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 2250 20 2350 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 280 -30 330 330 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 890 -30 940 250 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1450 -30 1500 330 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1770 -30 1820 260 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 2260 -30 2310 330 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 0 -30 2600 90 1 VSS
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 -30 2600 1590
string GDS_END 242606
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 216576
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
