magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 407 2326 870
rect -86 352 575 407
rect 943 352 2326 407
<< pwell >>
rect 575 352 943 407
rect -86 -86 2326 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 1064 68 1184 176
rect 1288 68 1408 176
rect 1548 68 1668 232
rect 1772 68 1892 232
rect 1996 68 2116 232
<< mvpmos >>
rect 172 527 272 716
rect 376 527 476 716
rect 660 527 760 716
rect 1130 514 1230 716
rect 1334 514 1434 716
rect 1574 481 1674 716
rect 1778 481 1878 716
rect 1982 481 2082 716
<< mvndiff >>
rect 752 274 824 287
rect 752 232 765 274
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 128 348 232
rect 244 82 273 128
rect 319 82 348 128
rect 244 68 348 82
rect 468 169 572 232
rect 468 123 497 169
rect 543 123 572 169
rect 468 68 572 123
rect 692 228 765 232
rect 811 228 824 274
rect 692 68 824 228
rect 1468 176 1548 232
rect 932 95 1064 176
rect 932 49 945 95
rect 991 68 1064 95
rect 1184 163 1288 176
rect 1184 117 1213 163
rect 1259 117 1288 163
rect 1184 68 1288 117
rect 1408 127 1548 176
rect 1408 81 1455 127
rect 1501 81 1548 127
rect 1408 68 1548 81
rect 1668 219 1772 232
rect 1668 173 1697 219
rect 1743 173 1772 219
rect 1668 68 1772 173
rect 1892 127 1996 232
rect 1892 81 1921 127
rect 1967 81 1996 127
rect 1892 68 1996 81
rect 2116 219 2204 232
rect 2116 173 2145 219
rect 2191 173 2204 219
rect 2116 68 2204 173
rect 991 49 1004 68
rect 932 36 1004 49
<< mvpdiff >>
rect 84 602 172 716
rect 84 556 97 602
rect 143 556 172 602
rect 84 527 172 556
rect 272 698 376 716
rect 272 652 301 698
rect 347 652 376 698
rect 272 527 376 652
rect 476 678 660 716
rect 476 632 585 678
rect 631 632 660 678
rect 476 527 660 632
rect 760 586 848 716
rect 760 540 789 586
rect 835 540 848 586
rect 760 527 848 540
rect 1042 703 1130 716
rect 1042 657 1055 703
rect 1101 657 1130 703
rect 1042 514 1130 657
rect 1230 667 1334 716
rect 1230 527 1259 667
rect 1305 527 1334 667
rect 1230 514 1334 527
rect 1434 703 1574 716
rect 1434 657 1463 703
rect 1509 657 1574 703
rect 1434 514 1574 657
rect 1494 481 1574 514
rect 1674 667 1778 716
rect 1674 527 1703 667
rect 1749 527 1778 667
rect 1674 481 1778 527
rect 1878 703 1982 716
rect 1878 657 1907 703
rect 1953 657 1982 703
rect 1878 481 1982 657
rect 2082 667 2170 716
rect 2082 527 2111 667
rect 2157 527 2170 667
rect 2082 481 2170 527
<< mvndiffc >>
rect 49 173 95 219
rect 273 82 319 128
rect 497 123 543 169
rect 765 228 811 274
rect 945 49 991 95
rect 1213 117 1259 163
rect 1455 81 1501 127
rect 1697 173 1743 219
rect 1921 81 1967 127
rect 2145 173 2191 219
<< mvpdiffc >>
rect 97 556 143 602
rect 301 652 347 698
rect 585 632 631 678
rect 789 540 835 586
rect 1055 657 1101 703
rect 1259 527 1305 667
rect 1463 657 1509 703
rect 1703 527 1749 667
rect 1907 657 1953 703
rect 2111 527 2157 667
<< polysilicon >>
rect 172 716 272 760
rect 376 716 476 760
rect 660 716 760 760
rect 1130 716 1230 760
rect 1334 716 1434 760
rect 1574 716 1674 760
rect 1778 716 1878 760
rect 1982 716 2082 760
rect 172 413 272 527
rect 376 413 476 527
rect 660 493 760 527
rect 660 447 673 493
rect 719 447 760 493
rect 660 434 760 447
rect 1130 415 1230 514
rect 124 412 612 413
rect 124 366 185 412
rect 231 373 612 412
rect 1130 399 1157 415
rect 231 366 244 373
rect 124 232 244 366
rect 348 311 468 324
rect 348 265 385 311
rect 431 265 468 311
rect 348 232 468 265
rect 572 288 612 373
rect 1064 369 1157 399
rect 1203 399 1230 415
rect 1334 415 1434 514
rect 1334 399 1361 415
rect 1203 369 1361 399
rect 1407 369 1434 415
rect 1574 439 1674 481
rect 1574 393 1601 439
rect 1647 420 1674 439
rect 1778 439 1878 481
rect 1778 420 1805 439
rect 1647 393 1805 420
rect 1851 420 1878 439
rect 1982 439 2082 481
rect 1982 420 2009 439
rect 1851 393 2009 420
rect 2055 393 2082 439
rect 1574 380 2082 393
rect 1064 349 1434 369
rect 572 232 692 288
rect 1064 176 1184 349
rect 1288 176 1408 349
rect 1548 319 2116 332
rect 1548 273 1585 319
rect 1631 292 1809 319
rect 1631 273 1668 292
rect 1548 232 1668 273
rect 1772 273 1809 292
rect 1855 292 2033 319
rect 1855 273 1892 292
rect 1772 232 1892 273
rect 1996 273 2033 292
rect 2079 273 2116 319
rect 1996 232 2116 273
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1064 24 1184 68
rect 1288 24 1408 68
rect 1548 24 1668 68
rect 1772 24 1892 68
rect 1996 24 2116 68
<< polycontact >>
rect 673 447 719 493
rect 185 366 231 412
rect 385 265 431 311
rect 1157 369 1203 415
rect 1361 369 1407 415
rect 1601 393 1647 439
rect 1805 393 1851 439
rect 2009 393 2055 439
rect 1585 273 1631 319
rect 1809 273 1855 319
rect 2033 273 2079 319
<< metal1 >>
rect 0 724 2240 844
rect 290 698 358 724
rect 290 652 301 698
rect 347 652 358 698
rect 1044 703 1112 724
rect 574 632 585 678
rect 631 632 965 678
rect 1044 657 1055 703
rect 1101 657 1112 703
rect 1452 703 1520 724
rect 1248 667 1316 678
rect 84 556 97 602
rect 143 556 431 602
rect 385 504 431 556
rect 778 540 789 586
rect 835 540 846 586
rect 385 493 730 504
rect 385 447 673 493
rect 719 447 730 493
rect 109 412 326 437
rect 109 366 185 412
rect 231 366 326 412
rect 109 355 326 366
rect 385 311 431 447
rect 778 401 846 540
rect 38 219 431 265
rect 497 355 846 401
rect 919 561 965 632
rect 1248 561 1259 667
rect 919 527 1259 561
rect 1305 561 1316 667
rect 1452 657 1463 703
rect 1509 657 1520 703
rect 1896 703 1964 724
rect 1692 667 1760 678
rect 1305 527 1571 561
rect 919 515 1571 527
rect 38 173 49 219
rect 95 173 106 219
rect 38 170 106 173
rect 497 169 543 355
rect 919 309 965 515
rect 1525 439 1571 515
rect 1692 527 1703 667
rect 1749 554 1760 667
rect 1896 657 1907 703
rect 1953 657 1964 703
rect 2100 667 2168 678
rect 2100 554 2111 667
rect 1749 527 2111 554
rect 2157 554 2168 667
rect 2157 527 2214 554
rect 1692 508 2214 527
rect 1018 415 1455 424
rect 1018 369 1157 415
rect 1203 369 1361 415
rect 1407 369 1455 415
rect 1525 393 1601 439
rect 1647 393 1805 439
rect 1851 393 2009 439
rect 2055 393 2074 439
rect 1018 360 1455 369
rect 754 274 965 309
rect 754 228 765 274
rect 811 263 965 274
rect 1557 273 1585 319
rect 1631 273 1809 319
rect 1855 273 2033 319
rect 2079 273 2098 319
rect 811 228 822 263
rect 1557 219 1603 273
rect 2148 227 2214 508
rect 1184 187 1603 219
rect 262 128 330 131
rect 262 82 273 128
rect 319 82 330 128
rect 843 173 1603 187
rect 1668 219 2214 227
rect 1668 173 1697 219
rect 1743 173 2145 219
rect 2191 173 2214 219
rect 843 163 1274 173
rect 843 152 1213 163
rect 543 141 1213 152
rect 543 123 888 141
rect 497 106 888 123
rect 1184 117 1213 141
rect 1259 117 1274 163
rect 262 60 330 82
rect 934 60 945 95
rect 0 49 945 60
rect 991 60 1002 95
rect 1444 81 1455 127
rect 1501 81 1512 127
rect 1444 60 1512 81
rect 1910 81 1921 127
rect 1967 81 1978 127
rect 1910 60 1978 81
rect 991 49 2240 60
rect 0 -60 2240 49
<< labels >>
flabel metal1 s 109 355 326 437 0 FreeSans 600 0 0 0 EN
port 1 nsew default input
flabel metal1 s 0 724 2240 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 262 127 330 131 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2100 554 2168 678 0 FreeSans 400 0 0 0 Z
port 3 nsew default output
flabel metal1 s 1018 360 1455 424 0 FreeSans 400 0 0 0 I
port 2 nsew default input
rlabel metal1 s 1692 554 1760 678 1 Z
port 3 nsew default output
rlabel metal1 s 1692 508 2214 554 1 Z
port 3 nsew default output
rlabel metal1 s 2148 227 2214 508 1 Z
port 3 nsew default output
rlabel metal1 s 1668 173 2214 227 1 Z
port 3 nsew default output
rlabel metal1 s 1896 657 1964 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1452 657 1520 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1044 657 1112 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 657 358 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1910 95 1978 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1444 95 1512 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 95 330 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1910 60 1978 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1444 60 1512 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2240 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2240 784
string GDS_END 1374566
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1368900
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
