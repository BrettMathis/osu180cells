magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 5889 11760 13827 16428
rect 6717 7412 7860 7872
rect 6493 7185 7860 7412
rect 542 6727 5430 7122
rect 542 6338 5654 6727
rect 4800 5991 5654 6338
rect 6234 5995 7860 7185
rect 10123 5152 10509 9334
rect -73 2245 8748 3429
rect 7919 852 8748 2245
rect 7137 -1400 8748 852
<< mvnmos >>
rect 9526 262 9646 4798
rect 9750 262 9870 4798
rect 9974 262 10094 4798
rect 10725 484 10845 4113
rect 10949 484 11069 4113
rect 11173 484 11293 4113
rect 11397 484 11517 4113
rect 12010 3205 12130 4113
rect 12233 3205 12353 4113
rect 12458 3205 12578 4113
rect 12681 3205 12801 4113
<< mvpmos >>
rect 5055 6131 5174 6587
rect 5279 6131 5398 6587
<< mvndiff >>
rect 9407 4752 9526 4798
rect 9407 4706 9451 4752
rect 9497 4706 9526 4752
rect 9407 4584 9526 4706
rect 9407 4538 9451 4584
rect 9497 4538 9526 4584
rect 9407 4417 9526 4538
rect 9407 4371 9451 4417
rect 9497 4371 9526 4417
rect 9407 4249 9526 4371
rect 9407 4203 9451 4249
rect 9497 4203 9526 4249
rect 9407 4081 9526 4203
rect 9407 4035 9451 4081
rect 9497 4035 9526 4081
rect 9407 3913 9526 4035
rect 9407 3867 9451 3913
rect 9497 3867 9526 3913
rect 9407 3746 9526 3867
rect 9407 3700 9451 3746
rect 9497 3700 9526 3746
rect 9407 3578 9526 3700
rect 9407 3532 9451 3578
rect 9497 3532 9526 3578
rect 9407 3410 9526 3532
rect 9407 3364 9451 3410
rect 9497 3364 9526 3410
rect 9407 3242 9526 3364
rect 9407 3196 9451 3242
rect 9497 3196 9526 3242
rect 9407 3075 9526 3196
rect 9407 3029 9451 3075
rect 9497 3029 9526 3075
rect 9407 2905 9526 3029
rect 9407 2859 9451 2905
rect 9497 2859 9526 2905
rect 9407 2735 9526 2859
rect 9407 2689 9451 2735
rect 9497 2689 9526 2735
rect 9407 2565 9526 2689
rect 9407 2519 9451 2565
rect 9497 2519 9526 2565
rect 9407 2395 9526 2519
rect 9407 2349 9451 2395
rect 9497 2349 9526 2395
rect 9407 2225 9526 2349
rect 9407 2179 9451 2225
rect 9497 2179 9526 2225
rect 9407 2055 9526 2179
rect 9407 2009 9451 2055
rect 9497 2009 9526 2055
rect 9407 1884 9526 2009
rect 9407 1838 9451 1884
rect 9497 1838 9526 1884
rect 9407 1714 9526 1838
rect 9407 1668 9451 1714
rect 9497 1668 9526 1714
rect 9407 1544 9526 1668
rect 9407 1498 9451 1544
rect 9497 1498 9526 1544
rect 9407 1374 9526 1498
rect 9407 1328 9451 1374
rect 9497 1328 9526 1374
rect 9407 1204 9526 1328
rect 9407 1158 9451 1204
rect 9497 1158 9526 1204
rect 9407 1034 9526 1158
rect 9407 988 9451 1034
rect 9497 988 9526 1034
rect 9407 864 9526 988
rect 9407 818 9451 864
rect 9497 818 9526 864
rect 9407 694 9526 818
rect 9407 648 9451 694
rect 9497 648 9526 694
rect 9407 524 9526 648
rect 9407 478 9451 524
rect 9497 478 9526 524
rect 9407 354 9526 478
rect 9407 308 9451 354
rect 9497 308 9526 354
rect 9407 262 9526 308
rect 9646 262 9750 4798
rect 9870 262 9974 4798
rect 10094 4584 10212 4798
rect 10094 4538 10123 4584
rect 10169 4538 10212 4584
rect 10094 4417 10212 4538
rect 10094 4371 10123 4417
rect 10169 4371 10212 4417
rect 10094 4249 10212 4371
rect 10094 4203 10123 4249
rect 10169 4203 10212 4249
rect 10094 4081 10212 4203
rect 10094 4035 10123 4081
rect 10169 4035 10212 4081
rect 10094 3913 10212 4035
rect 10094 3867 10123 3913
rect 10169 3867 10212 3913
rect 10094 3746 10212 3867
rect 10094 3700 10123 3746
rect 10169 3700 10212 3746
rect 10094 3578 10212 3700
rect 10094 3532 10123 3578
rect 10169 3532 10212 3578
rect 10094 3410 10212 3532
rect 10094 3364 10123 3410
rect 10169 3364 10212 3410
rect 10094 3242 10212 3364
rect 10094 3196 10123 3242
rect 10169 3196 10212 3242
rect 10094 3075 10212 3196
rect 10094 3029 10123 3075
rect 10169 3029 10212 3075
rect 10094 2905 10212 3029
rect 10094 2859 10123 2905
rect 10169 2859 10212 2905
rect 10094 2735 10212 2859
rect 10094 2689 10123 2735
rect 10169 2689 10212 2735
rect 10094 2565 10212 2689
rect 10094 2519 10123 2565
rect 10169 2519 10212 2565
rect 10094 2395 10212 2519
rect 10094 2349 10123 2395
rect 10169 2349 10212 2395
rect 10094 2225 10212 2349
rect 10094 2179 10123 2225
rect 10169 2179 10212 2225
rect 10094 2055 10212 2179
rect 10094 2009 10123 2055
rect 10169 2009 10212 2055
rect 10094 1884 10212 2009
rect 10094 1838 10123 1884
rect 10169 1838 10212 1884
rect 10094 1714 10212 1838
rect 10094 1668 10123 1714
rect 10169 1668 10212 1714
rect 10094 1544 10212 1668
rect 10094 1498 10123 1544
rect 10169 1498 10212 1544
rect 10094 1374 10212 1498
rect 10094 1328 10123 1374
rect 10169 1328 10212 1374
rect 10094 1204 10212 1328
rect 10094 1158 10123 1204
rect 10169 1158 10212 1204
rect 10094 1034 10212 1158
rect 10094 988 10123 1034
rect 10169 988 10212 1034
rect 10094 864 10212 988
rect 10094 818 10123 864
rect 10169 818 10212 864
rect 10094 694 10212 818
rect 10094 648 10123 694
rect 10169 648 10212 694
rect 10094 524 10212 648
rect 10094 478 10123 524
rect 10169 478 10212 524
rect 10606 4068 10725 4113
rect 10606 4022 10650 4068
rect 10696 4022 10725 4068
rect 10606 3900 10725 4022
rect 10606 3854 10650 3900
rect 10696 3854 10725 3900
rect 10606 3732 10725 3854
rect 10606 3686 10650 3732
rect 10696 3686 10725 3732
rect 10606 3564 10725 3686
rect 10606 3518 10650 3564
rect 10696 3518 10725 3564
rect 10606 3397 10725 3518
rect 10606 3351 10650 3397
rect 10696 3351 10725 3397
rect 10606 3229 10725 3351
rect 10606 3183 10650 3229
rect 10696 3183 10725 3229
rect 10606 3061 10725 3183
rect 10606 3015 10650 3061
rect 10696 3015 10725 3061
rect 10606 2893 10725 3015
rect 10606 2847 10650 2893
rect 10696 2847 10725 2893
rect 10606 2726 10725 2847
rect 10606 2680 10650 2726
rect 10696 2680 10725 2726
rect 10606 2558 10725 2680
rect 10606 2512 10650 2558
rect 10696 2512 10725 2558
rect 10606 2390 10725 2512
rect 10606 2344 10650 2390
rect 10696 2344 10725 2390
rect 10606 2220 10725 2344
rect 10606 2174 10650 2220
rect 10696 2174 10725 2220
rect 10606 2050 10725 2174
rect 10606 2004 10650 2050
rect 10696 2004 10725 2050
rect 10606 1880 10725 2004
rect 10606 1834 10650 1880
rect 10696 1834 10725 1880
rect 10606 1710 10725 1834
rect 10606 1664 10650 1710
rect 10696 1664 10725 1710
rect 10606 1540 10725 1664
rect 10606 1494 10650 1540
rect 10696 1494 10725 1540
rect 10606 1370 10725 1494
rect 10606 1324 10650 1370
rect 10696 1324 10725 1370
rect 10606 1200 10725 1324
rect 10606 1154 10650 1200
rect 10696 1154 10725 1200
rect 10606 1030 10725 1154
rect 10606 984 10650 1030
rect 10696 984 10725 1030
rect 10606 860 10725 984
rect 10606 814 10650 860
rect 10696 814 10725 860
rect 10606 690 10725 814
rect 10606 644 10650 690
rect 10696 644 10725 690
rect 10606 484 10725 644
rect 10845 484 10949 4113
rect 11069 4068 11173 4113
rect 11069 4022 11098 4068
rect 11144 4022 11173 4068
rect 11069 3900 11173 4022
rect 11069 3854 11098 3900
rect 11144 3854 11173 3900
rect 11069 3732 11173 3854
rect 11069 3686 11098 3732
rect 11144 3686 11173 3732
rect 11069 3564 11173 3686
rect 11069 3518 11098 3564
rect 11144 3518 11173 3564
rect 11069 3397 11173 3518
rect 11069 3351 11098 3397
rect 11144 3351 11173 3397
rect 11069 3229 11173 3351
rect 11069 3183 11098 3229
rect 11144 3183 11173 3229
rect 11069 3061 11173 3183
rect 11069 3015 11098 3061
rect 11144 3015 11173 3061
rect 11069 2893 11173 3015
rect 11069 2847 11098 2893
rect 11144 2847 11173 2893
rect 11069 2726 11173 2847
rect 11069 2680 11098 2726
rect 11144 2680 11173 2726
rect 11069 2558 11173 2680
rect 11069 2512 11098 2558
rect 11144 2512 11173 2558
rect 11069 2390 11173 2512
rect 11069 2344 11098 2390
rect 11144 2344 11173 2390
rect 11069 2220 11173 2344
rect 11069 2174 11098 2220
rect 11144 2174 11173 2220
rect 11069 2050 11173 2174
rect 11069 2004 11098 2050
rect 11144 2004 11173 2050
rect 11069 1880 11173 2004
rect 11069 1834 11098 1880
rect 11144 1834 11173 1880
rect 11069 1710 11173 1834
rect 11069 1664 11098 1710
rect 11144 1664 11173 1710
rect 11069 1540 11173 1664
rect 11069 1494 11098 1540
rect 11144 1494 11173 1540
rect 11069 1370 11173 1494
rect 11069 1324 11098 1370
rect 11144 1324 11173 1370
rect 11069 1200 11173 1324
rect 11069 1154 11098 1200
rect 11144 1154 11173 1200
rect 11069 1030 11173 1154
rect 11069 984 11098 1030
rect 11144 984 11173 1030
rect 11069 860 11173 984
rect 11069 814 11098 860
rect 11144 814 11173 860
rect 11069 690 11173 814
rect 11069 644 11098 690
rect 11144 644 11173 690
rect 11069 484 11173 644
rect 11293 484 11397 4113
rect 11517 4068 11635 4113
rect 11517 4022 11546 4068
rect 11592 4022 11635 4068
rect 11517 3900 11635 4022
rect 11517 3854 11546 3900
rect 11592 3854 11635 3900
rect 11517 3732 11635 3854
rect 11517 3686 11546 3732
rect 11592 3686 11635 3732
rect 11517 3564 11635 3686
rect 11517 3518 11546 3564
rect 11592 3518 11635 3564
rect 11517 3397 11635 3518
rect 11517 3351 11546 3397
rect 11592 3351 11635 3397
rect 11517 3229 11635 3351
rect 11517 3183 11546 3229
rect 11592 3183 11635 3229
rect 11891 4068 12010 4113
rect 11891 4022 11934 4068
rect 11980 4022 12010 4068
rect 11891 3900 12010 4022
rect 11891 3854 11934 3900
rect 11980 3854 12010 3900
rect 11891 3732 12010 3854
rect 11891 3686 11934 3732
rect 11980 3686 12010 3732
rect 11891 3564 12010 3686
rect 11891 3518 11934 3564
rect 11980 3518 12010 3564
rect 11891 3397 12010 3518
rect 11891 3351 11934 3397
rect 11980 3351 12010 3397
rect 11891 3205 12010 3351
rect 12130 3205 12233 4113
rect 12353 4068 12458 4113
rect 12353 4022 12382 4068
rect 12428 4022 12458 4068
rect 12353 3900 12458 4022
rect 12353 3854 12382 3900
rect 12428 3854 12458 3900
rect 12353 3732 12458 3854
rect 12353 3686 12382 3732
rect 12428 3686 12458 3732
rect 12353 3564 12458 3686
rect 12353 3518 12382 3564
rect 12428 3518 12458 3564
rect 12353 3397 12458 3518
rect 12353 3351 12382 3397
rect 12428 3351 12458 3397
rect 12353 3205 12458 3351
rect 12578 3205 12681 4113
rect 12801 4068 12920 4113
rect 12801 4022 12830 4068
rect 12876 4022 12920 4068
rect 12801 3732 12920 4022
rect 12801 3686 12830 3732
rect 12876 3686 12920 3732
rect 12801 3564 12920 3686
rect 12801 3518 12830 3564
rect 12876 3518 12920 3564
rect 12801 3397 12920 3518
rect 12801 3351 12830 3397
rect 12876 3351 12920 3397
rect 12801 3205 12920 3351
rect 11517 3061 11635 3183
rect 11517 3015 11546 3061
rect 11592 3015 11635 3061
rect 11517 2893 11635 3015
rect 11517 2847 11546 2893
rect 11592 2847 11635 2893
rect 11517 2726 11635 2847
rect 11517 2680 11546 2726
rect 11592 2680 11635 2726
rect 11517 2558 11635 2680
rect 11517 2512 11546 2558
rect 11592 2512 11635 2558
rect 11517 2390 11635 2512
rect 11517 2344 11546 2390
rect 11592 2344 11635 2390
rect 11517 2220 11635 2344
rect 11517 2174 11546 2220
rect 11592 2174 11635 2220
rect 11517 2050 11635 2174
rect 11517 2004 11546 2050
rect 11592 2004 11635 2050
rect 11517 1880 11635 2004
rect 11517 1834 11546 1880
rect 11592 1834 11635 1880
rect 11517 1710 11635 1834
rect 11517 1664 11546 1710
rect 11592 1664 11635 1710
rect 11517 1540 11635 1664
rect 11517 1494 11546 1540
rect 11592 1494 11635 1540
rect 11517 1370 11635 1494
rect 11517 1324 11546 1370
rect 11592 1324 11635 1370
rect 11517 1200 11635 1324
rect 11517 1154 11546 1200
rect 11592 1154 11635 1200
rect 11517 1030 11635 1154
rect 11517 984 11546 1030
rect 11592 984 11635 1030
rect 11517 860 11635 984
rect 11517 814 11546 860
rect 11592 814 11635 860
rect 11517 690 11635 814
rect 11517 644 11546 690
rect 11592 644 11635 690
rect 11517 484 11635 644
rect 10094 354 10212 478
rect 10094 308 10123 354
rect 10169 308 10212 354
rect 10094 262 10212 308
<< mvpdiff >>
rect 4936 6405 5055 6587
rect 4936 6359 4980 6405
rect 5026 6359 5055 6405
rect 4936 6224 5055 6359
rect 4936 6178 4980 6224
rect 5026 6178 5055 6224
rect 4936 6131 5055 6178
rect 5174 6131 5279 6587
rect 5398 6405 5517 6587
rect 5398 6359 5428 6405
rect 5474 6359 5517 6405
rect 5398 6224 5517 6359
rect 5398 6178 5428 6224
rect 5474 6178 5517 6224
rect 5398 6131 5517 6178
<< mvndiffc >>
rect 9451 4706 9497 4752
rect 9451 4538 9497 4584
rect 9451 4371 9497 4417
rect 9451 4203 9497 4249
rect 9451 4035 9497 4081
rect 9451 3867 9497 3913
rect 9451 3700 9497 3746
rect 9451 3532 9497 3578
rect 9451 3364 9497 3410
rect 9451 3196 9497 3242
rect 9451 3029 9497 3075
rect 9451 2859 9497 2905
rect 9451 2689 9497 2735
rect 9451 2519 9497 2565
rect 9451 2349 9497 2395
rect 9451 2179 9497 2225
rect 9451 2009 9497 2055
rect 9451 1838 9497 1884
rect 9451 1668 9497 1714
rect 9451 1498 9497 1544
rect 9451 1328 9497 1374
rect 9451 1158 9497 1204
rect 9451 988 9497 1034
rect 9451 818 9497 864
rect 9451 648 9497 694
rect 9451 478 9497 524
rect 9451 308 9497 354
rect 10123 4538 10169 4584
rect 10123 4371 10169 4417
rect 10123 4203 10169 4249
rect 10123 4035 10169 4081
rect 10123 3867 10169 3913
rect 10123 3700 10169 3746
rect 10123 3532 10169 3578
rect 10123 3364 10169 3410
rect 10123 3196 10169 3242
rect 10123 3029 10169 3075
rect 10123 2859 10169 2905
rect 10123 2689 10169 2735
rect 10123 2519 10169 2565
rect 10123 2349 10169 2395
rect 10123 2179 10169 2225
rect 10123 2009 10169 2055
rect 10123 1838 10169 1884
rect 10123 1668 10169 1714
rect 10123 1498 10169 1544
rect 10123 1328 10169 1374
rect 10123 1158 10169 1204
rect 10123 988 10169 1034
rect 10123 818 10169 864
rect 10123 648 10169 694
rect 10123 478 10169 524
rect 10650 4022 10696 4068
rect 10650 3854 10696 3900
rect 10650 3686 10696 3732
rect 10650 3518 10696 3564
rect 10650 3351 10696 3397
rect 10650 3183 10696 3229
rect 10650 3015 10696 3061
rect 10650 2847 10696 2893
rect 10650 2680 10696 2726
rect 10650 2512 10696 2558
rect 10650 2344 10696 2390
rect 10650 2174 10696 2220
rect 10650 2004 10696 2050
rect 10650 1834 10696 1880
rect 10650 1664 10696 1710
rect 10650 1494 10696 1540
rect 10650 1324 10696 1370
rect 10650 1154 10696 1200
rect 10650 984 10696 1030
rect 10650 814 10696 860
rect 10650 644 10696 690
rect 11098 4022 11144 4068
rect 11098 3854 11144 3900
rect 11098 3686 11144 3732
rect 11098 3518 11144 3564
rect 11098 3351 11144 3397
rect 11098 3183 11144 3229
rect 11098 3015 11144 3061
rect 11098 2847 11144 2893
rect 11098 2680 11144 2726
rect 11098 2512 11144 2558
rect 11098 2344 11144 2390
rect 11098 2174 11144 2220
rect 11098 2004 11144 2050
rect 11098 1834 11144 1880
rect 11098 1664 11144 1710
rect 11098 1494 11144 1540
rect 11098 1324 11144 1370
rect 11098 1154 11144 1200
rect 11098 984 11144 1030
rect 11098 814 11144 860
rect 11098 644 11144 690
rect 11546 4022 11592 4068
rect 11546 3854 11592 3900
rect 11546 3686 11592 3732
rect 11546 3518 11592 3564
rect 11546 3351 11592 3397
rect 11546 3183 11592 3229
rect 11934 4022 11980 4068
rect 11934 3854 11980 3900
rect 11934 3686 11980 3732
rect 11934 3518 11980 3564
rect 11934 3351 11980 3397
rect 12382 4022 12428 4068
rect 12382 3854 12428 3900
rect 12382 3686 12428 3732
rect 12382 3518 12428 3564
rect 12382 3351 12428 3397
rect 12830 4022 12876 4068
rect 12830 3686 12876 3732
rect 12830 3518 12876 3564
rect 12830 3351 12876 3397
rect 11546 3015 11592 3061
rect 11546 2847 11592 2893
rect 11546 2680 11592 2726
rect 11546 2512 11592 2558
rect 11546 2344 11592 2390
rect 11546 2174 11592 2220
rect 11546 2004 11592 2050
rect 11546 1834 11592 1880
rect 11546 1664 11592 1710
rect 11546 1494 11592 1540
rect 11546 1324 11592 1370
rect 11546 1154 11592 1200
rect 11546 984 11592 1030
rect 11546 814 11592 860
rect 11546 644 11592 690
rect 10123 308 10169 354
<< mvpdiffc >>
rect 4980 6359 5026 6405
rect 4980 6178 5026 6224
rect 5428 6359 5474 6405
rect 5428 6178 5474 6224
<< mvpsubdiff >>
rect 7991 11543 13744 11653
rect 7991 11536 8304 11543
rect 7990 11375 8304 11536
rect 7991 11227 8304 11375
rect 6339 5707 6473 5766
rect 6339 5661 6383 5707
rect 6429 5661 6473 5707
rect 6339 5543 6473 5661
rect 6339 5497 6383 5543
rect 6429 5497 6473 5543
rect 6339 5001 6473 5497
<< mvnsubdiff >>
rect 5994 16273 13722 16319
rect 5994 16227 6192 16273
rect 6238 16227 6350 16273
rect 6396 16227 6508 16273
rect 6554 16227 6666 16273
rect 6712 16227 6824 16273
rect 6870 16227 6982 16273
rect 7028 16227 7140 16273
rect 7186 16227 7298 16273
rect 7344 16227 7457 16273
rect 7503 16227 7615 16273
rect 7661 16227 7773 16273
rect 7819 16227 7931 16273
rect 7977 16227 8089 16273
rect 8135 16227 8247 16273
rect 8293 16227 8405 16273
rect 8451 16227 8563 16273
rect 8609 16227 8721 16273
rect 8767 16227 8880 16273
rect 8926 16227 9038 16273
rect 9084 16227 9196 16273
rect 9242 16227 9354 16273
rect 9400 16227 9512 16273
rect 9558 16227 9670 16273
rect 9716 16227 9828 16273
rect 9874 16227 9986 16273
rect 10032 16227 10144 16273
rect 10190 16227 10303 16273
rect 10349 16227 10461 16273
rect 10507 16227 10619 16273
rect 10665 16227 10777 16273
rect 10823 16227 10935 16273
rect 10981 16227 11093 16273
rect 11139 16227 11251 16273
rect 11297 16227 11409 16273
rect 11455 16227 11567 16273
rect 11613 16227 11726 16273
rect 11772 16227 11884 16273
rect 11930 16227 12042 16273
rect 12088 16227 12200 16273
rect 12246 16227 12358 16273
rect 12404 16227 12516 16273
rect 12562 16227 12674 16273
rect 12720 16227 12832 16273
rect 12878 16227 12990 16273
rect 13036 16227 13149 16273
rect 13195 16227 13307 16273
rect 13353 16227 13465 16273
rect 13511 16227 13722 16273
rect 5994 16181 13722 16227
rect 5994 16092 6128 16181
rect 5994 16046 6038 16092
rect 6084 16046 6128 16092
rect 5994 15928 6128 16046
rect 13588 16092 13722 16181
rect 13588 16046 13632 16092
rect 13678 16046 13722 16092
rect 5994 15882 6038 15928
rect 6084 15882 6128 15928
rect 5994 15765 6128 15882
rect 5994 15719 6038 15765
rect 6084 15719 6128 15765
rect 5994 15602 6128 15719
rect 5994 15556 6038 15602
rect 6084 15556 6128 15602
rect 5994 15439 6128 15556
rect 5994 15393 6038 15439
rect 6084 15393 6128 15439
rect 5994 15275 6128 15393
rect 5994 15229 6038 15275
rect 6084 15229 6128 15275
rect 5994 15112 6128 15229
rect 5994 15066 6038 15112
rect 6084 15066 6128 15112
rect 5994 14949 6128 15066
rect 5994 14903 6038 14949
rect 6084 14903 6128 14949
rect 5994 14786 6128 14903
rect 5994 14740 6038 14786
rect 6084 14740 6128 14786
rect 5994 14622 6128 14740
rect 5994 14576 6038 14622
rect 6084 14576 6128 14622
rect 5994 14459 6128 14576
rect 5994 14413 6038 14459
rect 6084 14413 6128 14459
rect 5994 14296 6128 14413
rect 5994 14250 6038 14296
rect 6084 14250 6128 14296
rect 5994 14133 6128 14250
rect 5994 14087 6038 14133
rect 6084 14087 6128 14133
rect 5994 13970 6128 14087
rect 5994 13924 6038 13970
rect 6084 13924 6128 13970
rect 5994 13806 6128 13924
rect 5994 13760 6038 13806
rect 6084 13760 6128 13806
rect 5994 13643 6128 13760
rect 5994 13597 6038 13643
rect 6084 13597 6128 13643
rect 5994 13480 6128 13597
rect 5994 13434 6038 13480
rect 6084 13434 6128 13480
rect 13588 15928 13722 16046
rect 13588 15882 13632 15928
rect 13678 15882 13722 15928
rect 13588 15765 13722 15882
rect 13588 15719 13632 15765
rect 13678 15719 13722 15765
rect 13588 15602 13722 15719
rect 13588 15556 13632 15602
rect 13678 15556 13722 15602
rect 13588 15439 13722 15556
rect 13588 15393 13632 15439
rect 13678 15393 13722 15439
rect 13588 15275 13722 15393
rect 13588 15229 13632 15275
rect 13678 15229 13722 15275
rect 13588 15112 13722 15229
rect 13588 15066 13632 15112
rect 13678 15066 13722 15112
rect 13588 14949 13722 15066
rect 13588 14903 13632 14949
rect 13678 14903 13722 14949
rect 13588 14786 13722 14903
rect 13588 14740 13632 14786
rect 13678 14740 13722 14786
rect 13588 14622 13722 14740
rect 13588 14576 13632 14622
rect 13678 14576 13722 14622
rect 13588 14459 13722 14576
rect 13588 14413 13632 14459
rect 13678 14413 13722 14459
rect 13588 14296 13722 14413
rect 13588 14250 13632 14296
rect 13678 14250 13722 14296
rect 13588 14133 13722 14250
rect 13588 14087 13632 14133
rect 13678 14087 13722 14133
rect 13588 13970 13722 14087
rect 13588 13924 13632 13970
rect 13678 13924 13722 13970
rect 13588 13806 13722 13924
rect 13588 13760 13632 13806
rect 13678 13760 13722 13806
rect 13588 13643 13722 13760
rect 13588 13597 13632 13643
rect 13678 13597 13722 13643
rect 13588 13480 13722 13597
rect 5994 13317 6128 13434
rect 13588 13434 13632 13480
rect 13678 13434 13722 13480
rect 13588 13317 13722 13434
rect 5994 13271 6038 13317
rect 6084 13271 6128 13317
rect 5994 13161 6128 13271
rect 13588 13271 13632 13317
rect 13678 13271 13722 13317
rect 5994 13153 8664 13161
rect 5994 13107 6038 13153
rect 6084 13107 8664 13153
rect 5994 12990 8664 13107
rect 5994 12944 6038 12990
rect 6084 12944 8664 12990
rect 5994 12827 8664 12944
rect 5994 12781 6038 12827
rect 6084 12781 8664 12827
rect 5994 12664 8664 12781
rect 5994 12618 6038 12664
rect 6084 12618 8664 12664
rect 5994 12501 8664 12618
rect 5994 12455 6038 12501
rect 6084 12455 8664 12501
rect 5994 12337 8664 12455
rect 5994 12291 6038 12337
rect 6084 12291 8664 12337
rect 5994 12174 8664 12291
rect 13588 13153 13722 13271
rect 13588 13107 13632 13153
rect 13678 13107 13722 13153
rect 13588 12990 13722 13107
rect 13588 12944 13632 12990
rect 13678 12944 13722 12990
rect 13588 12827 13722 12944
rect 13588 12781 13632 12827
rect 13678 12781 13722 12827
rect 13588 12664 13722 12781
rect 13588 12618 13632 12664
rect 13678 12618 13722 12664
rect 13588 12501 13722 12618
rect 13588 12455 13632 12501
rect 13678 12455 13722 12501
rect 13588 12337 13722 12455
rect 13588 12291 13632 12337
rect 13678 12291 13722 12337
rect 5994 12128 6038 12174
rect 6084 12128 8664 12174
rect 13588 12174 13722 12291
rect 5994 12011 8664 12128
rect 5994 11965 6038 12011
rect 6084 12007 8664 12011
rect 13588 12128 13632 12174
rect 13678 12128 13722 12174
rect 13588 12011 13722 12128
rect 13588 12007 13632 12011
rect 6084 11965 13632 12007
rect 13678 11965 13722 12011
rect 5994 11961 13722 11965
rect 5994 11915 6192 11961
rect 6238 11915 6350 11961
rect 6396 11915 6508 11961
rect 6554 11915 6666 11961
rect 6712 11915 6824 11961
rect 6870 11915 6982 11961
rect 7028 11915 7140 11961
rect 7186 11915 7298 11961
rect 7344 11915 7457 11961
rect 7503 11915 7615 11961
rect 7661 11915 7773 11961
rect 7819 11915 7931 11961
rect 7977 11915 8089 11961
rect 8135 11915 8247 11961
rect 8293 11915 8405 11961
rect 8451 11915 8563 11961
rect 8609 11915 8721 11961
rect 8767 11915 8880 11961
rect 8926 11915 9038 11961
rect 9084 11915 9196 11961
rect 9242 11915 9354 11961
rect 9400 11915 9512 11961
rect 9558 11915 9670 11961
rect 9716 11915 9828 11961
rect 9874 11915 9986 11961
rect 10032 11915 10144 11961
rect 10190 11915 10303 11961
rect 10349 11915 10461 11961
rect 10507 11915 10619 11961
rect 10665 11915 10777 11961
rect 10823 11915 10935 11961
rect 10981 11915 11093 11961
rect 11139 11915 11251 11961
rect 11297 11915 11409 11961
rect 11455 11915 11567 11961
rect 11613 11915 11726 11961
rect 11772 11915 11884 11961
rect 11930 11915 12042 11961
rect 12088 11915 12200 11961
rect 12246 11915 12358 11961
rect 12404 11915 12516 11961
rect 12562 11915 12674 11961
rect 12720 11915 12832 11961
rect 12878 11915 12990 11961
rect 13036 11915 13149 11961
rect 13195 11915 13307 11961
rect 13353 11915 13465 11961
rect 13511 11915 13722 11961
rect 5994 11869 13722 11915
rect 6339 6969 6473 7045
rect 6339 6923 6383 6969
rect 6429 6923 6473 6969
rect 6339 6777 6473 6923
rect 6339 6731 6383 6777
rect 6429 6731 6473 6777
rect 6339 6584 6473 6731
rect 6339 6538 6383 6584
rect 6429 6538 6473 6584
rect 6339 6421 6473 6538
rect 6339 6375 6383 6421
rect 6429 6375 6473 6421
rect 6339 6213 6473 6375
<< mvpsubdiffcont >>
rect 6383 5661 6429 5707
rect 6383 5497 6429 5543
<< mvnsubdiffcont >>
rect 6192 16227 6238 16273
rect 6350 16227 6396 16273
rect 6508 16227 6554 16273
rect 6666 16227 6712 16273
rect 6824 16227 6870 16273
rect 6982 16227 7028 16273
rect 7140 16227 7186 16273
rect 7298 16227 7344 16273
rect 7457 16227 7503 16273
rect 7615 16227 7661 16273
rect 7773 16227 7819 16273
rect 7931 16227 7977 16273
rect 8089 16227 8135 16273
rect 8247 16227 8293 16273
rect 8405 16227 8451 16273
rect 8563 16227 8609 16273
rect 8721 16227 8767 16273
rect 8880 16227 8926 16273
rect 9038 16227 9084 16273
rect 9196 16227 9242 16273
rect 9354 16227 9400 16273
rect 9512 16227 9558 16273
rect 9670 16227 9716 16273
rect 9828 16227 9874 16273
rect 9986 16227 10032 16273
rect 10144 16227 10190 16273
rect 10303 16227 10349 16273
rect 10461 16227 10507 16273
rect 10619 16227 10665 16273
rect 10777 16227 10823 16273
rect 10935 16227 10981 16273
rect 11093 16227 11139 16273
rect 11251 16227 11297 16273
rect 11409 16227 11455 16273
rect 11567 16227 11613 16273
rect 11726 16227 11772 16273
rect 11884 16227 11930 16273
rect 12042 16227 12088 16273
rect 12200 16227 12246 16273
rect 12358 16227 12404 16273
rect 12516 16227 12562 16273
rect 12674 16227 12720 16273
rect 12832 16227 12878 16273
rect 12990 16227 13036 16273
rect 13149 16227 13195 16273
rect 13307 16227 13353 16273
rect 13465 16227 13511 16273
rect 6038 16046 6084 16092
rect 13632 16046 13678 16092
rect 6038 15882 6084 15928
rect 6038 15719 6084 15765
rect 6038 15556 6084 15602
rect 6038 15393 6084 15439
rect 6038 15229 6084 15275
rect 6038 15066 6084 15112
rect 6038 14903 6084 14949
rect 6038 14740 6084 14786
rect 6038 14576 6084 14622
rect 6038 14413 6084 14459
rect 6038 14250 6084 14296
rect 6038 14087 6084 14133
rect 6038 13924 6084 13970
rect 6038 13760 6084 13806
rect 6038 13597 6084 13643
rect 6038 13434 6084 13480
rect 13632 15882 13678 15928
rect 13632 15719 13678 15765
rect 13632 15556 13678 15602
rect 13632 15393 13678 15439
rect 13632 15229 13678 15275
rect 13632 15066 13678 15112
rect 13632 14903 13678 14949
rect 13632 14740 13678 14786
rect 13632 14576 13678 14622
rect 13632 14413 13678 14459
rect 13632 14250 13678 14296
rect 13632 14087 13678 14133
rect 13632 13924 13678 13970
rect 13632 13760 13678 13806
rect 13632 13597 13678 13643
rect 13632 13434 13678 13480
rect 6038 13271 6084 13317
rect 13632 13271 13678 13317
rect 6038 13107 6084 13153
rect 6038 12944 6084 12990
rect 6038 12781 6084 12827
rect 6038 12618 6084 12664
rect 6038 12455 6084 12501
rect 6038 12291 6084 12337
rect 13632 13107 13678 13153
rect 13632 12944 13678 12990
rect 13632 12781 13678 12827
rect 13632 12618 13678 12664
rect 13632 12455 13678 12501
rect 13632 12291 13678 12337
rect 6038 12128 6084 12174
rect 6038 11965 6084 12011
rect 13632 12128 13678 12174
rect 13632 11965 13678 12011
rect 6192 11915 6238 11961
rect 6350 11915 6396 11961
rect 6508 11915 6554 11961
rect 6666 11915 6712 11961
rect 6824 11915 6870 11961
rect 6982 11915 7028 11961
rect 7140 11915 7186 11961
rect 7298 11915 7344 11961
rect 7457 11915 7503 11961
rect 7615 11915 7661 11961
rect 7773 11915 7819 11961
rect 7931 11915 7977 11961
rect 8089 11915 8135 11961
rect 8247 11915 8293 11961
rect 8405 11915 8451 11961
rect 8563 11915 8609 11961
rect 8721 11915 8767 11961
rect 8880 11915 8926 11961
rect 9038 11915 9084 11961
rect 9196 11915 9242 11961
rect 9354 11915 9400 11961
rect 9512 11915 9558 11961
rect 9670 11915 9716 11961
rect 9828 11915 9874 11961
rect 9986 11915 10032 11961
rect 10144 11915 10190 11961
rect 10303 11915 10349 11961
rect 10461 11915 10507 11961
rect 10619 11915 10665 11961
rect 10777 11915 10823 11961
rect 10935 11915 10981 11961
rect 11093 11915 11139 11961
rect 11251 11915 11297 11961
rect 11409 11915 11455 11961
rect 11567 11915 11613 11961
rect 11726 11915 11772 11961
rect 11884 11915 11930 11961
rect 12042 11915 12088 11961
rect 12200 11915 12246 11961
rect 12358 11915 12404 11961
rect 12516 11915 12562 11961
rect 12674 11915 12720 11961
rect 12832 11915 12878 11961
rect 12990 11915 13036 11961
rect 13149 11915 13195 11961
rect 13307 11915 13353 11961
rect 13465 11915 13511 11961
rect 6383 6923 6429 6969
rect 6383 6731 6429 6777
rect 6383 6538 6429 6584
rect 6383 6375 6429 6421
<< polysilicon >>
rect 6408 15956 6527 16028
rect 6632 15956 6751 16028
rect 6856 15956 6975 16028
rect 7080 15956 7199 16028
rect 7304 15956 7423 16028
rect 7528 15956 7647 16028
rect 7752 15956 7871 16028
rect 7976 15956 8095 16028
rect 8200 15956 8319 16028
rect 8424 15956 8543 16028
rect 6408 13317 6528 13461
rect 6632 13317 6752 13461
rect 6856 13317 6976 13461
rect 7080 13317 7200 13461
rect 7304 13317 7424 13461
rect 7528 13317 7648 13461
rect 7752 13317 7872 13461
rect 7976 13317 8096 13461
rect 8200 13317 8320 13461
rect 8424 13317 8544 13461
rect 8937 12223 9057 12282
rect 9161 12223 9281 12276
rect 9385 12223 9505 12276
rect 9609 12223 9729 12276
rect 9833 12223 9953 12276
rect 10057 12223 10177 12276
rect 10281 12223 10401 12276
rect 10505 12223 10625 12276
rect 10729 12223 10849 12276
rect 10953 12223 11073 12276
rect 11177 12223 11297 12276
rect 11401 12223 11521 12276
rect 11625 12223 11745 12276
rect 11849 12223 11969 12276
rect 12073 12223 12193 12276
rect 12297 12223 12417 12276
rect 12521 12223 12641 12276
rect 12745 12223 12865 12276
rect 12969 12223 13089 12276
rect 13193 12223 13313 12276
rect 8937 12139 13313 12223
rect 8937 11302 9057 11389
rect 9161 11302 9281 11389
rect 9385 11302 9505 11389
rect 9609 11302 9729 11389
rect 9833 11302 9953 11389
rect 10057 11302 10177 11389
rect 10281 11302 10401 11389
rect 10505 11302 10625 11389
rect 10729 11302 10849 11389
rect 10953 11302 11073 11389
rect 11177 11302 11297 11389
rect 11401 11302 11521 11389
rect 11625 11302 11745 11389
rect 11849 11302 11969 11389
rect 12073 11302 12193 11389
rect 12297 11302 12417 11389
rect 12521 11302 12641 11389
rect 12745 11302 12865 11389
rect 12969 11302 13089 11389
rect 13193 11302 13313 11389
rect 6700 11033 6820 11179
rect 6924 11033 7044 11179
rect 7148 11033 7268 11179
rect 7372 11033 7492 11179
rect 7596 11033 7716 11179
rect 5055 7680 5174 7911
rect 6972 7761 7092 7981
rect 7486 7961 7606 7993
rect 7755 7985 7947 8031
rect 7755 7961 7828 7985
rect 7486 7939 7828 7961
rect 7874 7939 7947 7985
rect 7486 7896 7947 7939
rect 7755 7821 7947 7896
rect 7755 7775 7828 7821
rect 7874 7775 7947 7821
rect 7755 7729 7947 7775
rect 7486 7477 7606 7509
rect 6166 7394 7092 7454
rect 7486 7432 7723 7477
rect 6166 7393 6519 7394
rect 6166 7391 6518 7393
rect 6166 7345 6240 7391
rect 6286 7345 6398 7391
rect 6444 7345 6518 7391
rect 6166 7299 6518 7345
rect 7486 7386 7604 7432
rect 7650 7386 7723 7432
rect 7486 7340 7723 7386
rect 5055 7123 5175 7151
rect 5055 7078 5376 7123
rect 5055 7032 5256 7078
rect 5302 7032 5376 7078
rect 5055 6986 5376 7032
rect 7791 6978 7911 7729
rect 7486 6891 7911 6978
rect 5055 6587 5174 6659
rect 5279 6587 5398 6659
rect 5055 6069 5174 6131
rect 4981 6024 5174 6069
rect 4981 5978 5054 6024
rect 5100 5978 5174 6024
rect 4981 5932 5174 5978
rect 5055 5718 5174 5932
rect 5279 5857 5398 6131
rect 6748 6063 6868 6136
rect 6972 6063 7092 6136
rect 6748 6017 7254 6063
rect 6748 5971 7134 6017
rect 7180 5971 7254 6017
rect 7719 6033 7912 6078
rect 7719 6002 7793 6033
rect 6748 5925 7254 5971
rect 7486 5987 7793 6002
rect 7839 5987 7912 6033
rect 7486 5941 7912 5987
rect 6748 5886 6868 5925
rect 6972 5886 7092 5925
rect 5279 5811 5867 5857
rect 7486 5855 7606 5941
rect 5279 5765 5788 5811
rect 5834 5765 5867 5811
rect 5279 5734 5867 5765
rect 5279 5718 5399 5734
rect 9526 5095 9646 5263
rect 9526 4955 9568 5095
rect 9614 4955 9646 5095
rect 9526 4798 9646 4955
rect 9750 5095 9870 5263
rect 9750 4955 9791 5095
rect 9837 4955 9870 5095
rect 9750 4798 9870 4955
rect 9974 5095 10094 5263
rect 9974 4955 10015 5095
rect 10061 4955 10094 5095
rect 9974 4798 10094 4955
rect 6467 3790 6469 3823
rect 5157 3603 5397 3762
rect 5157 3557 5623 3603
rect 6235 3602 6475 3762
rect 6954 3602 7154 3797
rect 7600 3760 7719 3790
rect 7600 3602 7720 3760
rect 8114 3603 8234 3760
rect 8114 3602 8458 3603
rect 5157 3511 5345 3557
rect 5391 3511 5503 3557
rect 5549 3511 5623 3557
rect 5157 3465 5623 3511
rect 6109 3557 6475 3602
rect 6109 3511 6183 3557
rect 6229 3511 6475 3557
rect 6109 3465 6475 3511
rect 6833 3557 7154 3602
rect 6833 3511 6907 3557
rect 6953 3511 7154 3557
rect 6833 3465 7154 3511
rect 7473 3557 7720 3602
rect 7473 3511 7547 3557
rect 7593 3511 7720 3557
rect 7473 3465 7720 3511
rect 7991 3557 8458 3602
rect 7991 3511 8065 3557
rect 8111 3511 8458 3557
rect 7991 3465 8458 3511
rect 5157 3261 5397 3465
rect 6235 3261 6475 3465
rect 6954 3291 7154 3465
rect 7600 3291 7720 3465
rect 8114 3291 8234 3465
rect 8338 3291 8458 3465
rect 7600 3261 7719 3291
rect 7600 2810 7719 2883
rect 10725 4537 10845 4628
rect 10725 4491 10763 4537
rect 10809 4491 10845 4537
rect 10725 4113 10845 4491
rect 10949 4338 11069 4628
rect 11173 4338 11293 4628
rect 10949 4319 11293 4338
rect 10949 4273 11049 4319
rect 11189 4273 11293 4319
rect 10949 4254 11293 4273
rect 10949 4113 11069 4254
rect 11173 4113 11293 4254
rect 11397 4537 11517 4628
rect 11397 4491 11434 4537
rect 11480 4491 11517 4537
rect 11397 4113 11517 4491
rect 12010 4288 12130 4628
rect 12234 4525 12354 4628
rect 12458 4525 12578 4628
rect 12010 4242 12046 4288
rect 12092 4242 12130 4288
rect 12010 4113 12130 4242
rect 12233 4506 12578 4525
rect 12233 4460 12294 4506
rect 12528 4460 12578 4506
rect 12233 4441 12578 4460
rect 12233 4113 12353 4441
rect 12458 4113 12578 4441
rect 12682 4307 12802 4628
rect 12681 4288 12802 4307
rect 12681 4242 12718 4288
rect 12764 4242 12802 4288
rect 12681 4223 12802 4242
rect 12681 4113 12801 4223
rect 12010 3132 12130 3205
rect 12233 3132 12353 3205
rect 12458 3132 12578 3205
rect 12681 3132 12801 3205
rect 10725 412 10845 484
rect 10949 412 11069 484
rect 11173 412 11293 484
rect 11397 412 11517 484
rect 9526 190 9646 262
rect 9750 190 9870 262
rect 9974 190 10094 262
<< polycontact >>
rect 7828 7939 7874 7985
rect 7828 7775 7874 7821
rect 6240 7345 6286 7391
rect 6398 7345 6444 7391
rect 7604 7386 7650 7432
rect 5256 7032 5302 7078
rect 5054 5978 5100 6024
rect 7134 5971 7180 6017
rect 7793 5987 7839 6033
rect 5788 5765 5834 5811
rect 9568 4955 9614 5095
rect 9791 4955 9837 5095
rect 10015 4955 10061 5095
rect 5345 3511 5391 3557
rect 5503 3511 5549 3557
rect 6183 3511 6229 3557
rect 6907 3511 6953 3557
rect 7547 3511 7593 3557
rect 8065 3511 8111 3557
rect 10763 4491 10809 4537
rect 11049 4273 11189 4319
rect 11434 4491 11480 4537
rect 12046 4242 12092 4288
rect 12294 4460 12528 4506
rect 12718 4242 12764 4288
<< metal1 >>
rect 6003 16273 13713 16310
rect 6003 16227 6192 16273
rect 6238 16227 6350 16273
rect 6396 16227 6508 16273
rect 6554 16227 6666 16273
rect 6712 16227 6824 16273
rect 6870 16227 6982 16273
rect 7028 16227 7140 16273
rect 7186 16227 7298 16273
rect 7344 16227 7457 16273
rect 7503 16227 7615 16273
rect 7661 16227 7773 16273
rect 7819 16227 7931 16273
rect 7977 16227 8089 16273
rect 8135 16227 8247 16273
rect 8293 16227 8405 16273
rect 8451 16227 8563 16273
rect 8609 16227 8721 16273
rect 8767 16227 8880 16273
rect 8926 16227 9038 16273
rect 9084 16227 9196 16273
rect 9242 16227 9354 16273
rect 9400 16227 9512 16273
rect 9558 16227 9670 16273
rect 9716 16227 9828 16273
rect 9874 16227 9986 16273
rect 10032 16227 10144 16273
rect 10190 16227 10303 16273
rect 10349 16227 10461 16273
rect 10507 16227 10619 16273
rect 10665 16227 10777 16273
rect 10823 16227 10935 16273
rect 10981 16227 11093 16273
rect 11139 16227 11251 16273
rect 11297 16227 11409 16273
rect 11455 16227 11567 16273
rect 11613 16227 11726 16273
rect 11772 16227 11884 16273
rect 11930 16227 12042 16273
rect 12088 16227 12200 16273
rect 12246 16227 12358 16273
rect 12404 16227 12516 16273
rect 12562 16227 12674 16273
rect 12720 16227 12832 16273
rect 12878 16227 12990 16273
rect 13036 16227 13149 16273
rect 13195 16227 13307 16273
rect 13353 16227 13465 16273
rect 13511 16227 13713 16273
rect 6003 16190 13713 16227
rect 6003 16092 6413 16190
rect 6003 16046 6038 16092
rect 6084 16046 6413 16092
rect 6003 15928 6413 16046
rect 6003 15882 6038 15928
rect 6084 15882 6413 15928
rect 6003 15765 6413 15882
rect 6003 15719 6038 15765
rect 6084 15719 6413 15765
rect 6003 15602 6413 15719
rect 6003 15556 6038 15602
rect 6084 15556 6413 15602
rect 6003 15439 6413 15556
rect 6003 15393 6038 15439
rect 6084 15393 6413 15439
rect 6003 15275 6413 15393
rect 6003 15229 6038 15275
rect 6084 15229 6413 15275
rect 6003 15112 6413 15229
rect 6003 15066 6038 15112
rect 6084 15066 6413 15112
rect 6003 14949 6413 15066
rect 6003 14903 6038 14949
rect 6084 14903 6413 14949
rect 6003 14786 6413 14903
rect 6003 14740 6038 14786
rect 6084 14740 6413 14786
rect 6003 14622 6413 14740
rect 6003 14576 6038 14622
rect 6084 14576 6413 14622
rect 6003 14459 6413 14576
rect 13301 16092 13713 16190
rect 13301 16046 13632 16092
rect 13678 16046 13713 16092
rect 13301 15928 13713 16046
rect 13301 15882 13632 15928
rect 13678 15882 13713 15928
rect 13301 15765 13713 15882
rect 13301 15719 13632 15765
rect 13678 15719 13713 15765
rect 13301 15602 13713 15719
rect 13301 15556 13632 15602
rect 13678 15556 13713 15602
rect 13301 15439 13713 15556
rect 13301 15393 13632 15439
rect 13678 15393 13713 15439
rect 13301 15275 13713 15393
rect 13301 15229 13632 15275
rect 13678 15229 13713 15275
rect 13301 15112 13713 15229
rect 13301 15066 13632 15112
rect 13678 15066 13713 15112
rect 13301 14949 13713 15066
rect 13301 14903 13632 14949
rect 13678 14903 13713 14949
rect 13301 14786 13713 14903
rect 13301 14740 13632 14786
rect 13678 14740 13713 14786
rect 13301 14622 13713 14740
rect 13301 14576 13632 14622
rect 13678 14576 13713 14622
rect 6003 14413 6038 14459
rect 6084 14413 6413 14459
rect 6003 14296 6413 14413
rect 6003 14250 6038 14296
rect 6084 14250 6413 14296
rect 6003 14133 6413 14250
rect 6003 14087 6038 14133
rect 6084 14087 6413 14133
rect 6003 13970 6413 14087
rect 6003 13924 6038 13970
rect 6084 13924 6413 13970
rect 6003 13806 6413 13924
rect 6003 13760 6038 13806
rect 6084 13760 6413 13806
rect 6003 13643 6413 13760
rect 6003 13597 6038 13643
rect 6084 13597 6413 13643
rect 6003 13480 6413 13597
rect 6003 13434 6038 13480
rect 6084 13470 6413 13480
rect 6513 14433 6640 14474
rect 6513 14381 6551 14433
rect 6603 14381 6640 14433
rect 6513 14216 6640 14381
rect 6513 14164 6551 14216
rect 6603 14164 6640 14216
rect 6513 13998 6640 14164
rect 6513 13946 6551 13998
rect 6603 13946 6640 13998
rect 6513 13780 6640 13946
rect 6513 13728 6551 13780
rect 6603 13728 6640 13780
rect 6513 13563 6640 13728
rect 6513 13511 6551 13563
rect 6603 13511 6640 13563
rect 6513 13470 6640 13511
rect 6961 14433 7088 14474
rect 6961 14381 6999 14433
rect 7051 14381 7088 14433
rect 6961 14216 7088 14381
rect 6961 14164 6999 14216
rect 7051 14164 7088 14216
rect 6961 13998 7088 14164
rect 6961 13946 6999 13998
rect 7051 13946 7088 13998
rect 6961 13780 7088 13946
rect 6961 13728 6999 13780
rect 7051 13728 7088 13780
rect 6961 13563 7088 13728
rect 6961 13511 6999 13563
rect 7051 13511 7088 13563
rect 6961 13470 7088 13511
rect 7409 14433 7536 14474
rect 7409 14381 7447 14433
rect 7499 14381 7536 14433
rect 7409 14216 7536 14381
rect 7409 14164 7447 14216
rect 7499 14164 7536 14216
rect 7409 13998 7536 14164
rect 7409 13946 7447 13998
rect 7499 13946 7536 13998
rect 7409 13780 7536 13946
rect 7409 13728 7447 13780
rect 7499 13728 7536 13780
rect 7409 13563 7536 13728
rect 7409 13511 7447 13563
rect 7499 13511 7536 13563
rect 7409 13470 7536 13511
rect 7857 14433 7984 14474
rect 7857 14381 7895 14433
rect 7947 14381 7984 14433
rect 7857 14216 7984 14381
rect 7857 14164 7895 14216
rect 7947 14164 7984 14216
rect 7857 13998 7984 14164
rect 7857 13946 7895 13998
rect 7947 13946 7984 13998
rect 7857 13780 7984 13946
rect 7857 13728 7895 13780
rect 7947 13728 7984 13780
rect 7857 13563 7984 13728
rect 7857 13511 7895 13563
rect 7947 13511 7984 13563
rect 7857 13470 7984 13511
rect 8305 14433 8432 14474
rect 8305 14381 8343 14433
rect 8395 14381 8432 14433
rect 8305 14216 8432 14381
rect 8305 14164 8343 14216
rect 8395 14164 8432 14216
rect 8305 13998 8432 14164
rect 8305 13946 8343 13998
rect 8395 13946 8432 13998
rect 8305 13780 8432 13946
rect 8305 13728 8343 13780
rect 8395 13728 8432 13780
rect 8305 13563 8432 13728
rect 8305 13511 8343 13563
rect 8395 13511 8432 13563
rect 8305 13470 8432 13511
rect 13301 14459 13713 14576
rect 13301 14413 13632 14459
rect 13678 14413 13713 14459
rect 13301 14296 13713 14413
rect 13301 14250 13632 14296
rect 13678 14250 13713 14296
rect 13301 14133 13713 14250
rect 13301 14087 13632 14133
rect 13678 14087 13713 14133
rect 13301 13970 13713 14087
rect 13301 13924 13632 13970
rect 13678 13924 13713 13970
rect 13301 13806 13713 13924
rect 13301 13760 13632 13806
rect 13678 13760 13713 13806
rect 13301 13643 13713 13760
rect 13301 13597 13632 13643
rect 13678 13597 13713 13643
rect 13301 13480 13713 13597
rect 6084 13434 6119 13470
rect 6003 13317 6119 13434
rect 13301 13434 13632 13480
rect 13678 13434 13713 13480
rect 6003 13271 6038 13317
rect 6084 13271 6119 13317
rect 6003 13153 6119 13271
rect 6539 13336 7301 13376
rect 6539 13284 6577 13336
rect 6629 13284 6788 13336
rect 6840 13284 7000 13336
rect 7052 13284 7211 13336
rect 7263 13284 7301 13336
rect 6539 13243 7301 13284
rect 13301 13317 13713 13434
rect 13301 13271 13632 13317
rect 13678 13271 13713 13317
rect 6003 13107 6038 13153
rect 6084 13141 6119 13153
rect 13301 13153 13713 13271
rect 6084 13107 8645 13141
rect 6003 12990 8645 13107
rect 6003 12944 6038 12990
rect 6084 12944 8645 12990
rect 6003 12827 8645 12944
rect 6003 12781 6038 12827
rect 6084 12781 8645 12827
rect 6003 12664 8645 12781
rect 6003 12618 6038 12664
rect 6084 12618 8645 12664
rect 6003 12501 8645 12618
rect 6003 12455 6038 12501
rect 6084 12455 8645 12501
rect 6003 12337 8645 12455
rect 6003 12291 6038 12337
rect 6084 12291 8645 12337
rect 13301 13107 13632 13153
rect 13678 13107 13713 13153
rect 13301 12990 13713 13107
rect 13301 12944 13632 12990
rect 13678 12944 13713 12990
rect 13301 12827 13713 12944
rect 13301 12781 13632 12827
rect 13678 12781 13713 12827
rect 13301 12664 13713 12781
rect 13301 12618 13632 12664
rect 13678 12618 13713 12664
rect 13301 12501 13713 12618
rect 13301 12455 13632 12501
rect 13678 12455 13713 12501
rect 13301 12337 13713 12455
rect 13301 12291 13632 12337
rect 13678 12291 13713 12337
rect 6003 12174 8645 12291
rect 6003 12128 6038 12174
rect 6084 12128 8645 12174
rect 6003 12011 8645 12128
rect 6003 11965 6038 12011
rect 6084 11998 8645 12011
rect 13597 12174 13713 12291
rect 13597 12128 13632 12174
rect 13678 12128 13713 12174
rect 13597 12011 13713 12128
rect 13597 11998 13632 12011
rect 6084 11965 13632 11998
rect 13678 11965 13713 12011
rect 6003 11961 13713 11965
rect 6003 11915 6192 11961
rect 6238 11915 6350 11961
rect 6396 11915 6508 11961
rect 6554 11915 6666 11961
rect 6712 11915 6824 11961
rect 6870 11915 6982 11961
rect 7028 11915 7140 11961
rect 7186 11915 7298 11961
rect 7344 11915 7457 11961
rect 7503 11915 7615 11961
rect 7661 11915 7773 11961
rect 7819 11915 7931 11961
rect 7977 11915 8089 11961
rect 8135 11915 8247 11961
rect 8293 11915 8405 11961
rect 8451 11915 8563 11961
rect 8609 11915 8721 11961
rect 8767 11915 8880 11961
rect 8926 11915 9038 11961
rect 9084 11915 9196 11961
rect 9242 11915 9354 11961
rect 9400 11915 9512 11961
rect 9558 11915 9670 11961
rect 9716 11915 9828 11961
rect 9874 11915 9986 11961
rect 10032 11915 10144 11961
rect 10190 11915 10303 11961
rect 10349 11915 10461 11961
rect 10507 11915 10619 11961
rect 10665 11915 10777 11961
rect 10823 11915 10935 11961
rect 10981 11915 11093 11961
rect 11139 11915 11251 11961
rect 11297 11915 11409 11961
rect 11455 11915 11567 11961
rect 11613 11915 11726 11961
rect 11772 11915 11884 11961
rect 11930 11915 12042 11961
rect 12088 11915 12200 11961
rect 12246 11915 12358 11961
rect 12404 11915 12516 11961
rect 12562 11915 12674 11961
rect 12720 11915 12832 11961
rect 12878 11915 12990 11961
rect 13036 11915 13149 11961
rect 13195 11915 13307 11961
rect 13353 11915 13465 11961
rect 13511 11915 13713 11961
rect 6003 11878 13713 11915
rect 6283 11333 6397 11334
rect 6276 11332 6401 11333
rect 6276 11293 6404 11332
rect 6276 11241 6314 11293
rect 6366 11241 6404 11293
rect 6276 11075 6404 11241
rect 6569 11200 7331 11240
rect 8010 11227 8284 11515
rect 6569 11148 6607 11200
rect 6659 11148 6818 11200
rect 6870 11148 7030 11200
rect 7082 11148 7241 11200
rect 7293 11148 7331 11200
rect 6569 11107 7331 11148
rect 9045 11195 9173 11236
rect 9045 11143 9083 11195
rect 9135 11143 9173 11195
rect 6276 11023 6314 11075
rect 6366 11025 6404 11075
rect 6366 11023 6705 11025
rect 6276 10858 6705 11023
rect 9045 10978 9173 11143
rect 6815 10955 6929 10956
rect 7262 10955 7376 10956
rect 7710 10955 7824 10956
rect 6276 10806 6314 10858
rect 6366 10806 6705 10858
rect 6276 10640 6705 10806
rect 6276 10588 6314 10640
rect 6366 10588 6705 10640
rect 6276 10422 6705 10588
rect 6276 10370 6314 10422
rect 6366 10370 6705 10422
rect 6276 10205 6705 10370
rect 6276 10153 6314 10205
rect 6366 10153 6705 10205
rect 6276 9987 6705 10153
rect 6276 9935 6314 9987
rect 6366 9935 6705 9987
rect 6276 9895 6705 9935
rect 6289 9047 6705 9895
rect 6808 10954 6933 10955
rect 7255 10954 7380 10955
rect 7703 10954 7828 10955
rect 6808 10915 6936 10954
rect 6808 10863 6846 10915
rect 6898 10863 6936 10915
rect 6808 10697 6936 10863
rect 6808 10645 6846 10697
rect 6898 10645 6936 10697
rect 6808 10480 6936 10645
rect 6808 10428 6846 10480
rect 6898 10428 6936 10480
rect 6808 10262 6936 10428
rect 7255 10915 7383 10954
rect 7255 10863 7293 10915
rect 7345 10863 7383 10915
rect 7255 10697 7383 10863
rect 7255 10645 7293 10697
rect 7345 10645 7383 10697
rect 7255 10480 7383 10645
rect 7255 10428 7293 10480
rect 7345 10428 7383 10480
rect 6808 10210 6846 10262
rect 6898 10210 6936 10262
rect 6808 10044 6936 10210
rect 6808 9992 6846 10044
rect 6898 9992 6936 10044
rect 6808 9827 6936 9992
rect 6808 9775 6846 9827
rect 6898 9775 6936 9827
rect 6808 9609 6936 9775
rect 6808 9557 6846 9609
rect 6898 9557 6936 9609
rect 6808 9517 6936 9557
rect 6821 9516 6936 9517
rect 7032 10262 7160 10302
rect 7032 10210 7070 10262
rect 7122 10210 7160 10262
rect 7032 10044 7160 10210
rect 7032 9992 7070 10044
rect 7122 9992 7160 10044
rect 7032 9826 7160 9992
rect 7032 9774 7070 9826
rect 7122 9774 7160 9826
rect 7032 9608 7160 9774
rect 7032 9556 7070 9608
rect 7122 9556 7160 9608
rect 7032 9516 7160 9556
rect 7255 10262 7383 10428
rect 7703 10915 7831 10954
rect 7703 10863 7741 10915
rect 7793 10863 7831 10915
rect 7703 10697 7831 10863
rect 7703 10645 7741 10697
rect 7793 10645 7831 10697
rect 7703 10480 7831 10645
rect 9045 10926 9083 10978
rect 9135 10926 9173 10978
rect 9045 10760 9173 10926
rect 9045 10708 9083 10760
rect 9135 10708 9173 10760
rect 7703 10428 7741 10480
rect 7793 10428 7831 10480
rect 7255 10210 7293 10262
rect 7345 10210 7383 10262
rect 7255 10044 7383 10210
rect 7255 9992 7293 10044
rect 7345 9992 7383 10044
rect 7255 9827 7383 9992
rect 7255 9775 7293 9827
rect 7345 9775 7383 9827
rect 7255 9609 7383 9775
rect 7255 9557 7293 9609
rect 7345 9557 7383 9609
rect 7255 9517 7383 9557
rect 7268 9516 7383 9517
rect 7479 10262 7607 10302
rect 7479 10210 7517 10262
rect 7569 10210 7607 10262
rect 7479 10044 7607 10210
rect 7479 9992 7517 10044
rect 7569 9992 7607 10044
rect 7479 9826 7607 9992
rect 7479 9774 7517 9826
rect 7569 9774 7607 9826
rect 7479 9608 7607 9774
rect 7479 9556 7517 9608
rect 7569 9556 7607 9608
rect 7479 9516 7607 9556
rect 7703 10262 7831 10428
rect 7703 10210 7741 10262
rect 7793 10210 7831 10262
rect 7703 10044 7831 10210
rect 7703 9992 7741 10044
rect 7793 9992 7831 10044
rect 7703 9827 7831 9992
rect 8823 10593 8951 10633
rect 8823 10541 8861 10593
rect 8913 10541 8951 10593
rect 8823 10375 8951 10541
rect 8823 10323 8861 10375
rect 8913 10323 8951 10375
rect 8823 10157 8951 10323
rect 8823 10105 8861 10157
rect 8913 10105 8951 10157
rect 8823 9939 8951 10105
rect 9045 10542 9173 10708
rect 9493 11195 9621 11236
rect 9493 11143 9531 11195
rect 9583 11143 9621 11195
rect 9493 10978 9621 11143
rect 9493 10926 9531 10978
rect 9583 10926 9621 10978
rect 9493 10760 9621 10926
rect 9493 10708 9531 10760
rect 9583 10708 9621 10760
rect 9045 10490 9083 10542
rect 9135 10490 9173 10542
rect 9045 10324 9173 10490
rect 9045 10272 9083 10324
rect 9135 10272 9173 10324
rect 9045 10107 9173 10272
rect 9045 10055 9083 10107
rect 9135 10055 9173 10107
rect 9045 10015 9173 10055
rect 9271 10593 9399 10633
rect 9271 10541 9309 10593
rect 9361 10541 9399 10593
rect 9271 10375 9399 10541
rect 9271 10323 9309 10375
rect 9361 10323 9399 10375
rect 9271 10157 9399 10323
rect 9271 10105 9309 10157
rect 9361 10105 9399 10157
rect 9051 10014 9167 10015
rect 8823 9887 8861 9939
rect 8913 9887 8951 9939
rect 8823 9847 8951 9887
rect 9271 9939 9399 10105
rect 9493 10542 9621 10708
rect 9941 11195 10069 11236
rect 9941 11143 9979 11195
rect 10031 11143 10069 11195
rect 9941 10978 10069 11143
rect 9941 10926 9979 10978
rect 10031 10926 10069 10978
rect 9941 10760 10069 10926
rect 9941 10708 9979 10760
rect 10031 10708 10069 10760
rect 9493 10490 9531 10542
rect 9583 10490 9621 10542
rect 9493 10324 9621 10490
rect 9493 10272 9531 10324
rect 9583 10272 9621 10324
rect 9493 10107 9621 10272
rect 9493 10055 9531 10107
rect 9583 10055 9621 10107
rect 9493 10015 9621 10055
rect 9719 10593 9847 10633
rect 9719 10541 9757 10593
rect 9809 10541 9847 10593
rect 9719 10375 9847 10541
rect 9719 10323 9757 10375
rect 9809 10323 9847 10375
rect 9719 10157 9847 10323
rect 9719 10105 9757 10157
rect 9809 10105 9847 10157
rect 9499 10014 9615 10015
rect 9271 9887 9309 9939
rect 9361 9887 9399 9939
rect 9271 9847 9399 9887
rect 9719 9939 9847 10105
rect 9941 10542 10069 10708
rect 10389 11195 10517 11236
rect 10389 11143 10427 11195
rect 10479 11143 10517 11195
rect 10389 10978 10517 11143
rect 10389 10926 10427 10978
rect 10479 10926 10517 10978
rect 10389 10760 10517 10926
rect 10389 10708 10427 10760
rect 10479 10708 10517 10760
rect 9941 10490 9979 10542
rect 10031 10490 10069 10542
rect 9941 10324 10069 10490
rect 9941 10272 9979 10324
rect 10031 10272 10069 10324
rect 9941 10107 10069 10272
rect 9941 10055 9979 10107
rect 10031 10055 10069 10107
rect 9941 10015 10069 10055
rect 10167 10593 10295 10633
rect 10167 10541 10205 10593
rect 10257 10541 10295 10593
rect 10167 10375 10295 10541
rect 10167 10323 10205 10375
rect 10257 10323 10295 10375
rect 10167 10157 10295 10323
rect 10167 10105 10205 10157
rect 10257 10105 10295 10157
rect 9947 10014 10063 10015
rect 9719 9887 9757 9939
rect 9809 9887 9847 9939
rect 9719 9847 9847 9887
rect 10167 9939 10295 10105
rect 10389 10542 10517 10708
rect 10837 11195 10965 11236
rect 10837 11143 10875 11195
rect 10927 11143 10965 11195
rect 10837 10978 10965 11143
rect 10837 10926 10875 10978
rect 10927 10926 10965 10978
rect 10837 10760 10965 10926
rect 10837 10708 10875 10760
rect 10927 10708 10965 10760
rect 10389 10490 10427 10542
rect 10479 10490 10517 10542
rect 10389 10324 10517 10490
rect 10389 10272 10427 10324
rect 10479 10272 10517 10324
rect 10389 10107 10517 10272
rect 10389 10055 10427 10107
rect 10479 10055 10517 10107
rect 10389 10015 10517 10055
rect 10615 10593 10743 10633
rect 10615 10541 10653 10593
rect 10705 10541 10743 10593
rect 10615 10375 10743 10541
rect 10615 10323 10653 10375
rect 10705 10323 10743 10375
rect 10615 10157 10743 10323
rect 10615 10105 10653 10157
rect 10705 10105 10743 10157
rect 10395 10014 10511 10015
rect 10167 9887 10205 9939
rect 10257 9887 10295 9939
rect 10167 9847 10295 9887
rect 10615 9939 10743 10105
rect 10837 10542 10965 10708
rect 11285 11195 11413 11236
rect 11285 11143 11323 11195
rect 11375 11143 11413 11195
rect 11285 10978 11413 11143
rect 11285 10926 11323 10978
rect 11375 10926 11413 10978
rect 11285 10760 11413 10926
rect 11285 10708 11323 10760
rect 11375 10708 11413 10760
rect 10837 10490 10875 10542
rect 10927 10490 10965 10542
rect 10837 10324 10965 10490
rect 10837 10272 10875 10324
rect 10927 10272 10965 10324
rect 10837 10107 10965 10272
rect 10837 10055 10875 10107
rect 10927 10055 10965 10107
rect 10837 10015 10965 10055
rect 11063 10593 11191 10633
rect 11063 10541 11101 10593
rect 11153 10541 11191 10593
rect 11063 10375 11191 10541
rect 11063 10323 11101 10375
rect 11153 10323 11191 10375
rect 11063 10157 11191 10323
rect 11063 10105 11101 10157
rect 11153 10105 11191 10157
rect 10843 10014 10959 10015
rect 10615 9887 10653 9939
rect 10705 9887 10743 9939
rect 10615 9847 10743 9887
rect 11063 9939 11191 10105
rect 11285 10542 11413 10708
rect 11733 11195 11861 11236
rect 11733 11143 11771 11195
rect 11823 11143 11861 11195
rect 11733 10978 11861 11143
rect 11733 10926 11771 10978
rect 11823 10926 11861 10978
rect 11733 10760 11861 10926
rect 11733 10708 11771 10760
rect 11823 10708 11861 10760
rect 11285 10490 11323 10542
rect 11375 10490 11413 10542
rect 11285 10324 11413 10490
rect 11285 10272 11323 10324
rect 11375 10272 11413 10324
rect 11285 10107 11413 10272
rect 11285 10055 11323 10107
rect 11375 10055 11413 10107
rect 11285 10015 11413 10055
rect 11511 10593 11639 10633
rect 11511 10541 11549 10593
rect 11601 10541 11639 10593
rect 11511 10375 11639 10541
rect 11511 10323 11549 10375
rect 11601 10323 11639 10375
rect 11511 10157 11639 10323
rect 11511 10105 11549 10157
rect 11601 10105 11639 10157
rect 11291 10014 11407 10015
rect 11063 9887 11101 9939
rect 11153 9887 11191 9939
rect 11063 9847 11191 9887
rect 11511 9939 11639 10105
rect 11733 10542 11861 10708
rect 12181 11195 12309 11236
rect 12181 11143 12219 11195
rect 12271 11143 12309 11195
rect 12181 10978 12309 11143
rect 12181 10926 12219 10978
rect 12271 10926 12309 10978
rect 12181 10760 12309 10926
rect 12181 10708 12219 10760
rect 12271 10708 12309 10760
rect 11733 10490 11771 10542
rect 11823 10490 11861 10542
rect 11733 10324 11861 10490
rect 11733 10272 11771 10324
rect 11823 10272 11861 10324
rect 11733 10107 11861 10272
rect 11733 10055 11771 10107
rect 11823 10055 11861 10107
rect 11733 10015 11861 10055
rect 11959 10593 12087 10633
rect 11959 10541 11997 10593
rect 12049 10541 12087 10593
rect 11959 10375 12087 10541
rect 11959 10323 11997 10375
rect 12049 10323 12087 10375
rect 11959 10157 12087 10323
rect 11959 10105 11997 10157
rect 12049 10105 12087 10157
rect 11739 10014 11855 10015
rect 11511 9887 11549 9939
rect 11601 9887 11639 9939
rect 11511 9847 11639 9887
rect 11959 9939 12087 10105
rect 12181 10542 12309 10708
rect 12629 11195 12757 11236
rect 12629 11143 12667 11195
rect 12719 11143 12757 11195
rect 12629 10978 12757 11143
rect 12629 10926 12667 10978
rect 12719 10926 12757 10978
rect 12629 10760 12757 10926
rect 12629 10708 12667 10760
rect 12719 10708 12757 10760
rect 12181 10490 12219 10542
rect 12271 10490 12309 10542
rect 12181 10324 12309 10490
rect 12181 10272 12219 10324
rect 12271 10272 12309 10324
rect 12181 10107 12309 10272
rect 12181 10055 12219 10107
rect 12271 10055 12309 10107
rect 12181 10015 12309 10055
rect 12407 10593 12535 10633
rect 12407 10541 12445 10593
rect 12497 10541 12535 10593
rect 12407 10375 12535 10541
rect 12407 10323 12445 10375
rect 12497 10323 12535 10375
rect 12407 10157 12535 10323
rect 12407 10105 12445 10157
rect 12497 10105 12535 10157
rect 12187 10014 12303 10015
rect 11959 9887 11997 9939
rect 12049 9887 12087 9939
rect 11959 9847 12087 9887
rect 12407 9939 12535 10105
rect 12629 10542 12757 10708
rect 13077 11195 13205 11236
rect 13077 11143 13115 11195
rect 13167 11143 13205 11195
rect 13077 10978 13205 11143
rect 13077 10926 13115 10978
rect 13167 10926 13205 10978
rect 13077 10760 13205 10926
rect 13077 10708 13115 10760
rect 13167 10708 13205 10760
rect 12629 10490 12667 10542
rect 12719 10490 12757 10542
rect 12629 10324 12757 10490
rect 12629 10272 12667 10324
rect 12719 10272 12757 10324
rect 12629 10107 12757 10272
rect 12629 10055 12667 10107
rect 12719 10055 12757 10107
rect 12629 10015 12757 10055
rect 12855 10593 12983 10633
rect 12855 10541 12893 10593
rect 12945 10541 12983 10593
rect 12855 10375 12983 10541
rect 12855 10323 12893 10375
rect 12945 10323 12983 10375
rect 12855 10157 12983 10323
rect 12855 10105 12893 10157
rect 12945 10105 12983 10157
rect 12635 10014 12751 10015
rect 12407 9887 12445 9939
rect 12497 9887 12535 9939
rect 12407 9847 12535 9887
rect 12855 9939 12983 10105
rect 13077 10542 13205 10708
rect 13077 10490 13115 10542
rect 13167 10490 13205 10542
rect 13077 10324 13205 10490
rect 13077 10272 13115 10324
rect 13167 10272 13205 10324
rect 13077 10107 13205 10272
rect 13077 10055 13115 10107
rect 13167 10055 13205 10107
rect 13077 10015 13205 10055
rect 13301 10667 13724 11304
rect 13301 10627 13730 10667
rect 13301 10593 13640 10627
rect 13301 10541 13339 10593
rect 13391 10575 13640 10593
rect 13692 10575 13730 10627
rect 13391 10541 13730 10575
rect 13301 10409 13730 10541
rect 13301 10375 13640 10409
rect 13301 10323 13339 10375
rect 13391 10357 13640 10375
rect 13692 10357 13730 10409
rect 13391 10323 13730 10357
rect 13301 10191 13730 10323
rect 13301 10157 13640 10191
rect 13301 10105 13339 10157
rect 13391 10139 13640 10157
rect 13692 10139 13730 10191
rect 13391 10105 13730 10139
rect 13083 10014 13199 10015
rect 12855 9887 12893 9939
rect 12945 9887 12983 9939
rect 12855 9847 12983 9887
rect 13301 9973 13730 10105
rect 13301 9939 13640 9973
rect 13301 9887 13339 9939
rect 13391 9921 13640 9939
rect 13692 9921 13730 9973
rect 13391 9887 13730 9921
rect 13301 9881 13730 9887
rect 13301 9847 13724 9881
rect 7703 9775 7741 9827
rect 7793 9775 7831 9827
rect 7703 9609 7831 9775
rect 7703 9557 7741 9609
rect 7793 9557 7831 9609
rect 7703 9517 7831 9557
rect 7716 9516 7831 9517
rect 6289 8668 6405 8915
rect 355 7730 4292 8668
rect 4944 8543 5061 8663
rect 6288 8566 6405 8668
rect 7905 8548 8284 8668
rect 4945 7949 5061 8543
rect 6862 8287 7702 8391
rect 5169 7970 5285 8124
rect 5169 7913 5713 7970
rect 5169 7861 5411 7913
rect 5463 7861 5623 7913
rect 5675 7861 5713 7913
rect 5169 7786 5713 7861
rect 4945 7106 5061 7641
rect 5169 7204 5285 7786
rect 6638 7444 6754 7616
rect 6862 7548 6978 8287
rect 7082 8153 7206 8193
rect 7082 8101 7118 8153
rect 7170 8101 7206 8153
rect 7082 7935 7206 8101
rect 7082 7883 7118 7935
rect 7170 7883 7206 7935
rect 7082 7843 7206 7883
rect 7086 7444 7202 7616
rect 6154 7391 6494 7432
rect 6154 7339 6192 7391
rect 6286 7345 6398 7391
rect 6244 7339 6404 7345
rect 6456 7339 6494 7391
rect 6638 7342 7202 7444
rect 6154 7298 6494 7339
rect 6858 7222 6982 7262
rect 6858 7170 6894 7222
rect 6946 7170 6982 7222
rect 4944 7104 5061 7106
rect 4938 7065 5066 7104
rect 4938 7013 4976 7065
rect 5028 7013 5066 7065
rect 4938 6847 5066 7013
rect 5221 7078 5509 7115
rect 5221 7032 5256 7078
rect 5302 7032 5509 7078
rect 5221 6993 5509 7032
rect 4938 6795 4976 6847
rect 5028 6795 5066 6847
rect 4938 6629 5066 6795
rect 4938 6577 4976 6629
rect 5028 6577 5066 6629
rect 4938 6537 5066 6577
rect 5393 6770 5509 6993
rect 6348 6969 6754 7036
rect 6348 6923 6383 6969
rect 6429 6923 6754 6969
rect 6348 6857 6754 6923
rect 6858 7004 6982 7170
rect 7086 7115 7202 7342
rect 6858 6952 6894 7004
rect 6946 6952 6982 7004
rect 6858 6912 6982 6952
rect 7080 7075 7208 7115
rect 7080 7023 7118 7075
rect 7170 7023 7208 7075
rect 6348 6805 6386 6857
rect 6438 6805 6754 6857
rect 6348 6777 6754 6805
rect 5393 6730 5519 6770
rect 5393 6678 5431 6730
rect 5483 6678 5519 6730
rect 4945 6405 5061 6537
rect 4945 6359 4980 6405
rect 5026 6359 5061 6405
rect 4945 6224 5061 6359
rect 4945 6178 4980 6224
rect 5026 6178 5061 6224
rect 4945 6140 5061 6178
rect 5393 6512 5519 6678
rect 5393 6460 5431 6512
rect 5483 6460 5519 6512
rect 5393 6420 5519 6460
rect 6348 6731 6383 6777
rect 6429 6731 6754 6777
rect 6348 6639 6754 6731
rect 6348 6587 6386 6639
rect 6438 6587 6754 6639
rect 6348 6584 6754 6587
rect 6348 6538 6383 6584
rect 6429 6538 6754 6584
rect 6348 6421 6754 6538
rect 5393 6405 5509 6420
rect 5393 6359 5428 6405
rect 5474 6359 5509 6405
rect 5393 6224 5509 6359
rect 5393 6178 5428 6224
rect 5474 6178 5509 6224
rect 4802 6024 5142 6061
rect 4802 6020 5054 6024
rect 5100 6020 5142 6024
rect 4802 5968 4840 6020
rect 4892 5968 5052 6020
rect 5104 5968 5142 6020
rect 4802 5928 5142 5968
rect 5393 5848 5509 6178
rect 6348 6375 6383 6421
rect 6348 6369 6386 6375
rect 6438 6369 6754 6421
rect 6348 6145 6754 6369
rect 6862 6158 6978 6912
rect 7080 6857 7208 7023
rect 7080 6805 7118 6857
rect 7170 6805 7208 6857
rect 7080 6639 7208 6805
rect 7080 6587 7118 6639
rect 7170 6587 7208 6639
rect 7080 6421 7208 6587
rect 7080 6369 7118 6421
rect 7170 6369 7208 6421
rect 7080 6329 7208 6369
rect 6855 6118 6985 6158
rect 6855 6066 6894 6118
rect 6946 6066 6985 6118
rect 6350 5970 6474 6010
rect 6350 5918 6386 5970
rect 6438 5918 6474 5970
rect 6350 5848 6474 5918
rect 6855 5900 6985 6066
rect 7376 6054 7492 8051
rect 7600 7614 7702 8287
rect 7795 8083 7919 8123
rect 7795 8031 7831 8083
rect 7883 8031 7919 8083
rect 7795 7985 7919 8031
rect 7795 7939 7828 7985
rect 7874 7939 7919 7985
rect 7795 7865 7919 7939
rect 7795 7821 7831 7865
rect 7795 7775 7828 7821
rect 7883 7813 7919 7865
rect 7874 7775 7919 7813
rect 7795 7773 7919 7775
rect 7795 7738 7907 7773
rect 7569 7468 7874 7469
rect 7569 7432 7919 7468
rect 7569 7386 7604 7432
rect 7650 7428 7919 7432
rect 7650 7386 7831 7428
rect 7569 7376 7831 7386
rect 7883 7376 7919 7428
rect 7569 7349 7919 7376
rect 7793 7210 7919 7349
rect 7793 7158 7831 7210
rect 7883 7158 7919 7210
rect 7793 7118 7919 7158
rect 7099 6017 7492 6054
rect 7099 5971 7134 6017
rect 7180 5971 7492 6017
rect 7099 5934 7492 5971
rect 6855 5848 6894 5900
rect 6946 5848 6985 5900
rect 4945 5746 5509 5848
rect 4945 5639 5061 5746
rect 5164 5626 5288 5666
rect 5164 5574 5200 5626
rect 5252 5574 5288 5626
rect 5393 5621 5509 5746
rect 5751 5811 5880 5848
rect 5751 5765 5788 5811
rect 5834 5807 5880 5811
rect 5751 5755 5789 5765
rect 5841 5755 5880 5807
rect 5164 5408 5288 5574
rect 5751 5589 5880 5755
rect 5751 5537 5789 5589
rect 5841 5537 5880 5589
rect 5751 5497 5880 5537
rect 6348 5752 6754 5848
rect 6855 5807 6985 5848
rect 6348 5707 6386 5752
rect 6348 5661 6383 5707
rect 6438 5700 6754 5752
rect 6862 5737 6978 5807
rect 7376 5759 7492 5934
rect 6429 5661 6754 5700
rect 6348 5543 6754 5661
rect 6348 5497 6383 5543
rect 6429 5501 6754 5543
rect 6429 5497 6464 5501
rect 5164 5356 5200 5408
rect 5252 5356 5288 5408
rect 5164 5316 5288 5356
rect 5168 5315 5285 5316
rect 5169 5165 5285 5315
rect 6348 5165 6464 5497
rect 7086 5165 7202 5757
rect 7569 5716 7680 6831
rect 7793 6069 7874 7118
rect 7758 6033 7874 6069
rect 7758 5987 7793 6033
rect 7839 5987 7874 6033
rect 7758 5950 7874 5987
rect 7569 5596 8811 5716
rect 8948 5658 9532 9452
rect 9863 9412 9980 9482
rect 10838 9412 10955 9482
rect 11286 9412 11403 9482
rect 12123 9412 12239 9482
rect 9864 9126 9980 9412
rect 10155 9030 10300 9193
rect 10839 9126 10955 9412
rect 11287 9126 11403 9412
rect 12124 9126 12239 9412
rect 12571 9126 12687 9482
rect 9636 8990 9760 9030
rect 9636 8938 9672 8990
rect 9724 8938 9760 8990
rect 9636 8772 9760 8938
rect 9636 8720 9672 8772
rect 9724 8720 9760 8772
rect 9636 8680 9760 8720
rect 10086 8990 10300 9030
rect 10086 8938 10122 8990
rect 10174 8938 10300 8990
rect 10086 8772 10300 8938
rect 10086 8720 10122 8772
rect 10174 8720 10300 8772
rect 10086 8680 10300 8720
rect 9416 5657 9532 5658
rect 7569 5410 7680 5596
rect 8696 5249 8811 5596
rect 10155 5293 10300 8680
rect 8585 5208 8925 5249
rect 67 4191 8120 5165
rect 8585 5156 8623 5208
rect 8675 5156 8835 5208
rect 8887 5156 8925 5208
rect 9752 5201 9868 5202
rect 9978 5201 10094 5202
rect 8585 5115 8925 5156
rect 9745 5161 9875 5201
rect 9745 5109 9784 5161
rect 9836 5109 9875 5161
rect 9557 5095 9625 5106
rect 9557 5002 9568 5095
rect 8228 4955 9568 5002
rect 9614 4955 9625 5095
rect 8228 4882 9625 4955
rect 9745 5095 9875 5109
rect 9745 4955 9791 5095
rect 9837 4955 9875 5095
rect 9745 4943 9875 4955
rect 9745 4891 9784 4943
rect 9836 4891 9875 4943
rect 8228 4281 8344 4882
rect 9745 4850 9875 4891
rect 9971 5161 10101 5201
rect 9971 5109 10010 5161
rect 10062 5109 10101 5161
rect 9971 5095 10101 5109
rect 9971 4955 10015 5095
rect 10061 4955 10101 5095
rect 9971 4943 10101 4955
rect 9971 4891 10010 4943
rect 10062 4891 10101 4943
rect 9971 4850 10101 4891
rect 8878 4752 9532 4789
rect 8878 4706 9451 4752
rect 9497 4706 9532 4752
rect 8878 4584 9532 4706
rect 10184 4696 10300 5293
rect 8878 4538 9451 4584
rect 9497 4538 9532 4584
rect 8878 4417 9532 4538
rect 8878 4371 9451 4417
rect 9497 4371 9532 4417
rect 5082 3832 5128 4191
rect 5386 3772 5859 3892
rect 6127 3772 6242 4191
rect 5324 3594 5664 3599
rect 5310 3558 5664 3594
rect 5310 3557 5362 3558
rect 5414 3557 5574 3558
rect 5310 3511 5345 3557
rect 5414 3511 5503 3557
rect 5549 3511 5574 3557
rect 5310 3506 5362 3511
rect 5414 3506 5574 3511
rect 5626 3506 5664 3558
rect 5310 3474 5664 3506
rect 5324 3466 5664 3474
rect 5743 3594 5859 3772
rect 6504 3594 6619 3918
rect 6848 3777 6925 4191
rect 7183 3594 7299 3918
rect 7490 3789 7606 4191
rect 7749 3594 7795 3941
rect 8004 3789 8120 4191
rect 8878 4249 9532 4371
rect 8878 4203 9451 4249
rect 9497 4203 9532 4249
rect 8878 4081 9532 4203
rect 8878 4035 9451 4081
rect 9497 4035 9532 4081
rect 5743 3557 6264 3594
rect 5743 3511 6183 3557
rect 6229 3511 6264 3557
rect 5743 3474 6264 3511
rect 6504 3557 6987 3594
rect 6504 3511 6907 3557
rect 6953 3511 6987 3557
rect 6504 3474 6987 3511
rect 7183 3593 7598 3594
rect 7183 3557 7627 3593
rect 7183 3511 7547 3557
rect 7593 3511 7627 3557
rect 7183 3474 7627 3511
rect 7749 3557 8146 3594
rect 7749 3511 8065 3557
rect 8111 3511 8146 3557
rect 7749 3474 8146 3511
rect 5743 3260 5859 3474
rect 5082 2477 5128 3108
rect 5426 3080 5859 3260
rect 6117 2543 6233 3260
rect 6504 3252 6619 3474
rect 6503 3050 6619 3252
rect 6841 2543 6957 3260
rect 7183 3080 7299 3474
rect 7490 2751 7606 3260
rect 7749 3132 7795 3474
rect 7003 2335 7606 2751
rect 8004 3063 8120 3260
rect 8263 3132 8309 3921
rect 8878 3913 9532 4035
rect 8878 3867 9451 3913
rect 9497 3867 9532 3913
rect 8878 3746 9532 3867
rect 8878 3700 9451 3746
rect 9497 3700 9532 3746
rect 8878 3578 9532 3700
rect 8878 3532 9451 3578
rect 9497 3532 9532 3578
rect 8878 3410 9532 3532
rect 8878 3364 9451 3410
rect 9497 3364 9532 3410
rect 8004 2699 8036 3063
rect 8088 2699 8120 3063
rect 8004 2543 8120 2699
rect 8452 3063 8568 3260
rect 8452 2699 8484 3063
rect 8536 2699 8568 3063
rect 8452 2543 8568 2699
rect 8878 3242 9532 3364
rect 8878 3196 9451 3242
rect 9497 3196 9532 3242
rect 8878 3075 9532 3196
rect 8878 3029 9451 3075
rect 9497 3029 9532 3075
rect 8878 2905 9532 3029
rect 8878 2859 9451 2905
rect 9497 2859 9532 2905
rect 8878 2735 9532 2859
rect 8878 2689 9451 2735
rect 9497 2689 9532 2735
rect 8878 2565 9532 2689
rect 8878 2519 9451 2565
rect 9497 2519 9532 2565
rect 8878 2395 9532 2519
rect 8878 2349 9451 2395
rect 9497 2349 9532 2395
rect 8878 2225 9532 2349
rect 8878 2179 9451 2225
rect 9497 2179 9532 2225
rect 8878 2055 9532 2179
rect 8878 2009 9451 2055
rect 9497 2009 9532 2055
rect 8878 1884 9532 2009
rect 8878 1838 9451 1884
rect 9497 1838 9532 1884
rect 8878 1714 9532 1838
rect 8878 1668 9451 1714
rect 9497 1668 9532 1714
rect 8878 1544 9532 1668
rect 8878 1498 9451 1544
rect 9497 1498 9532 1544
rect 8878 1374 9532 1498
rect 8878 1328 9451 1374
rect 9497 1328 9532 1374
rect 8878 1204 9532 1328
rect 8878 1158 9451 1204
rect 9497 1158 9532 1204
rect 8878 1034 9532 1158
rect 8878 988 9451 1034
rect 9497 988 9532 1034
rect 8878 864 9532 988
rect 8878 818 9451 864
rect 9497 818 9532 864
rect 8878 694 9532 818
rect 8878 648 9451 694
rect 9497 648 9532 694
rect 8878 524 9532 648
rect 8878 478 9451 524
rect 9497 478 9532 524
rect 8878 354 9532 478
rect 8878 308 9451 354
rect 9497 308 9532 354
rect 8878 -110 9532 308
rect 10088 4584 10300 4696
rect 10088 4538 10123 4584
rect 10169 4538 10300 4584
rect 11893 5413 12021 5453
rect 11893 5361 11931 5413
rect 11983 5361 12021 5413
rect 11893 5195 12021 5361
rect 11893 5143 11931 5195
rect 11983 5143 12021 5195
rect 11893 4977 12021 5143
rect 11893 4925 11931 4977
rect 11983 4925 12021 4977
rect 11893 4759 12021 4925
rect 11893 4707 11931 4759
rect 11983 4712 12021 4759
rect 12341 5413 12469 5453
rect 12341 5361 12379 5413
rect 12431 5361 12469 5413
rect 12341 5195 12469 5361
rect 12341 5143 12379 5195
rect 12431 5143 12469 5195
rect 12341 4977 12469 5143
rect 12341 4925 12379 4977
rect 12431 4925 12469 4977
rect 12341 4759 12469 4925
rect 11983 4707 12022 4712
rect 11893 4574 12022 4707
rect 12341 4707 12379 4759
rect 12431 4707 12469 4759
rect 12341 4667 12469 4707
rect 12789 5413 12917 5453
rect 12789 5361 12827 5413
rect 12879 5361 12917 5413
rect 12789 5195 12917 5361
rect 12789 5143 12827 5195
rect 12879 5143 12917 5195
rect 12789 4977 12917 5143
rect 12789 4925 12827 4977
rect 12879 4925 12917 4977
rect 12789 4759 12917 4925
rect 12789 4707 12827 4759
rect 12879 4707 12917 4759
rect 12789 4667 12917 4707
rect 10088 4417 10300 4538
rect 10727 4537 12022 4574
rect 12595 4540 12935 4553
rect 10727 4491 10763 4537
rect 10809 4491 11434 4537
rect 11480 4491 12022 4537
rect 10727 4454 12022 4491
rect 12268 4512 12935 4540
rect 12268 4506 12633 4512
rect 12268 4460 12294 4506
rect 12528 4460 12633 4506
rect 12685 4460 12845 4512
rect 12897 4460 12935 4512
rect 12268 4420 12935 4460
rect 10088 4371 10123 4417
rect 10169 4371 10300 4417
rect 10088 4356 10300 4371
rect 10088 4319 11258 4356
rect 10088 4273 11049 4319
rect 11189 4273 11258 4319
rect 10088 4249 11258 4273
rect 10088 4203 10123 4249
rect 10169 4236 11258 4249
rect 11557 4324 11897 4331
rect 11557 4290 12799 4324
rect 11557 4238 11595 4290
rect 11647 4238 11807 4290
rect 11859 4288 12799 4290
rect 11859 4242 12046 4288
rect 12092 4242 12718 4288
rect 12764 4242 12799 4288
rect 11859 4238 12799 4242
rect 10169 4203 10300 4236
rect 10088 4081 10300 4203
rect 11557 4204 12799 4238
rect 11557 4198 11897 4204
rect 10088 4035 10123 4081
rect 10169 4035 10300 4081
rect 10088 3913 10300 4035
rect 10615 4068 10731 4104
rect 10615 4032 10650 4068
rect 10088 3867 10123 3913
rect 10169 3867 10300 3913
rect 10088 3746 10300 3867
rect 10088 3700 10123 3746
rect 10169 3700 10300 3746
rect 10088 3578 10300 3700
rect 10088 3532 10123 3578
rect 10169 3532 10300 3578
rect 10088 3410 10300 3532
rect 10088 3364 10123 3410
rect 10169 3364 10300 3410
rect 10088 3242 10300 3364
rect 10088 3196 10123 3242
rect 10169 3196 10300 3242
rect 10088 3075 10300 3196
rect 10088 3029 10123 3075
rect 10169 3029 10300 3075
rect 10088 2905 10300 3029
rect 10088 2859 10123 2905
rect 10169 2859 10300 2905
rect 10088 2735 10300 2859
rect 10088 2689 10123 2735
rect 10169 2689 10300 2735
rect 10088 2565 10300 2689
rect 10088 2519 10123 2565
rect 10169 2519 10300 2565
rect 10088 2395 10300 2519
rect 10088 2349 10123 2395
rect 10169 2349 10300 2395
rect 10088 2225 10300 2349
rect 10088 2179 10123 2225
rect 10169 2179 10300 2225
rect 10088 2055 10300 2179
rect 10088 2009 10123 2055
rect 10169 2009 10300 2055
rect 10088 1884 10300 2009
rect 10088 1838 10123 1884
rect 10169 1838 10300 1884
rect 10088 1714 10300 1838
rect 10088 1668 10123 1714
rect 10169 1668 10300 1714
rect 10088 1544 10300 1668
rect 10088 1498 10123 1544
rect 10169 1498 10300 1544
rect 10088 1374 10300 1498
rect 10088 1328 10123 1374
rect 10169 1328 10300 1374
rect 10088 1204 10300 1328
rect 10088 1158 10123 1204
rect 10169 1158 10300 1204
rect 10088 1034 10300 1158
rect 10088 988 10123 1034
rect 10169 988 10300 1034
rect 10088 864 10300 988
rect 10088 818 10123 864
rect 10169 818 10300 864
rect 10088 694 10300 818
rect 10088 648 10123 694
rect 10169 648 10300 694
rect 10088 524 10300 648
rect 10088 478 10123 524
rect 10169 478 10300 524
rect 10088 354 10300 478
rect 10088 308 10123 354
rect 10169 308 10300 354
rect 10088 271 10300 308
rect 10614 4022 10650 4032
rect 10696 4022 10731 4068
rect 10614 3900 10731 4022
rect 10614 3854 10650 3900
rect 10696 3854 10731 3900
rect 10614 3732 10731 3854
rect 10614 3686 10650 3732
rect 10696 3686 10731 3732
rect 10614 3564 10731 3686
rect 10614 3518 10650 3564
rect 10696 3518 10731 3564
rect 10614 3397 10731 3518
rect 10614 3351 10650 3397
rect 10696 3351 10731 3397
rect 10614 3229 10731 3351
rect 10614 3183 10650 3229
rect 10696 3183 10731 3229
rect 10614 3061 10731 3183
rect 10614 3015 10650 3061
rect 10696 3015 10731 3061
rect 10614 2893 10731 3015
rect 10614 2847 10650 2893
rect 10696 2847 10731 2893
rect 10614 2726 10731 2847
rect 10614 2680 10650 2726
rect 10696 2680 10731 2726
rect 10614 2558 10731 2680
rect 10614 2512 10650 2558
rect 10696 2512 10731 2558
rect 10614 2390 10731 2512
rect 10614 2344 10650 2390
rect 10696 2344 10731 2390
rect 10614 2220 10731 2344
rect 11062 4068 11179 4104
rect 11062 4022 11098 4068
rect 11144 4022 11179 4068
rect 11511 4068 11627 4104
rect 11511 4032 11546 4068
rect 11062 3900 11179 4022
rect 11062 3854 11098 3900
rect 11144 3854 11179 3900
rect 11062 3732 11179 3854
rect 11062 3686 11098 3732
rect 11144 3686 11179 3732
rect 11062 3564 11179 3686
rect 11062 3518 11098 3564
rect 11144 3518 11179 3564
rect 11062 3397 11179 3518
rect 11062 3351 11098 3397
rect 11144 3351 11179 3397
rect 11062 3229 11179 3351
rect 11062 3183 11098 3229
rect 11144 3183 11179 3229
rect 11062 3061 11179 3183
rect 11062 3015 11098 3061
rect 11144 3015 11179 3061
rect 11062 2893 11179 3015
rect 11062 2847 11098 2893
rect 11144 2847 11179 2893
rect 11062 2726 11179 2847
rect 11062 2680 11098 2726
rect 11144 2680 11179 2726
rect 11062 2558 11179 2680
rect 11062 2512 11098 2558
rect 11144 2512 11179 2558
rect 11062 2390 11179 2512
rect 11062 2344 11098 2390
rect 11144 2344 11179 2390
rect 11062 2230 11179 2344
rect 10614 2174 10650 2220
rect 10696 2174 10731 2220
rect 10614 2050 10731 2174
rect 10614 2004 10650 2050
rect 10696 2004 10731 2050
rect 10614 1880 10731 2004
rect 10614 1834 10650 1880
rect 10696 1834 10731 1880
rect 10614 1710 10731 1834
rect 10614 1664 10650 1710
rect 10696 1664 10731 1710
rect 10614 1540 10731 1664
rect 10614 1494 10650 1540
rect 10696 1494 10731 1540
rect 10614 1370 10731 1494
rect 10614 1324 10650 1370
rect 10696 1324 10731 1370
rect 10614 1200 10731 1324
rect 10614 1154 10650 1200
rect 10696 1154 10731 1200
rect 10614 1030 10731 1154
rect 10614 984 10650 1030
rect 10696 984 10731 1030
rect 10614 860 10731 984
rect 10614 814 10650 860
rect 10696 814 10731 860
rect 10614 690 10731 814
rect 10614 644 10650 690
rect 10696 644 10731 690
rect 10614 199 10731 644
rect 11063 2220 11179 2230
rect 11063 2174 11098 2220
rect 11144 2174 11179 2220
rect 11063 2050 11179 2174
rect 11063 2004 11098 2050
rect 11144 2004 11179 2050
rect 11063 1880 11179 2004
rect 11063 1834 11098 1880
rect 11144 1834 11179 1880
rect 11063 1710 11179 1834
rect 11063 1664 11098 1710
rect 11144 1664 11179 1710
rect 11063 1540 11179 1664
rect 11063 1494 11098 1540
rect 11144 1494 11179 1540
rect 11063 1370 11179 1494
rect 11063 1324 11098 1370
rect 11144 1324 11179 1370
rect 11063 1200 11179 1324
rect 11063 1154 11098 1200
rect 11144 1154 11179 1200
rect 11063 1030 11179 1154
rect 11063 984 11098 1030
rect 11144 984 11179 1030
rect 11063 860 11179 984
rect 11063 814 11098 860
rect 11144 814 11179 860
rect 11063 690 11179 814
rect 11063 644 11098 690
rect 11144 644 11179 690
rect 11063 493 11179 644
rect 11510 4022 11546 4032
rect 11592 4022 11627 4068
rect 11900 4068 12015 4104
rect 11900 4032 11934 4068
rect 11510 3900 11627 4022
rect 11510 3854 11546 3900
rect 11592 3854 11627 3900
rect 11510 3732 11627 3854
rect 11510 3686 11546 3732
rect 11592 3686 11627 3732
rect 11510 3564 11627 3686
rect 11510 3518 11546 3564
rect 11592 3518 11627 3564
rect 11510 3397 11627 3518
rect 11510 3351 11546 3397
rect 11592 3351 11627 3397
rect 11510 3229 11627 3351
rect 11510 3183 11546 3229
rect 11592 3183 11627 3229
rect 11510 3061 11627 3183
rect 11510 3015 11546 3061
rect 11592 3015 11627 3061
rect 11510 2893 11627 3015
rect 11510 2847 11546 2893
rect 11592 2847 11627 2893
rect 11510 2726 11627 2847
rect 11510 2680 11546 2726
rect 11592 2680 11627 2726
rect 11510 2558 11627 2680
rect 11510 2512 11546 2558
rect 11592 2512 11627 2558
rect 11510 2390 11627 2512
rect 11510 2344 11546 2390
rect 11592 2344 11627 2390
rect 11510 2220 11627 2344
rect 11510 2174 11546 2220
rect 11592 2174 11627 2220
rect 11510 2050 11627 2174
rect 11510 2004 11546 2050
rect 11592 2004 11627 2050
rect 11510 1880 11627 2004
rect 11510 1834 11546 1880
rect 11592 1834 11627 1880
rect 11510 1710 11627 1834
rect 11510 1664 11546 1710
rect 11592 1664 11627 1710
rect 11510 1540 11627 1664
rect 11510 1494 11546 1540
rect 11592 1494 11627 1540
rect 11510 1370 11627 1494
rect 11510 1324 11546 1370
rect 11592 1324 11627 1370
rect 11510 1200 11627 1324
rect 11510 1154 11546 1200
rect 11592 1154 11627 1200
rect 11510 1030 11627 1154
rect 11510 984 11546 1030
rect 11592 984 11627 1030
rect 11510 860 11627 984
rect 11510 814 11546 860
rect 11592 814 11627 860
rect 11510 690 11627 814
rect 11510 644 11546 690
rect 11592 644 11627 690
rect 11510 199 11627 644
rect 11899 4022 11934 4032
rect 11980 4022 12015 4068
rect 11899 3900 12015 4022
rect 11899 3854 11934 3900
rect 11980 3854 12015 3900
rect 11899 3732 12015 3854
rect 11899 3686 11934 3732
rect 11980 3686 12015 3732
rect 11899 3564 12015 3686
rect 11899 3518 11934 3564
rect 11980 3518 12015 3564
rect 11899 3397 12015 3518
rect 11899 3351 11934 3397
rect 11980 3351 12015 3397
rect 11899 199 12015 3351
rect 12347 4068 12463 4104
rect 12347 4022 12382 4068
rect 12428 4022 12463 4068
rect 12347 3900 12463 4022
rect 12347 3854 12382 3900
rect 12428 3854 12463 3900
rect 12347 3732 12463 3854
rect 12347 3686 12382 3732
rect 12428 3686 12463 3732
rect 12347 3564 12463 3686
rect 12347 3518 12382 3564
rect 12428 3518 12463 3564
rect 12347 3397 12463 3518
rect 12347 3351 12382 3397
rect 12428 3351 12463 3397
rect 12347 2230 12463 3351
rect 12795 4068 13605 4104
rect 12795 4022 12830 4068
rect 12876 4022 13605 4068
rect 12795 3732 13605 4022
rect 12795 3686 12830 3732
rect 12876 3686 13605 3732
rect 12795 3564 13605 3686
rect 12795 3518 12830 3564
rect 12876 3518 13605 3564
rect 12795 3397 13605 3518
rect 12795 3351 12830 3397
rect 12876 3351 13605 3397
rect 10615 37 10731 199
rect 11511 37 11627 199
rect 11900 37 12015 199
rect 10614 -67 10731 37
rect 11510 -110 11627 37
rect 11899 -58 12015 37
rect 12795 -37 13605 3351
rect 8999 -477 13686 -384
rect 8999 -529 10253 -477
rect 10305 -529 10465 -477
rect 10517 -529 12976 -477
rect 13028 -529 13188 -477
rect 13240 -529 13686 -477
rect 8999 -695 13686 -529
rect 8999 -747 10253 -695
rect 10305 -747 10465 -695
rect 10517 -747 12976 -695
rect 13028 -747 13188 -695
rect 13240 -747 13686 -695
rect 8999 -840 13686 -747
<< via1 >>
rect 6551 14381 6603 14433
rect 6551 14164 6603 14216
rect 6551 13946 6603 13998
rect 6551 13728 6603 13780
rect 6551 13511 6603 13563
rect 6999 14381 7051 14433
rect 6999 14164 7051 14216
rect 6999 13946 7051 13998
rect 6999 13728 7051 13780
rect 6999 13511 7051 13563
rect 7447 14381 7499 14433
rect 7447 14164 7499 14216
rect 7447 13946 7499 13998
rect 7447 13728 7499 13780
rect 7447 13511 7499 13563
rect 7895 14381 7947 14433
rect 7895 14164 7947 14216
rect 7895 13946 7947 13998
rect 7895 13728 7947 13780
rect 7895 13511 7947 13563
rect 8343 14381 8395 14433
rect 8343 14164 8395 14216
rect 8343 13946 8395 13998
rect 8343 13728 8395 13780
rect 8343 13511 8395 13563
rect 6577 13284 6629 13336
rect 6788 13284 6840 13336
rect 7000 13284 7052 13336
rect 7211 13284 7263 13336
rect 6314 11241 6366 11293
rect 6607 11148 6659 11200
rect 6818 11148 6870 11200
rect 7030 11148 7082 11200
rect 7241 11148 7293 11200
rect 9083 11143 9135 11195
rect 6314 11023 6366 11075
rect 6314 10806 6366 10858
rect 6314 10588 6366 10640
rect 6314 10370 6366 10422
rect 6314 10153 6366 10205
rect 6314 9935 6366 9987
rect 6846 10863 6898 10915
rect 6846 10645 6898 10697
rect 6846 10428 6898 10480
rect 7293 10863 7345 10915
rect 7293 10645 7345 10697
rect 7293 10428 7345 10480
rect 6846 10210 6898 10262
rect 6846 9992 6898 10044
rect 6846 9775 6898 9827
rect 6846 9557 6898 9609
rect 7070 10210 7122 10262
rect 7070 9992 7122 10044
rect 7070 9774 7122 9826
rect 7070 9556 7122 9608
rect 7741 10863 7793 10915
rect 7741 10645 7793 10697
rect 9083 10926 9135 10978
rect 9083 10708 9135 10760
rect 7741 10428 7793 10480
rect 7293 10210 7345 10262
rect 7293 9992 7345 10044
rect 7293 9775 7345 9827
rect 7293 9557 7345 9609
rect 7517 10210 7569 10262
rect 7517 9992 7569 10044
rect 7517 9774 7569 9826
rect 7517 9556 7569 9608
rect 7741 10210 7793 10262
rect 7741 9992 7793 10044
rect 8861 10541 8913 10593
rect 8861 10323 8913 10375
rect 8861 10105 8913 10157
rect 9531 11143 9583 11195
rect 9531 10926 9583 10978
rect 9531 10708 9583 10760
rect 9083 10490 9135 10542
rect 9083 10272 9135 10324
rect 9083 10055 9135 10107
rect 9309 10541 9361 10593
rect 9309 10323 9361 10375
rect 9309 10105 9361 10157
rect 8861 9887 8913 9939
rect 9979 11143 10031 11195
rect 9979 10926 10031 10978
rect 9979 10708 10031 10760
rect 9531 10490 9583 10542
rect 9531 10272 9583 10324
rect 9531 10055 9583 10107
rect 9757 10541 9809 10593
rect 9757 10323 9809 10375
rect 9757 10105 9809 10157
rect 9309 9887 9361 9939
rect 10427 11143 10479 11195
rect 10427 10926 10479 10978
rect 10427 10708 10479 10760
rect 9979 10490 10031 10542
rect 9979 10272 10031 10324
rect 9979 10055 10031 10107
rect 10205 10541 10257 10593
rect 10205 10323 10257 10375
rect 10205 10105 10257 10157
rect 9757 9887 9809 9939
rect 10875 11143 10927 11195
rect 10875 10926 10927 10978
rect 10875 10708 10927 10760
rect 10427 10490 10479 10542
rect 10427 10272 10479 10324
rect 10427 10055 10479 10107
rect 10653 10541 10705 10593
rect 10653 10323 10705 10375
rect 10653 10105 10705 10157
rect 10205 9887 10257 9939
rect 11323 11143 11375 11195
rect 11323 10926 11375 10978
rect 11323 10708 11375 10760
rect 10875 10490 10927 10542
rect 10875 10272 10927 10324
rect 10875 10055 10927 10107
rect 11101 10541 11153 10593
rect 11101 10323 11153 10375
rect 11101 10105 11153 10157
rect 10653 9887 10705 9939
rect 11771 11143 11823 11195
rect 11771 10926 11823 10978
rect 11771 10708 11823 10760
rect 11323 10490 11375 10542
rect 11323 10272 11375 10324
rect 11323 10055 11375 10107
rect 11549 10541 11601 10593
rect 11549 10323 11601 10375
rect 11549 10105 11601 10157
rect 11101 9887 11153 9939
rect 12219 11143 12271 11195
rect 12219 10926 12271 10978
rect 12219 10708 12271 10760
rect 11771 10490 11823 10542
rect 11771 10272 11823 10324
rect 11771 10055 11823 10107
rect 11997 10541 12049 10593
rect 11997 10323 12049 10375
rect 11997 10105 12049 10157
rect 11549 9887 11601 9939
rect 12667 11143 12719 11195
rect 12667 10926 12719 10978
rect 12667 10708 12719 10760
rect 12219 10490 12271 10542
rect 12219 10272 12271 10324
rect 12219 10055 12271 10107
rect 12445 10541 12497 10593
rect 12445 10323 12497 10375
rect 12445 10105 12497 10157
rect 11997 9887 12049 9939
rect 13115 11143 13167 11195
rect 13115 10926 13167 10978
rect 13115 10708 13167 10760
rect 12667 10490 12719 10542
rect 12667 10272 12719 10324
rect 12667 10055 12719 10107
rect 12893 10541 12945 10593
rect 12893 10323 12945 10375
rect 12893 10105 12945 10157
rect 12445 9887 12497 9939
rect 13115 10490 13167 10542
rect 13115 10272 13167 10324
rect 13115 10055 13167 10107
rect 13339 10541 13391 10593
rect 13640 10575 13692 10627
rect 13339 10323 13391 10375
rect 13640 10357 13692 10409
rect 13339 10105 13391 10157
rect 13640 10139 13692 10191
rect 12893 9887 12945 9939
rect 13339 9887 13391 9939
rect 13640 9921 13692 9973
rect 7741 9775 7793 9827
rect 7741 9557 7793 9609
rect 5411 7861 5463 7913
rect 5623 7861 5675 7913
rect 7118 8101 7170 8153
rect 7118 7883 7170 7935
rect 6192 7345 6240 7391
rect 6240 7345 6244 7391
rect 6404 7345 6444 7391
rect 6444 7345 6456 7391
rect 6192 7339 6244 7345
rect 6404 7339 6456 7345
rect 6894 7170 6946 7222
rect 4976 7013 5028 7065
rect 4976 6795 5028 6847
rect 4976 6577 5028 6629
rect 6894 6952 6946 7004
rect 7118 7023 7170 7075
rect 6386 6805 6438 6857
rect 5431 6678 5483 6730
rect 5431 6460 5483 6512
rect 6386 6587 6438 6639
rect 4840 5968 4892 6020
rect 5052 5978 5054 6020
rect 5054 5978 5100 6020
rect 5100 5978 5104 6020
rect 5052 5968 5104 5978
rect 6386 6375 6429 6421
rect 6429 6375 6438 6421
rect 6386 6369 6438 6375
rect 7118 6805 7170 6857
rect 7118 6587 7170 6639
rect 7118 6369 7170 6421
rect 6894 6066 6946 6118
rect 6386 5918 6438 5970
rect 7831 8031 7883 8083
rect 7831 7821 7883 7865
rect 7831 7813 7874 7821
rect 7874 7813 7883 7821
rect 7831 7376 7883 7428
rect 7831 7158 7883 7210
rect 6894 5848 6946 5900
rect 5200 5574 5252 5626
rect 5789 5765 5834 5807
rect 5834 5765 5841 5807
rect 5789 5755 5841 5765
rect 5789 5537 5841 5589
rect 6386 5707 6438 5752
rect 6386 5700 6429 5707
rect 6429 5700 6438 5707
rect 5200 5356 5252 5408
rect 9672 8938 9724 8990
rect 9672 8720 9724 8772
rect 10122 8938 10174 8990
rect 10122 8720 10174 8772
rect 8623 5156 8675 5208
rect 8835 5156 8887 5208
rect 9784 5109 9836 5161
rect 9784 4891 9836 4943
rect 10010 5109 10062 5161
rect 10010 4891 10062 4943
rect 5362 3557 5414 3558
rect 5362 3511 5391 3557
rect 5391 3511 5414 3557
rect 5362 3506 5414 3511
rect 5574 3506 5626 3558
rect 8036 2699 8088 3063
rect 8484 2699 8536 3063
rect 11931 5361 11983 5413
rect 11931 5143 11983 5195
rect 11931 4925 11983 4977
rect 11931 4707 11983 4759
rect 12379 5361 12431 5413
rect 12379 5143 12431 5195
rect 12379 4925 12431 4977
rect 12379 4707 12431 4759
rect 12827 5361 12879 5413
rect 12827 5143 12879 5195
rect 12827 4925 12879 4977
rect 12827 4707 12879 4759
rect 12633 4460 12685 4512
rect 12845 4460 12897 4512
rect 11595 4238 11647 4290
rect 11807 4238 11859 4290
rect 10253 -529 10305 -477
rect 10465 -529 10517 -477
rect 12976 -529 13028 -477
rect 13188 -529 13240 -477
rect 10253 -747 10305 -695
rect 10465 -747 10517 -695
rect 12976 -747 13028 -695
rect 13188 -747 13240 -695
<< metal2 >>
rect 6225 14621 13430 16278
rect 6513 14433 8434 14474
rect 6513 14381 6551 14433
rect 6603 14381 6999 14433
rect 7051 14381 7447 14433
rect 7499 14381 7895 14433
rect 7947 14381 8343 14433
rect 8395 14381 8434 14433
rect 6513 14216 8434 14381
rect 6513 14164 6551 14216
rect 6603 14164 6999 14216
rect 7051 14164 7447 14216
rect 7499 14164 7895 14216
rect 7947 14164 8343 14216
rect 8395 14164 8434 14216
rect 6513 13998 8434 14164
rect 6513 13946 6551 13998
rect 6603 13946 6999 13998
rect 7051 13946 7447 13998
rect 7499 13946 7895 13998
rect 7947 13946 8343 13998
rect 8395 13946 8434 13998
rect 6513 13780 8434 13946
rect 6513 13728 6551 13780
rect 6603 13728 6999 13780
rect 7051 13728 7447 13780
rect 7499 13728 7895 13780
rect 7947 13728 8343 13780
rect 8395 13728 8434 13780
rect 6513 13563 8434 13728
rect 6513 13511 6551 13563
rect 6603 13511 6999 13563
rect 7051 13511 7447 13563
rect 7499 13511 7895 13563
rect 7947 13511 8343 13563
rect 8395 13511 8434 13563
rect 6513 13470 8434 13511
rect 6497 13336 7364 13376
rect 6497 13284 6577 13336
rect 6629 13284 6788 13336
rect 6840 13284 7000 13336
rect 7052 13284 7211 13336
rect 7263 13284 7364 13336
rect 6276 11295 6404 11332
rect 6276 11239 6312 11295
rect 6368 11239 6404 11295
rect 6276 11077 6404 11239
rect 6276 11021 6312 11077
rect 6368 11021 6404 11077
rect 6276 10860 6404 11021
rect 6276 10804 6312 10860
rect 6368 10804 6404 10860
rect 6276 10642 6404 10804
rect 6276 10586 6312 10642
rect 6368 10586 6404 10642
rect 6276 10424 6404 10586
rect 6276 10368 6312 10424
rect 6368 10368 6404 10424
rect 6276 10207 6404 10368
rect 6276 10151 6312 10207
rect 6368 10151 6404 10207
rect 6276 9989 6404 10151
rect 6276 9933 6312 9989
rect 6368 9933 6404 9989
rect 6276 9895 6404 9933
rect 6497 11200 7364 13284
rect 6497 11148 6607 11200
rect 6659 11148 6818 11200
rect 6870 11148 7030 11200
rect 7082 11148 7241 11200
rect 7293 11148 7364 11200
rect 6497 11107 7364 11148
rect 7591 12211 8192 13470
rect 9045 12502 13206 14376
rect 7591 11384 11159 12211
rect 6497 9258 6725 11107
rect 7591 10955 8192 11384
rect 11555 11282 13206 12502
rect 6838 10954 8192 10955
rect 6808 10915 8192 10954
rect 6808 10863 6846 10915
rect 6898 10863 7293 10915
rect 7345 10863 7741 10915
rect 7793 10863 8192 10915
rect 6808 10697 8192 10863
rect 6808 10645 6846 10697
rect 6898 10656 7293 10697
rect 6898 10645 6936 10656
rect 6808 10480 6936 10645
rect 6808 10428 6846 10480
rect 6898 10428 6936 10480
rect 6808 10262 6936 10428
rect 7255 10645 7293 10656
rect 7345 10656 7741 10697
rect 7345 10645 7383 10656
rect 7255 10480 7383 10645
rect 7255 10428 7293 10480
rect 7345 10428 7383 10480
rect 6808 10210 6846 10262
rect 6898 10210 6936 10262
rect 6808 10044 6936 10210
rect 6808 9992 6846 10044
rect 6898 9992 6936 10044
rect 6808 9827 6936 9992
rect 6808 9775 6846 9827
rect 6898 9775 6936 9827
rect 6808 9609 6936 9775
rect 6808 9557 6846 9609
rect 6898 9557 6936 9609
rect 6808 9517 6936 9557
rect 7032 10264 7160 10301
rect 7032 10208 7068 10264
rect 7124 10208 7160 10264
rect 7032 10046 7160 10208
rect 7032 9990 7068 10046
rect 7124 9990 7160 10046
rect 7032 9828 7160 9990
rect 7032 9772 7068 9828
rect 7124 9772 7160 9828
rect 7032 9610 7160 9772
rect 7032 9554 7068 9610
rect 7124 9554 7160 9610
rect 7032 9516 7160 9554
rect 7255 10262 7383 10428
rect 7703 10645 7741 10656
rect 7793 10656 8192 10697
rect 8428 11195 13206 11282
rect 8428 11143 9083 11195
rect 9135 11143 9531 11195
rect 9583 11143 9979 11195
rect 10031 11143 10427 11195
rect 10479 11143 10875 11195
rect 10927 11143 11323 11195
rect 11375 11143 11771 11195
rect 11823 11143 12219 11195
rect 12271 11143 12667 11195
rect 12719 11143 13115 11195
rect 13167 11143 13206 11195
rect 8428 10978 13206 11143
rect 8428 10926 9083 10978
rect 9135 10926 9531 10978
rect 9583 10926 9979 10978
rect 10031 10926 10427 10978
rect 10479 10926 10875 10978
rect 10927 10926 11323 10978
rect 11375 10926 11771 10978
rect 11823 10926 12219 10978
rect 12271 10926 12667 10978
rect 12719 10926 13115 10978
rect 13167 10926 13206 10978
rect 8428 10760 13206 10926
rect 8428 10731 9083 10760
rect 7793 10645 7831 10656
rect 7703 10480 7831 10645
rect 7703 10428 7741 10480
rect 7793 10428 7831 10480
rect 7255 10210 7293 10262
rect 7345 10210 7383 10262
rect 7255 10044 7383 10210
rect 7255 9992 7293 10044
rect 7345 9992 7383 10044
rect 7255 9827 7383 9992
rect 7255 9775 7293 9827
rect 7345 9775 7383 9827
rect 7255 9609 7383 9775
rect 7255 9557 7293 9609
rect 7345 9557 7383 9609
rect 7255 9517 7383 9557
rect 7479 10264 7607 10301
rect 7479 10208 7515 10264
rect 7571 10208 7607 10264
rect 7479 10046 7607 10208
rect 7479 9990 7515 10046
rect 7571 9990 7607 10046
rect 7479 9828 7607 9990
rect 7479 9772 7515 9828
rect 7571 9772 7607 9828
rect 7479 9610 7607 9772
rect 7479 9554 7515 9610
rect 7571 9554 7607 9610
rect 7479 9516 7607 9554
rect 7703 10262 7831 10428
rect 7703 10210 7741 10262
rect 7793 10210 7831 10262
rect 7703 10044 7831 10210
rect 7703 9992 7741 10044
rect 7793 9992 7831 10044
rect 7703 9827 7831 9992
rect 7703 9775 7741 9827
rect 7793 9775 7831 9827
rect 7703 9609 7831 9775
rect 7703 9557 7741 9609
rect 7793 9557 7831 9609
rect 7703 9517 7831 9557
rect 8428 9736 8719 10731
rect 9045 10708 9083 10731
rect 9135 10731 9531 10760
rect 9135 10708 9174 10731
rect 8823 10595 8951 10632
rect 8823 10539 8859 10595
rect 8915 10539 8951 10595
rect 8823 10377 8951 10539
rect 8823 10321 8859 10377
rect 8915 10321 8951 10377
rect 8823 10159 8951 10321
rect 8823 10103 8859 10159
rect 8915 10103 8951 10159
rect 8823 9941 8951 10103
rect 8823 9885 8859 9941
rect 8915 9885 8951 9941
rect 8823 9847 8951 9885
rect 9045 10542 9174 10708
rect 9493 10708 9531 10731
rect 9583 10731 9979 10760
rect 9583 10708 9622 10731
rect 9045 10490 9083 10542
rect 9135 10490 9174 10542
rect 9045 10324 9174 10490
rect 9045 10272 9083 10324
rect 9135 10272 9174 10324
rect 9045 10107 9174 10272
rect 9045 10055 9083 10107
rect 9135 10055 9174 10107
rect 9045 9736 9174 10055
rect 9271 10595 9399 10632
rect 9271 10539 9307 10595
rect 9363 10539 9399 10595
rect 9271 10377 9399 10539
rect 9271 10321 9307 10377
rect 9363 10321 9399 10377
rect 9271 10159 9399 10321
rect 9271 10103 9307 10159
rect 9363 10103 9399 10159
rect 9271 9941 9399 10103
rect 9271 9885 9307 9941
rect 9363 9885 9399 9941
rect 9271 9847 9399 9885
rect 9493 10542 9622 10708
rect 9941 10708 9979 10731
rect 10031 10731 10427 10760
rect 10031 10708 10070 10731
rect 9493 10490 9531 10542
rect 9583 10490 9622 10542
rect 9493 10324 9622 10490
rect 9493 10272 9531 10324
rect 9583 10272 9622 10324
rect 9493 10107 9622 10272
rect 9493 10055 9531 10107
rect 9583 10055 9622 10107
rect 9493 9736 9622 10055
rect 9719 10595 9847 10632
rect 9719 10539 9755 10595
rect 9811 10539 9847 10595
rect 9719 10377 9847 10539
rect 9719 10321 9755 10377
rect 9811 10321 9847 10377
rect 9719 10159 9847 10321
rect 9719 10103 9755 10159
rect 9811 10103 9847 10159
rect 9719 9941 9847 10103
rect 9719 9885 9755 9941
rect 9811 9885 9847 9941
rect 9719 9847 9847 9885
rect 9941 10542 10070 10708
rect 10389 10708 10427 10731
rect 10479 10731 10875 10760
rect 10479 10708 10518 10731
rect 9941 10490 9979 10542
rect 10031 10490 10070 10542
rect 9941 10324 10070 10490
rect 9941 10272 9979 10324
rect 10031 10272 10070 10324
rect 9941 10107 10070 10272
rect 9941 10055 9979 10107
rect 10031 10055 10070 10107
rect 9941 9736 10070 10055
rect 10167 10595 10295 10632
rect 10167 10539 10203 10595
rect 10259 10539 10295 10595
rect 10167 10377 10295 10539
rect 10167 10321 10203 10377
rect 10259 10321 10295 10377
rect 10167 10159 10295 10321
rect 10167 10103 10203 10159
rect 10259 10103 10295 10159
rect 10167 9941 10295 10103
rect 10167 9885 10203 9941
rect 10259 9885 10295 9941
rect 10167 9847 10295 9885
rect 10389 10542 10518 10708
rect 10837 10708 10875 10731
rect 10927 10731 11323 10760
rect 10927 10708 10966 10731
rect 10389 10490 10427 10542
rect 10479 10490 10518 10542
rect 10389 10324 10518 10490
rect 10389 10272 10427 10324
rect 10479 10272 10518 10324
rect 10389 10107 10518 10272
rect 10389 10055 10427 10107
rect 10479 10055 10518 10107
rect 10389 9736 10518 10055
rect 10615 10595 10743 10632
rect 10615 10539 10651 10595
rect 10707 10539 10743 10595
rect 10615 10377 10743 10539
rect 10615 10321 10651 10377
rect 10707 10321 10743 10377
rect 10615 10159 10743 10321
rect 10615 10103 10651 10159
rect 10707 10103 10743 10159
rect 10615 9941 10743 10103
rect 10615 9885 10651 9941
rect 10707 9885 10743 9941
rect 10615 9847 10743 9885
rect 10837 10542 10966 10708
rect 11285 10708 11323 10731
rect 11375 10731 11771 10760
rect 11375 10708 11414 10731
rect 10837 10490 10875 10542
rect 10927 10490 10966 10542
rect 10837 10324 10966 10490
rect 10837 10272 10875 10324
rect 10927 10272 10966 10324
rect 10837 10107 10966 10272
rect 10837 10055 10875 10107
rect 10927 10055 10966 10107
rect 10837 9736 10966 10055
rect 11063 10595 11191 10632
rect 11063 10539 11099 10595
rect 11155 10539 11191 10595
rect 11063 10377 11191 10539
rect 11063 10321 11099 10377
rect 11155 10321 11191 10377
rect 11063 10159 11191 10321
rect 11063 10103 11099 10159
rect 11155 10103 11191 10159
rect 11063 9941 11191 10103
rect 11063 9885 11099 9941
rect 11155 9885 11191 9941
rect 11063 9847 11191 9885
rect 11285 10542 11414 10708
rect 11733 10708 11771 10731
rect 11823 10731 12219 10760
rect 11823 10708 11862 10731
rect 11285 10490 11323 10542
rect 11375 10490 11414 10542
rect 11285 10324 11414 10490
rect 11285 10272 11323 10324
rect 11375 10272 11414 10324
rect 11285 10107 11414 10272
rect 11285 10055 11323 10107
rect 11375 10055 11414 10107
rect 11285 9736 11414 10055
rect 11511 10595 11639 10632
rect 11511 10539 11547 10595
rect 11603 10539 11639 10595
rect 11511 10377 11639 10539
rect 11511 10321 11547 10377
rect 11603 10321 11639 10377
rect 11511 10159 11639 10321
rect 11511 10103 11547 10159
rect 11603 10103 11639 10159
rect 11511 9941 11639 10103
rect 11511 9885 11547 9941
rect 11603 9885 11639 9941
rect 11511 9847 11639 9885
rect 11733 10542 11862 10708
rect 12181 10708 12219 10731
rect 12271 10731 12667 10760
rect 12271 10708 12310 10731
rect 11733 10490 11771 10542
rect 11823 10490 11862 10542
rect 11733 10324 11862 10490
rect 11733 10272 11771 10324
rect 11823 10272 11862 10324
rect 11733 10107 11862 10272
rect 11733 10055 11771 10107
rect 11823 10055 11862 10107
rect 11733 9736 11862 10055
rect 11959 10595 12087 10632
rect 11959 10539 11995 10595
rect 12051 10539 12087 10595
rect 11959 10377 12087 10539
rect 11959 10321 11995 10377
rect 12051 10321 12087 10377
rect 11959 10159 12087 10321
rect 11959 10103 11995 10159
rect 12051 10103 12087 10159
rect 11959 9941 12087 10103
rect 11959 9885 11995 9941
rect 12051 9885 12087 9941
rect 11959 9847 12087 9885
rect 12181 10542 12310 10708
rect 12629 10708 12667 10731
rect 12719 10731 13115 10760
rect 12719 10708 12758 10731
rect 12181 10490 12219 10542
rect 12271 10490 12310 10542
rect 12181 10324 12310 10490
rect 12181 10272 12219 10324
rect 12271 10272 12310 10324
rect 12181 10107 12310 10272
rect 12181 10055 12219 10107
rect 12271 10055 12310 10107
rect 12181 9736 12310 10055
rect 12407 10595 12535 10632
rect 12407 10539 12443 10595
rect 12499 10539 12535 10595
rect 12407 10377 12535 10539
rect 12407 10321 12443 10377
rect 12499 10321 12535 10377
rect 12407 10159 12535 10321
rect 12407 10103 12443 10159
rect 12499 10103 12535 10159
rect 12407 9941 12535 10103
rect 12407 9885 12443 9941
rect 12499 9885 12535 9941
rect 12407 9847 12535 9885
rect 12629 10542 12758 10708
rect 13077 10708 13115 10731
rect 13167 10708 13206 10760
rect 12629 10490 12667 10542
rect 12719 10490 12758 10542
rect 12629 10324 12758 10490
rect 12629 10272 12667 10324
rect 12719 10272 12758 10324
rect 12629 10107 12758 10272
rect 12629 10055 12667 10107
rect 12719 10055 12758 10107
rect 12629 9736 12758 10055
rect 12855 10595 12983 10632
rect 12855 10539 12891 10595
rect 12947 10539 12983 10595
rect 12855 10377 12983 10539
rect 12855 10321 12891 10377
rect 12947 10321 12983 10377
rect 12855 10159 12983 10321
rect 12855 10103 12891 10159
rect 12947 10103 12983 10159
rect 12855 9941 12983 10103
rect 12855 9885 12891 9941
rect 12947 9885 12983 9941
rect 12855 9847 12983 9885
rect 13077 10542 13206 10708
rect 13077 10490 13115 10542
rect 13167 10490 13206 10542
rect 13077 10324 13206 10490
rect 13077 10272 13115 10324
rect 13167 10272 13206 10324
rect 13077 10107 13206 10272
rect 13077 10055 13115 10107
rect 13167 10055 13206 10107
rect 13077 9736 13206 10055
rect 13301 10595 13429 10632
rect 13301 10539 13337 10595
rect 13393 10539 13429 10595
rect 13301 10377 13429 10539
rect 13301 10321 13337 10377
rect 13393 10321 13429 10377
rect 13301 10159 13429 10321
rect 13301 10103 13337 10159
rect 13393 10103 13429 10159
rect 13301 9941 13429 10103
rect 13301 9885 13337 9941
rect 13393 9885 13429 9941
rect 13301 9847 13429 9885
rect 13602 10629 13730 10666
rect 13602 10573 13638 10629
rect 13694 10573 13730 10629
rect 13602 10411 13730 10573
rect 13602 10355 13638 10411
rect 13694 10355 13730 10411
rect 13602 10193 13730 10355
rect 13602 10137 13638 10193
rect 13694 10137 13730 10193
rect 13602 9975 13730 10137
rect 13602 9919 13638 9975
rect 13694 9919 13730 9975
rect 13602 9881 13730 9919
rect 8428 9355 13206 9736
rect 6497 9257 6768 9258
rect 6497 9219 6888 9257
rect 6497 9163 6584 9219
rect 6640 9163 6796 9219
rect 6852 9163 6888 9219
rect 6497 9001 6888 9163
rect 6497 8945 6584 9001
rect 6640 8945 6796 9001
rect 6852 8945 6888 9001
rect 6497 8906 6888 8945
rect 8428 8808 8719 9355
rect 4611 8760 8719 8808
rect 4611 8704 4647 8760
rect 4703 8704 4859 8760
rect 4915 8704 8719 8760
rect 4611 8659 8719 8704
rect 9633 8990 10212 9030
rect 9633 8938 9672 8990
rect 9724 8938 10122 8990
rect 10174 8938 10212 8990
rect 9633 8772 10212 8938
rect 9633 8720 9672 8772
rect 9724 8720 10122 8772
rect 10174 8720 10212 8772
rect 9633 8679 10212 8720
rect -319 7396 21 7435
rect -319 7340 -283 7396
rect -227 7340 -71 7396
rect -15 7340 21 7396
rect -319 7301 21 7340
rect -279 -2007 -146 7301
rect 4714 6061 4848 8659
rect 5474 8565 5713 8566
rect 7897 8565 8027 8566
rect 5374 8527 5713 8565
rect 5374 8471 5409 8527
rect 5465 8471 5621 8527
rect 5677 8471 5713 8527
rect 5374 8432 5713 8471
rect 7688 8527 8027 8565
rect 7688 8471 7723 8527
rect 7779 8471 7935 8527
rect 7991 8471 8027 8527
rect 7688 8432 8027 8471
rect 5474 7954 5603 8432
rect 7081 8155 7206 8194
rect 7081 8099 7116 8155
rect 7172 8099 7206 8155
rect 5373 7913 5713 7954
rect 5373 7861 5411 7913
rect 5463 7861 5623 7913
rect 5675 7861 5713 7913
rect 5373 7820 5713 7861
rect 7081 7937 7206 8099
rect 7081 7881 7116 7937
rect 7172 7881 7206 7937
rect 7081 7843 7206 7881
rect 7793 8083 7922 8432
rect 7793 8031 7831 8083
rect 7883 8031 7922 8083
rect 7793 7865 7922 8031
rect 7793 7813 7831 7865
rect 7883 7813 7922 7865
rect 7793 7773 7922 7813
rect 5391 7528 7926 7666
rect 4938 7067 5066 7104
rect 4938 7011 4974 7067
rect 5030 7011 5066 7067
rect 4938 6849 5066 7011
rect 4938 6793 4974 6849
rect 5030 6793 5066 6849
rect 4938 6631 5066 6793
rect 4938 6575 4974 6631
rect 5030 6575 5066 6631
rect 4938 6537 5066 6575
rect 5391 6730 5524 7528
rect 5641 7396 5981 7435
rect 5641 7340 5677 7396
rect 5733 7340 5889 7396
rect 5945 7340 5981 7396
rect 5641 7301 5981 7340
rect 6154 7391 6494 7432
rect 6154 7339 6192 7391
rect 6244 7339 6404 7391
rect 6456 7339 6494 7391
rect 5391 6678 5431 6730
rect 5483 6678 5524 6730
rect 5391 6512 5524 6678
rect 5391 6460 5431 6512
rect 5483 6460 5524 6512
rect 5391 6451 5524 6460
rect 5395 6420 5519 6451
rect 4714 6020 5142 6061
rect 4714 5968 4840 6020
rect 4892 5968 5052 6020
rect 5104 5968 5142 6020
rect 4714 5928 5142 5968
rect 4714 5927 4848 5928
rect 5738 5807 5886 7301
rect 6154 7298 6494 7339
rect 7793 7428 7926 7528
rect 7793 7376 7831 7428
rect 7883 7376 7926 7428
rect 6273 7149 6407 7298
rect 6858 7222 6982 7262
rect 6858 7170 6894 7222
rect 6946 7170 6982 7222
rect 6858 7149 6982 7170
rect 6273 7011 6982 7149
rect 7793 7210 7926 7376
rect 7793 7158 7831 7210
rect 7883 7158 7926 7210
rect 7793 7117 7926 7158
rect 6858 7004 6982 7011
rect 6858 6952 6894 7004
rect 6946 6952 6982 7004
rect 6858 6912 6982 6952
rect 7080 7077 7208 7114
rect 7080 7021 7116 7077
rect 7172 7021 7208 7077
rect 6348 6859 6476 6896
rect 6348 6803 6384 6859
rect 6440 6803 6476 6859
rect 6348 6641 6476 6803
rect 6348 6585 6384 6641
rect 6440 6585 6476 6641
rect 6348 6423 6476 6585
rect 6348 6367 6384 6423
rect 6440 6367 6476 6423
rect 6348 6329 6476 6367
rect 7080 6859 7208 7021
rect 7080 6803 7116 6859
rect 7172 6803 7208 6859
rect 7080 6641 7208 6803
rect 7080 6585 7116 6641
rect 7172 6585 7208 6641
rect 7080 6423 7208 6585
rect 7080 6367 7116 6423
rect 7172 6367 7208 6423
rect 7080 6329 7208 6367
rect 6855 6118 6985 6158
rect 6855 6066 6894 6118
rect 6946 6066 6985 6118
rect 6855 6063 6985 6066
rect 5738 5755 5789 5807
rect 5841 5755 5886 5807
rect 5164 5628 5289 5667
rect 5164 5572 5198 5628
rect 5254 5572 5289 5628
rect 5164 5410 5289 5572
rect 5164 5354 5198 5410
rect 5254 5354 5289 5410
rect 5164 5316 5289 5354
rect 5738 5589 5886 5755
rect 6349 5972 6474 6011
rect 6349 5916 6384 5972
rect 6440 5916 6474 5972
rect 6349 5754 6474 5916
rect 6855 5930 10100 6063
rect 6855 5900 6985 5930
rect 6855 5848 6894 5900
rect 6946 5848 6985 5900
rect 6855 5807 6985 5848
rect 6349 5698 6384 5754
rect 6440 5698 6474 5754
rect 6349 5660 6474 5698
rect 5738 5537 5789 5589
rect 5841 5537 5886 5589
rect 5738 5496 5886 5537
rect 5738 5363 9874 5496
rect 5738 3599 5886 5363
rect 8585 5208 8925 5249
rect 8585 5156 8623 5208
rect 8675 5156 8835 5208
rect 8887 5156 8925 5208
rect 8585 5115 8925 5156
rect 9745 5201 9874 5363
rect 9971 5201 10100 5930
rect 9745 5161 9875 5201
rect 5325 3558 5886 3599
rect 5325 3506 5362 3558
rect 5414 3506 5574 3558
rect 5626 3506 5886 3558
rect 5325 3466 5886 3506
rect 8024 3065 8100 3075
rect 8024 2697 8034 3065
rect 8090 2697 8100 3065
rect 8024 2687 8100 2697
rect 8472 3065 8548 3075
rect 8472 2697 8482 3065
rect 8538 2697 8548 3065
rect 8472 2687 8548 2697
rect 8689 -253 8822 5115
rect 9745 5109 9784 5161
rect 9836 5109 9875 5161
rect 9745 4943 9875 5109
rect 9745 4891 9784 4943
rect 9836 4891 9875 4943
rect 9745 4850 9875 4891
rect 9971 5161 10101 5201
rect 9971 5109 10010 5161
rect 10062 5109 10101 5161
rect 9971 4943 10101 5109
rect 9971 4891 10010 4943
rect 10062 4891 10101 4943
rect 9971 4850 10101 4891
rect 10321 -436 10450 9355
rect 10607 9219 10732 9258
rect 10607 9163 10642 9219
rect 10698 9163 10732 9219
rect 10607 9001 10732 9163
rect 10607 8945 10642 9001
rect 10698 8945 10732 9001
rect 10607 8907 10732 8945
rect 11058 9219 11183 9258
rect 11058 9163 11093 9219
rect 11149 9163 11183 9219
rect 11058 9001 11183 9163
rect 11058 8945 11093 9001
rect 11149 8945 11183 9001
rect 11058 8907 11183 8945
rect 11506 9219 11631 9258
rect 11506 9163 11541 9219
rect 11597 9163 11631 9219
rect 11506 9001 11631 9163
rect 11506 8945 11541 9001
rect 11597 8945 11631 9001
rect 11506 8907 11631 8945
rect 11812 8555 13206 9355
rect 11062 5331 11179 8484
rect 11893 5413 12918 5453
rect 11893 5361 11931 5413
rect 11983 5361 12379 5413
rect 12431 5361 12827 5413
rect 12879 5361 12918 5413
rect 10608 4869 11633 5331
rect 11893 5195 12918 5361
rect 11893 5143 11931 5195
rect 11983 5143 12379 5195
rect 12431 5143 12827 5195
rect 12879 5143 12918 5195
rect 11893 4977 12918 5143
rect 11893 4925 11931 4977
rect 11983 4925 12379 4977
rect 12431 4925 12827 4977
rect 12879 4925 12918 4977
rect 11063 4331 11179 4869
rect 11893 4759 12918 4925
rect 11893 4707 11931 4759
rect 11983 4707 12379 4759
rect 12431 4707 12827 4759
rect 12879 4707 12918 4759
rect 11893 4667 12918 4707
rect 11063 4290 11897 4331
rect 11063 4238 11595 4290
rect 11647 4238 11807 4290
rect 11859 4238 11897 4290
rect 11063 4198 11897 4238
rect 11063 4104 11179 4198
rect 12348 4104 12463 4667
rect 12595 4514 12935 4553
rect 12595 4458 12631 4514
rect 12687 4458 12843 4514
rect 12899 4458 12935 4514
rect 12595 4419 12935 4458
rect 11062 3771 11179 4104
rect 12347 3771 12463 4104
rect 13044 -436 13173 8555
rect 10215 -477 10555 -436
rect 10215 -529 10253 -477
rect 10305 -529 10465 -477
rect 10517 -529 10555 -477
rect 10215 -695 10555 -529
rect 10215 -747 10253 -695
rect 10305 -747 10465 -695
rect 10517 -747 10555 -695
rect 10215 -787 10555 -747
rect 12938 -477 13278 -436
rect 12938 -529 12976 -477
rect 13028 -529 13188 -477
rect 13240 -529 13278 -477
rect 12938 -695 13278 -529
rect 12938 -747 12976 -695
rect 13028 -747 13188 -695
rect 13240 -747 13278 -695
rect 12938 -787 13278 -747
rect -383 -2046 -43 -2007
rect -383 -2102 -347 -2046
rect -291 -2102 -135 -2046
rect -79 -2102 -43 -2046
rect -383 -2140 -43 -2102
rect -280 -2141 -146 -2140
<< via2 >>
rect 6312 11293 6368 11295
rect 6312 11241 6314 11293
rect 6314 11241 6366 11293
rect 6366 11241 6368 11293
rect 6312 11239 6368 11241
rect 6312 11075 6368 11077
rect 6312 11023 6314 11075
rect 6314 11023 6366 11075
rect 6366 11023 6368 11075
rect 6312 11021 6368 11023
rect 6312 10858 6368 10860
rect 6312 10806 6314 10858
rect 6314 10806 6366 10858
rect 6366 10806 6368 10858
rect 6312 10804 6368 10806
rect 6312 10640 6368 10642
rect 6312 10588 6314 10640
rect 6314 10588 6366 10640
rect 6366 10588 6368 10640
rect 6312 10586 6368 10588
rect 6312 10422 6368 10424
rect 6312 10370 6314 10422
rect 6314 10370 6366 10422
rect 6366 10370 6368 10422
rect 6312 10368 6368 10370
rect 6312 10205 6368 10207
rect 6312 10153 6314 10205
rect 6314 10153 6366 10205
rect 6366 10153 6368 10205
rect 6312 10151 6368 10153
rect 6312 9987 6368 9989
rect 6312 9935 6314 9987
rect 6314 9935 6366 9987
rect 6366 9935 6368 9987
rect 6312 9933 6368 9935
rect 7068 10262 7124 10264
rect 7068 10210 7070 10262
rect 7070 10210 7122 10262
rect 7122 10210 7124 10262
rect 7068 10208 7124 10210
rect 7068 10044 7124 10046
rect 7068 9992 7070 10044
rect 7070 9992 7122 10044
rect 7122 9992 7124 10044
rect 7068 9990 7124 9992
rect 7068 9826 7124 9828
rect 7068 9774 7070 9826
rect 7070 9774 7122 9826
rect 7122 9774 7124 9826
rect 7068 9772 7124 9774
rect 7068 9608 7124 9610
rect 7068 9556 7070 9608
rect 7070 9556 7122 9608
rect 7122 9556 7124 9608
rect 7068 9554 7124 9556
rect 7515 10262 7571 10264
rect 7515 10210 7517 10262
rect 7517 10210 7569 10262
rect 7569 10210 7571 10262
rect 7515 10208 7571 10210
rect 7515 10044 7571 10046
rect 7515 9992 7517 10044
rect 7517 9992 7569 10044
rect 7569 9992 7571 10044
rect 7515 9990 7571 9992
rect 7515 9826 7571 9828
rect 7515 9774 7517 9826
rect 7517 9774 7569 9826
rect 7569 9774 7571 9826
rect 7515 9772 7571 9774
rect 7515 9608 7571 9610
rect 7515 9556 7517 9608
rect 7517 9556 7569 9608
rect 7569 9556 7571 9608
rect 7515 9554 7571 9556
rect 8859 10593 8915 10595
rect 8859 10541 8861 10593
rect 8861 10541 8913 10593
rect 8913 10541 8915 10593
rect 8859 10539 8915 10541
rect 8859 10375 8915 10377
rect 8859 10323 8861 10375
rect 8861 10323 8913 10375
rect 8913 10323 8915 10375
rect 8859 10321 8915 10323
rect 8859 10157 8915 10159
rect 8859 10105 8861 10157
rect 8861 10105 8913 10157
rect 8913 10105 8915 10157
rect 8859 10103 8915 10105
rect 8859 9939 8915 9941
rect 8859 9887 8861 9939
rect 8861 9887 8913 9939
rect 8913 9887 8915 9939
rect 8859 9885 8915 9887
rect 9307 10593 9363 10595
rect 9307 10541 9309 10593
rect 9309 10541 9361 10593
rect 9361 10541 9363 10593
rect 9307 10539 9363 10541
rect 9307 10375 9363 10377
rect 9307 10323 9309 10375
rect 9309 10323 9361 10375
rect 9361 10323 9363 10375
rect 9307 10321 9363 10323
rect 9307 10157 9363 10159
rect 9307 10105 9309 10157
rect 9309 10105 9361 10157
rect 9361 10105 9363 10157
rect 9307 10103 9363 10105
rect 9307 9939 9363 9941
rect 9307 9887 9309 9939
rect 9309 9887 9361 9939
rect 9361 9887 9363 9939
rect 9307 9885 9363 9887
rect 9755 10593 9811 10595
rect 9755 10541 9757 10593
rect 9757 10541 9809 10593
rect 9809 10541 9811 10593
rect 9755 10539 9811 10541
rect 9755 10375 9811 10377
rect 9755 10323 9757 10375
rect 9757 10323 9809 10375
rect 9809 10323 9811 10375
rect 9755 10321 9811 10323
rect 9755 10157 9811 10159
rect 9755 10105 9757 10157
rect 9757 10105 9809 10157
rect 9809 10105 9811 10157
rect 9755 10103 9811 10105
rect 9755 9939 9811 9941
rect 9755 9887 9757 9939
rect 9757 9887 9809 9939
rect 9809 9887 9811 9939
rect 9755 9885 9811 9887
rect 10203 10593 10259 10595
rect 10203 10541 10205 10593
rect 10205 10541 10257 10593
rect 10257 10541 10259 10593
rect 10203 10539 10259 10541
rect 10203 10375 10259 10377
rect 10203 10323 10205 10375
rect 10205 10323 10257 10375
rect 10257 10323 10259 10375
rect 10203 10321 10259 10323
rect 10203 10157 10259 10159
rect 10203 10105 10205 10157
rect 10205 10105 10257 10157
rect 10257 10105 10259 10157
rect 10203 10103 10259 10105
rect 10203 9939 10259 9941
rect 10203 9887 10205 9939
rect 10205 9887 10257 9939
rect 10257 9887 10259 9939
rect 10203 9885 10259 9887
rect 10651 10593 10707 10595
rect 10651 10541 10653 10593
rect 10653 10541 10705 10593
rect 10705 10541 10707 10593
rect 10651 10539 10707 10541
rect 10651 10375 10707 10377
rect 10651 10323 10653 10375
rect 10653 10323 10705 10375
rect 10705 10323 10707 10375
rect 10651 10321 10707 10323
rect 10651 10157 10707 10159
rect 10651 10105 10653 10157
rect 10653 10105 10705 10157
rect 10705 10105 10707 10157
rect 10651 10103 10707 10105
rect 10651 9939 10707 9941
rect 10651 9887 10653 9939
rect 10653 9887 10705 9939
rect 10705 9887 10707 9939
rect 10651 9885 10707 9887
rect 11099 10593 11155 10595
rect 11099 10541 11101 10593
rect 11101 10541 11153 10593
rect 11153 10541 11155 10593
rect 11099 10539 11155 10541
rect 11099 10375 11155 10377
rect 11099 10323 11101 10375
rect 11101 10323 11153 10375
rect 11153 10323 11155 10375
rect 11099 10321 11155 10323
rect 11099 10157 11155 10159
rect 11099 10105 11101 10157
rect 11101 10105 11153 10157
rect 11153 10105 11155 10157
rect 11099 10103 11155 10105
rect 11099 9939 11155 9941
rect 11099 9887 11101 9939
rect 11101 9887 11153 9939
rect 11153 9887 11155 9939
rect 11099 9885 11155 9887
rect 11547 10593 11603 10595
rect 11547 10541 11549 10593
rect 11549 10541 11601 10593
rect 11601 10541 11603 10593
rect 11547 10539 11603 10541
rect 11547 10375 11603 10377
rect 11547 10323 11549 10375
rect 11549 10323 11601 10375
rect 11601 10323 11603 10375
rect 11547 10321 11603 10323
rect 11547 10157 11603 10159
rect 11547 10105 11549 10157
rect 11549 10105 11601 10157
rect 11601 10105 11603 10157
rect 11547 10103 11603 10105
rect 11547 9939 11603 9941
rect 11547 9887 11549 9939
rect 11549 9887 11601 9939
rect 11601 9887 11603 9939
rect 11547 9885 11603 9887
rect 11995 10593 12051 10595
rect 11995 10541 11997 10593
rect 11997 10541 12049 10593
rect 12049 10541 12051 10593
rect 11995 10539 12051 10541
rect 11995 10375 12051 10377
rect 11995 10323 11997 10375
rect 11997 10323 12049 10375
rect 12049 10323 12051 10375
rect 11995 10321 12051 10323
rect 11995 10157 12051 10159
rect 11995 10105 11997 10157
rect 11997 10105 12049 10157
rect 12049 10105 12051 10157
rect 11995 10103 12051 10105
rect 11995 9939 12051 9941
rect 11995 9887 11997 9939
rect 11997 9887 12049 9939
rect 12049 9887 12051 9939
rect 11995 9885 12051 9887
rect 12443 10593 12499 10595
rect 12443 10541 12445 10593
rect 12445 10541 12497 10593
rect 12497 10541 12499 10593
rect 12443 10539 12499 10541
rect 12443 10375 12499 10377
rect 12443 10323 12445 10375
rect 12445 10323 12497 10375
rect 12497 10323 12499 10375
rect 12443 10321 12499 10323
rect 12443 10157 12499 10159
rect 12443 10105 12445 10157
rect 12445 10105 12497 10157
rect 12497 10105 12499 10157
rect 12443 10103 12499 10105
rect 12443 9939 12499 9941
rect 12443 9887 12445 9939
rect 12445 9887 12497 9939
rect 12497 9887 12499 9939
rect 12443 9885 12499 9887
rect 12891 10593 12947 10595
rect 12891 10541 12893 10593
rect 12893 10541 12945 10593
rect 12945 10541 12947 10593
rect 12891 10539 12947 10541
rect 12891 10375 12947 10377
rect 12891 10323 12893 10375
rect 12893 10323 12945 10375
rect 12945 10323 12947 10375
rect 12891 10321 12947 10323
rect 12891 10157 12947 10159
rect 12891 10105 12893 10157
rect 12893 10105 12945 10157
rect 12945 10105 12947 10157
rect 12891 10103 12947 10105
rect 12891 9939 12947 9941
rect 12891 9887 12893 9939
rect 12893 9887 12945 9939
rect 12945 9887 12947 9939
rect 12891 9885 12947 9887
rect 13337 10593 13393 10595
rect 13337 10541 13339 10593
rect 13339 10541 13391 10593
rect 13391 10541 13393 10593
rect 13337 10539 13393 10541
rect 13337 10375 13393 10377
rect 13337 10323 13339 10375
rect 13339 10323 13391 10375
rect 13391 10323 13393 10375
rect 13337 10321 13393 10323
rect 13337 10157 13393 10159
rect 13337 10105 13339 10157
rect 13339 10105 13391 10157
rect 13391 10105 13393 10157
rect 13337 10103 13393 10105
rect 13337 9939 13393 9941
rect 13337 9887 13339 9939
rect 13339 9887 13391 9939
rect 13391 9887 13393 9939
rect 13337 9885 13393 9887
rect 13638 10627 13694 10629
rect 13638 10575 13640 10627
rect 13640 10575 13692 10627
rect 13692 10575 13694 10627
rect 13638 10573 13694 10575
rect 13638 10409 13694 10411
rect 13638 10357 13640 10409
rect 13640 10357 13692 10409
rect 13692 10357 13694 10409
rect 13638 10355 13694 10357
rect 13638 10191 13694 10193
rect 13638 10139 13640 10191
rect 13640 10139 13692 10191
rect 13692 10139 13694 10191
rect 13638 10137 13694 10139
rect 13638 9973 13694 9975
rect 13638 9921 13640 9973
rect 13640 9921 13692 9973
rect 13692 9921 13694 9973
rect 13638 9919 13694 9921
rect 6584 9163 6640 9219
rect 6796 9163 6852 9219
rect 6584 8945 6640 9001
rect 6796 8945 6852 9001
rect 4647 8704 4703 8760
rect 4859 8704 4915 8760
rect -283 7340 -227 7396
rect -71 7340 -15 7396
rect 5409 8471 5465 8527
rect 5621 8471 5677 8527
rect 7723 8471 7779 8527
rect 7935 8471 7991 8527
rect 7116 8153 7172 8155
rect 7116 8101 7118 8153
rect 7118 8101 7170 8153
rect 7170 8101 7172 8153
rect 7116 8099 7172 8101
rect 7116 7935 7172 7937
rect 7116 7883 7118 7935
rect 7118 7883 7170 7935
rect 7170 7883 7172 7935
rect 7116 7881 7172 7883
rect 4974 7065 5030 7067
rect 4974 7013 4976 7065
rect 4976 7013 5028 7065
rect 5028 7013 5030 7065
rect 4974 7011 5030 7013
rect 4974 6847 5030 6849
rect 4974 6795 4976 6847
rect 4976 6795 5028 6847
rect 5028 6795 5030 6847
rect 4974 6793 5030 6795
rect 4974 6629 5030 6631
rect 4974 6577 4976 6629
rect 4976 6577 5028 6629
rect 5028 6577 5030 6629
rect 4974 6575 5030 6577
rect 5677 7340 5733 7396
rect 5889 7340 5945 7396
rect 7116 7075 7172 7077
rect 7116 7023 7118 7075
rect 7118 7023 7170 7075
rect 7170 7023 7172 7075
rect 7116 7021 7172 7023
rect 6384 6857 6440 6859
rect 6384 6805 6386 6857
rect 6386 6805 6438 6857
rect 6438 6805 6440 6857
rect 6384 6803 6440 6805
rect 6384 6639 6440 6641
rect 6384 6587 6386 6639
rect 6386 6587 6438 6639
rect 6438 6587 6440 6639
rect 6384 6585 6440 6587
rect 6384 6421 6440 6423
rect 6384 6369 6386 6421
rect 6386 6369 6438 6421
rect 6438 6369 6440 6421
rect 6384 6367 6440 6369
rect 7116 6857 7172 6859
rect 7116 6805 7118 6857
rect 7118 6805 7170 6857
rect 7170 6805 7172 6857
rect 7116 6803 7172 6805
rect 7116 6639 7172 6641
rect 7116 6587 7118 6639
rect 7118 6587 7170 6639
rect 7170 6587 7172 6639
rect 7116 6585 7172 6587
rect 7116 6421 7172 6423
rect 7116 6369 7118 6421
rect 7118 6369 7170 6421
rect 7170 6369 7172 6421
rect 7116 6367 7172 6369
rect 5198 5626 5254 5628
rect 5198 5574 5200 5626
rect 5200 5574 5252 5626
rect 5252 5574 5254 5626
rect 5198 5572 5254 5574
rect 5198 5408 5254 5410
rect 5198 5356 5200 5408
rect 5200 5356 5252 5408
rect 5252 5356 5254 5408
rect 5198 5354 5254 5356
rect 6384 5970 6440 5972
rect 6384 5918 6386 5970
rect 6386 5918 6438 5970
rect 6438 5918 6440 5970
rect 6384 5916 6440 5918
rect 6384 5752 6440 5754
rect 6384 5700 6386 5752
rect 6386 5700 6438 5752
rect 6438 5700 6440 5752
rect 6384 5698 6440 5700
rect 8034 3063 8090 3065
rect 8034 2699 8036 3063
rect 8036 2699 8088 3063
rect 8088 2699 8090 3063
rect 8034 2697 8090 2699
rect 8482 3063 8538 3065
rect 8482 2699 8484 3063
rect 8484 2699 8536 3063
rect 8536 2699 8538 3063
rect 8482 2697 8538 2699
rect 10642 9163 10698 9219
rect 10642 8945 10698 9001
rect 11093 9163 11149 9219
rect 11093 8945 11149 9001
rect 11541 9163 11597 9219
rect 11541 8945 11597 9001
rect 12631 4512 12687 4514
rect 12631 4460 12633 4512
rect 12633 4460 12685 4512
rect 12685 4460 12687 4512
rect 12631 4458 12687 4460
rect 12843 4512 12899 4514
rect 12843 4460 12845 4512
rect 12845 4460 12897 4512
rect 12897 4460 12899 4512
rect 12843 4458 12899 4460
rect -347 -2102 -291 -2046
rect -135 -2102 -79 -2046
<< metal3 >>
rect 2733 14544 13946 16283
rect 5986 11295 13946 11359
rect 5986 11239 6312 11295
rect 6368 11239 13946 11295
rect 5986 11077 13946 11239
rect 5986 11021 6312 11077
rect 6368 11021 13946 11077
rect 5986 10860 13946 11021
rect 5986 10804 6312 10860
rect 6368 10804 13946 10860
rect 5986 10642 13946 10804
rect 5986 10586 6312 10642
rect 6368 10629 13946 10642
rect 6368 10595 13638 10629
rect 6368 10586 8859 10595
rect 5986 10539 8859 10586
rect 8915 10539 9307 10595
rect 9363 10539 9755 10595
rect 9811 10539 10203 10595
rect 10259 10539 10651 10595
rect 10707 10539 11099 10595
rect 11155 10539 11547 10595
rect 11603 10539 11995 10595
rect 12051 10539 12443 10595
rect 12499 10539 12891 10595
rect 12947 10539 13337 10595
rect 13393 10573 13638 10595
rect 13694 10573 13946 10629
rect 13393 10539 13946 10573
rect 5986 10424 13946 10539
rect 5986 10368 6312 10424
rect 6368 10411 13946 10424
rect 6368 10377 13638 10411
rect 6368 10368 8859 10377
rect 5986 10321 8859 10368
rect 8915 10321 9307 10377
rect 9363 10321 9755 10377
rect 9811 10321 10203 10377
rect 10259 10321 10651 10377
rect 10707 10321 11099 10377
rect 11155 10321 11547 10377
rect 11603 10321 11995 10377
rect 12051 10321 12443 10377
rect 12499 10321 12891 10377
rect 12947 10321 13337 10377
rect 13393 10355 13638 10377
rect 13694 10355 13946 10411
rect 13393 10321 13946 10355
rect 5986 10264 13946 10321
rect 5986 10208 7068 10264
rect 7124 10208 7515 10264
rect 7571 10208 13946 10264
rect 5986 10207 13946 10208
rect 5986 10151 6312 10207
rect 6368 10193 13946 10207
rect 6368 10159 13638 10193
rect 6368 10151 8859 10159
rect 5986 10103 8859 10151
rect 8915 10103 9307 10159
rect 9363 10103 9755 10159
rect 9811 10103 10203 10159
rect 10259 10103 10651 10159
rect 10707 10103 11099 10159
rect 11155 10103 11547 10159
rect 11603 10103 11995 10159
rect 12051 10103 12443 10159
rect 12499 10103 12891 10159
rect 12947 10103 13337 10159
rect 13393 10137 13638 10159
rect 13694 10137 13946 10193
rect 13393 10103 13946 10137
rect 5986 10046 13946 10103
rect 5986 9990 7068 10046
rect 7124 9990 7515 10046
rect 7571 9990 13946 10046
rect 5986 9989 13946 9990
rect 5986 9933 6312 9989
rect 6368 9975 13946 9989
rect 6368 9941 13638 9975
rect 6368 9933 8859 9941
rect 5986 9885 8859 9933
rect 8915 9885 9307 9941
rect 9363 9885 9755 9941
rect 9811 9885 10203 9941
rect 10259 9885 10651 9941
rect 10707 9885 11099 9941
rect 11155 9885 11547 9941
rect 11603 9885 11995 9941
rect 12051 9885 12443 9941
rect 12499 9885 12891 9941
rect 12947 9885 13337 9941
rect 13393 9919 13638 9941
rect 13694 9919 13946 9975
rect 13393 9885 13946 9919
rect 5986 9828 13946 9885
rect 5986 9772 7068 9828
rect 7124 9772 7515 9828
rect 7571 9772 13946 9828
rect 5986 9610 13946 9772
rect 5986 9554 7068 9610
rect 7124 9554 7515 9610
rect 7571 9554 13946 9610
rect 5986 9541 13946 9554
rect 5986 9511 10061 9541
rect 6548 9257 6888 9258
rect 10607 9257 10733 9258
rect 11058 9257 11184 9258
rect 11506 9257 11632 9258
rect 6497 9219 11632 9257
rect 6497 9163 6584 9219
rect 6640 9163 6796 9219
rect 6852 9163 10642 9219
rect 10698 9163 11093 9219
rect 11149 9163 11541 9219
rect 11597 9163 11632 9219
rect 6497 9001 11632 9163
rect 6497 8945 6584 9001
rect 6640 8945 6796 9001
rect 6852 8945 10642 9001
rect 10698 8945 11093 9001
rect 11149 8945 11541 9001
rect 11597 8945 11632 9001
rect 6497 8906 11632 8945
rect 4611 8760 4951 8799
rect 4611 8704 4647 8760
rect 4703 8704 4859 8760
rect 4915 8704 4951 8760
rect 4611 8665 4951 8704
rect 11812 8582 15246 9368
rect 5373 8527 8027 8566
rect 5373 8471 5409 8527
rect 5465 8471 5621 8527
rect 5677 8471 7723 8527
rect 7779 8471 7935 8527
rect 7991 8471 8027 8527
rect 5373 8428 8027 8471
rect -206 8155 8076 8335
rect -206 8099 7116 8155
rect 7172 8099 8076 8155
rect -206 7937 8076 8099
rect -206 7881 7116 7937
rect 7172 7881 8076 7937
rect -206 7653 8076 7881
rect -319 7396 5981 7435
rect -319 7340 -283 7396
rect -227 7340 -71 7396
rect -15 7340 5677 7396
rect 5733 7340 5889 7396
rect 5945 7340 5981 7396
rect -319 7301 5981 7340
rect 8529 7149 13873 8441
rect 24 7077 13873 7149
rect 24 7067 7116 7077
rect 24 7011 4974 7067
rect 5030 7021 7116 7067
rect 7172 7021 13873 7077
rect 5030 7011 13873 7021
rect 24 6859 13873 7011
rect 24 6849 6384 6859
rect 24 6793 4974 6849
rect 5030 6803 6384 6849
rect 6440 6803 7116 6859
rect 7172 6803 13873 6859
rect 5030 6793 13873 6803
rect 24 6641 13873 6793
rect 24 6631 6384 6641
rect 24 6575 4974 6631
rect 5030 6585 6384 6631
rect 6440 6585 7116 6641
rect 7172 6585 13873 6641
rect 5030 6575 13873 6585
rect 24 6423 13873 6575
rect 24 6367 6384 6423
rect 6440 6367 7116 6423
rect 7172 6367 13873 6423
rect 24 6272 13873 6367
rect 562 5972 13878 6102
rect 562 5916 6384 5972
rect 6440 5916 13878 5972
rect 562 5754 13878 5916
rect 562 5698 6384 5754
rect 6440 5698 13878 5754
rect 562 5628 13878 5698
rect 562 5572 5198 5628
rect 5254 5572 13878 5628
rect 562 5410 13878 5572
rect 562 5354 5198 5410
rect 5254 5354 13878 5410
rect 562 5315 13878 5354
rect 158 4077 9731 4995
rect 12595 4514 12935 4553
rect 12595 4458 12631 4514
rect 12687 4458 12843 4514
rect 12899 4458 12935 4514
rect 12595 4419 12935 4458
rect 12596 4352 12935 4419
rect 12596 4256 17136 4352
rect 158 3740 13783 4077
rect 71 3065 8829 3327
rect 71 2697 8034 3065
rect 8090 2697 8482 3065
rect 8538 2697 8829 3065
rect 71 2265 8829 2697
rect 9223 1450 13783 3740
rect -930 1167 13783 1450
rect 9223 180 13783 1167
rect -930 -109 8587 175
rect -17790 -1261 17624 -806
rect -17790 -1901 15799 -1550
rect -383 -2008 -43 -2007
rect -14200 -2046 15799 -2008
rect -14200 -2102 -347 -2046
rect -291 -2102 -135 -2046
rect -79 -2102 15799 -2046
rect -14200 -2141 15799 -2102
use CON_128x8m81  CON_128x8m81_0
timestamp 1669390400
transform 1 0 6373 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_1
timestamp 1669390400
transform 1 0 6531 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_2
timestamp 1669390400
transform 1 0 6689 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_3
timestamp 1669390400
transform 1 0 6689 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_4
timestamp 1669390400
transform 1 0 6215 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_5
timestamp 1669390400
transform 1 0 6373 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_6
timestamp 1669390400
transform 1 0 6531 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_7
timestamp 1669390400
transform 1 0 6061 0 1 11988
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_8
timestamp 1669390400
transform 1 0 6061 0 1 12151
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_9
timestamp 1669390400
transform 1 0 6061 0 1 12314
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_10
timestamp 1669390400
transform 1 0 6061 0 1 12478
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_11
timestamp 1669390400
transform 1 0 6061 0 1 12641
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_12
timestamp 1669390400
transform 1 0 6061 0 1 12804
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_13
timestamp 1669390400
transform 1 0 6061 0 1 12967
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_14
timestamp 1669390400
transform 1 0 6061 0 1 13130
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_15
timestamp 1669390400
transform 1 0 6061 0 1 13294
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_16
timestamp 1669390400
transform 1 0 6061 0 1 13457
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_17
timestamp 1669390400
transform 1 0 6061 0 1 13620
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_18
timestamp 1669390400
transform 1 0 6061 0 1 13783
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_19
timestamp 1669390400
transform 1 0 6061 0 1 13947
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_20
timestamp 1669390400
transform 1 0 6061 0 1 14110
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_21
timestamp 1669390400
transform 1 0 6061 0 1 14273
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_22
timestamp 1669390400
transform 1 0 6061 0 1 14436
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_23
timestamp 1669390400
transform 1 0 6061 0 1 14599
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_24
timestamp 1669390400
transform 1 0 6061 0 1 14763
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_25
timestamp 1669390400
transform 1 0 6061 0 1 14926
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_26
timestamp 1669390400
transform 1 0 6061 0 1 15089
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_27
timestamp 1669390400
transform 1 0 6061 0 1 15252
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_28
timestamp 1669390400
transform 1 0 6061 0 1 15416
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_29
timestamp 1669390400
transform 1 0 6061 0 1 15579
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_30
timestamp 1669390400
transform 1 0 6061 0 1 15742
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_31
timestamp 1669390400
transform 1 0 6061 0 1 15905
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_32
timestamp 1669390400
transform 1 0 6061 0 1 16069
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_33
timestamp 1669390400
transform 1 0 6215 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_34
timestamp 1669390400
transform 1 0 6847 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_35
timestamp 1669390400
transform 1 0 7005 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_36
timestamp 1669390400
transform 1 0 7163 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_37
timestamp 1669390400
transform 1 0 7321 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_38
timestamp 1669390400
transform 1 0 7480 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_39
timestamp 1669390400
transform 1 0 7638 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_40
timestamp 1669390400
transform 1 0 7796 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_41
timestamp 1669390400
transform 1 0 7954 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_42
timestamp 1669390400
transform 1 0 8112 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_43
timestamp 1669390400
transform 1 0 8270 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_44
timestamp 1669390400
transform 1 0 8428 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_45
timestamp 1669390400
transform 1 0 8586 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_46
timestamp 1669390400
transform 1 0 8744 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_47
timestamp 1669390400
transform 1 0 8903 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_48
timestamp 1669390400
transform 1 0 9061 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_49
timestamp 1669390400
transform 1 0 9219 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_50
timestamp 1669390400
transform 1 0 9377 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_51
timestamp 1669390400
transform 1 0 9535 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_52
timestamp 1669390400
transform 1 0 9693 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_53
timestamp 1669390400
transform 1 0 9851 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_54
timestamp 1669390400
transform 1 0 10009 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_55
timestamp 1669390400
transform 1 0 10167 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_56
timestamp 1669390400
transform 1 0 6847 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_57
timestamp 1669390400
transform 1 0 7005 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_58
timestamp 1669390400
transform 1 0 7163 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_59
timestamp 1669390400
transform 1 0 7321 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_60
timestamp 1669390400
transform 1 0 7480 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_61
timestamp 1669390400
transform 1 0 7638 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_62
timestamp 1669390400
transform 1 0 7796 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_63
timestamp 1669390400
transform 1 0 7954 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_64
timestamp 1669390400
transform 1 0 8112 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_65
timestamp 1669390400
transform 1 0 8270 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_66
timestamp 1669390400
transform 1 0 8428 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_67
timestamp 1669390400
transform 1 0 8586 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_68
timestamp 1669390400
transform 1 0 8744 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_69
timestamp 1669390400
transform 1 0 8903 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_70
timestamp 1669390400
transform 1 0 9061 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_71
timestamp 1669390400
transform 1 0 9219 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_72
timestamp 1669390400
transform 1 0 9377 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_73
timestamp 1669390400
transform 1 0 9535 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_74
timestamp 1669390400
transform 1 0 9693 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_75
timestamp 1669390400
transform 1 0 9851 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_76
timestamp 1669390400
transform 1 0 10009 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_77
timestamp 1669390400
transform 1 0 10167 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_78
timestamp 1669390400
transform 1 0 13655 0 1 11988
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_79
timestamp 1669390400
transform 1 0 13655 0 1 12151
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_80
timestamp 1669390400
transform 1 0 13655 0 1 12314
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_81
timestamp 1669390400
transform 1 0 13655 0 1 12478
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_82
timestamp 1669390400
transform 1 0 13655 0 1 12641
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_83
timestamp 1669390400
transform 1 0 13655 0 1 12804
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_84
timestamp 1669390400
transform 1 0 13655 0 1 12967
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_85
timestamp 1669390400
transform 1 0 13655 0 1 13130
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_86
timestamp 1669390400
transform 1 0 13655 0 1 13294
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_87
timestamp 1669390400
transform 1 0 13655 0 1 13457
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_88
timestamp 1669390400
transform 1 0 13655 0 1 13620
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_89
timestamp 1669390400
transform 1 0 13655 0 1 13783
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_90
timestamp 1669390400
transform 1 0 13655 0 1 13947
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_91
timestamp 1669390400
transform 1 0 13655 0 1 14110
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_92
timestamp 1669390400
transform 1 0 13655 0 1 14273
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_93
timestamp 1669390400
transform 1 0 13655 0 1 14436
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_94
timestamp 1669390400
transform 1 0 13655 0 1 14599
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_95
timestamp 1669390400
transform 1 0 13655 0 1 14763
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_96
timestamp 1669390400
transform 1 0 13655 0 1 14926
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_97
timestamp 1669390400
transform 1 0 13655 0 1 15089
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_98
timestamp 1669390400
transform 1 0 13655 0 1 15252
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_99
timestamp 1669390400
transform 1 0 13655 0 1 15416
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_100
timestamp 1669390400
transform 1 0 13655 0 1 15579
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_101
timestamp 1669390400
transform 1 0 13655 0 1 15742
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_102
timestamp 1669390400
transform 1 0 13655 0 1 15905
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_103
timestamp 1669390400
transform 1 0 13655 0 1 16069
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_104
timestamp 1669390400
transform 1 0 10326 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_105
timestamp 1669390400
transform 1 0 10484 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_106
timestamp 1669390400
transform 1 0 10642 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_107
timestamp 1669390400
transform 1 0 10800 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_108
timestamp 1669390400
transform 1 0 10958 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_109
timestamp 1669390400
transform 1 0 11116 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_110
timestamp 1669390400
transform 1 0 11274 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_111
timestamp 1669390400
transform 1 0 11432 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_112
timestamp 1669390400
transform 1 0 11590 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_113
timestamp 1669390400
transform 1 0 11749 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_114
timestamp 1669390400
transform 1 0 11907 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_115
timestamp 1669390400
transform 1 0 12065 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_116
timestamp 1669390400
transform 1 0 12223 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_117
timestamp 1669390400
transform 1 0 12381 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_118
timestamp 1669390400
transform 1 0 12539 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_119
timestamp 1669390400
transform 1 0 12697 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_120
timestamp 1669390400
transform 1 0 12855 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_121
timestamp 1669390400
transform 1 0 13013 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_122
timestamp 1669390400
transform 1 0 13172 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_123
timestamp 1669390400
transform 1 0 13330 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_124
timestamp 1669390400
transform 1 0 13488 0 1 11938
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_125
timestamp 1669390400
transform 1 0 10326 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_126
timestamp 1669390400
transform 1 0 10484 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_127
timestamp 1669390400
transform 1 0 10642 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_128
timestamp 1669390400
transform 1 0 10800 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_129
timestamp 1669390400
transform 1 0 10958 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_130
timestamp 1669390400
transform 1 0 11116 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_131
timestamp 1669390400
transform 1 0 11274 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_132
timestamp 1669390400
transform 1 0 11432 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_133
timestamp 1669390400
transform 1 0 11590 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_134
timestamp 1669390400
transform 1 0 11749 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_135
timestamp 1669390400
transform 1 0 11907 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_136
timestamp 1669390400
transform 1 0 12065 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_137
timestamp 1669390400
transform 1 0 12223 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_138
timestamp 1669390400
transform 1 0 12381 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_139
timestamp 1669390400
transform 1 0 12539 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_140
timestamp 1669390400
transform 1 0 12697 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_141
timestamp 1669390400
transform 1 0 12855 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_142
timestamp 1669390400
transform 1 0 13013 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_143
timestamp 1669390400
transform 1 0 13172 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_144
timestamp 1669390400
transform 1 0 13330 0 1 16250
box 0 0 1 1
use CON_128x8m81  CON_128x8m81_145
timestamp 1669390400
transform 1 0 13488 0 1 16250
box 0 0 1 1
use M1_NACTIVE4310590548762_128x8m81  M1_NACTIVE4310590548762_128x8m81_0
timestamp 1669390400
transform 1 0 5593 0 1 2510
box -1840 -228 1840 228
use M1_NWELL$$47635500_R90_128x8m81  M1_NWELL$$47635500_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 9084 1 0 7595
box -2105 -300 2105 299
use M1_NWELL$$48078892_128x8m81  M1_NWELL$$48078892_128x8m81_0
timestamp 1669390400
transform -1 0 11140 0 -1 9472
box -2355 -227 2354 228
use M1_NWELL$$48079916_R90_128x8m81  M1_NWELL$$48079916_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 13354 1 0 7187
box -2512 -300 2513 300
use M1_NWELL$$48080940_128x8m81  M1_NWELL$$48080940_128x8m81_0
timestamp 1669390400
transform 1 0 7479 0 1 12591
box -1327 -717 1327 717
use M1_NWELL$$169758764_128x8m81  M1_NWELL$$169758764_128x8m81_0
timestamp 1669390400
transform 1 0 2580 0 1 6728
box -2038 -390 2039 391
use M1_PACTIVE$$48070_R90_128x8m81  M1_PACTIVE$$48070_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 6346 1 0 10149
box -1386 -78 1386 77
use M1_PACTIVE$$48071_R90_128x8m81  M1_PACTIVE$$48071_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 13666 1 0 10757
box -896 -78 896 78
use M1_PACTIVE$$48073_128x8m81  M1_PACTIVE$$48073_128x8m81_0
timestamp 1669390400
transform 0 -1 8147 1 0 9914
box -1386 -157 1386 157
use M1_PACTIVE$$48067628_128x8m81  M1_PACTIVE$$48067628_128x8m81_0
timestamp 1669390400
transform 1 0 4139 0 1 8608
box -3793 -80 3793 80
use M1_PACTIVE$$48072748_128x8m81  M1_PACTIVE$$48072748_128x8m81_0
timestamp 1669390400
transform -1 0 7216 0 -1 11455
box -947 -80 947 80
use M1_PACTIVE$$169762860_128x8m81  M1_PACTIVE$$169762860_128x8m81_0
timestamp 1669390400
transform 1 0 2580 0 1 5745
box -1895 -244 1896 243
use M1_PACTIVE4310590548767_128x8m81  M1_PACTIVE4310590548767_128x8m81_0
timestamp 1669390400
transform 1 0 4037 0 1 4674
box -3742 -342 3742 342
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_0
timestamp 1669390400
transform 1 0 7816 0 1 6010
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_1
timestamp 1669390400
transform 1 0 8088 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_2
timestamp 1669390400
transform 1 0 7570 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_3
timestamp 1669390400
transform 1 0 6930 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_4
timestamp 1669390400
transform 1 0 7157 0 1 5994
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_5
timestamp 1669390400
transform -1 0 5077 0 1 6001
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_6
timestamp 1669390400
transform 1 0 6206 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_7
timestamp 1669390400
transform 1 0 5279 0 1 7055
box 0 0 1 1
use M1_POLY2$$44753964_128x8m81  M1_POLY2$$44753964_128x8m81_8
timestamp 1669390400
transform 1 0 7627 0 1 7409
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_0
timestamp 1669390400
transform 1 0 7851 0 1 7880
box 0 0 1 1
use M1_POLY2$$46559276_128x8m81_0  M1_POLY2$$46559276_128x8m81_0_0
timestamp 1669390400
transform 1 0 5447 0 1 3534
box 0 0 1 1
use M1_POLY2$$46559276_128x8m81_0  M1_POLY2$$46559276_128x8m81_0_1
timestamp 1669390400
transform 1 0 6342 0 1 7368
box 0 0 1 1
use M1_POLY24310590548731_128x8m81  M1_POLY24310590548731_128x8m81_0
timestamp 1669390400
transform 1 0 12411 0 1 4483
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1669390400
transform 1 0 12741 0 1 4265
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1669390400
transform 1 0 12069 0 1 4265
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_2
timestamp 1669390400
transform 1 0 11457 0 1 4514
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_3
timestamp 1669390400
transform 1 0 10786 0 1 4514
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_4
timestamp 1669390400
transform 1 0 5811 0 1 5788
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_0
timestamp 1669390400
transform 1 0 11119 0 1 4296
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1669390400
transform 1 0 9814 0 1 5025
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1669390400
transform 1 0 9591 0 1 5025
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1669390400
transform 1 0 10038 0 1 5025
box 0 0 1 1
use M1_POLY24310590548760_128x8m81  M1_POLY24310590548760_128x8m81_0
timestamp 1669390400
transform 1 0 11141 0 1 12181
box -2157 -42 2157 42
use M1_POLY24310590548761_128x8m81  M1_POLY24310590548761_128x8m81_0
timestamp 1669390400
transform 1 0 11109 0 1 11415
box -2204 -42 2204 42
use M1_POLY24310590548765_128x8m81  M1_POLY24310590548765_128x8m81_0
timestamp 1669390400
transform 1 0 7484 0 1 13359
box -1029 -42 1029 42
use M1_POLY24310590548766_128x8m81  M1_POLY24310590548766_128x8m81_0
timestamp 1669390400
transform 1 0 7212 0 1 11137
box -465 -42 465 42
use M1_PSUB$$48310316_R90_128x8m81  M1_PSUB$$48310316_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 13455 1 0 2086
box -2205 -159 2204 159
use M1_PSUB$$48311340_R90_128x8m81  M1_PSUB$$48311340_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 9028 1 0 2330
box -2449 -159 2449 159
use M1_PSUB$$48312364_128x8m81  M1_PSUB$$48312364_128x8m81_0
timestamp 1669390400
transform 1 0 11321 0 1 -37
box -2294 -83 2294 83
use M1_PSUB$$169764908_128x8m81  M1_PSUB$$169764908_128x8m81_0
timestamp 1669390400
transform -1 0 2323 0 1 8120
box -1977 -245 1977 246
use M2_M1$$34864172_128x8m81  M2_M1$$34864172_128x8m81_0
timestamp 1669390400
transform 1 0 11727 0 1 4264
box 0 0 1 1
use M2_M1$$34864172_128x8m81  M2_M1$$34864172_128x8m81_1
timestamp 1669390400
transform 1 0 12765 0 1 4486
box 0 0 1 1
use M2_M1$$34864172_128x8m81  M2_M1$$34864172_128x8m81_2
timestamp 1669390400
transform 1 0 4972 0 1 5994
box 0 0 1 1
use M2_M1$$34864172_128x8m81  M2_M1$$34864172_128x8m81_3
timestamp 1669390400
transform 1 0 5494 0 1 3532
box 0 0 1 1
use M2_M1$$34864172_R90_128x8m81  M2_M1$$34864172_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 10036 1 0 5026
box 0 0 1 1
use M2_M1$$34864172_R90_128x8m81  M2_M1$$34864172_R90_128x8m81_1
timestamp 1669390400
transform 0 -1 9810 1 0 5026
box 0 0 1 1
use M2_M1$$34864172_R90_128x8m81  M2_M1$$34864172_R90_128x8m81_2
timestamp 1669390400
transform 0 -1 6920 1 0 5983
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1669390400
transform 1 0 6412 0 1 5835
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1669390400
transform -1 0 5457 0 1 6595
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1669390400
transform -1 0 5226 0 1 5491
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_3
timestamp 1669390400
transform 1 0 10148 0 1 8855
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_4
timestamp 1669390400
transform 1 0 7144 0 1 8018
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_5
timestamp 1669390400
transform 1 0 7857 0 1 7293
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_6
timestamp 1669390400
transform 1 0 7857 0 1 7948
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_7
timestamp 1669390400
transform 1 0 9698 0 1 8855
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_8
timestamp 1669390400
transform 1 0 6920 0 1 7087
box 0 0 1 1
use M2_M1$$43375660_R90_128x8m81  M2_M1$$43375660_R90_128x8m81_0
timestamp 1669390400
transform 0 -1 8755 1 0 5182
box 0 0 1 1
use M2_M1$$43375660_R90_128x8m81  M2_M1$$43375660_R90_128x8m81_1
timestamp 1669390400
transform 0 -1 6324 1 0 7365
box 0 0 1 1
use M2_M1$$43375660_R270_128x8m81  M2_M1$$43375660_R270_128x8m81_0
timestamp 1669390400
transform 0 -1 5543 -1 0 7887
box 0 0 1 1
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_0
timestamp 1669390400
transform 1 0 6355 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_1
timestamp 1669390400
transform 1 0 8885 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_2
timestamp 1669390400
transform 1 0 8595 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_3
timestamp 1669390400
transform 1 0 6803 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_4
timestamp 1669390400
transform 1 0 7251 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_5
timestamp 1669390400
transform 1 0 7699 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_6
timestamp 1669390400
transform 1 0 8147 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_7
timestamp 1669390400
transform 1 0 9781 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_8
timestamp 1669390400
transform 1 0 9333 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_9
timestamp 1669390400
transform 1 0 11573 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_10
timestamp 1669390400
transform 1 0 11125 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_11
timestamp 1669390400
transform 1 0 10677 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_12
timestamp 1669390400
transform 1 0 13365 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_13
timestamp 1669390400
transform 1 0 12917 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_14
timestamp 1669390400
transform 1 0 12469 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_15
timestamp 1669390400
transform 1 0 12021 0 1 15450
box -63 -828 64 828
use M2_M1$$43376684_128x8m81  M2_M1$$43376684_128x8m81_16
timestamp 1669390400
transform 1 0 10229 0 1 15450
box -63 -828 64 828
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_0
timestamp 1669390400
transform 1 0 12245 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_1
timestamp 1669390400
transform 1 0 11797 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_2
timestamp 1669390400
transform 1 0 13141 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_3
timestamp 1669390400
transform 1 0 11349 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_4
timestamp 1669390400
transform 1 0 10901 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_5
timestamp 1669390400
transform 1 0 10453 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_6
timestamp 1669390400
transform 1 0 12693 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_7
timestamp 1669390400
transform 1 0 10005 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_8
timestamp 1669390400
transform 1 0 9109 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_9
timestamp 1669390400
transform 1 0 9557 0 1 10625
box 0 0 1 1
use M2_M1$$43378732_128x8m81  M2_M1$$43378732_128x8m81_0
timestamp 1669390400
transform 1 0 6577 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_128x8m81  M2_M1$$43378732_128x8m81_1
timestamp 1669390400
transform 1 0 7921 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_128x8m81  M2_M1$$43378732_128x8m81_2
timestamp 1669390400
transform 1 0 8369 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_128x8m81  M2_M1$$43378732_128x8m81_3
timestamp 1669390400
transform 1 0 7473 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_128x8m81  M2_M1$$43378732_128x8m81_4
timestamp 1669390400
transform 1 0 7025 0 1 13972
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_0
timestamp 1669390400
transform 1 0 12853 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_1
timestamp 1669390400
transform 1 0 11957 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_2
timestamp 1669390400
transform 1 0 12405 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_3
timestamp 1669390400
transform 1 0 13365 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_4
timestamp 1669390400
transform 1 0 12919 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_5
timestamp 1669390400
transform 1 0 11575 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_6
timestamp 1669390400
transform 1 0 12023 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_7
timestamp 1669390400
transform 1 0 12471 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_8
timestamp 1669390400
transform 1 0 13666 0 1 10274
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_9
timestamp 1669390400
transform 1 0 10679 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_10
timestamp 1669390400
transform 1 0 11127 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_11
timestamp 1669390400
transform 1 0 7543 0 1 9909
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_12
timestamp 1669390400
transform 1 0 9783 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_13
timestamp 1669390400
transform 1 0 9335 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_14
timestamp 1669390400
transform 1 0 8887 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_15
timestamp 1669390400
transform 1 0 7096 0 1 9909
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_16
timestamp 1669390400
transform 1 0 10231 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_17
timestamp 1669390400
transform 1 0 7144 0 1 6722
box 0 0 1 1
use M2_M1$$43380780_128x8m81  M2_M1$$43380780_128x8m81_0
timestamp 1669390400
transform 1 0 6412 0 1 6613
box 0 0 1 1
use M2_M1$$43380780_128x8m81  M2_M1$$43380780_128x8m81_1
timestamp 1669390400
transform -1 0 5002 0 1 6821
box 0 0 1 1
use M2_M1$$45013036_128x8m81  M2_M1$$45013036_128x8m81_0
timestamp 1669390400
transform 1 0 6920 0 1 13310
box 0 0 1 1
use M2_M1$$45013036_128x8m81  M2_M1$$45013036_128x8m81_1
timestamp 1669390400
transform 1 0 6950 0 1 11174
box 0 0 1 1
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_0
timestamp 1669390400
transform 1 0 13426 0 1 7395
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_1
timestamp 1669390400
transform 1 0 12179 0 1 7395
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_2
timestamp 1669390400
transform 1 0 12627 0 1 7395
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_3
timestamp 1669390400
transform 1 0 9922 0 1 7390
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_4
timestamp 1669390400
transform 1 0 9474 0 1 7390
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_5
timestamp 1669390400
transform 1 0 11345 0 1 7381
box -64 -1046 64 1046
use M2_M1$$47500332_128x8m81  M2_M1$$47500332_128x8m81_6
timestamp 1669390400
transform 1 0 10897 0 1 7381
box -64 -1046 64 1046
use M2_M1$$47515692_128x8m81  M2_M1$$47515692_128x8m81_0
timestamp 1669390400
transform 1 0 6340 0 1 10614
box 0 0 1 1
use M2_M1$$47515692_128x8m81  M2_M1$$47515692_128x8m81_1
timestamp 1669390400
transform 1 0 7767 0 1 10236
box 0 0 1 1
use M2_M1$$47515692_128x8m81  M2_M1$$47515692_128x8m81_2
timestamp 1669390400
transform 1 0 7319 0 1 10236
box 0 0 1 1
use M2_M1$$47515692_128x8m81  M2_M1$$47515692_128x8m81_3
timestamp 1669390400
transform 1 0 6872 0 1 10236
box 0 0 1 1
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_0
timestamp 1669390400
transform 1 0 11121 0 1 3167
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_1
timestamp 1669390400
transform 1 0 12405 0 1 3167
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_2
timestamp 1669390400
transform 1 0 10005 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_3
timestamp 1669390400
transform 1 0 9557 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_4
timestamp 1669390400
transform 1 0 9109 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_5
timestamp 1669390400
transform 1 0 13141 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_6
timestamp 1669390400
transform 1 0 11797 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_7
timestamp 1669390400
transform 1 0 12245 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_8
timestamp 1669390400
transform 1 0 12693 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_9
timestamp 1669390400
transform 1 0 10453 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_10
timestamp 1669390400
transform 1 0 10901 0 1 13439
box -64 -937 65 937
use M2_M1$$48217132_128x8m81  M2_M1$$48217132_128x8m81_11
timestamp 1669390400
transform 1 0 11349 0 1 13439
box -64 -937 65 937
use M2_M1$$48218156_128x8m81  M2_M1$$48218156_128x8m81_0
timestamp 1669390400
transform 1 0 10117 0 1 12144
box -1013 -67 1013 67
use M2_M1$$48218156_128x8m81  M2_M1$$48218156_128x8m81_1
timestamp 1669390400
transform 1 0 10117 0 1 11451
box -1013 -67 1013 67
use M2_M1$$48219180_128x8m81  M2_M1$$48219180_128x8m81_0
timestamp 1669390400
transform 1 0 9113 0 1 4348
box -170 -393 170 393
use M2_M1$$48220204_128x8m81  M2_M1$$48220204_128x8m81_0
timestamp 1669390400
transform 1 0 9109 0 1 7390
box -170 -1046 170 1046
use M2_M1$$48221228_128x8m81  M2_M1$$48221228_128x8m81_0
timestamp 1669390400
transform 1 0 13541 0 1 2115
box -64 -1917 65 1917
use M2_M1$$48221228_128x8m81  M2_M1$$48221228_128x8m81_1
timestamp 1669390400
transform 1 0 11569 0 1 2115
box -64 -1917 65 1917
use M2_M1$$48221228_128x8m81  M2_M1$$48221228_128x8m81_2
timestamp 1669390400
transform 1 0 11957 0 1 2115
box -64 -1917 65 1917
use M2_M1$$48221228_128x8m81  M2_M1$$48221228_128x8m81_3
timestamp 1669390400
transform 1 0 12853 0 1 2115
box -64 -1917 65 1917
use M2_M1$$48221228_128x8m81  M2_M1$$48221228_128x8m81_4
timestamp 1669390400
transform 1 0 10673 0 1 2115
box -64 -1917 65 1917
use M2_M1$$48222252_128x8m81  M2_M1$$48222252_128x8m81_0
timestamp 1669390400
transform 1 0 11569 0 1 7003
box -65 -2134 65 2134
use M2_M1$$48222252_128x8m81  M2_M1$$48222252_128x8m81_1
timestamp 1669390400
transform 1 0 10673 0 1 7003
box -65 -2134 65 2134
use M2_M1$$48222252_128x8m81  M2_M1$$48222252_128x8m81_2
timestamp 1669390400
transform 1 0 11121 0 1 7003
box -65 -2134 65 2134
use M2_M1$$48224300_128x8m81  M2_M1$$48224300_128x8m81_0
timestamp 1669390400
transform 1 0 8149 0 1 10013
box -169 -502 170 502
use M2_M1$$48316460_128x8m81  M2_M1$$48316460_128x8m81_0
timestamp 1669390400
transform 1 0 9480 0 1 2532
box -65 -2243 65 2243
use M2_M1$$168351788_128x8m81  M2_M1$$168351788_128x8m81_0
timestamp 1669390400
transform 1 0 5815 0 1 5672
box 0 0 1 1
use M2_M1$$170061868_128x8m81  M2_M1$$170061868_128x8m81_0
timestamp 1669390400
transform 1 0 2811 0 1 4584
box -2594 -393 2594 393
use M2_M1$$170063916_128x8m81  M2_M1$$170063916_128x8m81_0
timestamp 1669390400
transform -1 0 2275 0 1 8014
box -1857 -284 1857 284
use M2_M1$$170064940_128x8m81  M2_M1$$170064940_128x8m81_0
timestamp 1669390400
transform -1 0 2561 0 1 5742
box -1857 -176 1857 176
use M2_M1$$170064940_128x8m81  M2_M1$$170064940_128x8m81_1
timestamp 1669390400
transform -1 0 2561 0 1 6726
box -1857 -176 1857 176
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_0
timestamp 1669390400
transform 1 0 13108 0 1 -612
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_1
timestamp 1669390400
transform 1 0 10385 0 1 -612
box 0 0 1 1
use M2_M14310590548726_128x8m81  M2_M14310590548726_128x8m81_0
timestamp 1669390400
transform 1 0 8062 0 1 2881
box 0 0 1 1
use M2_M14310590548726_128x8m81  M2_M14310590548726_128x8m81_1
timestamp 1669390400
transform 1 0 8510 0 1 2881
box 0 0 1 1
use M2_M14310590548764_128x8m81  M2_M14310590548764_128x8m81_0
timestamp 1669390400
transform 1 0 5060 0 1 2506
box -2546 -236 2546 236
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_0
timestamp 1669390400
transform 1 0 6412 0 1 5835
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_1
timestamp 1669390400
transform -1 0 5226 0 1 5491
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_2
timestamp 1669390400
transform 1 0 11569 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_3
timestamp 1669390400
transform 1 0 11121 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_4
timestamp 1669390400
transform 1 0 10670 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_5
timestamp 1669390400
transform 1 0 7144 0 1 8018
box 0 0 1 1
use M3_M2$$43368492_R270_128x8m81  M3_M2$$43368492_R270_128x8m81_0
timestamp 1669390400
transform 0 -1 5543 -1 0 8499
box 0 0 1 1
use M3_M2$$43368492_R270_128x8m81  M3_M2$$43368492_R270_128x8m81_1
timestamp 1669390400
transform 0 -1 7857 -1 0 8499
box 0 0 1 1
use M3_M2$$43371564_128x8m81  M3_M2$$43371564_128x8m81_0
timestamp 1669390400
transform 1 0 12765 0 1 4486
box 0 0 1 1
use M3_M2$$43371564_128x8m81  M3_M2$$43371564_128x8m81_1
timestamp 1669390400
transform 1 0 -149 0 1 7368
box 0 0 1 1
use M3_M2$$43371564_128x8m81  M3_M2$$43371564_128x8m81_2
timestamp 1669390400
transform 1 0 4781 0 1 8732
box 0 0 1 1
use M3_M2$$43371564_128x8m81  M3_M2$$43371564_128x8m81_3
timestamp 1669390400
transform 1 0 5811 0 1 7368
box 0 0 1 1
use M3_M2$$45008940_128x8m81  M3_M2$$45008940_128x8m81_0
timestamp 1669390400
transform 1 0 6718 0 1 9082
box 0 0 1 1
use M3_M2$$47108140_128x8m81  M3_M2$$47108140_128x8m81_0
timestamp 1669390400
transform 1 0 6412 0 1 6613
box 0 0 1 1
use M3_M2$$47108140_128x8m81  M3_M2$$47108140_128x8m81_1
timestamp 1669390400
transform -1 0 5002 0 1 6821
box 0 0 1 1
use M3_M2$$47115308_128x8m81  M3_M2$$47115308_128x8m81_0
timestamp 1669390400
transform 1 0 9113 0 1 4348
box -170 -393 170 393
use M3_M2$$47332396_128x8m81  M3_M2$$47332396_128x8m81_0
timestamp 1669390400
transform 1 0 6340 0 1 10614
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_0
timestamp 1669390400
transform 1 0 12023 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_1
timestamp 1669390400
transform 1 0 11575 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_2
timestamp 1669390400
transform 1 0 12919 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_3
timestamp 1669390400
transform 1 0 13365 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_4
timestamp 1669390400
transform 1 0 13666 0 1 10274
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_5
timestamp 1669390400
transform 1 0 11127 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_6
timestamp 1669390400
transform 1 0 10679 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_7
timestamp 1669390400
transform 1 0 12471 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_8
timestamp 1669390400
transform 1 0 9783 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_9
timestamp 1669390400
transform 1 0 7096 0 1 9909
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_10
timestamp 1669390400
transform 1 0 7543 0 1 9909
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_11
timestamp 1669390400
transform 1 0 8887 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_12
timestamp 1669390400
transform 1 0 9335 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_13
timestamp 1669390400
transform 1 0 10231 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_14
timestamp 1669390400
transform 1 0 7144 0 1 6722
box 0 0 1 1
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_0
timestamp 1669390400
transform 1 0 12179 0 1 7395
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_1
timestamp 1669390400
transform 1 0 12627 0 1 7395
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_2
timestamp 1669390400
transform 1 0 9922 0 1 7390
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_3
timestamp 1669390400
transform 1 0 9474 0 1 7390
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_4
timestamp 1669390400
transform 1 0 11345 0 1 7381
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_5
timestamp 1669390400
transform 1 0 10897 0 1 7381
box -65 -1046 65 1046
use M3_M2$$47644716_128x8m81  M3_M2$$47644716_128x8m81_6
timestamp 1669390400
transform 1 0 13426 0 1 7395
box -65 -1046 65 1046
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_0
timestamp 1669390400
transform 1 0 6355 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_1
timestamp 1669390400
transform 1 0 8595 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_2
timestamp 1669390400
transform 1 0 6803 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_3
timestamp 1669390400
transform 1 0 7251 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_4
timestamp 1669390400
transform 1 0 7699 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_5
timestamp 1669390400
transform 1 0 8147 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_6
timestamp 1669390400
transform 1 0 9333 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_7
timestamp 1669390400
transform 1 0 8885 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_8
timestamp 1669390400
transform 1 0 9781 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_9
timestamp 1669390400
transform 1 0 10677 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_10
timestamp 1669390400
transform 1 0 13365 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_11
timestamp 1669390400
transform 1 0 12917 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_12
timestamp 1669390400
transform 1 0 12469 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_13
timestamp 1669390400
transform 1 0 12021 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_14
timestamp 1669390400
transform 1 0 11573 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_15
timestamp 1669390400
transform 1 0 11125 0 1 15450
box -65 -828 65 828
use M3_M2$$47645740_128x8m81  M3_M2$$47645740_128x8m81_16
timestamp 1669390400
transform 1 0 10229 0 1 15450
box -65 -828 65 828
use M3_M2$$48066604_128x8m81  M3_M2$$48066604_128x8m81_0
timestamp 1669390400
transform 1 0 12508 0 1 8975
box -697 -393 697 393
use M3_M2$$48227372_128x8m81  M3_M2$$48227372_128x8m81_0
timestamp 1669390400
transform 1 0 9480 0 1 2532
box -65 -2243 65 2243
use M3_M2$$48228396_128x8m81  M3_M2$$48228396_128x8m81_0
timestamp 1669390400
transform 1 0 9109 0 1 7390
box -170 -1046 170 1046
use M3_M2$$48229420_128x8m81  M3_M2$$48229420_128x8m81_0
timestamp 1669390400
transform 1 0 11569 0 1 2115
box -65 -1917 65 1917
use M3_M2$$48229420_128x8m81  M3_M2$$48229420_128x8m81_1
timestamp 1669390400
transform 1 0 11957 0 1 2115
box -65 -1917 65 1917
use M3_M2$$48229420_128x8m81  M3_M2$$48229420_128x8m81_2
timestamp 1669390400
transform 1 0 12853 0 1 2115
box -65 -1917 65 1917
use M3_M2$$48229420_128x8m81  M3_M2$$48229420_128x8m81_3
timestamp 1669390400
transform 1 0 10673 0 1 2115
box -65 -1917 65 1917
use M3_M2$$48229420_128x8m81  M3_M2$$48229420_128x8m81_4
timestamp 1669390400
transform 1 0 13541 0 1 2115
box -65 -1917 65 1917
use M3_M2$$48231468_128x8m81  M3_M2$$48231468_128x8m81_0
timestamp 1669390400
transform 1 0 8149 0 1 10013
box -170 -502 170 502
use M3_M2$$169753644_128x8m81  M3_M2$$169753644_128x8m81_0
timestamp 1669390400
transform 1 0 2811 0 1 4584
box -2594 -393 2594 393
use M3_M2$$169755692_128x8m81  M3_M2$$169755692_128x8m81_0
timestamp 1669390400
transform -1 0 2275 0 1 8014
box -1857 -284 1857 284
use M3_M2$$169756716_128x8m81  M3_M2$$169756716_128x8m81_0
timestamp 1669390400
transform -1 0 2561 0 1 6726
box -1857 -176 1857 176
use M3_M2$$169756716_128x8m81  M3_M2$$169756716_128x8m81_1
timestamp 1669390400
transform -1 0 2561 0 1 5742
box -1857 -176 1857 176
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_0
timestamp 1669390400
transform 1 0 -213 0 1 -2074
box 0 0 1 1
use M3_M24310590548727_128x8m81  M3_M24310590548727_128x8m81_0
timestamp 1669390400
transform 1 0 8062 0 1 2881
box 0 0 1 1
use M3_M24310590548727_128x8m81  M3_M24310590548727_128x8m81_1
timestamp 1669390400
transform 1 0 8510 0 1 2881
box 0 0 1 1
use M3_M24310590548763_128x8m81  M3_M24310590548763_128x8m81_0
timestamp 1669390400
transform 1 0 5060 0 1 2506
box -2546 -236 2546 236
use nmos_1p2$$46551084_128x8m81  nmos_1p2$$46551084_128x8m81_0
timestamp 1669390400
transform 1 0 7517 0 1 5402
box -119 -73 177 527
use nmos_1p2$$46563372_128x8m81  nmos_1p2$$46563372_128x8m81_0
timestamp 1669390400
transform 1 0 5086 0 1 7941
box -119 -74 177 264
use nmos_1p2$$46563372_128x8m81  nmos_1p2$$46563372_128x8m81_1
timestamp 1669390400
transform 1 0 7517 0 -1 8213
box -119 -74 177 264
use nmos_1p2$$46563372_128x8m81  nmos_1p2$$46563372_128x8m81_2
timestamp 1669390400
transform 1 0 7003 0 -1 8213
box -119 -74 177 264
use nmos_1p2$$47342636_128x8m81  nmos_1p2$$47342636_128x8m81_0
timestamp 1669390400
transform 1 0 5310 0 1 5402
box -119 -73 177 316
use nmos_1p2$$47342636_128x8m81  nmos_1p2$$47342636_128x8m81_1
timestamp 1669390400
transform 1 0 5086 0 1 5402
box -119 -73 177 316
use nmos_1p2$$48302124_128x8m81  nmos_1p2$$48302124_128x8m81_0
timestamp 1669390400
transform 1 0 8145 0 -1 4393
box -119 -74 177 677
use nmos_1p2$$48306220_128x8m81  nmos_1p2$$48306220_128x8m81_0
timestamp 1669390400
transform 1 0 6731 0 1 9039
box -119 -74 1073 2040
use nmos_1p2$$48308268_128x8m81  nmos_1p2$$48308268_128x8m81_0
timestamp 1669390400
transform 1 0 8968 0 1 9839
box -119 -44 4433 1518
use nmos_1p2$$48629804_128x8m81  nmos_1p2$$48629804_128x8m81_0
timestamp 1669390400
transform 1 0 6779 0 1 5402
box -119 -73 401 527
use nmos_5p04310590548787_128x8m81  nmos_5p04310590548787_128x8m81_0
timestamp 1669390400
transform 1 0 7600 0 -1 3940
box -88 -44 208 194
use nmos_5p04310590548794_128x8m81  nmos_5p04310590548794_128x8m81_0
timestamp 1669390400
transform 1 0 6954 0 -1 3897
box -88 -44 288 164
use nmos_5p04310590548797_128x8m81  nmos_5p04310590548797_128x8m81_0
timestamp 1669390400
transform 1 0 5157 0 -1 3892
box -88 -44 328 164
use nmos_5p04310590548797_128x8m81  nmos_5p04310590548797_128x8m81_1
timestamp 1669390400
transform 1 0 6235 0 -1 3892
box -88 -44 328 164
use pmos_1p2$$46273580_128x8m81  pmos_1p2$$46273580_128x8m81_0
timestamp 1669390400
transform 1 0 6779 0 -1 7742
box -286 -142 568 348
use pmos_1p2$$46285868_128x8m81  pmos_1p2$$46285868_128x8m81_0
timestamp 1669390400
transform 1 0 5086 0 1 7195
box -286 -142 344 595
use pmos_1p2$$46285868_128x8m81  pmos_1p2$$46285868_128x8m81_1
timestamp 1669390400
transform 1 0 7517 0 1 6377
box -286 -142 344 595
use pmos_1p2$$47330348_128x8m81  pmos_1p2$$47330348_128x8m81_0
timestamp 1669390400
transform 1 0 7517 0 -1 7742
box -286 -141 344 332
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_0
timestamp 1669390400
transform 1 0 12489 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_1
timestamp 1669390400
transform 1 0 12713 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_2
timestamp 1669390400
transform 1 0 12265 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_3
timestamp 1669390400
transform 1 0 12041 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_4
timestamp 1669390400
transform 1 0 11428 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_5
timestamp 1669390400
transform 1 0 10980 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_6
timestamp 1669390400
transform 1 0 10756 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$47815724_128x8m81  pmos_1p2$$47815724_128x8m81_7
timestamp 1669390400
transform 1 0 11204 0 1 4659
box -286 -141 344 4676
use pmos_1p2$$48623660_128x8m81  pmos_1p2$$48623660_128x8m81_0
timestamp 1669390400
transform 1 0 8145 0 -1 3260
box -286 -142 568 894
use pmos_1p2$$48624684_128x8m81  pmos_1p2$$48624684_128x8m81_0
timestamp 1669390400
transform 1 0 10005 0 1 5293
box -286 -141 344 4041
use pmos_1p2$$48624684_128x8m81  pmos_1p2$$48624684_128x8m81_1
timestamp 1669390400
transform 1 0 9557 0 1 5293
box -286 -141 344 4041
use pmos_1p2$$48624684_128x8m81  pmos_1p2$$48624684_128x8m81_2
timestamp 1669390400
transform 1 0 9781 0 1 5293
box -286 -141 344 4041
use pmos_5p04310590548751_128x8m81  pmos_5p04310590548751_128x8m81_0
timestamp 1669390400
transform 1 0 6748 0 1 6137
box -208 -120 552 1254
use pmos_5p04310590548778_128x8m81  pmos_5p04310590548778_128x8m81_0
timestamp 1669390400
transform 1 0 5157 0 -1 3260
box -208 -120 448 300
use pmos_5p04310590548778_128x8m81  pmos_5p04310590548778_128x8m81_1
timestamp 1669390400
transform 1 0 6235 0 -1 3260
box -208 -120 448 300
use pmos_5p04310590548792_128x8m81  pmos_5p04310590548792_128x8m81_0
timestamp 1669390400
transform 1 0 6408 0 1 13461
box -208 -120 2344 2616
use pmos_5p04310590548793_128x8m81  pmos_5p04310590548793_128x8m81_0
timestamp 1669390400
transform 1 0 8937 0 1 12283
box -208 -120 4584 3794
use pmos_5p04310590548796_128x8m81  pmos_5p04310590548796_128x8m81_0
timestamp 1669390400
transform 1 0 6954 0 -1 3260
box -208 -120 408 300
use pmos_5p04310590548798_128x8m81  pmos_5p04310590548798_128x8m81_0
timestamp 1669390400
transform 1 0 7600 0 -1 3260
box -208 -120 328 498
use wen_v2_128x8m81  wen_v2_128x8m81_0
timestamp 1669390400
transform 1 0 -16 0 1 -2104
box -27 -266 7407 3658
<< labels >>
flabel metal3 s 847 5774 847 5774 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
flabel metal3 s 320 4011 320 4011 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
flabel metal3 s 429 6678 429 6678 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal3 s 847 8050 847 8050 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
flabel metal3 s -445 -1708 -445 -1708 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
rlabel metal3 s 12652 4305 12652 4305 4 tblhl
port 3 nsew
flabel metal3 s 6414 10067 6414 10067 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
flabel metal3 s -445 -1060 -445 -1060 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal3 s -445 -26 -445 -26 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal3 s 344 2456 344 2456 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6414 15414 6414 15414 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal3 s -445 1250 -445 1250 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
rlabel metal2 s 8753 -181 8753 -181 4 cen
port 4 nsew
rlabel metal2 s -215 7409 -215 7409 4 clk
port 5 nsew
rlabel metal2 s 12456 13280 12456 13280 4 men
port 6 nsew
flabel metal1 s 529 -493 529 -493 0 FreeSans 1000 0 0 0 WEN
port 7 nsew
flabel metal1 s 6616 1004 6616 1004 0 FreeSans 1000 0 0 0 GWE
port 8 nsew
<< properties >>
string GDS_END 1566384
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1519784
string path 25.525 19.160 25.525 21.230 
<< end >>
