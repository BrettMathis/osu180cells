magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 4100 1230
<< nmos >>
rect 190 190 250 360
rect 540 190 600 360
rect 710 190 770 360
rect 820 190 880 360
rect 1220 190 1280 360
rect 1430 190 1490 360
rect 1660 190 1720 360
rect 1770 190 1830 360
rect 1940 190 2000 360
rect 2050 190 2110 360
rect 2280 190 2340 360
rect 2490 190 2550 360
rect 2660 190 2720 360
rect 3040 190 3100 360
rect 3150 190 3210 360
rect 3320 190 3380 360
rect 3670 190 3730 360
rect 3840 190 3900 360
<< pmos >>
rect 190 700 250 1040
rect 510 700 570 1040
rect 680 700 740 1040
rect 850 700 910 1040
rect 1220 700 1280 1040
rect 1430 700 1490 1040
rect 1660 700 1720 1040
rect 1770 700 1830 1040
rect 1940 700 2000 1040
rect 2050 700 2110 1040
rect 2280 700 2340 1040
rect 2490 700 2550 1040
rect 2660 700 2720 1040
rect 3010 700 3070 1040
rect 3180 700 3240 1040
rect 3350 700 3410 1040
rect 3670 700 3730 1040
rect 3840 700 3900 1040
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 350 360
rect 250 252 282 298
rect 328 252 350 298
rect 250 190 350 252
rect 440 258 540 360
rect 440 212 462 258
rect 508 212 540 258
rect 440 190 540 212
rect 600 283 710 360
rect 600 237 632 283
rect 678 237 710 283
rect 600 190 710 237
rect 770 190 820 360
rect 880 263 980 360
rect 880 217 912 263
rect 958 217 980 263
rect 880 190 980 217
rect 1120 263 1220 360
rect 1120 217 1142 263
rect 1188 217 1220 263
rect 1120 190 1220 217
rect 1280 190 1430 360
rect 1490 263 1660 360
rect 1490 217 1552 263
rect 1598 217 1660 263
rect 1490 190 1660 217
rect 1720 190 1770 360
rect 1830 258 1940 360
rect 1830 212 1862 258
rect 1908 212 1940 258
rect 1830 190 1940 212
rect 2000 190 2050 360
rect 2110 258 2280 360
rect 2110 212 2172 258
rect 2218 212 2280 258
rect 2110 190 2280 212
rect 2340 190 2490 360
rect 2550 283 2660 360
rect 2550 237 2582 283
rect 2628 237 2660 283
rect 2550 190 2660 237
rect 2720 298 2820 360
rect 2720 252 2752 298
rect 2798 252 2820 298
rect 2720 190 2820 252
rect 2940 298 3040 360
rect 2940 252 2962 298
rect 3008 252 3040 298
rect 2940 190 3040 252
rect 3100 190 3150 360
rect 3210 273 3320 360
rect 3210 227 3242 273
rect 3288 227 3320 273
rect 3210 190 3320 227
rect 3380 258 3480 360
rect 3380 212 3412 258
rect 3458 212 3480 258
rect 3380 190 3480 212
rect 3570 298 3670 360
rect 3570 252 3592 298
rect 3638 252 3670 298
rect 3570 190 3670 252
rect 3730 278 3840 360
rect 3730 232 3762 278
rect 3808 232 3840 278
rect 3730 190 3840 232
rect 3900 298 4000 360
rect 3900 252 3932 298
rect 3978 252 4000 298
rect 3900 190 4000 252
<< pdiff >>
rect 90 987 190 1040
rect 90 753 112 987
rect 158 753 190 987
rect 90 700 190 753
rect 250 987 350 1040
rect 250 753 282 987
rect 328 753 350 987
rect 250 700 350 753
rect 410 1020 510 1040
rect 410 880 432 1020
rect 478 880 510 1020
rect 410 700 510 880
rect 570 1015 680 1040
rect 570 875 602 1015
rect 648 875 680 1015
rect 570 700 680 875
rect 740 1015 850 1040
rect 740 875 772 1015
rect 818 875 850 1015
rect 740 700 850 875
rect 910 1015 1010 1040
rect 910 875 942 1015
rect 988 875 1010 1015
rect 910 700 1010 875
rect 1120 1018 1220 1040
rect 1120 972 1142 1018
rect 1188 972 1220 1018
rect 1120 700 1220 972
rect 1280 700 1430 1040
rect 1490 1010 1660 1040
rect 1490 870 1552 1010
rect 1598 870 1660 1010
rect 1490 700 1660 870
rect 1720 700 1770 1040
rect 1830 1000 1940 1040
rect 1830 860 1862 1000
rect 1908 860 1940 1000
rect 1830 700 1940 860
rect 2000 700 2050 1040
rect 2110 1007 2280 1040
rect 2110 773 2172 1007
rect 2218 773 2280 1007
rect 2110 700 2280 773
rect 2340 700 2490 1040
rect 2550 1018 2660 1040
rect 2550 972 2582 1018
rect 2628 972 2660 1018
rect 2550 700 2660 972
rect 2720 997 2820 1040
rect 2720 763 2752 997
rect 2798 763 2820 997
rect 2720 700 2820 763
rect 2910 1015 3010 1040
rect 2910 875 2932 1015
rect 2978 875 3010 1015
rect 2910 700 3010 875
rect 3070 1015 3180 1040
rect 3070 875 3102 1015
rect 3148 875 3180 1015
rect 3070 700 3180 875
rect 3240 1015 3350 1040
rect 3240 875 3272 1015
rect 3318 875 3350 1015
rect 3240 700 3350 875
rect 3410 1020 3510 1040
rect 3410 880 3442 1020
rect 3488 880 3510 1020
rect 3410 700 3510 880
rect 3570 992 3670 1040
rect 3570 758 3592 992
rect 3638 758 3670 992
rect 3570 700 3670 758
rect 3730 995 3840 1040
rect 3730 855 3762 995
rect 3808 855 3840 995
rect 3730 700 3840 855
rect 3900 987 4000 1040
rect 3900 753 3932 987
rect 3978 753 4000 987
rect 3900 700 4000 753
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 462 212 508 258
rect 632 237 678 283
rect 912 217 958 263
rect 1142 217 1188 263
rect 1552 217 1598 263
rect 1862 212 1908 258
rect 2172 212 2218 258
rect 2582 237 2628 283
rect 2752 252 2798 298
rect 2962 252 3008 298
rect 3242 227 3288 273
rect 3412 212 3458 258
rect 3592 252 3638 298
rect 3762 232 3808 278
rect 3932 252 3978 298
<< pdiffc >>
rect 112 753 158 987
rect 282 753 328 987
rect 432 880 478 1020
rect 602 875 648 1015
rect 772 875 818 1015
rect 942 875 988 1015
rect 1142 972 1188 1018
rect 1552 870 1598 1010
rect 1862 860 1908 1000
rect 2172 773 2218 1007
rect 2582 972 2628 1018
rect 2752 763 2798 997
rect 2932 875 2978 1015
rect 3102 875 3148 1015
rect 3272 875 3318 1015
rect 3442 880 3488 1020
rect 3592 758 3638 992
rect 3762 855 3808 995
rect 3932 753 3978 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 340 98 430 120
rect 340 52 362 98
rect 408 52 430 98
rect 340 30 430 52
rect 580 98 670 120
rect 580 52 602 98
rect 648 52 670 98
rect 580 30 670 52
rect 820 98 910 120
rect 820 52 842 98
rect 888 52 910 98
rect 820 30 910 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
rect 2730 98 2820 120
rect 2730 52 2752 98
rect 2798 52 2820 98
rect 2730 30 2820 52
rect 2970 98 3060 120
rect 2970 52 2992 98
rect 3038 52 3060 98
rect 2970 30 3060 52
rect 3210 98 3300 120
rect 3210 52 3232 98
rect 3278 52 3300 98
rect 3210 30 3300 52
rect 3450 98 3540 120
rect 3450 52 3472 98
rect 3518 52 3540 98
rect 3450 30 3540 52
rect 3690 98 3780 120
rect 3690 52 3712 98
rect 3758 52 3780 98
rect 3690 30 3780 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 340 1178 430 1200
rect 340 1132 362 1178
rect 408 1132 430 1178
rect 340 1110 430 1132
rect 580 1178 670 1200
rect 580 1132 602 1178
rect 648 1132 670 1178
rect 580 1110 670 1132
rect 820 1178 910 1200
rect 820 1132 842 1178
rect 888 1132 910 1178
rect 820 1110 910 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
rect 1290 1178 1380 1200
rect 1290 1132 1312 1178
rect 1358 1132 1380 1178
rect 1290 1110 1380 1132
rect 1530 1178 1620 1200
rect 1530 1132 1552 1178
rect 1598 1132 1620 1178
rect 1530 1110 1620 1132
rect 1770 1178 1860 1200
rect 1770 1132 1792 1178
rect 1838 1132 1860 1178
rect 1770 1110 1860 1132
rect 2010 1178 2100 1200
rect 2010 1132 2032 1178
rect 2078 1132 2100 1178
rect 2010 1110 2100 1132
rect 2250 1178 2340 1200
rect 2250 1132 2272 1178
rect 2318 1132 2340 1178
rect 2250 1110 2340 1132
rect 2490 1178 2580 1200
rect 2490 1132 2512 1178
rect 2558 1132 2580 1178
rect 2490 1110 2580 1132
rect 2730 1178 2820 1200
rect 2730 1132 2752 1178
rect 2798 1132 2820 1178
rect 2730 1110 2820 1132
rect 2970 1178 3060 1200
rect 2970 1132 2992 1178
rect 3038 1132 3060 1178
rect 2970 1110 3060 1132
rect 3210 1178 3300 1200
rect 3210 1132 3232 1178
rect 3278 1132 3300 1178
rect 3210 1110 3300 1132
rect 3450 1178 3540 1200
rect 3450 1132 3472 1178
rect 3518 1132 3540 1178
rect 3450 1110 3540 1132
rect 3690 1178 3780 1200
rect 3690 1132 3712 1178
rect 3758 1132 3780 1178
rect 3690 1110 3780 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 362 52 408 98
rect 602 52 648 98
rect 842 52 888 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
rect 2752 52 2798 98
rect 2992 52 3038 98
rect 3232 52 3278 98
rect 3472 52 3518 98
rect 3712 52 3758 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 362 1132 408 1178
rect 602 1132 648 1178
rect 842 1132 888 1178
rect 1072 1132 1118 1178
rect 1312 1132 1358 1178
rect 1552 1132 1598 1178
rect 1792 1132 1838 1178
rect 2032 1132 2078 1178
rect 2272 1132 2318 1178
rect 2512 1132 2558 1178
rect 2752 1132 2798 1178
rect 2992 1132 3038 1178
rect 3232 1132 3278 1178
rect 3472 1132 3518 1178
rect 3712 1132 3758 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 510 1040 570 1090
rect 680 1040 740 1090
rect 850 1040 910 1090
rect 1220 1040 1280 1090
rect 1430 1040 1490 1090
rect 1660 1040 1720 1090
rect 1770 1040 1830 1090
rect 1940 1040 2000 1090
rect 2050 1040 2110 1090
rect 2280 1040 2340 1090
rect 2490 1040 2550 1090
rect 2660 1040 2720 1090
rect 3010 1040 3070 1090
rect 3180 1040 3240 1090
rect 3350 1040 3410 1090
rect 3670 1040 3730 1090
rect 3840 1040 3900 1090
rect 190 650 250 700
rect 140 623 250 650
rect 140 577 167 623
rect 213 577 250 623
rect 140 550 250 577
rect 190 360 250 550
rect 510 520 570 700
rect 680 680 740 700
rect 850 680 910 700
rect 680 653 800 680
rect 680 607 707 653
rect 753 607 800 653
rect 680 580 800 607
rect 850 653 990 680
rect 850 607 907 653
rect 953 607 990 653
rect 1220 650 1280 700
rect 1430 680 1490 700
rect 1360 653 1490 680
rect 850 580 990 607
rect 1200 623 1310 650
rect 510 493 630 520
rect 510 447 557 493
rect 603 447 630 493
rect 510 420 630 447
rect 680 430 740 580
rect 850 430 910 580
rect 1200 577 1237 623
rect 1283 577 1310 623
rect 1360 607 1387 653
rect 1433 650 1490 653
rect 1433 607 1460 650
rect 1360 580 1460 607
rect 1660 600 1720 700
rect 1770 680 1830 700
rect 1940 680 2000 700
rect 1770 610 2000 680
rect 2050 610 2110 700
rect 2280 680 2340 700
rect 2280 653 2400 680
rect 2280 650 2327 653
rect 1200 550 1310 577
rect 1510 550 1720 600
rect 540 360 600 420
rect 680 380 770 430
rect 710 360 770 380
rect 820 390 910 430
rect 820 360 880 390
rect 1220 360 1280 550
rect 1510 510 1570 550
rect 1390 483 1570 510
rect 1390 437 1427 483
rect 1473 437 1570 483
rect 1390 410 1570 437
rect 1620 478 1720 500
rect 1850 480 1910 610
rect 2050 560 2250 610
rect 2300 607 2327 650
rect 2373 607 2400 653
rect 2300 580 2400 607
rect 2490 570 2550 700
rect 2660 650 2720 700
rect 2660 623 2760 650
rect 2660 577 2687 623
rect 2733 577 2760 623
rect 2200 530 2250 560
rect 2470 543 2570 570
rect 1620 432 1647 478
rect 1693 432 1720 478
rect 1620 410 1720 432
rect 1430 360 1490 410
rect 1660 360 1720 410
rect 1770 460 1910 480
rect 2050 488 2150 510
rect 1770 453 2000 460
rect 1770 407 1807 453
rect 1853 407 2000 453
rect 1770 380 2000 407
rect 1770 360 1830 380
rect 1940 360 2000 380
rect 2050 442 2077 488
rect 2123 442 2150 488
rect 2200 503 2370 530
rect 2200 460 2287 503
rect 2050 420 2150 442
rect 2260 457 2287 460
rect 2333 457 2370 503
rect 2470 497 2497 543
rect 2543 497 2570 543
rect 2470 470 2570 497
rect 2660 550 2760 577
rect 2260 430 2370 457
rect 2050 360 2110 420
rect 2280 360 2340 430
rect 2490 360 2550 470
rect 2660 360 2720 550
rect 3010 490 3070 700
rect 2910 463 3070 490
rect 2910 417 2947 463
rect 2993 460 3070 463
rect 3180 650 3240 700
rect 3180 623 3280 650
rect 3180 577 3207 623
rect 3253 577 3280 623
rect 3180 550 3280 577
rect 2993 417 3100 460
rect 3180 430 3240 550
rect 3350 500 3410 700
rect 3670 590 3730 700
rect 3840 670 3900 700
rect 2910 390 3100 417
rect 3040 360 3100 390
rect 3150 380 3240 430
rect 3300 478 3410 500
rect 3620 563 3730 590
rect 3790 648 3900 670
rect 3790 602 3812 648
rect 3858 602 3900 648
rect 3790 580 3900 602
rect 3620 517 3647 563
rect 3693 517 3730 563
rect 3620 490 3730 517
rect 3300 432 3327 478
rect 3373 432 3410 478
rect 3300 410 3410 432
rect 3150 360 3210 380
rect 3320 360 3380 410
rect 3670 360 3730 490
rect 3840 360 3900 580
rect 190 140 250 190
rect 540 140 600 190
rect 710 140 770 190
rect 820 140 880 190
rect 1220 140 1280 190
rect 1430 140 1490 190
rect 1660 140 1720 190
rect 1770 140 1830 190
rect 1940 140 2000 190
rect 2050 140 2110 190
rect 2280 140 2340 190
rect 2490 140 2550 190
rect 2660 140 2720 190
rect 3040 140 3100 190
rect 3150 140 3210 190
rect 3320 140 3380 190
rect 3670 140 3730 190
rect 3840 140 3900 190
<< polycontact >>
rect 167 577 213 623
rect 707 607 753 653
rect 907 607 953 653
rect 557 447 603 493
rect 1237 577 1283 623
rect 1387 607 1433 653
rect 1427 437 1473 483
rect 2327 607 2373 653
rect 2687 577 2733 623
rect 1647 432 1693 478
rect 1807 407 1853 453
rect 2077 442 2123 488
rect 2287 457 2333 503
rect 2497 497 2543 543
rect 2947 417 2993 463
rect 3207 577 3253 623
rect 3812 602 3858 648
rect 3647 517 3693 563
rect 3327 432 3373 478
<< metal1 >>
rect 0 1178 4100 1230
rect 0 1132 112 1178
rect 158 1176 362 1178
rect 408 1176 602 1178
rect 648 1176 842 1178
rect 0 1124 114 1132
rect 166 1124 354 1176
rect 408 1132 594 1176
rect 648 1132 834 1176
rect 888 1132 1072 1178
rect 1118 1176 1312 1178
rect 1358 1176 1552 1178
rect 1598 1176 1792 1178
rect 1838 1176 2032 1178
rect 2078 1176 2272 1178
rect 2318 1176 2512 1178
rect 2558 1176 2752 1178
rect 2798 1176 2992 1178
rect 3038 1176 3232 1178
rect 3278 1176 3472 1178
rect 3518 1176 3712 1178
rect 3758 1176 4100 1178
rect 1126 1132 1312 1176
rect 1366 1132 1552 1176
rect 1606 1132 1792 1176
rect 1846 1132 2032 1176
rect 2086 1132 2272 1176
rect 2326 1132 2512 1176
rect 2566 1132 2752 1176
rect 2806 1132 2992 1176
rect 3046 1132 3232 1176
rect 3286 1132 3472 1176
rect 3526 1132 3712 1176
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1314 1132
rect 1366 1124 1554 1132
rect 1606 1124 1794 1132
rect 1846 1124 2034 1132
rect 2086 1124 2274 1132
rect 2326 1124 2514 1132
rect 2566 1124 2754 1132
rect 2806 1124 2994 1132
rect 3046 1124 3234 1132
rect 3286 1124 3474 1132
rect 3526 1124 3714 1132
rect 3766 1124 4100 1176
rect 0 1110 4100 1124
rect 110 987 160 1110
rect 110 753 112 987
rect 158 753 160 987
rect 110 700 160 753
rect 280 987 330 1040
rect 280 753 282 987
rect 328 753 330 987
rect 160 626 220 650
rect 160 574 164 626
rect 216 574 220 626
rect 160 550 220 574
rect 280 510 330 753
rect 430 1020 480 1040
rect 430 880 432 1020
rect 478 880 480 1020
rect 280 500 340 510
rect 280 496 360 500
rect 280 444 284 496
rect 336 444 360 496
rect 280 440 360 444
rect 280 380 340 440
rect 430 380 480 880
rect 600 1015 650 1040
rect 600 875 602 1015
rect 648 875 650 1015
rect 600 800 650 875
rect 770 1015 820 1110
rect 770 875 772 1015
rect 818 875 820 1015
rect 770 850 820 875
rect 940 1015 990 1040
rect 940 875 942 1015
rect 988 875 990 1015
rect 1140 1018 1190 1110
rect 1140 972 1142 1018
rect 1188 972 1190 1018
rect 1140 950 1190 972
rect 1520 1010 1630 1040
rect 1520 900 1552 1010
rect 940 800 990 875
rect 600 750 990 800
rect 1080 870 1552 900
rect 1598 870 1630 1010
rect 1080 840 1630 870
rect 1860 1000 1910 1110
rect 1860 860 1862 1000
rect 1908 860 1910 1000
rect 1080 660 1140 840
rect 1860 820 1910 860
rect 2140 1007 2250 1040
rect 2140 786 2172 1007
rect 2140 734 2144 786
rect 2218 773 2250 1007
rect 2580 1018 2630 1110
rect 2580 972 2582 1018
rect 2628 972 2630 1018
rect 2580 950 2630 972
rect 2750 997 2800 1040
rect 2470 896 2570 900
rect 2470 844 2494 896
rect 2546 844 2570 896
rect 2470 840 2570 844
rect 2490 820 2550 840
rect 2196 740 2250 773
rect 2750 763 2752 997
rect 2798 770 2800 997
rect 2930 1015 2980 1040
rect 2930 875 2932 1015
rect 2978 875 2980 1015
rect 2930 800 2980 875
rect 3100 1015 3150 1110
rect 3100 875 3102 1015
rect 3148 875 3150 1015
rect 3100 850 3150 875
rect 3270 1015 3320 1040
rect 3270 875 3272 1015
rect 3318 875 3320 1015
rect 3270 800 3320 875
rect 2798 763 2860 770
rect 2196 734 2200 740
rect 2140 710 2200 734
rect 2750 720 2860 763
rect 2930 750 3320 800
rect 3440 1020 3490 1040
rect 3440 880 3442 1020
rect 3488 880 3490 1020
rect 3440 820 3490 880
rect 3590 992 3640 1040
rect 3440 770 3500 820
rect 680 656 780 660
rect 680 604 704 656
rect 756 604 780 656
rect 680 600 780 604
rect 880 656 1140 660
rect 880 604 904 656
rect 956 604 1140 656
rect 1360 653 2740 660
rect 880 600 1140 604
rect 1080 500 1140 600
rect 1210 626 1310 630
rect 1210 574 1234 626
rect 1286 574 1310 626
rect 1360 607 1387 653
rect 1433 607 2327 653
rect 2373 630 2740 653
rect 2373 626 2760 630
rect 2373 607 2684 626
rect 1360 600 2684 607
rect 1210 570 1310 574
rect 530 496 630 500
rect 530 444 554 496
rect 606 444 630 496
rect 530 440 630 444
rect 1080 440 1310 500
rect 1640 490 1700 600
rect 2070 490 2130 600
rect 2660 574 2684 600
rect 2736 574 2760 626
rect 2660 570 2760 574
rect 2470 546 2570 550
rect 2280 506 2340 540
rect 770 436 1030 440
rect 770 384 954 436
rect 1006 384 1030 436
rect 770 380 1030 384
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 380
rect 430 330 820 380
rect 280 252 282 298
rect 328 252 330 298
rect 630 320 820 330
rect 1250 330 1310 440
rect 1400 486 1500 490
rect 1400 434 1424 486
rect 1476 434 1500 486
rect 1400 430 1500 434
rect 1620 478 1720 490
rect 1620 432 1647 478
rect 1693 432 1720 478
rect 2050 488 2150 490
rect 1800 460 1860 470
rect 1620 430 1720 432
rect 1780 456 1880 460
rect 1780 404 1804 456
rect 1856 404 1880 456
rect 2050 442 2077 488
rect 2123 442 2150 488
rect 2050 440 2150 442
rect 2280 454 2284 506
rect 2336 454 2340 506
rect 2470 494 2494 546
rect 2546 494 2570 546
rect 2810 500 2860 720
rect 2910 626 3130 630
rect 2910 574 2934 626
rect 2986 574 3130 626
rect 2910 570 3130 574
rect 3180 626 3280 630
rect 3180 574 3204 626
rect 3256 574 3280 626
rect 3180 570 3280 574
rect 3450 570 3500 770
rect 3590 758 3592 992
rect 3638 760 3640 992
rect 3760 995 3810 1110
rect 3760 855 3762 995
rect 3808 855 3810 995
rect 3930 987 3980 1040
rect 3930 910 3932 987
rect 3760 810 3810 855
rect 3920 886 3932 910
rect 3920 834 3924 886
rect 3920 810 3932 834
rect 3638 758 3880 760
rect 3590 756 3880 758
rect 3590 704 3804 756
rect 3856 704 3880 756
rect 3590 700 3880 704
rect 3930 753 3932 810
rect 3978 753 3980 987
rect 3800 690 3860 700
rect 3810 648 3860 690
rect 3810 602 3812 648
rect 3858 602 3860 648
rect 2470 490 2570 494
rect 2280 440 2340 454
rect 2750 440 2860 500
rect 2920 466 3020 470
rect 1780 400 1880 404
rect 2280 390 2800 440
rect 2920 414 2944 466
rect 2996 414 3020 466
rect 2920 410 3020 414
rect 2140 366 2200 390
rect 630 283 680 320
rect 280 190 330 252
rect 460 258 510 280
rect 460 212 462 258
rect 508 212 510 258
rect 460 120 510 212
rect 630 237 632 283
rect 678 237 680 283
rect 630 190 680 237
rect 910 263 960 290
rect 910 217 912 263
rect 958 217 960 263
rect 910 120 960 217
rect 1140 263 1190 300
rect 1250 280 1630 330
rect 2140 314 2144 366
rect 2196 330 2200 366
rect 2196 314 2250 330
rect 1140 217 1142 263
rect 1188 217 1190 263
rect 1140 120 1190 217
rect 1520 263 1630 280
rect 1520 217 1552 263
rect 1598 217 1630 263
rect 1520 190 1630 217
rect 1860 258 1910 280
rect 1860 212 1862 258
rect 1908 212 1910 258
rect 1860 120 1910 212
rect 2140 258 2250 314
rect 2140 212 2172 258
rect 2218 212 2250 258
rect 2140 190 2250 212
rect 2580 283 2630 340
rect 2580 237 2582 283
rect 2628 237 2630 283
rect 2580 120 2630 237
rect 2750 298 2800 390
rect 3070 380 3130 570
rect 3450 566 3720 570
rect 3450 514 3644 566
rect 3696 514 3720 566
rect 3450 510 3720 514
rect 3300 486 3400 490
rect 3300 434 3324 486
rect 3376 434 3400 486
rect 3300 432 3327 434
rect 3373 432 3400 434
rect 3300 430 3400 432
rect 3450 380 3500 510
rect 3810 420 3860 602
rect 2750 252 2752 298
rect 2798 252 2800 298
rect 2750 190 2800 252
rect 2960 298 3010 360
rect 3070 330 3500 380
rect 3590 370 3860 420
rect 2960 252 2962 298
rect 3008 252 3010 298
rect 2960 120 3010 252
rect 3240 273 3290 330
rect 3590 298 3640 370
rect 3240 227 3242 273
rect 3288 227 3290 273
rect 3240 190 3290 227
rect 3410 258 3460 280
rect 3410 212 3412 258
rect 3458 212 3460 258
rect 3410 120 3460 212
rect 3590 252 3592 298
rect 3638 252 3640 298
rect 3590 190 3640 252
rect 3760 278 3810 320
rect 3760 232 3762 278
rect 3808 232 3810 278
rect 3760 120 3810 232
rect 3930 298 3980 753
rect 3930 252 3932 298
rect 3978 252 3980 298
rect 3930 190 3980 252
rect 0 106 4100 120
rect 0 98 114 106
rect 0 52 112 98
rect 166 54 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 2566 98 2754 106
rect 2806 98 2994 106
rect 3046 98 3234 106
rect 3286 98 3474 106
rect 3526 98 3714 106
rect 408 54 594 98
rect 648 54 834 98
rect 158 52 362 54
rect 408 52 602 54
rect 648 52 842 54
rect 888 52 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2752 98
rect 2806 54 2992 98
rect 3046 54 3232 98
rect 3286 54 3472 98
rect 3526 54 3712 98
rect 3766 54 4100 106
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2752 54
rect 2798 52 2992 54
rect 3038 52 3232 54
rect 3278 52 3472 54
rect 3518 52 3712 54
rect 3758 52 4100 54
rect 0 0 4100 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 114 1124 166 1132
rect 354 1132 362 1176
rect 362 1132 406 1176
rect 594 1132 602 1176
rect 602 1132 646 1176
rect 834 1132 842 1176
rect 842 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 1314 1132 1358 1176
rect 1358 1132 1366 1176
rect 1554 1132 1598 1176
rect 1598 1132 1606 1176
rect 1794 1132 1838 1176
rect 1838 1132 1846 1176
rect 2034 1132 2078 1176
rect 2078 1132 2086 1176
rect 2274 1132 2318 1176
rect 2318 1132 2326 1176
rect 2514 1132 2558 1176
rect 2558 1132 2566 1176
rect 2754 1132 2798 1176
rect 2798 1132 2806 1176
rect 2994 1132 3038 1176
rect 3038 1132 3046 1176
rect 3234 1132 3278 1176
rect 3278 1132 3286 1176
rect 3474 1132 3518 1176
rect 3518 1132 3526 1176
rect 3714 1132 3758 1176
rect 3758 1132 3766 1176
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 1554 1124 1606 1132
rect 1794 1124 1846 1132
rect 2034 1124 2086 1132
rect 2274 1124 2326 1132
rect 2514 1124 2566 1132
rect 2754 1124 2806 1132
rect 2994 1124 3046 1132
rect 3234 1124 3286 1132
rect 3474 1124 3526 1132
rect 3714 1124 3766 1132
rect 164 623 216 626
rect 164 577 167 623
rect 167 577 213 623
rect 213 577 216 623
rect 164 574 216 577
rect 284 444 336 496
rect 2144 773 2172 786
rect 2172 773 2196 786
rect 2494 844 2546 896
rect 2144 734 2196 773
rect 704 653 756 656
rect 704 607 707 653
rect 707 607 753 653
rect 753 607 756 653
rect 704 604 756 607
rect 904 653 956 656
rect 904 607 907 653
rect 907 607 953 653
rect 953 607 956 653
rect 904 604 956 607
rect 1234 623 1286 626
rect 1234 577 1237 623
rect 1237 577 1283 623
rect 1283 577 1286 623
rect 1234 574 1286 577
rect 2684 623 2736 626
rect 554 493 606 496
rect 554 447 557 493
rect 557 447 603 493
rect 603 447 606 493
rect 554 444 606 447
rect 2684 577 2687 623
rect 2687 577 2733 623
rect 2733 577 2736 623
rect 2684 574 2736 577
rect 954 384 1006 436
rect 1424 483 1476 486
rect 1424 437 1427 483
rect 1427 437 1473 483
rect 1473 437 1476 483
rect 1424 434 1476 437
rect 1804 453 1856 456
rect 1804 407 1807 453
rect 1807 407 1853 453
rect 1853 407 1856 453
rect 1804 404 1856 407
rect 2284 503 2336 506
rect 2284 457 2287 503
rect 2287 457 2333 503
rect 2333 457 2336 503
rect 2284 454 2336 457
rect 2494 543 2546 546
rect 2494 497 2497 543
rect 2497 497 2543 543
rect 2543 497 2546 543
rect 2494 494 2546 497
rect 2934 574 2986 626
rect 3204 623 3256 626
rect 3204 577 3207 623
rect 3207 577 3253 623
rect 3253 577 3256 623
rect 3204 574 3256 577
rect 3924 834 3932 886
rect 3932 834 3976 886
rect 3804 704 3856 756
rect 2944 463 2996 466
rect 2944 417 2947 463
rect 2947 417 2993 463
rect 2993 417 2996 463
rect 2944 414 2996 417
rect 2144 314 2196 366
rect 3644 563 3696 566
rect 3644 517 3647 563
rect 3647 517 3693 563
rect 3693 517 3696 563
rect 3644 514 3696 517
rect 3324 478 3376 486
rect 3324 434 3327 478
rect 3327 434 3373 478
rect 3373 434 3376 478
rect 114 98 166 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 2754 98 2806 106
rect 2994 98 3046 106
rect 3234 98 3286 106
rect 3474 98 3526 106
rect 3714 98 3766 106
rect 354 54 362 98
rect 362 54 406 98
rect 594 54 602 98
rect 602 54 646 98
rect 834 54 842 98
rect 842 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
rect 2754 54 2798 98
rect 2798 54 2806 98
rect 2994 54 3038 98
rect 3038 54 3046 98
rect 3234 54 3278 98
rect 3278 54 3286 98
rect 3474 54 3518 98
rect 3518 54 3526 98
rect 3714 54 3758 98
rect 3758 54 3766 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 1540 1180 1620 1190
rect 1780 1180 1860 1190
rect 2020 1180 2100 1190
rect 2260 1180 2340 1190
rect 2500 1180 2580 1190
rect 2740 1180 2820 1190
rect 2980 1180 3060 1190
rect 3220 1180 3300 1190
rect 3460 1180 3540 1190
rect 3700 1180 3780 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 1530 1176 1630 1180
rect 1530 1124 1554 1176
rect 1606 1124 1630 1176
rect 1530 1120 1630 1124
rect 1770 1176 1870 1180
rect 1770 1124 1794 1176
rect 1846 1124 1870 1176
rect 1770 1120 1870 1124
rect 2010 1176 2110 1180
rect 2010 1124 2034 1176
rect 2086 1124 2110 1176
rect 2010 1120 2110 1124
rect 2250 1176 2350 1180
rect 2250 1124 2274 1176
rect 2326 1124 2350 1176
rect 2250 1120 2350 1124
rect 2490 1176 2590 1180
rect 2490 1124 2514 1176
rect 2566 1124 2590 1176
rect 2490 1120 2590 1124
rect 2730 1176 2830 1180
rect 2730 1124 2754 1176
rect 2806 1124 2830 1176
rect 2730 1120 2830 1124
rect 2970 1176 3070 1180
rect 2970 1124 2994 1176
rect 3046 1124 3070 1176
rect 2970 1120 3070 1124
rect 3210 1176 3310 1180
rect 3210 1124 3234 1176
rect 3286 1124 3310 1176
rect 3210 1120 3310 1124
rect 3450 1176 3550 1180
rect 3450 1124 3474 1176
rect 3526 1124 3550 1176
rect 3450 1120 3550 1124
rect 3690 1176 3790 1180
rect 3690 1124 3714 1176
rect 3766 1124 3790 1176
rect 3690 1120 3790 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 1540 1110 1620 1120
rect 1780 1110 1860 1120
rect 2020 1110 2100 1120
rect 2260 1110 2340 1120
rect 2500 1110 2580 1120
rect 2740 1110 2820 1120
rect 2980 1110 3060 1120
rect 3220 1110 3300 1120
rect 3460 1110 3540 1120
rect 3700 1110 3780 1120
rect 700 990 3260 1050
rect 700 670 760 990
rect 1420 870 2340 930
rect 2480 900 2560 910
rect 680 656 780 670
rect 150 630 230 640
rect 140 626 240 630
rect 140 574 164 626
rect 216 574 240 626
rect 680 604 704 656
rect 756 604 780 656
rect 680 590 780 604
rect 880 656 980 670
rect 880 604 904 656
rect 956 604 980 656
rect 1210 630 1310 640
rect 880 590 980 604
rect 1200 626 1320 630
rect 140 570 240 574
rect 1200 574 1234 626
rect 1286 574 1320 626
rect 1200 570 1320 574
rect 150 560 230 570
rect 1210 560 1310 570
rect 270 500 350 510
rect 530 500 630 510
rect 1420 500 1480 870
rect 2140 800 2200 810
rect 2130 786 2210 800
rect 2130 734 2144 786
rect 2196 734 2210 786
rect 2130 720 2210 734
rect 260 496 630 500
rect 260 444 284 496
rect 336 444 554 496
rect 606 444 630 496
rect 1410 490 1500 500
rect 1400 486 1500 490
rect 260 440 630 444
rect 270 430 350 440
rect 530 430 630 440
rect 930 440 1030 450
rect 930 436 1320 440
rect 550 240 610 430
rect 930 384 954 436
rect 1006 384 1320 436
rect 1400 434 1424 486
rect 1476 434 1500 486
rect 1800 470 1860 480
rect 1400 430 1500 434
rect 1410 420 1500 430
rect 1790 460 1870 470
rect 1790 456 1880 460
rect 930 380 1320 384
rect 930 370 1030 380
rect 1260 360 1320 380
rect 1790 404 1804 456
rect 1856 404 1880 456
rect 1790 400 1880 404
rect 1790 390 1870 400
rect 1790 360 1860 390
rect 2140 380 2200 720
rect 2280 520 2340 870
rect 2470 896 2900 900
rect 2470 844 2494 896
rect 2546 844 2900 896
rect 2470 840 2900 844
rect 2480 830 2560 840
rect 2490 560 2550 830
rect 2840 640 2900 840
rect 3200 640 3260 990
rect 3910 890 3990 900
rect 3900 886 4000 890
rect 3900 834 3924 886
rect 3976 834 4000 886
rect 3900 830 4000 834
rect 3910 820 3990 830
rect 3790 760 3870 770
rect 3780 756 3880 760
rect 3780 704 3804 756
rect 3856 704 3880 756
rect 3780 700 3880 704
rect 3790 690 3870 700
rect 2670 630 2750 640
rect 2660 626 2760 630
rect 2660 574 2684 626
rect 2736 574 2760 626
rect 2660 570 2760 574
rect 2840 626 3010 640
rect 2840 574 2934 626
rect 2986 574 3010 626
rect 2840 570 3010 574
rect 2670 560 2750 570
rect 2910 560 3010 570
rect 3180 626 3280 640
rect 3180 574 3204 626
rect 3256 574 3280 626
rect 3180 560 3280 574
rect 3630 570 3710 580
rect 3600 566 3720 570
rect 2480 550 2560 560
rect 2470 546 2570 550
rect 2270 506 2350 520
rect 2270 454 2284 506
rect 2336 454 2350 506
rect 2470 494 2494 546
rect 2546 494 2570 546
rect 3600 514 3644 566
rect 3696 514 3720 566
rect 3600 510 3720 514
rect 3320 500 3380 510
rect 3630 500 3710 510
rect 2470 490 2570 494
rect 2480 480 2560 490
rect 3310 486 3390 500
rect 2270 440 2350 454
rect 2920 466 3020 480
rect 2280 430 2340 440
rect 2920 414 2944 466
rect 2996 414 3020 466
rect 2920 400 3020 414
rect 3310 434 3324 486
rect 3376 434 3390 486
rect 3310 410 3390 434
rect 2130 370 2210 380
rect 2920 370 3000 400
rect 1260 300 1860 360
rect 2120 366 3000 370
rect 2120 314 2144 366
rect 2196 314 3000 366
rect 2120 310 3000 314
rect 2130 300 2210 310
rect 3310 240 3370 410
rect 550 180 3370 240
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 2740 110 2820 120
rect 2980 110 3060 120
rect 3220 110 3300 120
rect 3460 110 3540 120
rect 3700 110 3780 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 50 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 50 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 50 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 50 2590 54
rect 2730 106 2830 110
rect 2730 54 2754 106
rect 2806 54 2830 106
rect 2730 50 2830 54
rect 2970 106 3070 110
rect 2970 54 2994 106
rect 3046 54 3070 106
rect 2970 50 3070 54
rect 3210 106 3310 110
rect 3210 54 3234 106
rect 3286 54 3310 106
rect 3210 50 3310 54
rect 3450 106 3550 110
rect 3450 54 3474 106
rect 3526 54 3550 106
rect 3450 50 3550 54
rect 3690 106 3790 110
rect 3690 54 3714 106
rect 3766 54 3790 106
rect 3690 50 3790 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
rect 1780 40 1860 50
rect 2020 40 2100 50
rect 2260 40 2340 50
rect 2500 40 2580 50
rect 2740 40 2820 50
rect 2980 40 3060 50
rect 3220 40 3300 50
rect 3460 40 3540 50
rect 3700 40 3780 50
<< labels >>
rlabel metal2 s 100 40 180 120 4 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 100 1110 180 1190 4 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1210 560 1310 640 4 D
port 1 nsew signal input
rlabel metal2 s 3910 820 3990 900 4 Q
port 2 nsew signal output
rlabel metal2 s 3790 690 3870 770 4 QN
port 3 nsew signal output
rlabel metal2 s 2670 560 2750 640 4 CLK
port 4 nsew clock input
rlabel metal2 s 150 560 230 640 4 RN
port 5 nsew signal input
rlabel metal2 s 700 590 760 1050 4 SN
port 6 nsew signal output
rlabel metal2 s 2660 570 2760 630 1 CLK
port 4 nsew clock input
rlabel metal1 s 1640 430 1700 660 1 CLK
port 4 nsew clock input
rlabel metal1 s 1620 430 1720 490 1 CLK
port 4 nsew clock input
rlabel metal1 s 2070 440 2130 660 1 CLK
port 4 nsew clock input
rlabel metal1 s 2050 440 2150 490 1 CLK
port 4 nsew clock input
rlabel metal1 s 1360 600 2740 660 1 CLK
port 4 nsew clock input
rlabel metal1 s 2660 570 2760 630 1 CLK
port 4 nsew clock input
rlabel metal2 s 1200 570 1320 630 1 D
port 1 nsew signal input
rlabel metal1 s 1210 570 1310 630 1 D
port 1 nsew signal input
rlabel metal2 s 3900 830 4000 890 1 Q
port 2 nsew signal output
rlabel metal1 s 3920 810 3980 910 1 Q
port 2 nsew signal output
rlabel metal1 s 3930 190 3980 1040 1 Q
port 2 nsew signal output
rlabel metal2 s 3780 700 3880 760 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 190 3640 420 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 700 3640 1040 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 370 3860 420 1 QN
port 3 nsew signal output
rlabel metal1 s 3810 370 3860 760 1 QN
port 3 nsew signal output
rlabel metal1 s 3800 690 3860 760 1 QN
port 3 nsew signal output
rlabel metal1 s 3590 700 3880 760 1 QN
port 3 nsew signal output
rlabel metal2 s 140 570 240 630 1 RN
port 5 nsew signal input
rlabel metal1 s 160 550 220 650 1 RN
port 5 nsew signal input
rlabel metal2 s 680 590 780 670 1 SN
port 6 nsew signal output
rlabel metal2 s 3200 560 3260 1050 1 SN
port 6 nsew signal output
rlabel metal2 s 700 990 3260 1050 1 SN
port 6 nsew signal output
rlabel metal2 s 3180 560 3280 640 1 SN
port 6 nsew signal output
rlabel metal1 s 680 600 780 660 1 SN
port 6 nsew signal output
rlabel metal1 s 3180 570 3280 630 1 SN
port 6 nsew signal output
rlabel metal2 s 90 1120 190 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1540 1110 1620 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1530 1120 1630 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1780 1110 1860 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1770 1120 1870 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2020 1110 2100 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2010 1120 2110 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2260 1110 2340 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2250 1120 2350 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2500 1110 2580 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2490 1120 2590 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2740 1110 2820 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2730 1120 2830 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2980 1110 3060 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2970 1120 3070 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3220 1110 3300 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3210 1120 3310 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3460 1110 3540 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3450 1120 3550 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3700 1110 3780 1190 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 3690 1120 3790 1180 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 110 700 160 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 770 850 820 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 1140 950 1190 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 1860 820 1910 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 2580 950 2630 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 3100 850 3150 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 3760 810 3810 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 0 1110 4100 1230 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1780 40 1860 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1770 50 1870 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2020 40 2100 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2010 50 2110 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2260 40 2340 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2250 50 2350 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2500 40 2580 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2490 50 2590 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2740 40 2820 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2730 50 2830 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2980 40 3060 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2970 50 3070 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3220 40 3300 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3210 50 3310 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3460 40 3540 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3450 50 3550 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3700 40 3780 120 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 3690 50 3790 110 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 110 0 160 360 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 460 0 510 280 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 910 0 960 290 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 1140 0 1190 300 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 1860 0 1910 280 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 2580 0 2630 340 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 2960 0 3010 360 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 3410 0 3460 280 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 3760 0 3810 320 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 0 0 4100 120 1 VSS
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4100 1230
string GDS_END 316728
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 277374
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
