magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4006 1094
<< pwell >>
rect -86 -86 4006 453
<< mvnmos >>
rect 124 150 244 308
rect 348 150 468 308
rect 716 192 836 332
rect 940 192 1060 332
rect 1164 192 1284 332
rect 1332 192 1452 332
rect 1536 192 1656 332
rect 1864 192 1984 332
rect 2088 192 2208 332
rect 2312 192 2432 332
rect 2536 192 2656 332
rect 2760 192 2880 332
rect 3020 69 3140 333
rect 3388 69 3508 333
rect 3612 69 3732 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 720 573 820 773
rect 924 573 1024 773
rect 1128 573 1228 773
rect 1332 573 1432 773
rect 1536 573 1636 773
rect 1884 652 1984 852
rect 2088 652 2188 852
rect 2313 652 2413 852
rect 2532 652 2632 852
rect 2780 573 2880 939
rect 3040 573 3140 939
rect 3408 573 3508 939
rect 3612 573 3712 939
<< mvndiff >>
rect 2940 332 3020 333
rect 36 295 124 308
rect 36 249 49 295
rect 95 249 124 295
rect 36 150 124 249
rect 244 209 348 308
rect 244 163 273 209
rect 319 163 348 209
rect 244 150 348 163
rect 468 295 556 308
rect 468 249 497 295
rect 543 249 556 295
rect 468 150 556 249
rect 628 251 716 332
rect 628 205 641 251
rect 687 205 716 251
rect 628 192 716 205
rect 836 319 940 332
rect 836 273 865 319
rect 911 273 940 319
rect 836 192 940 273
rect 1060 319 1164 332
rect 1060 273 1089 319
rect 1135 273 1164 319
rect 1060 192 1164 273
rect 1284 192 1332 332
rect 1452 192 1536 332
rect 1656 251 1864 332
rect 1656 205 1685 251
rect 1731 205 1864 251
rect 1656 192 1864 205
rect 1984 319 2088 332
rect 1984 273 2013 319
rect 2059 273 2088 319
rect 1984 192 2088 273
rect 2208 319 2312 332
rect 2208 273 2237 319
rect 2283 273 2312 319
rect 2208 192 2312 273
rect 2432 319 2536 332
rect 2432 273 2461 319
rect 2507 273 2536 319
rect 2432 192 2536 273
rect 2656 251 2760 332
rect 2656 205 2685 251
rect 2731 205 2760 251
rect 2656 192 2760 205
rect 2880 192 3020 332
rect 2940 69 3020 192
rect 3140 320 3228 333
rect 3140 180 3169 320
rect 3215 180 3228 320
rect 3140 69 3228 180
rect 3300 222 3388 333
rect 3300 82 3313 222
rect 3359 82 3388 222
rect 3300 69 3388 82
rect 3508 320 3612 333
rect 3508 180 3537 320
rect 3583 180 3612 320
rect 3508 69 3612 180
rect 3732 222 3820 333
rect 3732 82 3761 222
rect 3807 82 3820 222
rect 3732 69 3820 82
<< mvpdiff >>
rect 56 726 144 849
rect 56 586 69 726
rect 115 586 144 726
rect 56 573 144 586
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 2692 926 2780 939
rect 2692 880 2705 926
rect 2751 880 2780 926
rect 2692 852 2780 880
rect 1796 839 1884 852
rect 448 586 477 726
rect 523 586 536 726
rect 448 573 536 586
rect 632 760 720 773
rect 632 620 645 760
rect 691 620 720 760
rect 632 573 720 620
rect 820 726 924 773
rect 820 586 849 726
rect 895 586 924 726
rect 820 573 924 586
rect 1024 726 1128 773
rect 1024 586 1053 726
rect 1099 586 1128 726
rect 1024 573 1128 586
rect 1228 735 1332 773
rect 1228 595 1257 735
rect 1303 595 1332 735
rect 1228 573 1332 595
rect 1432 760 1536 773
rect 1432 714 1461 760
rect 1507 714 1536 760
rect 1432 573 1536 714
rect 1636 735 1724 773
rect 1636 595 1665 735
rect 1711 595 1724 735
rect 1796 699 1809 839
rect 1855 699 1884 839
rect 1796 652 1884 699
rect 1984 805 2088 852
rect 1984 665 2013 805
rect 2059 665 2088 805
rect 1984 652 2088 665
rect 2188 805 2313 852
rect 2188 665 2238 805
rect 2284 665 2313 805
rect 2188 652 2313 665
rect 2413 711 2532 852
rect 2413 665 2457 711
rect 2503 665 2532 711
rect 2413 652 2532 665
rect 2632 652 2780 852
rect 1636 573 1724 595
rect 2700 573 2780 652
rect 2880 632 3040 939
rect 2880 586 2909 632
rect 2955 586 3040 632
rect 2880 573 3040 586
rect 3140 926 3228 939
rect 3140 786 3169 926
rect 3215 786 3228 926
rect 3140 573 3228 786
rect 3320 926 3408 939
rect 3320 786 3333 926
rect 3379 786 3408 926
rect 3320 573 3408 786
rect 3508 726 3612 939
rect 3508 586 3537 726
rect 3583 586 3612 726
rect 3508 573 3612 586
rect 3712 926 3800 939
rect 3712 786 3741 926
rect 3787 786 3800 926
rect 3712 573 3800 786
<< mvndiffc >>
rect 49 249 95 295
rect 273 163 319 209
rect 497 249 543 295
rect 641 205 687 251
rect 865 273 911 319
rect 1089 273 1135 319
rect 1685 205 1731 251
rect 2013 273 2059 319
rect 2237 273 2283 319
rect 2461 273 2507 319
rect 2685 205 2731 251
rect 3169 180 3215 320
rect 3313 82 3359 222
rect 3537 180 3583 320
rect 3761 82 3807 222
<< mvpdiffc >>
rect 69 586 115 726
rect 273 696 319 836
rect 2705 880 2751 926
rect 477 586 523 726
rect 645 620 691 760
rect 849 586 895 726
rect 1053 586 1099 726
rect 1257 595 1303 735
rect 1461 714 1507 760
rect 1665 595 1711 735
rect 1809 699 1855 839
rect 2013 665 2059 805
rect 2238 665 2284 805
rect 2457 665 2503 711
rect 2909 586 2955 632
rect 3169 786 3215 926
rect 3333 786 3379 926
rect 3537 586 3583 726
rect 3741 786 3787 926
<< polysilicon >>
rect 348 909 1024 949
rect 144 849 244 893
rect 348 849 448 909
rect 720 773 820 817
rect 924 773 1024 909
rect 1129 944 2188 984
rect 1129 865 1228 944
rect 1128 852 1228 865
rect 1884 852 1984 896
rect 2088 852 2188 944
rect 2780 939 2880 983
rect 3040 939 3140 983
rect 3408 939 3508 983
rect 3612 939 3712 983
rect 2313 852 2413 896
rect 2532 852 2632 896
rect 1128 806 1141 852
rect 1187 806 1228 852
rect 1128 773 1228 806
rect 1332 773 1432 817
rect 1536 773 1636 817
rect 144 411 244 573
rect 144 365 157 411
rect 203 365 244 411
rect 144 352 244 365
rect 124 308 244 352
rect 348 387 448 573
rect 348 341 361 387
rect 407 352 448 387
rect 720 411 820 573
rect 924 529 1024 573
rect 1128 481 1228 573
rect 720 376 733 411
rect 716 365 733 376
rect 779 376 820 411
rect 940 472 1228 481
rect 940 441 1167 472
rect 1332 446 1432 573
rect 779 365 836 376
rect 407 341 468 352
rect 348 308 468 341
rect 716 332 836 365
rect 940 332 1060 441
rect 1212 411 1284 424
rect 1212 376 1225 411
rect 1164 365 1225 376
rect 1271 365 1284 411
rect 1164 332 1284 365
rect 1332 400 1373 446
rect 1419 400 1432 446
rect 1332 376 1432 400
rect 1536 376 1636 573
rect 1884 538 1984 652
rect 1884 492 1897 538
rect 1943 492 1984 538
rect 1884 376 1984 492
rect 2088 512 2188 652
rect 2313 619 2413 652
rect 2313 573 2329 619
rect 2375 573 2413 619
rect 2313 560 2413 573
rect 2532 522 2632 652
rect 2088 472 2432 512
rect 1332 332 1452 376
rect 1536 332 1656 376
rect 1864 332 1984 376
rect 2088 411 2208 424
rect 2088 365 2105 411
rect 2151 365 2208 411
rect 2088 332 2208 365
rect 2312 332 2432 472
rect 2532 476 2573 522
rect 2619 476 2632 522
rect 2532 392 2632 476
rect 2780 411 2880 573
rect 2536 332 2656 392
rect 2780 376 2821 411
rect 2760 365 2821 376
rect 2867 365 2880 411
rect 3040 540 3140 573
rect 3040 494 3053 540
rect 3099 494 3140 540
rect 3040 377 3140 494
rect 3408 465 3508 573
rect 3612 465 3712 573
rect 3408 412 3712 465
rect 3408 377 3421 412
rect 2760 332 2880 365
rect 3020 333 3140 377
rect 3388 366 3421 377
rect 3467 393 3712 412
rect 3467 366 3508 393
rect 3388 333 3508 366
rect 3612 377 3712 393
rect 3612 333 3732 377
rect 124 106 244 150
rect 348 106 468 150
rect 716 148 836 192
rect 940 148 1060 192
rect 1164 148 1284 192
rect 1332 148 1452 192
rect 428 90 468 106
rect 1164 90 1204 148
rect 428 50 1204 90
rect 1536 100 1656 192
rect 1864 148 1984 192
rect 2088 148 2208 192
rect 2312 148 2432 192
rect 2536 148 2656 192
rect 2760 100 2880 192
rect 1536 60 2880 100
rect 3020 25 3140 69
rect 3388 25 3508 69
rect 3612 25 3732 69
<< polycontact >>
rect 1141 806 1187 852
rect 157 365 203 411
rect 361 341 407 387
rect 733 365 779 411
rect 1225 365 1271 411
rect 1373 400 1419 446
rect 1897 492 1943 538
rect 2329 573 2375 619
rect 2105 365 2151 411
rect 2573 476 2619 522
rect 2821 365 2867 411
rect 3053 494 3099 540
rect 3421 366 3467 412
<< metal1 >>
rect 0 926 3920 1098
rect 0 918 2705 926
rect 273 836 319 918
rect 69 726 115 737
rect 645 760 691 918
rect 273 685 319 696
rect 477 726 523 737
rect 115 586 407 621
rect 69 575 407 586
rect 142 411 315 449
rect 142 365 157 411
rect 203 365 315 411
rect 142 354 315 365
rect 361 387 407 575
rect 361 308 407 341
rect 49 295 407 308
rect 95 262 407 295
rect 645 609 691 620
rect 737 806 1141 852
rect 1187 806 1198 852
rect 477 563 523 586
rect 737 563 783 806
rect 1461 760 1507 918
rect 477 517 783 563
rect 849 726 911 737
rect 895 586 911 726
rect 477 295 543 517
rect 589 411 779 430
rect 589 365 733 411
rect 589 354 779 365
rect 49 238 95 249
rect 477 249 497 295
rect 849 319 911 586
rect 849 273 865 319
rect 849 262 911 273
rect 1053 726 1099 737
rect 1053 538 1099 586
rect 1257 735 1303 746
rect 1809 839 1855 918
rect 2751 918 3169 926
rect 2705 869 2751 880
rect 1461 703 1507 714
rect 1665 735 1711 746
rect 1303 595 1665 630
rect 1809 688 1855 699
rect 2013 805 2059 816
rect 1257 584 1711 595
rect 1053 492 1897 538
rect 1943 492 1954 538
rect 1053 319 1135 492
rect 2013 446 2059 665
rect 1214 365 1225 411
rect 1271 365 1316 411
rect 1362 400 1373 446
rect 1419 400 2059 446
rect 2237 805 3099 816
rect 2237 665 2238 805
rect 2284 770 3099 805
rect 3215 918 3333 926
rect 3169 775 3215 786
rect 3379 918 3741 926
rect 3333 775 3379 786
rect 3787 918 3920 926
rect 3741 775 3787 786
rect 2237 654 2284 665
rect 2457 711 2507 722
rect 2503 665 2507 711
rect 1053 273 1089 319
rect 1270 354 1316 365
rect 1270 308 1967 354
rect 1053 262 1135 273
rect 477 238 543 249
rect 641 251 687 262
rect 262 209 330 216
rect 262 163 273 209
rect 319 163 330 209
rect 262 90 330 163
rect 641 90 687 205
rect 1685 251 1731 262
rect 1685 90 1731 205
rect 1921 216 1967 308
rect 2013 319 2059 400
rect 2013 262 2059 273
rect 2105 411 2151 422
rect 2105 216 2151 365
rect 2237 319 2283 654
rect 2237 262 2283 273
rect 2329 619 2375 630
rect 2329 216 2375 573
rect 2457 319 2507 665
rect 2909 632 2955 643
rect 2909 522 2955 586
rect 3053 540 3099 770
rect 3502 726 3583 766
rect 3502 690 3537 726
rect 2562 476 2573 522
rect 2619 476 3007 522
rect 3053 483 3099 494
rect 2961 437 3007 476
rect 2676 411 2882 430
rect 2676 365 2821 411
rect 2867 365 2882 411
rect 2961 412 3478 437
rect 2961 391 3421 412
rect 2676 335 2882 365
rect 3169 366 3421 391
rect 3467 366 3478 412
rect 2457 273 2461 319
rect 2457 262 2507 273
rect 3169 320 3215 366
rect 1921 170 2375 216
rect 2685 251 2731 262
rect 2685 90 2731 205
rect 3537 320 3583 586
rect 3169 169 3215 180
rect 3313 222 3359 233
rect 0 82 3313 90
rect 3537 169 3583 180
rect 3761 222 3807 233
rect 3359 82 3761 90
rect 3807 82 3920 90
rect 0 -90 3920 82
<< labels >>
flabel metal1 s 142 354 315 449 0 FreeSans 200 0 0 0 CLKN
port 3 nsew clock input
flabel metal1 s 589 354 779 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3502 690 3583 766 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2676 335 2882 430 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 0 918 3920 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2685 233 2731 262 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3537 169 3583 690 1 Q
port 4 nsew default output
rlabel metal1 s 3741 869 3787 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3333 869 3379 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3169 869 3215 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2705 869 2751 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 869 1855 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 869 1507 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 869 691 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 869 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3741 775 3787 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3333 775 3379 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3169 775 3215 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 775 1855 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 775 1507 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 775 691 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 703 1855 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 703 1507 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 703 691 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 703 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 688 1855 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 688 691 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 688 319 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 685 691 688 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 688 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 609 691 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1685 233 1731 262 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 262 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3761 216 3807 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3313 216 3359 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2685 216 2731 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1685 216 1731 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 216 687 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3761 90 3807 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3313 90 3359 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2685 90 2731 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1685 90 1731 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3920 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 1008
string GDS_END 1499268
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1490096
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
