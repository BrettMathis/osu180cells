magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 1000
rect 224 0 344 1000
<< mvndiff >>
rect -88 987 0 1000
rect -88 941 -75 987
rect -29 941 0 987
rect -88 884 0 941
rect -88 838 -75 884
rect -29 838 0 884
rect -88 781 0 838
rect -88 735 -75 781
rect -29 735 0 781
rect -88 678 0 735
rect -88 632 -75 678
rect -29 632 0 678
rect -88 575 0 632
rect -88 529 -75 575
rect -29 529 0 575
rect -88 472 0 529
rect -88 426 -75 472
rect -29 426 0 472
rect -88 369 0 426
rect -88 323 -75 369
rect -29 323 0 369
rect -88 266 0 323
rect -88 220 -75 266
rect -29 220 0 266
rect -88 163 0 220
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 987 224 1000
rect 120 941 149 987
rect 195 941 224 987
rect 120 884 224 941
rect 120 838 149 884
rect 195 838 224 884
rect 120 781 224 838
rect 120 735 149 781
rect 195 735 224 781
rect 120 678 224 735
rect 120 632 149 678
rect 195 632 224 678
rect 120 575 224 632
rect 120 529 149 575
rect 195 529 224 575
rect 120 472 224 529
rect 120 426 149 472
rect 195 426 224 472
rect 120 369 224 426
rect 120 323 149 369
rect 195 323 224 369
rect 120 266 224 323
rect 120 220 149 266
rect 195 220 224 266
rect 120 163 224 220
rect 120 117 149 163
rect 195 117 224 163
rect 120 59 224 117
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 987 432 1000
rect 344 941 373 987
rect 419 941 432 987
rect 344 884 432 941
rect 344 838 373 884
rect 419 838 432 884
rect 344 781 432 838
rect 344 735 373 781
rect 419 735 432 781
rect 344 678 432 735
rect 344 632 373 678
rect 419 632 432 678
rect 344 575 432 632
rect 344 529 373 575
rect 419 529 432 575
rect 344 472 432 529
rect 344 426 373 472
rect 419 426 432 472
rect 344 369 432 426
rect 344 323 373 369
rect 419 323 432 369
rect 344 266 432 323
rect 344 220 373 266
rect 419 220 432 266
rect 344 163 432 220
rect 344 117 373 163
rect 419 117 432 163
rect 344 59 432 117
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvndiffc >>
rect -75 941 -29 987
rect -75 838 -29 884
rect -75 735 -29 781
rect -75 632 -29 678
rect -75 529 -29 575
rect -75 426 -29 472
rect -75 323 -29 369
rect -75 220 -29 266
rect -75 117 -29 163
rect -75 13 -29 59
rect 149 941 195 987
rect 149 838 195 884
rect 149 735 195 781
rect 149 632 195 678
rect 149 529 195 575
rect 149 426 195 472
rect 149 323 195 369
rect 149 220 195 266
rect 149 117 195 163
rect 149 13 195 59
rect 373 941 419 987
rect 373 838 419 884
rect 373 735 419 781
rect 373 632 419 678
rect 373 529 419 575
rect 373 426 419 472
rect 373 323 419 369
rect 373 220 419 266
rect 373 117 419 163
rect 373 13 419 59
<< polysilicon >>
rect 0 1000 120 1044
rect 224 1000 344 1044
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 987 -29 1000
rect -75 884 -29 941
rect -75 781 -29 838
rect -75 678 -29 735
rect -75 575 -29 632
rect -75 472 -29 529
rect -75 369 -29 426
rect -75 266 -29 323
rect -75 163 -29 220
rect -75 59 -29 117
rect -75 0 -29 13
rect 149 987 195 1000
rect 149 884 195 941
rect 149 781 195 838
rect 149 678 195 735
rect 149 575 195 632
rect 149 472 195 529
rect 149 369 195 426
rect 149 266 195 323
rect 149 163 195 220
rect 149 59 195 117
rect 149 0 195 13
rect 373 987 419 1000
rect 373 884 419 941
rect 373 781 419 838
rect 373 678 419 735
rect 373 575 419 632
rect 373 472 419 529
rect 373 369 419 426
rect 373 266 419 323
rect 373 163 419 220
rect 373 59 419 117
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 500 -52 500 0 FreeSans 200 0 0 0 S
flabel metal1 s 396 500 396 500 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 500 172 500 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 332774
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 329576
<< end >>
