magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< pwell >>
rect 2995 6633 5171 11633
rect 5431 6633 7607 11633
rect 7867 6633 10043 11633
rect 7867 621 10043 5621
<< mvnmos >>
rect 3083 6633 5083 11633
rect 5519 6633 7519 11633
rect 7955 6633 9955 11633
rect 7955 621 9955 5621
<< mvndiff >>
rect 2995 11596 3083 11633
rect 2995 6670 3008 11596
rect 3054 6670 3083 11596
rect 2995 6633 3083 6670
rect 5083 11596 5171 11633
rect 5083 6670 5112 11596
rect 5158 6670 5171 11596
rect 5083 6633 5171 6670
rect 5431 11596 5519 11633
rect 5431 6670 5444 11596
rect 5490 6670 5519 11596
rect 5431 6633 5519 6670
rect 7519 11596 7607 11633
rect 7519 6670 7548 11596
rect 7594 6670 7607 11596
rect 7519 6633 7607 6670
rect 7867 11596 7955 11633
rect 7867 6670 7880 11596
rect 7926 6670 7955 11596
rect 7867 6633 7955 6670
rect 9955 11596 10043 11633
rect 9955 6670 9984 11596
rect 10030 6670 10043 11596
rect 9955 6633 10043 6670
rect 7867 5584 7955 5621
rect 7867 658 7880 5584
rect 7926 658 7955 5584
rect 7867 621 7955 658
rect 9955 5584 10043 5621
rect 9955 658 9984 5584
rect 10030 658 10043 5584
rect 9955 621 10043 658
<< mvndiffc >>
rect 3008 6670 3054 11596
rect 5112 6670 5158 11596
rect 5444 6670 5490 11596
rect 7548 6670 7594 11596
rect 7880 6670 7926 11596
rect 9984 6670 10030 11596
rect 7880 658 7926 5584
rect 9984 658 10030 5584
<< psubdiff >>
rect 2285 12298 10576 12320
rect 2285 12252 2307 12298
rect 2353 12252 2421 12298
rect 2467 12252 2575 12298
rect 2621 12252 2689 12298
rect 2735 12252 2803 12298
rect 2849 12252 2917 12298
rect 2963 12252 3031 12298
rect 3077 12252 3145 12298
rect 3191 12252 3259 12298
rect 3305 12252 3373 12298
rect 3419 12252 3487 12298
rect 3533 12252 3601 12298
rect 3647 12252 3715 12298
rect 3761 12252 3829 12298
rect 3875 12252 3943 12298
rect 3989 12252 4057 12298
rect 4103 12252 4171 12298
rect 4217 12252 4285 12298
rect 4331 12252 4399 12298
rect 4445 12252 4513 12298
rect 4559 12252 4627 12298
rect 4673 12252 4741 12298
rect 4787 12252 4855 12298
rect 4901 12252 4969 12298
rect 5015 12252 5083 12298
rect 5129 12252 5197 12298
rect 5243 12252 5311 12298
rect 5357 12252 5425 12298
rect 5471 12252 5539 12298
rect 5585 12252 5653 12298
rect 5699 12252 5767 12298
rect 5813 12252 5881 12298
rect 5927 12252 5995 12298
rect 6041 12252 6109 12298
rect 6155 12252 6223 12298
rect 6269 12252 6337 12298
rect 6383 12252 6451 12298
rect 6497 12252 6565 12298
rect 6611 12252 6679 12298
rect 6725 12252 6793 12298
rect 6839 12252 6907 12298
rect 6953 12252 7021 12298
rect 7067 12252 7135 12298
rect 7181 12252 7249 12298
rect 7295 12252 7363 12298
rect 7409 12252 7477 12298
rect 7523 12252 7591 12298
rect 7637 12252 7705 12298
rect 7751 12252 7819 12298
rect 7865 12252 7933 12298
rect 7979 12252 8047 12298
rect 8093 12252 8161 12298
rect 8207 12252 8275 12298
rect 8321 12252 8389 12298
rect 8435 12252 8503 12298
rect 8549 12252 8617 12298
rect 8663 12252 8731 12298
rect 8777 12252 8845 12298
rect 8891 12252 8959 12298
rect 9005 12252 9073 12298
rect 9119 12252 9187 12298
rect 9233 12252 9301 12298
rect 9347 12252 9415 12298
rect 9461 12252 9529 12298
rect 9575 12252 9643 12298
rect 9689 12252 9757 12298
rect 9803 12252 9871 12298
rect 9917 12252 9985 12298
rect 10031 12252 10099 12298
rect 10145 12252 10213 12298
rect 10259 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10576 12298
rect 2285 12184 10576 12252
rect 2285 12138 2307 12184
rect 2353 12138 2421 12184
rect 2467 12138 2575 12184
rect 2621 12138 2689 12184
rect 2735 12138 2803 12184
rect 2849 12138 2917 12184
rect 2963 12138 3031 12184
rect 3077 12138 3145 12184
rect 3191 12138 3259 12184
rect 3305 12138 3373 12184
rect 3419 12138 3487 12184
rect 3533 12138 3601 12184
rect 3647 12138 3715 12184
rect 3761 12138 3829 12184
rect 3875 12138 3943 12184
rect 3989 12138 4057 12184
rect 4103 12138 4171 12184
rect 4217 12138 4285 12184
rect 4331 12138 4399 12184
rect 4445 12138 4513 12184
rect 4559 12138 4627 12184
rect 4673 12138 4741 12184
rect 4787 12138 4855 12184
rect 4901 12138 4969 12184
rect 5015 12138 5083 12184
rect 5129 12138 5197 12184
rect 5243 12138 5311 12184
rect 5357 12138 5425 12184
rect 5471 12138 5539 12184
rect 5585 12138 5653 12184
rect 5699 12138 5767 12184
rect 5813 12138 5881 12184
rect 5927 12138 5995 12184
rect 6041 12138 6109 12184
rect 6155 12138 6223 12184
rect 6269 12138 6337 12184
rect 6383 12138 6451 12184
rect 6497 12138 6565 12184
rect 6611 12138 6679 12184
rect 6725 12138 6793 12184
rect 6839 12138 6907 12184
rect 6953 12138 7021 12184
rect 7067 12138 7135 12184
rect 7181 12138 7249 12184
rect 7295 12138 7363 12184
rect 7409 12138 7477 12184
rect 7523 12138 7591 12184
rect 7637 12138 7705 12184
rect 7751 12138 7819 12184
rect 7865 12138 7933 12184
rect 7979 12138 8047 12184
rect 8093 12138 8161 12184
rect 8207 12138 8275 12184
rect 8321 12138 8389 12184
rect 8435 12138 8503 12184
rect 8549 12138 8617 12184
rect 8663 12138 8731 12184
rect 8777 12138 8845 12184
rect 8891 12138 8959 12184
rect 9005 12138 9073 12184
rect 9119 12138 9187 12184
rect 9233 12138 9301 12184
rect 9347 12138 9415 12184
rect 9461 12138 9529 12184
rect 9575 12138 9643 12184
rect 9689 12138 9757 12184
rect 9803 12138 9871 12184
rect 9917 12138 9985 12184
rect 10031 12138 10099 12184
rect 10145 12138 10213 12184
rect 10259 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10576 12184
rect 2285 12116 10576 12138
rect 2285 12070 2489 12116
rect 2285 12024 2307 12070
rect 2353 12024 2421 12070
rect 2467 12024 2489 12070
rect 2285 11500 2489 12024
rect 10372 12070 10576 12116
rect 10372 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10576 12070
rect 10372 11956 10576 12024
rect 10372 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10576 11956
rect 10372 11842 10576 11910
rect 10372 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10576 11842
rect 10372 11728 10576 11796
rect 10372 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10576 11728
rect 2285 11454 2307 11500
rect 2353 11454 2421 11500
rect 2467 11454 2489 11500
rect 2285 11386 2489 11454
rect 2285 11340 2307 11386
rect 2353 11340 2421 11386
rect 2467 11340 2489 11386
rect 2285 11272 2489 11340
rect 2285 11226 2307 11272
rect 2353 11226 2421 11272
rect 2467 11226 2489 11272
rect 2285 11158 2489 11226
rect 2285 11112 2307 11158
rect 2353 11112 2421 11158
rect 2467 11112 2489 11158
rect 2285 11044 2489 11112
rect 2285 10998 2307 11044
rect 2353 10998 2421 11044
rect 2467 10998 2489 11044
rect 2285 10930 2489 10998
rect 2285 10884 2307 10930
rect 2353 10884 2421 10930
rect 2467 10884 2489 10930
rect 2285 10816 2489 10884
rect 2285 10770 2307 10816
rect 2353 10770 2421 10816
rect 2467 10770 2489 10816
rect 2285 10702 2489 10770
rect 2285 10656 2307 10702
rect 2353 10656 2421 10702
rect 2467 10656 2489 10702
rect 2285 10588 2489 10656
rect 2285 10542 2307 10588
rect 2353 10542 2421 10588
rect 2467 10542 2489 10588
rect 2285 10474 2489 10542
rect 2285 10428 2307 10474
rect 2353 10428 2421 10474
rect 2467 10428 2489 10474
rect 2285 10360 2489 10428
rect 2285 10314 2307 10360
rect 2353 10314 2421 10360
rect 2467 10314 2489 10360
rect 2285 10246 2489 10314
rect 2285 10200 2307 10246
rect 2353 10200 2421 10246
rect 2467 10200 2489 10246
rect 2285 10132 2489 10200
rect 2285 10086 2307 10132
rect 2353 10086 2421 10132
rect 2467 10086 2489 10132
rect 2285 10018 2489 10086
rect 2285 9972 2307 10018
rect 2353 9972 2421 10018
rect 2467 9972 2489 10018
rect 2285 9904 2489 9972
rect 2285 9858 2307 9904
rect 2353 9858 2421 9904
rect 2467 9858 2489 9904
rect 2285 9790 2489 9858
rect 2285 9744 2307 9790
rect 2353 9744 2421 9790
rect 2467 9744 2489 9790
rect 2285 9676 2489 9744
rect 2285 9630 2307 9676
rect 2353 9630 2421 9676
rect 2467 9630 2489 9676
rect 2285 9562 2489 9630
rect 2285 9516 2307 9562
rect 2353 9516 2421 9562
rect 2467 9516 2489 9562
rect 2285 9448 2489 9516
rect 2285 9402 2307 9448
rect 2353 9402 2421 9448
rect 2467 9402 2489 9448
rect 2285 9334 2489 9402
rect 2285 9288 2307 9334
rect 2353 9288 2421 9334
rect 2467 9288 2489 9334
rect 2285 9220 2489 9288
rect 2285 9174 2307 9220
rect 2353 9174 2421 9220
rect 2467 9174 2489 9220
rect 2285 9106 2489 9174
rect 2285 9060 2307 9106
rect 2353 9060 2421 9106
rect 2467 9060 2489 9106
rect 2285 8992 2489 9060
rect 2285 8946 2307 8992
rect 2353 8946 2421 8992
rect 2467 8946 2489 8992
rect 2285 8878 2489 8946
rect 2285 8832 2307 8878
rect 2353 8832 2421 8878
rect 2467 8832 2489 8878
rect 2285 8764 2489 8832
rect 2285 8718 2307 8764
rect 2353 8718 2421 8764
rect 2467 8718 2489 8764
rect 2285 8650 2489 8718
rect 2285 8604 2307 8650
rect 2353 8604 2421 8650
rect 2467 8604 2489 8650
rect 2285 8536 2489 8604
rect 2285 8490 2307 8536
rect 2353 8490 2421 8536
rect 2467 8490 2489 8536
rect 2285 8422 2489 8490
rect 2285 8376 2307 8422
rect 2353 8376 2421 8422
rect 2467 8376 2489 8422
rect 2285 8308 2489 8376
rect 2285 8262 2307 8308
rect 2353 8262 2421 8308
rect 2467 8262 2489 8308
rect 2285 8194 2489 8262
rect 2285 8148 2307 8194
rect 2353 8148 2421 8194
rect 2467 8148 2489 8194
rect 2285 8080 2489 8148
rect 2285 8034 2307 8080
rect 2353 8034 2421 8080
rect 2467 8034 2489 8080
rect 2285 7966 2489 8034
rect 2285 7920 2307 7966
rect 2353 7920 2421 7966
rect 2467 7920 2489 7966
rect 2285 7852 2489 7920
rect 2285 7806 2307 7852
rect 2353 7806 2421 7852
rect 2467 7806 2489 7852
rect 2285 7738 2489 7806
rect 2285 7692 2307 7738
rect 2353 7692 2421 7738
rect 2467 7692 2489 7738
rect 2285 7624 2489 7692
rect 2285 7578 2307 7624
rect 2353 7578 2421 7624
rect 2467 7578 2489 7624
rect 2285 7510 2489 7578
rect 2285 7464 2307 7510
rect 2353 7464 2421 7510
rect 2467 7464 2489 7510
rect 2285 7396 2489 7464
rect 2285 7350 2307 7396
rect 2353 7350 2421 7396
rect 2467 7350 2489 7396
rect 2285 7282 2489 7350
rect 2285 7236 2307 7282
rect 2353 7236 2421 7282
rect 2467 7236 2489 7282
rect 2285 7168 2489 7236
rect 2285 7122 2307 7168
rect 2353 7122 2421 7168
rect 2467 7122 2489 7168
rect 2285 7054 2489 7122
rect 2285 7008 2307 7054
rect 2353 7008 2421 7054
rect 2467 7008 2489 7054
rect 2285 6940 2489 7008
rect 2285 6894 2307 6940
rect 2353 6894 2421 6940
rect 2467 6894 2489 6940
rect 2285 6826 2489 6894
rect 2285 6780 2307 6826
rect 2353 6780 2421 6826
rect 2467 6780 2489 6826
rect 2285 6712 2489 6780
rect 2285 6666 2307 6712
rect 2353 6666 2421 6712
rect 2467 6666 2489 6712
rect 2285 6598 2489 6666
rect 10372 11614 10576 11682
rect 10372 11568 10394 11614
rect 10440 11568 10508 11614
rect 10554 11568 10576 11614
rect 10372 11500 10576 11568
rect 10372 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10576 11500
rect 10372 11386 10576 11454
rect 10372 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10576 11386
rect 10372 11272 10576 11340
rect 10372 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10576 11272
rect 10372 11158 10576 11226
rect 10372 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10576 11158
rect 10372 11044 10576 11112
rect 10372 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10576 11044
rect 10372 10930 10576 10998
rect 10372 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10576 10930
rect 10372 10816 10576 10884
rect 10372 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10576 10816
rect 10372 10702 10576 10770
rect 10372 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10576 10702
rect 10372 10588 10576 10656
rect 10372 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10576 10588
rect 10372 10474 10576 10542
rect 10372 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10576 10474
rect 10372 10360 10576 10428
rect 10372 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10576 10360
rect 10372 10246 10576 10314
rect 10372 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10576 10246
rect 10372 10132 10576 10200
rect 10372 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10576 10132
rect 10372 10018 10576 10086
rect 10372 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10576 10018
rect 10372 9904 10576 9972
rect 10372 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10576 9904
rect 10372 9790 10576 9858
rect 10372 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10576 9790
rect 10372 9676 10576 9744
rect 10372 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10576 9676
rect 10372 9562 10576 9630
rect 10372 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10576 9562
rect 10372 9448 10576 9516
rect 10372 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10576 9448
rect 10372 9334 10576 9402
rect 10372 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10576 9334
rect 10372 9220 10576 9288
rect 10372 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10576 9220
rect 10372 9106 10576 9174
rect 10372 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10576 9106
rect 10372 8992 10576 9060
rect 10372 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10576 8992
rect 10372 8878 10576 8946
rect 10372 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10576 8878
rect 10372 8764 10576 8832
rect 10372 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10576 8764
rect 10372 8650 10576 8718
rect 10372 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10576 8650
rect 10372 8536 10576 8604
rect 10372 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10576 8536
rect 10372 8422 10576 8490
rect 10372 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10576 8422
rect 10372 8308 10576 8376
rect 10372 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10576 8308
rect 10372 8194 10576 8262
rect 10372 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10576 8194
rect 10372 8080 10576 8148
rect 10372 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10576 8080
rect 10372 7966 10576 8034
rect 10372 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10576 7966
rect 10372 7852 10576 7920
rect 10372 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10576 7852
rect 10372 7738 10576 7806
rect 10372 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10576 7738
rect 10372 7624 10576 7692
rect 10372 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10576 7624
rect 10372 7510 10576 7578
rect 10372 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10576 7510
rect 10372 7396 10576 7464
rect 10372 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10576 7396
rect 10372 7282 10576 7350
rect 10372 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10576 7282
rect 10372 7168 10576 7236
rect 10372 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10576 7168
rect 10372 7054 10576 7122
rect 10372 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10576 7054
rect 10372 6940 10576 7008
rect 10372 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10576 6940
rect 10372 6826 10576 6894
rect 10372 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10576 6826
rect 10372 6712 10576 6780
rect 10372 6666 10394 6712
rect 10440 6666 10508 6712
rect 10554 6666 10576 6712
rect 2285 6552 2307 6598
rect 2353 6552 2421 6598
rect 2467 6552 2489 6598
rect 2285 6484 2489 6552
rect 10372 6598 10576 6666
rect 10372 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10576 6598
rect 2285 6438 2307 6484
rect 2353 6438 2421 6484
rect 2467 6438 2489 6484
rect 2285 6370 2489 6438
rect 2285 6324 2307 6370
rect 2353 6324 2421 6370
rect 2467 6324 2489 6370
rect 2285 6229 2489 6324
rect 10372 6484 10576 6552
rect 10372 6438 10394 6484
rect 10440 6438 10508 6484
rect 10554 6438 10576 6484
rect 10372 6370 10576 6438
rect 10372 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10576 6370
rect 10372 6256 10576 6324
rect 10372 6229 10394 6256
rect 2285 6210 10394 6229
rect 10440 6210 10508 6256
rect 10554 6210 10576 6256
rect 2285 6207 10576 6210
rect 2285 6161 2540 6207
rect 2586 6161 2654 6207
rect 2700 6161 2768 6207
rect 2814 6161 2882 6207
rect 2928 6161 2996 6207
rect 3042 6161 3110 6207
rect 3156 6161 3224 6207
rect 3270 6161 3338 6207
rect 3384 6161 3452 6207
rect 3498 6161 3566 6207
rect 3612 6161 3680 6207
rect 3726 6161 3794 6207
rect 3840 6161 3908 6207
rect 3954 6161 4022 6207
rect 4068 6161 4136 6207
rect 4182 6161 4250 6207
rect 4296 6161 4364 6207
rect 4410 6161 4478 6207
rect 4524 6161 4592 6207
rect 4638 6161 4706 6207
rect 4752 6161 4820 6207
rect 4866 6161 4934 6207
rect 4980 6161 5048 6207
rect 5094 6161 5162 6207
rect 5208 6161 5276 6207
rect 5322 6161 5390 6207
rect 5436 6161 5504 6207
rect 5550 6161 5618 6207
rect 5664 6161 5732 6207
rect 5778 6161 5846 6207
rect 5892 6161 5960 6207
rect 6006 6161 6074 6207
rect 6120 6161 6188 6207
rect 6234 6161 6302 6207
rect 6348 6161 6416 6207
rect 6462 6161 6530 6207
rect 6576 6161 6644 6207
rect 6690 6161 6758 6207
rect 6804 6161 6872 6207
rect 6918 6161 6986 6207
rect 7032 6161 7100 6207
rect 7146 6161 7214 6207
rect 7260 6161 7328 6207
rect 7374 6161 7442 6207
rect 7488 6161 7556 6207
rect 7602 6161 7670 6207
rect 7716 6161 7784 6207
rect 7830 6161 7898 6207
rect 7944 6161 8012 6207
rect 8058 6161 8126 6207
rect 8172 6161 8240 6207
rect 8286 6161 8354 6207
rect 8400 6161 8468 6207
rect 8514 6161 8582 6207
rect 8628 6161 8696 6207
rect 8742 6161 8810 6207
rect 8856 6161 8924 6207
rect 8970 6161 9038 6207
rect 9084 6161 9152 6207
rect 9198 6161 9266 6207
rect 9312 6161 9380 6207
rect 9426 6161 9494 6207
rect 9540 6161 9608 6207
rect 9654 6161 9722 6207
rect 9768 6161 9836 6207
rect 9882 6161 9950 6207
rect 9996 6161 10064 6207
rect 10110 6161 10178 6207
rect 10224 6161 10292 6207
rect 10338 6161 10576 6207
rect 2285 6142 10576 6161
rect 2285 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10576 6142
rect 2285 6093 10576 6096
rect 2285 6047 2540 6093
rect 2586 6047 2654 6093
rect 2700 6047 2768 6093
rect 2814 6047 2882 6093
rect 2928 6047 2996 6093
rect 3042 6047 3110 6093
rect 3156 6047 3224 6093
rect 3270 6047 3338 6093
rect 3384 6047 3452 6093
rect 3498 6047 3566 6093
rect 3612 6047 3680 6093
rect 3726 6047 3794 6093
rect 3840 6047 3908 6093
rect 3954 6047 4022 6093
rect 4068 6047 4136 6093
rect 4182 6047 4250 6093
rect 4296 6047 4364 6093
rect 4410 6047 4478 6093
rect 4524 6047 4592 6093
rect 4638 6047 4706 6093
rect 4752 6047 4820 6093
rect 4866 6047 4934 6093
rect 4980 6047 5048 6093
rect 5094 6047 5162 6093
rect 5208 6047 5276 6093
rect 5322 6047 5390 6093
rect 5436 6047 5504 6093
rect 5550 6047 5618 6093
rect 5664 6047 5732 6093
rect 5778 6047 5846 6093
rect 5892 6047 5960 6093
rect 6006 6047 6074 6093
rect 6120 6047 6188 6093
rect 6234 6047 6302 6093
rect 6348 6047 6416 6093
rect 6462 6047 6530 6093
rect 6576 6047 6644 6093
rect 6690 6047 6758 6093
rect 6804 6047 6872 6093
rect 6918 6047 6986 6093
rect 7032 6047 7100 6093
rect 7146 6047 7214 6093
rect 7260 6047 7328 6093
rect 7374 6047 7442 6093
rect 7488 6047 7556 6093
rect 7602 6047 7670 6093
rect 7716 6047 7784 6093
rect 7830 6047 7898 6093
rect 7944 6047 8012 6093
rect 8058 6047 8126 6093
rect 8172 6047 8240 6093
rect 8286 6047 8354 6093
rect 8400 6047 8468 6093
rect 8514 6047 8582 6093
rect 8628 6047 8696 6093
rect 8742 6047 8810 6093
rect 8856 6047 8924 6093
rect 8970 6047 9038 6093
rect 9084 6047 9152 6093
rect 9198 6047 9266 6093
rect 9312 6047 9380 6093
rect 9426 6047 9494 6093
rect 9540 6047 9608 6093
rect 9654 6047 9722 6093
rect 9768 6047 9836 6093
rect 9882 6047 9950 6093
rect 9996 6047 10064 6093
rect 10110 6047 10178 6093
rect 10224 6047 10292 6093
rect 10338 6047 10576 6093
rect 2285 6028 10576 6047
rect 2285 6025 10394 6028
rect 7260 5951 7474 6025
rect 7260 5905 7282 5951
rect 7328 5905 7406 5951
rect 7452 5905 7474 5951
rect 7260 5827 7474 5905
rect 7260 5781 7282 5827
rect 7328 5781 7406 5827
rect 7452 5781 7474 5827
rect 7260 5703 7474 5781
rect 10372 5982 10394 6025
rect 10440 5982 10508 6028
rect 10554 5982 10576 6028
rect 10372 5914 10576 5982
rect 10372 5868 10394 5914
rect 10440 5868 10508 5914
rect 10554 5868 10576 5914
rect 10372 5800 10576 5868
rect 10372 5754 10394 5800
rect 10440 5754 10508 5800
rect 10554 5754 10576 5800
rect 7260 5657 7282 5703
rect 7328 5657 7406 5703
rect 7452 5657 7474 5703
rect 7260 5579 7474 5657
rect 10372 5686 10576 5754
rect 10372 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10576 5686
rect 7260 5533 7282 5579
rect 7328 5533 7406 5579
rect 7452 5533 7474 5579
rect 7260 5455 7474 5533
rect 7260 5409 7282 5455
rect 7328 5409 7406 5455
rect 7452 5409 7474 5455
rect 7260 5331 7474 5409
rect 7260 5285 7282 5331
rect 7328 5285 7406 5331
rect 7452 5285 7474 5331
rect 7260 5207 7474 5285
rect 7260 5161 7282 5207
rect 7328 5161 7406 5207
rect 7452 5161 7474 5207
rect 7260 5083 7474 5161
rect 7260 5037 7282 5083
rect 7328 5037 7406 5083
rect 7452 5037 7474 5083
rect 7260 4959 7474 5037
rect 7260 4913 7282 4959
rect 7328 4913 7406 4959
rect 7452 4913 7474 4959
rect 7260 4835 7474 4913
rect 7260 4789 7282 4835
rect 7328 4789 7406 4835
rect 7452 4789 7474 4835
rect 7260 4711 7474 4789
rect 7260 4665 7282 4711
rect 7328 4665 7406 4711
rect 7452 4665 7474 4711
rect 7260 4587 7474 4665
rect 7260 4541 7282 4587
rect 7328 4541 7406 4587
rect 7452 4541 7474 4587
rect 7260 4463 7474 4541
rect 7260 4417 7282 4463
rect 7328 4417 7406 4463
rect 7452 4417 7474 4463
rect 7260 4339 7474 4417
rect 7260 4293 7282 4339
rect 7328 4293 7406 4339
rect 7452 4293 7474 4339
rect 7260 4215 7474 4293
rect 7260 4169 7282 4215
rect 7328 4169 7406 4215
rect 7452 4169 7474 4215
rect 7260 4091 7474 4169
rect 7260 4045 7282 4091
rect 7328 4045 7406 4091
rect 7452 4045 7474 4091
rect 7260 3967 7474 4045
rect 7260 3921 7282 3967
rect 7328 3921 7406 3967
rect 7452 3921 7474 3967
rect 7260 3843 7474 3921
rect 7260 3797 7282 3843
rect 7328 3797 7406 3843
rect 7452 3797 7474 3843
rect 7260 3719 7474 3797
rect 7260 3673 7282 3719
rect 7328 3673 7406 3719
rect 7452 3673 7474 3719
rect 7260 3595 7474 3673
rect 7260 3549 7282 3595
rect 7328 3549 7406 3595
rect 7452 3549 7474 3595
rect 7260 3471 7474 3549
rect 7260 3425 7282 3471
rect 7328 3425 7406 3471
rect 7452 3425 7474 3471
rect 7260 3347 7474 3425
rect 7260 3301 7282 3347
rect 7328 3301 7406 3347
rect 7452 3301 7474 3347
rect 7260 3223 7474 3301
rect 7260 3177 7282 3223
rect 7328 3177 7406 3223
rect 7452 3177 7474 3223
rect 7260 3099 7474 3177
rect 7260 3053 7282 3099
rect 7328 3053 7406 3099
rect 7452 3053 7474 3099
rect 7260 2975 7474 3053
rect 7260 2929 7282 2975
rect 7328 2929 7406 2975
rect 7452 2929 7474 2975
rect 7260 2851 7474 2929
rect 7260 2805 7282 2851
rect 7328 2805 7406 2851
rect 7452 2805 7474 2851
rect 7260 2727 7474 2805
rect 7260 2681 7282 2727
rect 7328 2681 7406 2727
rect 7452 2681 7474 2727
rect 7260 2603 7474 2681
rect 7260 2557 7282 2603
rect 7328 2557 7406 2603
rect 7452 2557 7474 2603
rect 7260 2479 7474 2557
rect 7260 2433 7282 2479
rect 7328 2433 7406 2479
rect 7452 2433 7474 2479
rect 7260 2355 7474 2433
rect 7260 2309 7282 2355
rect 7328 2309 7406 2355
rect 7452 2309 7474 2355
rect 7260 2231 7474 2309
rect 7260 2185 7282 2231
rect 7328 2185 7406 2231
rect 7452 2185 7474 2231
rect 7260 2107 7474 2185
rect 7260 2061 7282 2107
rect 7328 2061 7406 2107
rect 7452 2061 7474 2107
rect 7260 1983 7474 2061
rect 7260 1937 7282 1983
rect 7328 1937 7406 1983
rect 7452 1937 7474 1983
rect 7260 1859 7474 1937
rect 7260 1813 7282 1859
rect 7328 1813 7406 1859
rect 7452 1813 7474 1859
rect 7260 1735 7474 1813
rect 7260 1689 7282 1735
rect 7328 1689 7406 1735
rect 7452 1689 7474 1735
rect 7260 1611 7474 1689
rect 7260 1565 7282 1611
rect 7328 1565 7406 1611
rect 7452 1565 7474 1611
rect 7260 1487 7474 1565
rect 7260 1441 7282 1487
rect 7328 1441 7406 1487
rect 7452 1441 7474 1487
rect 7260 1363 7474 1441
rect 7260 1317 7282 1363
rect 7328 1317 7406 1363
rect 7452 1317 7474 1363
rect 7260 1239 7474 1317
rect 7260 1193 7282 1239
rect 7328 1193 7406 1239
rect 7452 1193 7474 1239
rect 7260 1115 7474 1193
rect 7260 1069 7282 1115
rect 7328 1069 7406 1115
rect 7452 1069 7474 1115
rect 7260 991 7474 1069
rect 7260 945 7282 991
rect 7328 945 7406 991
rect 7452 945 7474 991
rect 7260 867 7474 945
rect 7260 821 7282 867
rect 7328 821 7406 867
rect 7452 821 7474 867
rect 7260 743 7474 821
rect 7260 697 7282 743
rect 7328 697 7406 743
rect 7452 697 7474 743
rect 7260 619 7474 697
rect 10372 5572 10576 5640
rect 10372 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10576 5572
rect 10372 5458 10576 5526
rect 10372 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10576 5458
rect 10372 5344 10576 5412
rect 10372 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10576 5344
rect 10372 5230 10576 5298
rect 10372 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10576 5230
rect 10372 5116 10576 5184
rect 10372 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10576 5116
rect 10372 5002 10576 5070
rect 10372 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10576 5002
rect 10372 4888 10576 4956
rect 10372 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10576 4888
rect 10372 4774 10576 4842
rect 10372 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10576 4774
rect 10372 4660 10576 4728
rect 10372 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10576 4660
rect 10372 4546 10576 4614
rect 10372 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10576 4546
rect 10372 4432 10576 4500
rect 10372 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10576 4432
rect 10372 4318 10576 4386
rect 10372 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10576 4318
rect 10372 4204 10576 4272
rect 10372 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10576 4204
rect 10372 4090 10576 4158
rect 10372 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10576 4090
rect 10372 3976 10576 4044
rect 10372 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10576 3976
rect 10372 3862 10576 3930
rect 10372 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10576 3862
rect 10372 3748 10576 3816
rect 10372 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10576 3748
rect 10372 3634 10576 3702
rect 10372 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10576 3634
rect 10372 3520 10576 3588
rect 10372 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10576 3520
rect 10372 3406 10576 3474
rect 10372 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10576 3406
rect 10372 3292 10576 3360
rect 10372 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10576 3292
rect 10372 3178 10576 3246
rect 10372 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10576 3178
rect 10372 3064 10576 3132
rect 10372 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10576 3064
rect 10372 2950 10576 3018
rect 10372 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10576 2950
rect 10372 2836 10576 2904
rect 10372 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10576 2836
rect 10372 2722 10576 2790
rect 10372 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10576 2722
rect 10372 2608 10576 2676
rect 10372 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10576 2608
rect 10372 2494 10576 2562
rect 10372 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10576 2494
rect 10372 2380 10576 2448
rect 10372 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10576 2380
rect 10372 2266 10576 2334
rect 10372 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10576 2266
rect 10372 2152 10576 2220
rect 10372 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10576 2152
rect 10372 2038 10576 2106
rect 10372 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10576 2038
rect 10372 1924 10576 1992
rect 10372 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10576 1924
rect 10372 1810 10576 1878
rect 10372 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10576 1810
rect 10372 1696 10576 1764
rect 10372 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10576 1696
rect 10372 1582 10576 1650
rect 10372 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10576 1582
rect 10372 1468 10576 1536
rect 10372 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10576 1468
rect 10372 1354 10576 1422
rect 10372 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10576 1354
rect 10372 1240 10576 1308
rect 10372 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10576 1240
rect 10372 1126 10576 1194
rect 10372 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10576 1126
rect 10372 1012 10576 1080
rect 10372 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10576 1012
rect 10372 898 10576 966
rect 10372 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10576 898
rect 10372 784 10576 852
rect 10372 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10576 784
rect 10372 670 10576 738
rect 10372 624 10394 670
rect 10440 624 10508 670
rect 10554 624 10576 670
rect 7260 573 7282 619
rect 7328 573 7406 619
rect 7452 573 7474 619
rect 7260 495 7474 573
rect 10372 556 10576 624
rect 7260 449 7282 495
rect 7328 449 7406 495
rect 7452 449 7474 495
rect 7260 371 7474 449
rect 7260 325 7282 371
rect 7328 325 7406 371
rect 7452 325 7474 371
rect 7260 247 7474 325
rect 7260 201 7282 247
rect 7328 201 7406 247
rect 7452 236 7474 247
rect 10372 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10576 556
rect 10372 442 10576 510
rect 10372 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10576 442
rect 10372 328 10576 396
rect 10372 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10576 328
rect 10372 236 10576 282
rect 7452 214 10576 236
rect 7452 201 7612 214
rect 7260 168 7612 201
rect 7658 168 7726 214
rect 7772 168 7840 214
rect 7886 168 7954 214
rect 8000 168 8068 214
rect 8114 168 8182 214
rect 8228 168 8296 214
rect 8342 168 8410 214
rect 8456 168 8524 214
rect 8570 168 8638 214
rect 8684 168 8752 214
rect 8798 168 8866 214
rect 8912 168 8980 214
rect 9026 168 9094 214
rect 9140 168 9208 214
rect 9254 168 9322 214
rect 9368 168 9436 214
rect 9482 168 9550 214
rect 9596 168 9664 214
rect 9710 168 9778 214
rect 9824 168 9892 214
rect 9938 168 10006 214
rect 10052 168 10120 214
rect 10166 168 10234 214
rect 10280 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10576 214
rect 7260 123 10576 168
rect 7260 77 7282 123
rect 7328 77 7406 123
rect 7452 100 10576 123
rect 7452 77 7612 100
rect 7260 54 7612 77
rect 7658 54 7726 100
rect 7772 54 7840 100
rect 7886 54 7954 100
rect 8000 54 8068 100
rect 8114 54 8182 100
rect 8228 54 8296 100
rect 8342 54 8410 100
rect 8456 54 8524 100
rect 8570 54 8638 100
rect 8684 54 8752 100
rect 8798 54 8866 100
rect 8912 54 8980 100
rect 9026 54 9094 100
rect 9140 54 9208 100
rect 9254 54 9322 100
rect 9368 54 9436 100
rect 9482 54 9550 100
rect 9596 54 9664 100
rect 9710 54 9778 100
rect 9824 54 9892 100
rect 9938 54 10006 100
rect 10052 54 10120 100
rect 10166 54 10234 100
rect 10280 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10576 100
rect 7260 32 10576 54
<< psubdiffcont >>
rect 2307 12252 2353 12298
rect 2421 12252 2467 12298
rect 2575 12252 2621 12298
rect 2689 12252 2735 12298
rect 2803 12252 2849 12298
rect 2917 12252 2963 12298
rect 3031 12252 3077 12298
rect 3145 12252 3191 12298
rect 3259 12252 3305 12298
rect 3373 12252 3419 12298
rect 3487 12252 3533 12298
rect 3601 12252 3647 12298
rect 3715 12252 3761 12298
rect 3829 12252 3875 12298
rect 3943 12252 3989 12298
rect 4057 12252 4103 12298
rect 4171 12252 4217 12298
rect 4285 12252 4331 12298
rect 4399 12252 4445 12298
rect 4513 12252 4559 12298
rect 4627 12252 4673 12298
rect 4741 12252 4787 12298
rect 4855 12252 4901 12298
rect 4969 12252 5015 12298
rect 5083 12252 5129 12298
rect 5197 12252 5243 12298
rect 5311 12252 5357 12298
rect 5425 12252 5471 12298
rect 5539 12252 5585 12298
rect 5653 12252 5699 12298
rect 5767 12252 5813 12298
rect 5881 12252 5927 12298
rect 5995 12252 6041 12298
rect 6109 12252 6155 12298
rect 6223 12252 6269 12298
rect 6337 12252 6383 12298
rect 6451 12252 6497 12298
rect 6565 12252 6611 12298
rect 6679 12252 6725 12298
rect 6793 12252 6839 12298
rect 6907 12252 6953 12298
rect 7021 12252 7067 12298
rect 7135 12252 7181 12298
rect 7249 12252 7295 12298
rect 7363 12252 7409 12298
rect 7477 12252 7523 12298
rect 7591 12252 7637 12298
rect 7705 12252 7751 12298
rect 7819 12252 7865 12298
rect 7933 12252 7979 12298
rect 8047 12252 8093 12298
rect 8161 12252 8207 12298
rect 8275 12252 8321 12298
rect 8389 12252 8435 12298
rect 8503 12252 8549 12298
rect 8617 12252 8663 12298
rect 8731 12252 8777 12298
rect 8845 12252 8891 12298
rect 8959 12252 9005 12298
rect 9073 12252 9119 12298
rect 9187 12252 9233 12298
rect 9301 12252 9347 12298
rect 9415 12252 9461 12298
rect 9529 12252 9575 12298
rect 9643 12252 9689 12298
rect 9757 12252 9803 12298
rect 9871 12252 9917 12298
rect 9985 12252 10031 12298
rect 10099 12252 10145 12298
rect 10213 12252 10259 12298
rect 10394 12252 10440 12298
rect 10508 12252 10554 12298
rect 2307 12138 2353 12184
rect 2421 12138 2467 12184
rect 2575 12138 2621 12184
rect 2689 12138 2735 12184
rect 2803 12138 2849 12184
rect 2917 12138 2963 12184
rect 3031 12138 3077 12184
rect 3145 12138 3191 12184
rect 3259 12138 3305 12184
rect 3373 12138 3419 12184
rect 3487 12138 3533 12184
rect 3601 12138 3647 12184
rect 3715 12138 3761 12184
rect 3829 12138 3875 12184
rect 3943 12138 3989 12184
rect 4057 12138 4103 12184
rect 4171 12138 4217 12184
rect 4285 12138 4331 12184
rect 4399 12138 4445 12184
rect 4513 12138 4559 12184
rect 4627 12138 4673 12184
rect 4741 12138 4787 12184
rect 4855 12138 4901 12184
rect 4969 12138 5015 12184
rect 5083 12138 5129 12184
rect 5197 12138 5243 12184
rect 5311 12138 5357 12184
rect 5425 12138 5471 12184
rect 5539 12138 5585 12184
rect 5653 12138 5699 12184
rect 5767 12138 5813 12184
rect 5881 12138 5927 12184
rect 5995 12138 6041 12184
rect 6109 12138 6155 12184
rect 6223 12138 6269 12184
rect 6337 12138 6383 12184
rect 6451 12138 6497 12184
rect 6565 12138 6611 12184
rect 6679 12138 6725 12184
rect 6793 12138 6839 12184
rect 6907 12138 6953 12184
rect 7021 12138 7067 12184
rect 7135 12138 7181 12184
rect 7249 12138 7295 12184
rect 7363 12138 7409 12184
rect 7477 12138 7523 12184
rect 7591 12138 7637 12184
rect 7705 12138 7751 12184
rect 7819 12138 7865 12184
rect 7933 12138 7979 12184
rect 8047 12138 8093 12184
rect 8161 12138 8207 12184
rect 8275 12138 8321 12184
rect 8389 12138 8435 12184
rect 8503 12138 8549 12184
rect 8617 12138 8663 12184
rect 8731 12138 8777 12184
rect 8845 12138 8891 12184
rect 8959 12138 9005 12184
rect 9073 12138 9119 12184
rect 9187 12138 9233 12184
rect 9301 12138 9347 12184
rect 9415 12138 9461 12184
rect 9529 12138 9575 12184
rect 9643 12138 9689 12184
rect 9757 12138 9803 12184
rect 9871 12138 9917 12184
rect 9985 12138 10031 12184
rect 10099 12138 10145 12184
rect 10213 12138 10259 12184
rect 10394 12138 10440 12184
rect 10508 12138 10554 12184
rect 2307 12024 2353 12070
rect 2421 12024 2467 12070
rect 10394 12024 10440 12070
rect 10508 12024 10554 12070
rect 10394 11910 10440 11956
rect 10508 11910 10554 11956
rect 10394 11796 10440 11842
rect 10508 11796 10554 11842
rect 10394 11682 10440 11728
rect 10508 11682 10554 11728
rect 2307 11454 2353 11500
rect 2421 11454 2467 11500
rect 2307 11340 2353 11386
rect 2421 11340 2467 11386
rect 2307 11226 2353 11272
rect 2421 11226 2467 11272
rect 2307 11112 2353 11158
rect 2421 11112 2467 11158
rect 2307 10998 2353 11044
rect 2421 10998 2467 11044
rect 2307 10884 2353 10930
rect 2421 10884 2467 10930
rect 2307 10770 2353 10816
rect 2421 10770 2467 10816
rect 2307 10656 2353 10702
rect 2421 10656 2467 10702
rect 2307 10542 2353 10588
rect 2421 10542 2467 10588
rect 2307 10428 2353 10474
rect 2421 10428 2467 10474
rect 2307 10314 2353 10360
rect 2421 10314 2467 10360
rect 2307 10200 2353 10246
rect 2421 10200 2467 10246
rect 2307 10086 2353 10132
rect 2421 10086 2467 10132
rect 2307 9972 2353 10018
rect 2421 9972 2467 10018
rect 2307 9858 2353 9904
rect 2421 9858 2467 9904
rect 2307 9744 2353 9790
rect 2421 9744 2467 9790
rect 2307 9630 2353 9676
rect 2421 9630 2467 9676
rect 2307 9516 2353 9562
rect 2421 9516 2467 9562
rect 2307 9402 2353 9448
rect 2421 9402 2467 9448
rect 2307 9288 2353 9334
rect 2421 9288 2467 9334
rect 2307 9174 2353 9220
rect 2421 9174 2467 9220
rect 2307 9060 2353 9106
rect 2421 9060 2467 9106
rect 2307 8946 2353 8992
rect 2421 8946 2467 8992
rect 2307 8832 2353 8878
rect 2421 8832 2467 8878
rect 2307 8718 2353 8764
rect 2421 8718 2467 8764
rect 2307 8604 2353 8650
rect 2421 8604 2467 8650
rect 2307 8490 2353 8536
rect 2421 8490 2467 8536
rect 2307 8376 2353 8422
rect 2421 8376 2467 8422
rect 2307 8262 2353 8308
rect 2421 8262 2467 8308
rect 2307 8148 2353 8194
rect 2421 8148 2467 8194
rect 2307 8034 2353 8080
rect 2421 8034 2467 8080
rect 2307 7920 2353 7966
rect 2421 7920 2467 7966
rect 2307 7806 2353 7852
rect 2421 7806 2467 7852
rect 2307 7692 2353 7738
rect 2421 7692 2467 7738
rect 2307 7578 2353 7624
rect 2421 7578 2467 7624
rect 2307 7464 2353 7510
rect 2421 7464 2467 7510
rect 2307 7350 2353 7396
rect 2421 7350 2467 7396
rect 2307 7236 2353 7282
rect 2421 7236 2467 7282
rect 2307 7122 2353 7168
rect 2421 7122 2467 7168
rect 2307 7008 2353 7054
rect 2421 7008 2467 7054
rect 2307 6894 2353 6940
rect 2421 6894 2467 6940
rect 2307 6780 2353 6826
rect 2421 6780 2467 6826
rect 2307 6666 2353 6712
rect 2421 6666 2467 6712
rect 10394 11568 10440 11614
rect 10508 11568 10554 11614
rect 10394 11454 10440 11500
rect 10508 11454 10554 11500
rect 10394 11340 10440 11386
rect 10508 11340 10554 11386
rect 10394 11226 10440 11272
rect 10508 11226 10554 11272
rect 10394 11112 10440 11158
rect 10508 11112 10554 11158
rect 10394 10998 10440 11044
rect 10508 10998 10554 11044
rect 10394 10884 10440 10930
rect 10508 10884 10554 10930
rect 10394 10770 10440 10816
rect 10508 10770 10554 10816
rect 10394 10656 10440 10702
rect 10508 10656 10554 10702
rect 10394 10542 10440 10588
rect 10508 10542 10554 10588
rect 10394 10428 10440 10474
rect 10508 10428 10554 10474
rect 10394 10314 10440 10360
rect 10508 10314 10554 10360
rect 10394 10200 10440 10246
rect 10508 10200 10554 10246
rect 10394 10086 10440 10132
rect 10508 10086 10554 10132
rect 10394 9972 10440 10018
rect 10508 9972 10554 10018
rect 10394 9858 10440 9904
rect 10508 9858 10554 9904
rect 10394 9744 10440 9790
rect 10508 9744 10554 9790
rect 10394 9630 10440 9676
rect 10508 9630 10554 9676
rect 10394 9516 10440 9562
rect 10508 9516 10554 9562
rect 10394 9402 10440 9448
rect 10508 9402 10554 9448
rect 10394 9288 10440 9334
rect 10508 9288 10554 9334
rect 10394 9174 10440 9220
rect 10508 9174 10554 9220
rect 10394 9060 10440 9106
rect 10508 9060 10554 9106
rect 10394 8946 10440 8992
rect 10508 8946 10554 8992
rect 10394 8832 10440 8878
rect 10508 8832 10554 8878
rect 10394 8718 10440 8764
rect 10508 8718 10554 8764
rect 10394 8604 10440 8650
rect 10508 8604 10554 8650
rect 10394 8490 10440 8536
rect 10508 8490 10554 8536
rect 10394 8376 10440 8422
rect 10508 8376 10554 8422
rect 10394 8262 10440 8308
rect 10508 8262 10554 8308
rect 10394 8148 10440 8194
rect 10508 8148 10554 8194
rect 10394 8034 10440 8080
rect 10508 8034 10554 8080
rect 10394 7920 10440 7966
rect 10508 7920 10554 7966
rect 10394 7806 10440 7852
rect 10508 7806 10554 7852
rect 10394 7692 10440 7738
rect 10508 7692 10554 7738
rect 10394 7578 10440 7624
rect 10508 7578 10554 7624
rect 10394 7464 10440 7510
rect 10508 7464 10554 7510
rect 10394 7350 10440 7396
rect 10508 7350 10554 7396
rect 10394 7236 10440 7282
rect 10508 7236 10554 7282
rect 10394 7122 10440 7168
rect 10508 7122 10554 7168
rect 10394 7008 10440 7054
rect 10508 7008 10554 7054
rect 10394 6894 10440 6940
rect 10508 6894 10554 6940
rect 10394 6780 10440 6826
rect 10508 6780 10554 6826
rect 10394 6666 10440 6712
rect 10508 6666 10554 6712
rect 2307 6552 2353 6598
rect 2421 6552 2467 6598
rect 10394 6552 10440 6598
rect 10508 6552 10554 6598
rect 2307 6438 2353 6484
rect 2421 6438 2467 6484
rect 2307 6324 2353 6370
rect 2421 6324 2467 6370
rect 10394 6438 10440 6484
rect 10508 6438 10554 6484
rect 10394 6324 10440 6370
rect 10508 6324 10554 6370
rect 10394 6210 10440 6256
rect 10508 6210 10554 6256
rect 2540 6161 2586 6207
rect 2654 6161 2700 6207
rect 2768 6161 2814 6207
rect 2882 6161 2928 6207
rect 2996 6161 3042 6207
rect 3110 6161 3156 6207
rect 3224 6161 3270 6207
rect 3338 6161 3384 6207
rect 3452 6161 3498 6207
rect 3566 6161 3612 6207
rect 3680 6161 3726 6207
rect 3794 6161 3840 6207
rect 3908 6161 3954 6207
rect 4022 6161 4068 6207
rect 4136 6161 4182 6207
rect 4250 6161 4296 6207
rect 4364 6161 4410 6207
rect 4478 6161 4524 6207
rect 4592 6161 4638 6207
rect 4706 6161 4752 6207
rect 4820 6161 4866 6207
rect 4934 6161 4980 6207
rect 5048 6161 5094 6207
rect 5162 6161 5208 6207
rect 5276 6161 5322 6207
rect 5390 6161 5436 6207
rect 5504 6161 5550 6207
rect 5618 6161 5664 6207
rect 5732 6161 5778 6207
rect 5846 6161 5892 6207
rect 5960 6161 6006 6207
rect 6074 6161 6120 6207
rect 6188 6161 6234 6207
rect 6302 6161 6348 6207
rect 6416 6161 6462 6207
rect 6530 6161 6576 6207
rect 6644 6161 6690 6207
rect 6758 6161 6804 6207
rect 6872 6161 6918 6207
rect 6986 6161 7032 6207
rect 7100 6161 7146 6207
rect 7214 6161 7260 6207
rect 7328 6161 7374 6207
rect 7442 6161 7488 6207
rect 7556 6161 7602 6207
rect 7670 6161 7716 6207
rect 7784 6161 7830 6207
rect 7898 6161 7944 6207
rect 8012 6161 8058 6207
rect 8126 6161 8172 6207
rect 8240 6161 8286 6207
rect 8354 6161 8400 6207
rect 8468 6161 8514 6207
rect 8582 6161 8628 6207
rect 8696 6161 8742 6207
rect 8810 6161 8856 6207
rect 8924 6161 8970 6207
rect 9038 6161 9084 6207
rect 9152 6161 9198 6207
rect 9266 6161 9312 6207
rect 9380 6161 9426 6207
rect 9494 6161 9540 6207
rect 9608 6161 9654 6207
rect 9722 6161 9768 6207
rect 9836 6161 9882 6207
rect 9950 6161 9996 6207
rect 10064 6161 10110 6207
rect 10178 6161 10224 6207
rect 10292 6161 10338 6207
rect 10394 6096 10440 6142
rect 10508 6096 10554 6142
rect 2540 6047 2586 6093
rect 2654 6047 2700 6093
rect 2768 6047 2814 6093
rect 2882 6047 2928 6093
rect 2996 6047 3042 6093
rect 3110 6047 3156 6093
rect 3224 6047 3270 6093
rect 3338 6047 3384 6093
rect 3452 6047 3498 6093
rect 3566 6047 3612 6093
rect 3680 6047 3726 6093
rect 3794 6047 3840 6093
rect 3908 6047 3954 6093
rect 4022 6047 4068 6093
rect 4136 6047 4182 6093
rect 4250 6047 4296 6093
rect 4364 6047 4410 6093
rect 4478 6047 4524 6093
rect 4592 6047 4638 6093
rect 4706 6047 4752 6093
rect 4820 6047 4866 6093
rect 4934 6047 4980 6093
rect 5048 6047 5094 6093
rect 5162 6047 5208 6093
rect 5276 6047 5322 6093
rect 5390 6047 5436 6093
rect 5504 6047 5550 6093
rect 5618 6047 5664 6093
rect 5732 6047 5778 6093
rect 5846 6047 5892 6093
rect 5960 6047 6006 6093
rect 6074 6047 6120 6093
rect 6188 6047 6234 6093
rect 6302 6047 6348 6093
rect 6416 6047 6462 6093
rect 6530 6047 6576 6093
rect 6644 6047 6690 6093
rect 6758 6047 6804 6093
rect 6872 6047 6918 6093
rect 6986 6047 7032 6093
rect 7100 6047 7146 6093
rect 7214 6047 7260 6093
rect 7328 6047 7374 6093
rect 7442 6047 7488 6093
rect 7556 6047 7602 6093
rect 7670 6047 7716 6093
rect 7784 6047 7830 6093
rect 7898 6047 7944 6093
rect 8012 6047 8058 6093
rect 8126 6047 8172 6093
rect 8240 6047 8286 6093
rect 8354 6047 8400 6093
rect 8468 6047 8514 6093
rect 8582 6047 8628 6093
rect 8696 6047 8742 6093
rect 8810 6047 8856 6093
rect 8924 6047 8970 6093
rect 9038 6047 9084 6093
rect 9152 6047 9198 6093
rect 9266 6047 9312 6093
rect 9380 6047 9426 6093
rect 9494 6047 9540 6093
rect 9608 6047 9654 6093
rect 9722 6047 9768 6093
rect 9836 6047 9882 6093
rect 9950 6047 9996 6093
rect 10064 6047 10110 6093
rect 10178 6047 10224 6093
rect 10292 6047 10338 6093
rect 7282 5905 7328 5951
rect 7406 5905 7452 5951
rect 7282 5781 7328 5827
rect 7406 5781 7452 5827
rect 10394 5982 10440 6028
rect 10508 5982 10554 6028
rect 10394 5868 10440 5914
rect 10508 5868 10554 5914
rect 10394 5754 10440 5800
rect 10508 5754 10554 5800
rect 7282 5657 7328 5703
rect 7406 5657 7452 5703
rect 10394 5640 10440 5686
rect 10508 5640 10554 5686
rect 7282 5533 7328 5579
rect 7406 5533 7452 5579
rect 7282 5409 7328 5455
rect 7406 5409 7452 5455
rect 7282 5285 7328 5331
rect 7406 5285 7452 5331
rect 7282 5161 7328 5207
rect 7406 5161 7452 5207
rect 7282 5037 7328 5083
rect 7406 5037 7452 5083
rect 7282 4913 7328 4959
rect 7406 4913 7452 4959
rect 7282 4789 7328 4835
rect 7406 4789 7452 4835
rect 7282 4665 7328 4711
rect 7406 4665 7452 4711
rect 7282 4541 7328 4587
rect 7406 4541 7452 4587
rect 7282 4417 7328 4463
rect 7406 4417 7452 4463
rect 7282 4293 7328 4339
rect 7406 4293 7452 4339
rect 7282 4169 7328 4215
rect 7406 4169 7452 4215
rect 7282 4045 7328 4091
rect 7406 4045 7452 4091
rect 7282 3921 7328 3967
rect 7406 3921 7452 3967
rect 7282 3797 7328 3843
rect 7406 3797 7452 3843
rect 7282 3673 7328 3719
rect 7406 3673 7452 3719
rect 7282 3549 7328 3595
rect 7406 3549 7452 3595
rect 7282 3425 7328 3471
rect 7406 3425 7452 3471
rect 7282 3301 7328 3347
rect 7406 3301 7452 3347
rect 7282 3177 7328 3223
rect 7406 3177 7452 3223
rect 7282 3053 7328 3099
rect 7406 3053 7452 3099
rect 7282 2929 7328 2975
rect 7406 2929 7452 2975
rect 7282 2805 7328 2851
rect 7406 2805 7452 2851
rect 7282 2681 7328 2727
rect 7406 2681 7452 2727
rect 7282 2557 7328 2603
rect 7406 2557 7452 2603
rect 7282 2433 7328 2479
rect 7406 2433 7452 2479
rect 7282 2309 7328 2355
rect 7406 2309 7452 2355
rect 7282 2185 7328 2231
rect 7406 2185 7452 2231
rect 7282 2061 7328 2107
rect 7406 2061 7452 2107
rect 7282 1937 7328 1983
rect 7406 1937 7452 1983
rect 7282 1813 7328 1859
rect 7406 1813 7452 1859
rect 7282 1689 7328 1735
rect 7406 1689 7452 1735
rect 7282 1565 7328 1611
rect 7406 1565 7452 1611
rect 7282 1441 7328 1487
rect 7406 1441 7452 1487
rect 7282 1317 7328 1363
rect 7406 1317 7452 1363
rect 7282 1193 7328 1239
rect 7406 1193 7452 1239
rect 7282 1069 7328 1115
rect 7406 1069 7452 1115
rect 7282 945 7328 991
rect 7406 945 7452 991
rect 7282 821 7328 867
rect 7406 821 7452 867
rect 7282 697 7328 743
rect 7406 697 7452 743
rect 10394 5526 10440 5572
rect 10508 5526 10554 5572
rect 10394 5412 10440 5458
rect 10508 5412 10554 5458
rect 10394 5298 10440 5344
rect 10508 5298 10554 5344
rect 10394 5184 10440 5230
rect 10508 5184 10554 5230
rect 10394 5070 10440 5116
rect 10508 5070 10554 5116
rect 10394 4956 10440 5002
rect 10508 4956 10554 5002
rect 10394 4842 10440 4888
rect 10508 4842 10554 4888
rect 10394 4728 10440 4774
rect 10508 4728 10554 4774
rect 10394 4614 10440 4660
rect 10508 4614 10554 4660
rect 10394 4500 10440 4546
rect 10508 4500 10554 4546
rect 10394 4386 10440 4432
rect 10508 4386 10554 4432
rect 10394 4272 10440 4318
rect 10508 4272 10554 4318
rect 10394 4158 10440 4204
rect 10508 4158 10554 4204
rect 10394 4044 10440 4090
rect 10508 4044 10554 4090
rect 10394 3930 10440 3976
rect 10508 3930 10554 3976
rect 10394 3816 10440 3862
rect 10508 3816 10554 3862
rect 10394 3702 10440 3748
rect 10508 3702 10554 3748
rect 10394 3588 10440 3634
rect 10508 3588 10554 3634
rect 10394 3474 10440 3520
rect 10508 3474 10554 3520
rect 10394 3360 10440 3406
rect 10508 3360 10554 3406
rect 10394 3246 10440 3292
rect 10508 3246 10554 3292
rect 10394 3132 10440 3178
rect 10508 3132 10554 3178
rect 10394 3018 10440 3064
rect 10508 3018 10554 3064
rect 10394 2904 10440 2950
rect 10508 2904 10554 2950
rect 10394 2790 10440 2836
rect 10508 2790 10554 2836
rect 10394 2676 10440 2722
rect 10508 2676 10554 2722
rect 10394 2562 10440 2608
rect 10508 2562 10554 2608
rect 10394 2448 10440 2494
rect 10508 2448 10554 2494
rect 10394 2334 10440 2380
rect 10508 2334 10554 2380
rect 10394 2220 10440 2266
rect 10508 2220 10554 2266
rect 10394 2106 10440 2152
rect 10508 2106 10554 2152
rect 10394 1992 10440 2038
rect 10508 1992 10554 2038
rect 10394 1878 10440 1924
rect 10508 1878 10554 1924
rect 10394 1764 10440 1810
rect 10508 1764 10554 1810
rect 10394 1650 10440 1696
rect 10508 1650 10554 1696
rect 10394 1536 10440 1582
rect 10508 1536 10554 1582
rect 10394 1422 10440 1468
rect 10508 1422 10554 1468
rect 10394 1308 10440 1354
rect 10508 1308 10554 1354
rect 10394 1194 10440 1240
rect 10508 1194 10554 1240
rect 10394 1080 10440 1126
rect 10508 1080 10554 1126
rect 10394 966 10440 1012
rect 10508 966 10554 1012
rect 10394 852 10440 898
rect 10508 852 10554 898
rect 10394 738 10440 784
rect 10508 738 10554 784
rect 10394 624 10440 670
rect 10508 624 10554 670
rect 7282 573 7328 619
rect 7406 573 7452 619
rect 7282 449 7328 495
rect 7406 449 7452 495
rect 7282 325 7328 371
rect 7406 325 7452 371
rect 7282 201 7328 247
rect 7406 201 7452 247
rect 10394 510 10440 556
rect 10508 510 10554 556
rect 10394 396 10440 442
rect 10508 396 10554 442
rect 10394 282 10440 328
rect 10508 282 10554 328
rect 7612 168 7658 214
rect 7726 168 7772 214
rect 7840 168 7886 214
rect 7954 168 8000 214
rect 8068 168 8114 214
rect 8182 168 8228 214
rect 8296 168 8342 214
rect 8410 168 8456 214
rect 8524 168 8570 214
rect 8638 168 8684 214
rect 8752 168 8798 214
rect 8866 168 8912 214
rect 8980 168 9026 214
rect 9094 168 9140 214
rect 9208 168 9254 214
rect 9322 168 9368 214
rect 9436 168 9482 214
rect 9550 168 9596 214
rect 9664 168 9710 214
rect 9778 168 9824 214
rect 9892 168 9938 214
rect 10006 168 10052 214
rect 10120 168 10166 214
rect 10234 168 10280 214
rect 10394 168 10440 214
rect 10508 168 10554 214
rect 7282 77 7328 123
rect 7406 77 7452 123
rect 7612 54 7658 100
rect 7726 54 7772 100
rect 7840 54 7886 100
rect 7954 54 8000 100
rect 8068 54 8114 100
rect 8182 54 8228 100
rect 8296 54 8342 100
rect 8410 54 8456 100
rect 8524 54 8570 100
rect 8638 54 8684 100
rect 8752 54 8798 100
rect 8866 54 8912 100
rect 8980 54 9026 100
rect 9094 54 9140 100
rect 9208 54 9254 100
rect 9322 54 9368 100
rect 9436 54 9482 100
rect 9550 54 9596 100
rect 9664 54 9710 100
rect 9778 54 9824 100
rect 9892 54 9938 100
rect 10006 54 10052 100
rect 10120 54 10166 100
rect 10234 54 10280 100
rect 10394 54 10440 100
rect 10508 54 10554 100
<< polysilicon >>
rect 3083 11712 5083 11725
rect 3083 11666 3136 11712
rect 5030 11666 5083 11712
rect 3083 11633 5083 11666
rect 5519 11712 7519 11725
rect 5519 11666 5572 11712
rect 7466 11666 7519 11712
rect 5519 11633 7519 11666
rect 7955 11712 9955 11725
rect 7955 11666 8008 11712
rect 9902 11666 9955 11712
rect 7955 11633 9955 11666
rect 3083 6600 5083 6633
rect 3083 6554 3136 6600
rect 5030 6554 5083 6600
rect 3083 6541 5083 6554
rect 5519 6600 7519 6633
rect 5519 6554 5572 6600
rect 7466 6554 7519 6600
rect 5519 6541 7519 6554
rect 7955 6600 9955 6633
rect 7955 6554 8008 6600
rect 9902 6554 9955 6600
rect 7955 6541 9955 6554
rect 7955 5700 9955 5713
rect 7955 5654 8008 5700
rect 9902 5654 9955 5700
rect 7955 5621 9955 5654
rect 7955 588 9955 621
rect 7955 542 8008 588
rect 9902 542 9955 588
rect 7955 529 9955 542
<< polycontact >>
rect 3136 11666 5030 11712
rect 5572 11666 7466 11712
rect 8008 11666 9902 11712
rect 3136 6554 5030 6600
rect 5572 6554 7466 6600
rect 8008 6554 9902 6600
rect 8008 5654 9902 5700
rect 8008 542 9902 588
<< metal1 >>
rect 2296 12298 10565 12310
rect 2296 12252 2307 12298
rect 2353 12252 2421 12298
rect 2467 12252 2575 12298
rect 2621 12252 2689 12298
rect 2735 12252 2803 12298
rect 2849 12252 2917 12298
rect 2963 12252 3031 12298
rect 3077 12252 3145 12298
rect 3191 12252 3259 12298
rect 3305 12252 3373 12298
rect 3419 12252 3487 12298
rect 3533 12252 3601 12298
rect 3647 12252 3715 12298
rect 3761 12252 3829 12298
rect 3875 12252 3943 12298
rect 3989 12252 4057 12298
rect 4103 12252 4171 12298
rect 4217 12252 4285 12298
rect 4331 12252 4399 12298
rect 4445 12252 4513 12298
rect 4559 12252 4627 12298
rect 4673 12252 4741 12298
rect 4787 12252 4855 12298
rect 4901 12252 4969 12298
rect 5015 12252 5083 12298
rect 5129 12252 5197 12298
rect 5243 12252 5311 12298
rect 5357 12252 5425 12298
rect 5471 12252 5539 12298
rect 5585 12252 5653 12298
rect 5699 12252 5767 12298
rect 5813 12252 5881 12298
rect 5927 12252 5995 12298
rect 6041 12252 6109 12298
rect 6155 12252 6223 12298
rect 6269 12252 6337 12298
rect 6383 12252 6451 12298
rect 6497 12252 6565 12298
rect 6611 12252 6679 12298
rect 6725 12252 6793 12298
rect 6839 12252 6907 12298
rect 6953 12252 7021 12298
rect 7067 12252 7135 12298
rect 7181 12252 7249 12298
rect 7295 12252 7363 12298
rect 7409 12252 7477 12298
rect 7523 12252 7591 12298
rect 7637 12252 7705 12298
rect 7751 12252 7819 12298
rect 7865 12252 7933 12298
rect 7979 12252 8047 12298
rect 8093 12252 8161 12298
rect 8207 12252 8275 12298
rect 8321 12252 8389 12298
rect 8435 12252 8503 12298
rect 8549 12252 8617 12298
rect 8663 12252 8731 12298
rect 8777 12252 8845 12298
rect 8891 12252 8959 12298
rect 9005 12252 9073 12298
rect 9119 12252 9187 12298
rect 9233 12252 9301 12298
rect 9347 12252 9415 12298
rect 9461 12252 9529 12298
rect 9575 12252 9643 12298
rect 9689 12252 9757 12298
rect 9803 12252 9871 12298
rect 9917 12252 9985 12298
rect 10031 12252 10099 12298
rect 10145 12252 10213 12298
rect 10259 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10565 12298
rect 2296 12184 10565 12252
rect 2296 12138 2307 12184
rect 2353 12138 2421 12184
rect 2467 12138 2575 12184
rect 2621 12138 2689 12184
rect 2735 12138 2803 12184
rect 2849 12138 2917 12184
rect 2963 12138 3031 12184
rect 3077 12138 3145 12184
rect 3191 12138 3259 12184
rect 3305 12138 3373 12184
rect 3419 12138 3487 12184
rect 3533 12138 3601 12184
rect 3647 12138 3715 12184
rect 3761 12138 3829 12184
rect 3875 12138 3943 12184
rect 3989 12138 4057 12184
rect 4103 12138 4171 12184
rect 4217 12138 4285 12184
rect 4331 12138 4399 12184
rect 4445 12138 4513 12184
rect 4559 12138 4627 12184
rect 4673 12138 4741 12184
rect 4787 12138 4855 12184
rect 4901 12138 4969 12184
rect 5015 12138 5083 12184
rect 5129 12138 5197 12184
rect 5243 12138 5311 12184
rect 5357 12138 5425 12184
rect 5471 12138 5539 12184
rect 5585 12138 5653 12184
rect 5699 12138 5767 12184
rect 5813 12138 5881 12184
rect 5927 12138 5995 12184
rect 6041 12138 6109 12184
rect 6155 12138 6223 12184
rect 6269 12138 6337 12184
rect 6383 12138 6451 12184
rect 6497 12138 6565 12184
rect 6611 12138 6679 12184
rect 6725 12138 6793 12184
rect 6839 12138 6907 12184
rect 6953 12138 7021 12184
rect 7067 12138 7135 12184
rect 7181 12138 7249 12184
rect 7295 12138 7363 12184
rect 7409 12138 7477 12184
rect 7523 12138 7591 12184
rect 7637 12138 7705 12184
rect 7751 12138 7819 12184
rect 7865 12138 7933 12184
rect 7979 12138 8047 12184
rect 8093 12138 8161 12184
rect 8207 12138 8275 12184
rect 8321 12138 8389 12184
rect 8435 12138 8503 12184
rect 8549 12138 8617 12184
rect 8663 12138 8731 12184
rect 8777 12138 8845 12184
rect 8891 12138 8959 12184
rect 9005 12138 9073 12184
rect 9119 12138 9187 12184
rect 9233 12138 9301 12184
rect 9347 12138 9415 12184
rect 9461 12138 9529 12184
rect 9575 12138 9643 12184
rect 9689 12138 9757 12184
rect 9803 12138 9871 12184
rect 9917 12138 9985 12184
rect 10031 12138 10099 12184
rect 10145 12138 10213 12184
rect 10259 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10565 12184
rect 2296 12126 10565 12138
rect 2296 12070 2478 12126
rect 2296 12024 2307 12070
rect 2353 12024 2421 12070
rect 2467 12024 2478 12070
rect 2296 11633 2478 12024
rect 10383 12070 10565 12126
rect 10383 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10565 12070
rect 10383 11956 10565 12024
rect 10383 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10565 11956
rect 3125 11723 9913 11855
rect 3125 11712 5041 11723
rect 3125 11666 3136 11712
rect 5030 11666 5041 11712
rect 3125 11655 5041 11666
rect 5561 11712 7477 11723
rect 5561 11666 5572 11712
rect 7466 11666 7477 11712
rect 5561 11655 7477 11666
rect 7997 11712 9913 11723
rect 7997 11666 8008 11712
rect 9902 11666 9913 11712
rect 7997 11655 9913 11666
rect 10383 11842 10565 11910
rect 10383 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10565 11842
rect 10383 11728 10565 11796
rect 10383 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10565 11728
rect 2296 11596 3065 11633
rect 2296 11500 3008 11596
rect 2296 11454 2307 11500
rect 2353 11454 2421 11500
rect 2467 11454 3008 11500
rect 2296 11386 3008 11454
rect 2296 11340 2307 11386
rect 2353 11340 2421 11386
rect 2467 11340 3008 11386
rect 2296 11272 3008 11340
rect 2296 11226 2307 11272
rect 2353 11226 2421 11272
rect 2467 11226 3008 11272
rect 2296 11158 3008 11226
rect 2296 11112 2307 11158
rect 2353 11112 2421 11158
rect 2467 11112 3008 11158
rect 2296 11044 3008 11112
rect 2296 10998 2307 11044
rect 2353 10998 2421 11044
rect 2467 10998 3008 11044
rect 2296 10930 3008 10998
rect 2296 10884 2307 10930
rect 2353 10884 2421 10930
rect 2467 10884 3008 10930
rect 2296 10816 3008 10884
rect 2296 10770 2307 10816
rect 2353 10770 2421 10816
rect 2467 10770 3008 10816
rect 2296 10702 3008 10770
rect 2296 10656 2307 10702
rect 2353 10656 2421 10702
rect 2467 10656 3008 10702
rect 2296 10588 3008 10656
rect 2296 10542 2307 10588
rect 2353 10542 2421 10588
rect 2467 10542 3008 10588
rect 2296 10474 3008 10542
rect 2296 10428 2307 10474
rect 2353 10428 2421 10474
rect 2467 10428 3008 10474
rect 2296 10360 3008 10428
rect 2296 10314 2307 10360
rect 2353 10314 2421 10360
rect 2467 10314 3008 10360
rect 2296 10246 3008 10314
rect 2296 10200 2307 10246
rect 2353 10200 2421 10246
rect 2467 10200 3008 10246
rect 2296 10132 3008 10200
rect 2296 10086 2307 10132
rect 2353 10086 2421 10132
rect 2467 10086 3008 10132
rect 2296 10018 3008 10086
rect 2296 9972 2307 10018
rect 2353 9972 2421 10018
rect 2467 9972 3008 10018
rect 2296 9904 3008 9972
rect 2296 9858 2307 9904
rect 2353 9858 2421 9904
rect 2467 9858 3008 9904
rect 2296 9790 3008 9858
rect 2296 9744 2307 9790
rect 2353 9744 2421 9790
rect 2467 9744 3008 9790
rect 2296 9676 3008 9744
rect 2296 9630 2307 9676
rect 2353 9630 2421 9676
rect 2467 9630 3008 9676
rect 2296 9562 3008 9630
rect 2296 9516 2307 9562
rect 2353 9516 2421 9562
rect 2467 9516 3008 9562
rect 2296 9448 3008 9516
rect 2296 9402 2307 9448
rect 2353 9402 2421 9448
rect 2467 9402 3008 9448
rect 2296 9334 3008 9402
rect 2296 9288 2307 9334
rect 2353 9288 2421 9334
rect 2467 9288 3008 9334
rect 2296 9220 3008 9288
rect 2296 9174 2307 9220
rect 2353 9174 2421 9220
rect 2467 9174 3008 9220
rect 2296 9106 3008 9174
rect 2296 9060 2307 9106
rect 2353 9060 2421 9106
rect 2467 9060 3008 9106
rect 2296 8992 3008 9060
rect 2296 8946 2307 8992
rect 2353 8946 2421 8992
rect 2467 8946 3008 8992
rect 2296 8878 3008 8946
rect 2296 8832 2307 8878
rect 2353 8832 2421 8878
rect 2467 8832 3008 8878
rect 2296 8764 3008 8832
rect 2296 8718 2307 8764
rect 2353 8718 2421 8764
rect 2467 8718 3008 8764
rect 2296 8650 3008 8718
rect 2296 8604 2307 8650
rect 2353 8604 2421 8650
rect 2467 8604 3008 8650
rect 2296 8536 3008 8604
rect 2296 8490 2307 8536
rect 2353 8490 2421 8536
rect 2467 8490 3008 8536
rect 2296 8422 3008 8490
rect 2296 8376 2307 8422
rect 2353 8376 2421 8422
rect 2467 8376 3008 8422
rect 2296 8308 3008 8376
rect 2296 8262 2307 8308
rect 2353 8262 2421 8308
rect 2467 8262 3008 8308
rect 2296 8194 3008 8262
rect 2296 8148 2307 8194
rect 2353 8148 2421 8194
rect 2467 8148 3008 8194
rect 2296 8080 3008 8148
rect 2296 8034 2307 8080
rect 2353 8034 2421 8080
rect 2467 8034 3008 8080
rect 2296 7966 3008 8034
rect 2296 7920 2307 7966
rect 2353 7920 2421 7966
rect 2467 7920 3008 7966
rect 2296 7852 3008 7920
rect 2296 7806 2307 7852
rect 2353 7806 2421 7852
rect 2467 7806 3008 7852
rect 2296 7738 3008 7806
rect 2296 7692 2307 7738
rect 2353 7692 2421 7738
rect 2467 7692 3008 7738
rect 2296 7624 3008 7692
rect 2296 7578 2307 7624
rect 2353 7578 2421 7624
rect 2467 7578 3008 7624
rect 2296 7510 3008 7578
rect 2296 7464 2307 7510
rect 2353 7464 2421 7510
rect 2467 7464 3008 7510
rect 2296 7396 3008 7464
rect 2296 7350 2307 7396
rect 2353 7350 2421 7396
rect 2467 7350 3008 7396
rect 2296 7282 3008 7350
rect 2296 7236 2307 7282
rect 2353 7236 2421 7282
rect 2467 7236 3008 7282
rect 2296 7168 3008 7236
rect 2296 7122 2307 7168
rect 2353 7122 2421 7168
rect 2467 7122 3008 7168
rect 2296 7054 3008 7122
rect 2296 7008 2307 7054
rect 2353 7008 2421 7054
rect 2467 7008 3008 7054
rect 2296 6940 3008 7008
rect 2296 6894 2307 6940
rect 2353 6894 2421 6940
rect 2467 6894 3008 6940
rect 2296 6826 3008 6894
rect 2296 6780 2307 6826
rect 2353 6780 2421 6826
rect 2467 6780 3008 6826
rect 2296 6712 3008 6780
rect 2296 6666 2307 6712
rect 2353 6666 2421 6712
rect 2467 6670 3008 6712
rect 3054 6670 3065 11596
rect 2467 6666 3065 6670
rect 2296 6598 3065 6666
rect 3583 6611 4583 11655
rect 5101 11596 5501 11633
rect 5101 6670 5112 11596
rect 5158 6670 5444 11596
rect 5490 6670 5501 11596
rect 2296 6552 2307 6598
rect 2353 6552 2421 6598
rect 2467 6552 3065 6598
rect 2296 6484 3065 6552
rect 3125 6600 5041 6611
rect 3125 6554 3136 6600
rect 5030 6554 5041 6600
rect 3125 6543 5041 6554
rect 2296 6438 2307 6484
rect 2353 6438 2421 6484
rect 2467 6483 3065 6484
rect 5101 6483 5501 6670
rect 6019 6611 7019 11655
rect 7537 11596 7937 11633
rect 7537 6670 7548 11596
rect 7594 6670 7880 11596
rect 7926 6670 7937 11596
rect 5561 6600 7477 6611
rect 5561 6554 5572 6600
rect 7466 6554 7477 6600
rect 5561 6543 7477 6554
rect 7537 6483 7937 6670
rect 8455 6611 9455 11655
rect 10383 11633 10565 11682
rect 9973 11614 10565 11633
rect 9973 11596 10394 11614
rect 9973 6670 9984 11596
rect 10030 11568 10394 11596
rect 10440 11568 10508 11614
rect 10554 11568 10565 11614
rect 10030 11500 10565 11568
rect 10030 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10565 11500
rect 10030 11386 10565 11454
rect 10030 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10565 11386
rect 10030 11272 10565 11340
rect 10030 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10565 11272
rect 10030 11158 10565 11226
rect 10030 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10565 11158
rect 10030 11044 10565 11112
rect 10030 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10565 11044
rect 10030 10930 10565 10998
rect 10030 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10565 10930
rect 10030 10816 10565 10884
rect 10030 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10565 10816
rect 10030 10702 10565 10770
rect 10030 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10565 10702
rect 10030 10588 10565 10656
rect 10030 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10565 10588
rect 10030 10474 10565 10542
rect 10030 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10565 10474
rect 10030 10360 10565 10428
rect 10030 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10565 10360
rect 10030 10246 10565 10314
rect 10030 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10565 10246
rect 10030 10132 10565 10200
rect 10030 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10565 10132
rect 10030 10018 10565 10086
rect 10030 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10565 10018
rect 10030 9904 10565 9972
rect 10030 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10565 9904
rect 10030 9790 10565 9858
rect 10030 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10565 9790
rect 10030 9676 10565 9744
rect 10030 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10565 9676
rect 10030 9562 10565 9630
rect 10030 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10565 9562
rect 10030 9448 10565 9516
rect 10030 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10565 9448
rect 10030 9334 10565 9402
rect 10030 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10565 9334
rect 10030 9220 10565 9288
rect 10030 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10565 9220
rect 10030 9106 10565 9174
rect 10030 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10565 9106
rect 10030 8992 10565 9060
rect 10030 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10565 8992
rect 10030 8878 10565 8946
rect 10030 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10565 8878
rect 10030 8764 10565 8832
rect 10030 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10565 8764
rect 10030 8650 10565 8718
rect 10030 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10565 8650
rect 10030 8536 10565 8604
rect 10030 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10565 8536
rect 10030 8422 10565 8490
rect 10030 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10565 8422
rect 10030 8308 10565 8376
rect 10030 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10565 8308
rect 10030 8194 10565 8262
rect 10030 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10565 8194
rect 10030 8080 10565 8148
rect 10030 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10565 8080
rect 10030 7966 10565 8034
rect 10030 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10565 7966
rect 10030 7852 10565 7920
rect 10030 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10565 7852
rect 10030 7738 10565 7806
rect 10030 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10565 7738
rect 10030 7624 10565 7692
rect 10030 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10565 7624
rect 10030 7510 10565 7578
rect 10030 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10565 7510
rect 10030 7396 10565 7464
rect 10030 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10565 7396
rect 10030 7282 10565 7350
rect 10030 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10565 7282
rect 10030 7168 10565 7236
rect 10030 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10565 7168
rect 10030 7054 10565 7122
rect 10030 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10565 7054
rect 10030 6940 10565 7008
rect 10030 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10565 6940
rect 10030 6826 10565 6894
rect 10030 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10565 6826
rect 10030 6712 10565 6780
rect 10030 6670 10394 6712
rect 9973 6666 10394 6670
rect 10440 6666 10508 6712
rect 10554 6666 10565 6712
rect 7997 6600 9913 6611
rect 7997 6554 8008 6600
rect 9902 6554 9913 6600
rect 7997 6543 9913 6554
rect 9973 6598 10565 6666
rect 9973 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10565 6598
rect 9973 6484 10565 6552
rect 9973 6483 10394 6484
rect 2467 6438 10394 6483
rect 10440 6438 10508 6484
rect 10554 6438 10565 6484
rect 2296 6370 10565 6438
rect 2296 6324 2307 6370
rect 2353 6324 2421 6370
rect 2467 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10565 6370
rect 2296 6256 10565 6324
rect 2296 6210 10394 6256
rect 10440 6210 10508 6256
rect 10554 6210 10565 6256
rect 2296 6207 10565 6210
rect 2296 6161 2540 6207
rect 2586 6161 2654 6207
rect 2700 6161 2768 6207
rect 2814 6161 2882 6207
rect 2928 6161 2996 6207
rect 3042 6161 3110 6207
rect 3156 6161 3224 6207
rect 3270 6161 3338 6207
rect 3384 6161 3452 6207
rect 3498 6161 3566 6207
rect 3612 6161 3680 6207
rect 3726 6161 3794 6207
rect 3840 6161 3908 6207
rect 3954 6161 4022 6207
rect 4068 6161 4136 6207
rect 4182 6161 4250 6207
rect 4296 6161 4364 6207
rect 4410 6161 4478 6207
rect 4524 6161 4592 6207
rect 4638 6161 4706 6207
rect 4752 6161 4820 6207
rect 4866 6161 4934 6207
rect 4980 6161 5048 6207
rect 5094 6161 5162 6207
rect 5208 6161 5276 6207
rect 5322 6161 5390 6207
rect 5436 6161 5504 6207
rect 5550 6161 5618 6207
rect 5664 6161 5732 6207
rect 5778 6161 5846 6207
rect 5892 6161 5960 6207
rect 6006 6161 6074 6207
rect 6120 6161 6188 6207
rect 6234 6161 6302 6207
rect 6348 6161 6416 6207
rect 6462 6161 6530 6207
rect 6576 6161 6644 6207
rect 6690 6161 6758 6207
rect 6804 6161 6872 6207
rect 6918 6161 6986 6207
rect 7032 6161 7100 6207
rect 7146 6161 7214 6207
rect 7260 6161 7328 6207
rect 7374 6161 7442 6207
rect 7488 6161 7556 6207
rect 7602 6161 7670 6207
rect 7716 6161 7784 6207
rect 7830 6161 7898 6207
rect 7944 6161 8012 6207
rect 8058 6161 8126 6207
rect 8172 6161 8240 6207
rect 8286 6161 8354 6207
rect 8400 6161 8468 6207
rect 8514 6161 8582 6207
rect 8628 6161 8696 6207
rect 8742 6161 8810 6207
rect 8856 6161 8924 6207
rect 8970 6161 9038 6207
rect 9084 6161 9152 6207
rect 9198 6161 9266 6207
rect 9312 6161 9380 6207
rect 9426 6161 9494 6207
rect 9540 6161 9608 6207
rect 9654 6161 9722 6207
rect 9768 6161 9836 6207
rect 9882 6161 9950 6207
rect 9996 6161 10064 6207
rect 10110 6161 10178 6207
rect 10224 6161 10292 6207
rect 10338 6161 10565 6207
rect 2296 6142 10565 6161
rect 2296 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10565 6142
rect 2296 6093 10565 6096
rect 2296 6047 2540 6093
rect 2586 6047 2654 6093
rect 2700 6047 2768 6093
rect 2814 6047 2882 6093
rect 2928 6047 2996 6093
rect 3042 6047 3110 6093
rect 3156 6047 3224 6093
rect 3270 6047 3338 6093
rect 3384 6047 3452 6093
rect 3498 6047 3566 6093
rect 3612 6047 3680 6093
rect 3726 6047 3794 6093
rect 3840 6047 3908 6093
rect 3954 6047 4022 6093
rect 4068 6047 4136 6093
rect 4182 6047 4250 6093
rect 4296 6047 4364 6093
rect 4410 6047 4478 6093
rect 4524 6047 4592 6093
rect 4638 6047 4706 6093
rect 4752 6047 4820 6093
rect 4866 6047 4934 6093
rect 4980 6047 5048 6093
rect 5094 6047 5162 6093
rect 5208 6047 5276 6093
rect 5322 6047 5390 6093
rect 5436 6047 5504 6093
rect 5550 6047 5618 6093
rect 5664 6047 5732 6093
rect 5778 6047 5846 6093
rect 5892 6047 5960 6093
rect 6006 6047 6074 6093
rect 6120 6047 6188 6093
rect 6234 6047 6302 6093
rect 6348 6047 6416 6093
rect 6462 6047 6530 6093
rect 6576 6047 6644 6093
rect 6690 6047 6758 6093
rect 6804 6047 6872 6093
rect 6918 6047 6986 6093
rect 7032 6047 7100 6093
rect 7146 6047 7214 6093
rect 7260 6047 7328 6093
rect 7374 6047 7442 6093
rect 7488 6047 7556 6093
rect 7602 6047 7670 6093
rect 7716 6047 7784 6093
rect 7830 6047 7898 6093
rect 7944 6047 8012 6093
rect 8058 6047 8126 6093
rect 8172 6047 8240 6093
rect 8286 6047 8354 6093
rect 8400 6047 8468 6093
rect 8514 6047 8582 6093
rect 8628 6047 8696 6093
rect 8742 6047 8810 6093
rect 8856 6047 8924 6093
rect 8970 6047 9038 6093
rect 9084 6047 9152 6093
rect 9198 6047 9266 6093
rect 9312 6047 9380 6093
rect 9426 6047 9494 6093
rect 9540 6047 9608 6093
rect 9654 6047 9722 6093
rect 9768 6047 9836 6093
rect 9882 6047 9950 6093
rect 9996 6047 10064 6093
rect 10110 6047 10178 6093
rect 10224 6047 10292 6093
rect 10338 6047 10565 6093
rect 2296 6028 10565 6047
rect 2296 5982 10394 6028
rect 10440 5982 10508 6028
rect 10554 5982 10565 6028
rect 2296 5951 10565 5982
rect 2296 5905 7282 5951
rect 7328 5905 7406 5951
rect 7452 5914 10565 5951
rect 7452 5905 10394 5914
rect 2296 5868 10394 5905
rect 10440 5868 10508 5914
rect 10554 5868 10565 5914
rect 2296 5827 10565 5868
rect 2296 5781 7282 5827
rect 7328 5781 7406 5827
rect 7452 5800 10565 5827
rect 7452 5781 10394 5800
rect 2296 5771 10394 5781
rect 7271 5703 7937 5771
rect 9973 5754 10394 5771
rect 10440 5754 10508 5800
rect 10554 5754 10565 5800
rect 7271 5657 7282 5703
rect 7328 5657 7406 5703
rect 7452 5657 7937 5703
rect 7271 5584 7937 5657
rect 7997 5700 9913 5711
rect 7997 5654 8008 5700
rect 9902 5654 9913 5700
rect 7997 5643 9913 5654
rect 9973 5686 10565 5754
rect 7271 5579 7880 5584
rect 7271 5533 7282 5579
rect 7328 5533 7406 5579
rect 7452 5533 7880 5579
rect 7271 5455 7880 5533
rect 7271 5409 7282 5455
rect 7328 5409 7406 5455
rect 7452 5409 7880 5455
rect 7271 5331 7880 5409
rect 7271 5285 7282 5331
rect 7328 5285 7406 5331
rect 7452 5285 7880 5331
rect 7271 5207 7880 5285
rect 7271 5161 7282 5207
rect 7328 5161 7406 5207
rect 7452 5161 7880 5207
rect 7271 5083 7880 5161
rect 7271 5037 7282 5083
rect 7328 5037 7406 5083
rect 7452 5037 7880 5083
rect 7271 4959 7880 5037
rect 7271 4913 7282 4959
rect 7328 4913 7406 4959
rect 7452 4913 7880 4959
rect 7271 4835 7880 4913
rect 7271 4789 7282 4835
rect 7328 4789 7406 4835
rect 7452 4789 7880 4835
rect 7271 4711 7880 4789
rect 7271 4665 7282 4711
rect 7328 4665 7406 4711
rect 7452 4665 7880 4711
rect 7271 4587 7880 4665
rect 7271 4541 7282 4587
rect 7328 4541 7406 4587
rect 7452 4541 7880 4587
rect 7271 4463 7880 4541
rect 7271 4417 7282 4463
rect 7328 4417 7406 4463
rect 7452 4417 7880 4463
rect 7271 4339 7880 4417
rect 7271 4293 7282 4339
rect 7328 4293 7406 4339
rect 7452 4293 7880 4339
rect 7271 4215 7880 4293
rect 7271 4169 7282 4215
rect 7328 4169 7406 4215
rect 7452 4169 7880 4215
rect 7271 4091 7880 4169
rect 7271 4045 7282 4091
rect 7328 4045 7406 4091
rect 7452 4045 7880 4091
rect 7271 3967 7880 4045
rect 7271 3921 7282 3967
rect 7328 3921 7406 3967
rect 7452 3921 7880 3967
rect 7271 3843 7880 3921
rect 7271 3797 7282 3843
rect 7328 3797 7406 3843
rect 7452 3797 7880 3843
rect 7271 3719 7880 3797
rect 7271 3673 7282 3719
rect 7328 3673 7406 3719
rect 7452 3673 7880 3719
rect 7271 3595 7880 3673
rect 7271 3549 7282 3595
rect 7328 3549 7406 3595
rect 7452 3549 7880 3595
rect 7271 3471 7880 3549
rect 7271 3425 7282 3471
rect 7328 3425 7406 3471
rect 7452 3425 7880 3471
rect 7271 3347 7880 3425
rect 7271 3301 7282 3347
rect 7328 3301 7406 3347
rect 7452 3301 7880 3347
rect 7271 3223 7880 3301
rect 7271 3177 7282 3223
rect 7328 3177 7406 3223
rect 7452 3177 7880 3223
rect 7271 3099 7880 3177
rect 7271 3053 7282 3099
rect 7328 3053 7406 3099
rect 7452 3053 7880 3099
rect 7271 2975 7880 3053
rect 7271 2929 7282 2975
rect 7328 2929 7406 2975
rect 7452 2929 7880 2975
rect 7271 2851 7880 2929
rect 7271 2805 7282 2851
rect 7328 2805 7406 2851
rect 7452 2805 7880 2851
rect 7271 2727 7880 2805
rect 7271 2681 7282 2727
rect 7328 2681 7406 2727
rect 7452 2681 7880 2727
rect 7271 2603 7880 2681
rect 7271 2557 7282 2603
rect 7328 2557 7406 2603
rect 7452 2557 7880 2603
rect 7271 2479 7880 2557
rect 7271 2433 7282 2479
rect 7328 2433 7406 2479
rect 7452 2433 7880 2479
rect 7271 2355 7880 2433
rect 7271 2309 7282 2355
rect 7328 2309 7406 2355
rect 7452 2309 7880 2355
rect 7271 2231 7880 2309
rect 7271 2185 7282 2231
rect 7328 2185 7406 2231
rect 7452 2185 7880 2231
rect 7271 2107 7880 2185
rect 7271 2061 7282 2107
rect 7328 2061 7406 2107
rect 7452 2061 7880 2107
rect 7271 1983 7880 2061
rect 7271 1937 7282 1983
rect 7328 1937 7406 1983
rect 7452 1937 7880 1983
rect 7271 1859 7880 1937
rect 7271 1813 7282 1859
rect 7328 1813 7406 1859
rect 7452 1813 7880 1859
rect 7271 1735 7880 1813
rect 7271 1689 7282 1735
rect 7328 1689 7406 1735
rect 7452 1689 7880 1735
rect 7271 1611 7880 1689
rect 7271 1565 7282 1611
rect 7328 1565 7406 1611
rect 7452 1565 7880 1611
rect 7271 1487 7880 1565
rect 7271 1441 7282 1487
rect 7328 1441 7406 1487
rect 7452 1441 7880 1487
rect 7271 1363 7880 1441
rect 7271 1317 7282 1363
rect 7328 1317 7406 1363
rect 7452 1317 7880 1363
rect 7271 1239 7880 1317
rect 7271 1193 7282 1239
rect 7328 1193 7406 1239
rect 7452 1193 7880 1239
rect 7271 1115 7880 1193
rect 7271 1069 7282 1115
rect 7328 1069 7406 1115
rect 7452 1069 7880 1115
rect 7271 991 7880 1069
rect 7271 945 7282 991
rect 7328 945 7406 991
rect 7452 945 7880 991
rect 7271 867 7880 945
rect 7271 821 7282 867
rect 7328 821 7406 867
rect 7452 821 7880 867
rect 7271 743 7880 821
rect 7271 697 7282 743
rect 7328 697 7406 743
rect 7452 697 7880 743
rect 7271 658 7880 697
rect 7926 658 7937 5584
rect 7271 621 7937 658
rect 7271 619 7743 621
rect 7271 573 7282 619
rect 7328 573 7406 619
rect 7452 573 7743 619
rect 8455 599 9455 5643
rect 9973 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10565 5686
rect 9973 5584 10565 5640
rect 9973 658 9984 5584
rect 10030 5572 10565 5584
rect 10030 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10565 5572
rect 10030 5458 10565 5526
rect 10030 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10565 5458
rect 10030 5344 10565 5412
rect 10030 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10565 5344
rect 10030 5230 10565 5298
rect 10030 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10565 5230
rect 10030 5116 10565 5184
rect 10030 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10565 5116
rect 10030 5002 10565 5070
rect 10030 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10565 5002
rect 10030 4888 10565 4956
rect 10030 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10565 4888
rect 10030 4774 10565 4842
rect 10030 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10565 4774
rect 10030 4660 10565 4728
rect 10030 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10565 4660
rect 10030 4546 10565 4614
rect 10030 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10565 4546
rect 10030 4432 10565 4500
rect 10030 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10565 4432
rect 10030 4318 10565 4386
rect 10030 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10565 4318
rect 10030 4204 10565 4272
rect 10030 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10565 4204
rect 10030 4090 10565 4158
rect 10030 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10565 4090
rect 10030 3976 10565 4044
rect 10030 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10565 3976
rect 10030 3862 10565 3930
rect 10030 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10565 3862
rect 10030 3748 10565 3816
rect 10030 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10565 3748
rect 10030 3634 10565 3702
rect 10030 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10565 3634
rect 10030 3520 10565 3588
rect 10030 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10565 3520
rect 10030 3406 10565 3474
rect 10030 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10565 3406
rect 10030 3292 10565 3360
rect 10030 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10565 3292
rect 10030 3178 10565 3246
rect 10030 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10565 3178
rect 10030 3064 10565 3132
rect 10030 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10565 3064
rect 10030 2950 10565 3018
rect 10030 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10565 2950
rect 10030 2836 10565 2904
rect 10030 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10565 2836
rect 10030 2722 10565 2790
rect 10030 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10565 2722
rect 10030 2608 10565 2676
rect 10030 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10565 2608
rect 10030 2494 10565 2562
rect 10030 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10565 2494
rect 10030 2380 10565 2448
rect 10030 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10565 2380
rect 10030 2266 10565 2334
rect 10030 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10565 2266
rect 10030 2152 10565 2220
rect 10030 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10565 2152
rect 10030 2038 10565 2106
rect 10030 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10565 2038
rect 10030 1924 10565 1992
rect 10030 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10565 1924
rect 10030 1810 10565 1878
rect 10030 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10565 1810
rect 10030 1696 10565 1764
rect 10030 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10565 1696
rect 10030 1582 10565 1650
rect 10030 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10565 1582
rect 10030 1468 10565 1536
rect 10030 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10565 1468
rect 10030 1354 10565 1422
rect 10030 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10565 1354
rect 10030 1240 10565 1308
rect 10030 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10565 1240
rect 10030 1126 10565 1194
rect 10030 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10565 1126
rect 10030 1012 10565 1080
rect 10030 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10565 1012
rect 10030 898 10565 966
rect 10030 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10565 898
rect 10030 784 10565 852
rect 10030 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10565 784
rect 10030 670 10565 738
rect 10030 658 10394 670
rect 9973 624 10394 658
rect 10440 624 10508 670
rect 10554 624 10565 670
rect 9973 621 10565 624
rect 7271 495 7743 573
rect 7271 449 7282 495
rect 7328 449 7406 495
rect 7452 449 7743 495
rect 7271 371 7743 449
rect 7997 588 9913 599
rect 7997 542 8008 588
rect 9902 542 9913 588
rect 7997 399 9913 542
rect 10383 556 10565 621
rect 10383 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10565 556
rect 10383 442 10565 510
rect 7271 325 7282 371
rect 7328 325 7406 371
rect 7452 325 7743 371
rect 7271 247 7743 325
rect 7271 201 7282 247
rect 7328 201 7406 247
rect 7452 226 7743 247
rect 10383 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10565 442
rect 10383 328 10565 396
rect 10383 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10565 328
rect 10383 226 10565 282
rect 7452 214 10565 226
rect 7452 201 7612 214
rect 7271 168 7612 201
rect 7658 168 7726 214
rect 7772 168 7840 214
rect 7886 168 7954 214
rect 8000 168 8068 214
rect 8114 168 8182 214
rect 8228 168 8296 214
rect 8342 168 8410 214
rect 8456 168 8524 214
rect 8570 168 8638 214
rect 8684 168 8752 214
rect 8798 168 8866 214
rect 8912 168 8980 214
rect 9026 168 9094 214
rect 9140 168 9208 214
rect 9254 168 9322 214
rect 9368 168 9436 214
rect 9482 168 9550 214
rect 9596 168 9664 214
rect 9710 168 9778 214
rect 9824 168 9892 214
rect 9938 168 10006 214
rect 10052 168 10120 214
rect 10166 168 10234 214
rect 10280 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10565 214
rect 7271 123 10565 168
rect 7271 77 7282 123
rect 7328 77 7406 123
rect 7452 100 10565 123
rect 7452 77 7612 100
rect 7271 54 7612 77
rect 7658 54 7726 100
rect 7772 54 7840 100
rect 7886 54 7954 100
rect 8000 54 8068 100
rect 8114 54 8182 100
rect 8228 54 8296 100
rect 8342 54 8410 100
rect 8456 54 8524 100
rect 8570 54 8638 100
rect 8684 54 8752 100
rect 8798 54 8866 100
rect 8912 54 8980 100
rect 9026 54 9094 100
rect 9140 54 9208 100
rect 9254 54 9322 100
rect 9368 54 9436 100
rect 9482 54 9550 100
rect 9596 54 9664 100
rect 9710 54 9778 100
rect 9824 54 9892 100
rect 9938 54 10006 100
rect 10052 54 10120 100
rect 10166 54 10234 100
rect 10280 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10565 100
rect 7271 42 10565 54
use M1_PSUB_CDNS_40661954729136  M1_PSUB_CDNS_40661954729136_0
timestamp 1669390400
transform 1 0 10474 0 1 6176
box 0 0 1 1
use M1_PSUB_CDNS_40661954729141  M1_PSUB_CDNS_40661954729141_0
timestamp 1669390400
transform 0 -1 6417 1 0 12218
box 0 0 1 1
use M1_PSUB_CDNS_40661954729142  M1_PSUB_CDNS_40661954729142_0
timestamp 1669390400
transform 0 -1 8946 1 0 134
box 0 0 1 1
use M1_PSUB_CDNS_40661954729143  M1_PSUB_CDNS_40661954729143_0
timestamp 1669390400
transform 1 0 7367 0 1 3014
box 0 0 1 1
use M1_PSUB_CDNS_40661954729144  M1_PSUB_CDNS_40661954729144_0
timestamp 1669390400
transform 0 -1 6439 1 0 6127
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_0
timestamp 1669390400
transform 1 0 7955 0 -1 5621
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_1
timestamp 1669390400
transform 1 0 7955 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_2
timestamp 1669390400
transform 1 0 5519 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_3
timestamp 1669390400
transform 1 0 3083 0 1 6633
box 0 0 1 1
<< labels >>
rlabel metal1 s 5302 6126 5302 6126 4 VMINUS
port 1 nsew
<< properties >>
string GDS_END 4919486
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4911288
<< end >>
