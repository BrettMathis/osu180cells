magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 2800 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
rect 1550 190 1610 360
rect 1720 190 1780 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2230 190 2290 360
rect 2550 190 2610 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
rect 870 1090 930 1430
rect 1040 1090 1100 1430
rect 1210 1090 1270 1430
rect 1380 1090 1440 1430
rect 1550 1090 1610 1430
rect 1720 1090 1780 1430
rect 1890 1090 1950 1430
rect 2060 1090 2120 1430
rect 2230 1090 2290 1430
rect 2550 1090 2610 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 190 870 360
rect 930 298 1040 360
rect 930 252 962 298
rect 1008 252 1040 298
rect 930 190 1040 252
rect 1100 293 1210 360
rect 1100 247 1132 293
rect 1178 247 1210 293
rect 1100 190 1210 247
rect 1270 263 1380 360
rect 1270 217 1302 263
rect 1348 217 1380 263
rect 1270 190 1380 217
rect 1440 293 1550 360
rect 1440 247 1472 293
rect 1518 247 1550 293
rect 1440 190 1550 247
rect 1610 298 1720 360
rect 1610 252 1642 298
rect 1688 252 1720 298
rect 1610 190 1720 252
rect 1780 190 1890 360
rect 1950 190 2060 360
rect 2120 298 2230 360
rect 2120 252 2152 298
rect 2198 252 2230 298
rect 2120 190 2230 252
rect 2290 298 2390 360
rect 2290 252 2322 298
rect 2368 252 2390 298
rect 2290 190 2390 252
rect 2450 298 2550 360
rect 2450 252 2472 298
rect 2518 252 2550 298
rect 2450 190 2550 252
rect 2610 298 2710 360
rect 2610 252 2642 298
rect 2688 252 2710 298
rect 2610 190 2710 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1090 870 1430
rect 930 1377 1040 1430
rect 930 1143 962 1377
rect 1008 1143 1040 1377
rect 930 1090 1040 1143
rect 1100 1377 1210 1430
rect 1100 1143 1132 1377
rect 1178 1143 1210 1377
rect 1100 1090 1210 1143
rect 1270 1377 1380 1430
rect 1270 1143 1302 1377
rect 1348 1143 1380 1377
rect 1270 1090 1380 1143
rect 1440 1377 1550 1430
rect 1440 1143 1472 1377
rect 1518 1143 1550 1377
rect 1440 1090 1550 1143
rect 1610 1377 1720 1430
rect 1610 1143 1642 1377
rect 1688 1143 1720 1377
rect 1610 1090 1720 1143
rect 1780 1090 1890 1430
rect 1950 1090 2060 1430
rect 2120 1377 2230 1430
rect 2120 1143 2152 1377
rect 2198 1143 2230 1377
rect 2120 1090 2230 1143
rect 2290 1377 2390 1430
rect 2290 1143 2322 1377
rect 2368 1143 2390 1377
rect 2290 1090 2390 1143
rect 2450 1377 2550 1430
rect 2450 1143 2472 1377
rect 2518 1143 2550 1377
rect 2450 1090 2550 1143
rect 2610 1377 2710 1430
rect 2610 1143 2642 1377
rect 2688 1143 2710 1377
rect 2610 1090 2710 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 962 252 1008 298
rect 1132 247 1178 293
rect 1302 217 1348 263
rect 1472 247 1518 293
rect 1642 252 1688 298
rect 2152 252 2198 298
rect 2322 252 2368 298
rect 2472 252 2518 298
rect 2642 252 2688 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 962 1143 1008 1377
rect 1132 1143 1178 1377
rect 1302 1143 1348 1377
rect 1472 1143 1518 1377
rect 1642 1143 1688 1377
rect 2152 1143 2198 1377
rect 2322 1143 2368 1377
rect 2472 1143 2518 1377
rect 2642 1143 2688 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
rect 1290 1568 1380 1590
rect 1290 1522 1312 1568
rect 1358 1522 1380 1568
rect 1290 1500 1380 1522
rect 1530 1568 1620 1590
rect 1530 1522 1552 1568
rect 1598 1522 1620 1568
rect 1530 1500 1620 1522
rect 1770 1568 1860 1590
rect 1770 1522 1792 1568
rect 1838 1522 1860 1568
rect 1770 1500 1860 1522
rect 2010 1568 2100 1590
rect 2010 1522 2032 1568
rect 2078 1522 2100 1568
rect 2010 1500 2100 1522
rect 2250 1568 2340 1590
rect 2250 1522 2272 1568
rect 2318 1522 2340 1568
rect 2250 1500 2340 1522
rect 2490 1568 2580 1590
rect 2490 1522 2512 1568
rect 2558 1522 2580 1568
rect 2490 1500 2580 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
rect 1552 1522 1598 1568
rect 1792 1522 1838 1568
rect 2032 1522 2078 1568
rect 2272 1522 2318 1568
rect 2512 1522 2558 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 870 1430 930 1480
rect 1040 1430 1100 1480
rect 1210 1430 1270 1480
rect 1380 1430 1440 1480
rect 1550 1430 1610 1480
rect 1720 1430 1780 1480
rect 1890 1430 1950 1480
rect 2060 1430 2120 1480
rect 2230 1430 2290 1480
rect 2550 1430 2610 1480
rect 190 780 250 1090
rect 360 910 420 1090
rect 300 883 420 910
rect 300 837 327 883
rect 373 837 420 883
rect 300 810 420 837
rect 120 753 250 780
rect 120 707 147 753
rect 193 707 250 753
rect 120 680 250 707
rect 190 360 250 680
rect 360 360 420 810
rect 530 650 590 1090
rect 470 623 590 650
rect 470 577 497 623
rect 543 577 590 623
rect 470 550 590 577
rect 530 360 590 550
rect 700 910 760 1090
rect 870 1070 930 1090
rect 1040 1070 1100 1090
rect 870 1020 1100 1070
rect 700 883 820 910
rect 700 837 747 883
rect 793 837 820 883
rect 700 810 820 837
rect 700 360 760 810
rect 870 780 930 1020
rect 1210 910 1270 1090
rect 1150 883 1270 910
rect 1150 837 1177 883
rect 1223 837 1270 883
rect 1150 810 1270 837
rect 870 753 1020 780
rect 870 707 947 753
rect 993 707 1020 753
rect 870 680 1020 707
rect 870 430 930 680
rect 870 380 1100 430
rect 870 360 930 380
rect 1040 360 1100 380
rect 1210 360 1270 810
rect 1380 520 1440 1090
rect 1550 650 1610 1090
rect 1490 623 1610 650
rect 1490 577 1517 623
rect 1563 577 1610 623
rect 1490 550 1610 577
rect 1330 493 1440 520
rect 1330 447 1357 493
rect 1403 447 1440 493
rect 1330 420 1440 447
rect 1380 360 1440 420
rect 1550 360 1610 550
rect 1720 780 1780 1090
rect 1890 910 1950 1090
rect 1890 883 2010 910
rect 1890 837 1937 883
rect 1983 837 2010 883
rect 1890 810 2010 837
rect 1720 753 1840 780
rect 1720 707 1767 753
rect 1813 707 1840 753
rect 1720 680 1840 707
rect 1720 360 1780 680
rect 1890 360 1950 810
rect 2060 520 2120 1090
rect 2230 650 2290 1090
rect 2550 650 2610 1090
rect 2170 623 2290 650
rect 2170 577 2197 623
rect 2243 577 2290 623
rect 2170 550 2290 577
rect 2490 623 2610 650
rect 2490 577 2517 623
rect 2563 577 2610 623
rect 2490 550 2610 577
rect 2010 493 2120 520
rect 2010 447 2037 493
rect 2083 447 2120 493
rect 2010 420 2120 447
rect 2060 360 2120 420
rect 2230 360 2290 550
rect 2550 360 2610 550
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
rect 1550 140 1610 190
rect 1720 140 1780 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2230 140 2290 190
rect 2550 140 2610 190
<< polycontact >>
rect 327 837 373 883
rect 147 707 193 753
rect 497 577 543 623
rect 747 837 793 883
rect 1177 837 1223 883
rect 947 707 993 753
rect 1517 577 1563 623
rect 1357 447 1403 493
rect 1937 837 1983 883
rect 1767 707 1813 753
rect 2197 577 2243 623
rect 2517 577 2563 623
rect 2037 447 2083 493
<< metal1 >>
rect 0 1568 2800 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1552 1568
rect 1598 1566 1792 1568
rect 1838 1566 2032 1568
rect 2078 1566 2272 1568
rect 2318 1566 2512 1568
rect 2558 1566 2800 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 1366 1522 1552 1566
rect 1606 1522 1792 1566
rect 1846 1522 2032 1566
rect 2086 1522 2272 1566
rect 2326 1522 2512 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1794 1522
rect 1846 1514 2034 1522
rect 2086 1514 2274 1522
rect 2326 1514 2514 1522
rect 2566 1514 2800 1566
rect 0 1500 2800 1514
rect 110 1377 160 1430
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1040 160 1143
rect 280 1377 330 1500
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 1090 330 1143
rect 450 1377 500 1430
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1040 500 1143
rect 110 990 500 1040
rect 620 1377 670 1430
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 300 886 400 890
rect 300 834 324 886
rect 376 834 400 886
rect 300 830 400 834
rect 120 756 220 760
rect 120 704 144 756
rect 196 704 220 756
rect 120 700 220 704
rect 620 630 670 1143
rect 960 1377 1010 1500
rect 960 1143 962 1377
rect 1008 1143 1010 1377
rect 960 1090 1010 1143
rect 1130 1377 1180 1430
rect 1130 1143 1132 1377
rect 1178 1143 1180 1377
rect 1130 1040 1180 1143
rect 1300 1377 1350 1500
rect 1300 1143 1302 1377
rect 1348 1143 1350 1377
rect 1300 1090 1350 1143
rect 1470 1377 1520 1430
rect 1470 1143 1472 1377
rect 1518 1143 1520 1377
rect 1470 1040 1520 1143
rect 1130 990 1520 1040
rect 1640 1377 1690 1430
rect 1640 1143 1642 1377
rect 1688 1143 1690 1377
rect 720 886 1250 890
rect 720 834 744 886
rect 796 834 1174 886
rect 1226 834 1250 886
rect 720 830 1250 834
rect 920 756 1020 760
rect 920 704 944 756
rect 996 704 1020 756
rect 920 700 1020 704
rect 1640 630 1690 1143
rect 2150 1377 2200 1500
rect 2150 1143 2152 1377
rect 2198 1143 2200 1377
rect 2150 1090 2200 1143
rect 2320 1377 2370 1430
rect 2320 1143 2322 1377
rect 2368 1143 2370 1377
rect 2320 890 2370 1143
rect 2470 1377 2520 1500
rect 2470 1143 2472 1377
rect 2518 1143 2520 1377
rect 2470 1090 2520 1143
rect 2640 1377 2690 1430
rect 2640 1143 2642 1377
rect 2688 1143 2690 1377
rect 1910 886 2010 890
rect 1910 834 1934 886
rect 1986 834 2010 886
rect 1910 830 2010 834
rect 2320 886 2400 890
rect 2320 834 2324 886
rect 2376 834 2400 886
rect 2320 830 2400 834
rect 1740 756 1840 760
rect 1740 704 1764 756
rect 1816 704 1840 756
rect 1740 700 1840 704
rect 470 626 570 630
rect 470 574 494 626
rect 546 574 570 626
rect 470 570 570 574
rect 620 626 1590 630
rect 620 574 1514 626
rect 1566 574 1590 626
rect 620 570 1590 574
rect 1640 623 2270 630
rect 1640 577 2197 623
rect 2243 577 2270 623
rect 1640 570 2270 577
rect 110 410 500 460
rect 110 298 160 410
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 450 298 500 410
rect 450 252 452 298
rect 498 252 500 298
rect 450 190 500 252
rect 620 298 670 570
rect 1330 496 1430 500
rect 1330 444 1354 496
rect 1406 444 1430 496
rect 1330 440 1430 444
rect 620 252 622 298
rect 668 252 670 298
rect 620 190 670 252
rect 960 298 1010 360
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 120 1010 252
rect 1130 340 1520 390
rect 1130 293 1180 340
rect 1130 247 1132 293
rect 1178 247 1180 293
rect 1470 293 1520 340
rect 1130 190 1180 247
rect 1300 263 1350 290
rect 1300 217 1302 263
rect 1348 217 1350 263
rect 1300 120 1350 217
rect 1470 247 1472 293
rect 1518 247 1520 293
rect 1470 190 1520 247
rect 1640 298 1690 570
rect 2010 496 2110 500
rect 2010 444 2034 496
rect 2086 444 2110 496
rect 2010 440 2110 444
rect 1640 252 1642 298
rect 1688 252 1690 298
rect 1640 190 1690 252
rect 2150 298 2200 360
rect 2150 252 2152 298
rect 2198 252 2200 298
rect 2150 120 2200 252
rect 2320 298 2370 830
rect 2640 640 2690 1143
rect 2640 630 2720 640
rect 2490 626 2590 630
rect 2490 574 2514 626
rect 2566 574 2590 626
rect 2490 570 2590 574
rect 2640 626 2750 630
rect 2640 574 2674 626
rect 2726 574 2750 626
rect 2640 570 2750 574
rect 2640 560 2720 570
rect 2320 252 2322 298
rect 2368 252 2370 298
rect 2320 190 2370 252
rect 2470 298 2520 360
rect 2470 252 2472 298
rect 2518 252 2520 298
rect 2470 120 2520 252
rect 2640 298 2690 560
rect 2640 252 2642 298
rect 2688 252 2690 298
rect 2640 190 2690 252
rect 0 106 2800 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2800 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2800 54
rect 0 0 2800 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 1554 1522 1598 1566
rect 1598 1522 1606 1566
rect 1794 1522 1838 1566
rect 1838 1522 1846 1566
rect 2034 1522 2078 1566
rect 2078 1522 2086 1566
rect 2274 1522 2318 1566
rect 2318 1522 2326 1566
rect 2514 1522 2558 1566
rect 2558 1522 2566 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 1794 1514 1846 1522
rect 2034 1514 2086 1522
rect 2274 1514 2326 1522
rect 2514 1514 2566 1522
rect 324 883 376 886
rect 324 837 327 883
rect 327 837 373 883
rect 373 837 376 883
rect 324 834 376 837
rect 144 753 196 756
rect 144 707 147 753
rect 147 707 193 753
rect 193 707 196 753
rect 144 704 196 707
rect 744 883 796 886
rect 744 837 747 883
rect 747 837 793 883
rect 793 837 796 883
rect 744 834 796 837
rect 1174 883 1226 886
rect 1174 837 1177 883
rect 1177 837 1223 883
rect 1223 837 1226 883
rect 1174 834 1226 837
rect 944 753 996 756
rect 944 707 947 753
rect 947 707 993 753
rect 993 707 996 753
rect 944 704 996 707
rect 1934 883 1986 886
rect 1934 837 1937 883
rect 1937 837 1983 883
rect 1983 837 1986 883
rect 1934 834 1986 837
rect 2324 834 2376 886
rect 1764 753 1816 756
rect 1764 707 1767 753
rect 1767 707 1813 753
rect 1813 707 1816 753
rect 1764 704 1816 707
rect 494 623 546 626
rect 494 577 497 623
rect 497 577 543 623
rect 543 577 546 623
rect 494 574 546 577
rect 1514 623 1566 626
rect 1514 577 1517 623
rect 1517 577 1563 623
rect 1563 577 1566 623
rect 1514 574 1566 577
rect 1354 493 1406 496
rect 1354 447 1357 493
rect 1357 447 1403 493
rect 1403 447 1406 493
rect 1354 444 1406 447
rect 2034 493 2086 496
rect 2034 447 2037 493
rect 2037 447 2083 493
rect 2083 447 2086 493
rect 2034 444 2086 447
rect 2514 623 2566 626
rect 2514 577 2517 623
rect 2517 577 2563 623
rect 2563 577 2566 623
rect 2514 574 2566 577
rect 2674 574 2726 626
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect 1780 1570 1860 1580
rect 2020 1570 2100 1580
rect 2260 1570 2340 1580
rect 2500 1570 2580 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1510 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1510 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1510 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1510 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1510 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1510 1390 1514
rect 1530 1566 1630 1570
rect 1530 1514 1554 1566
rect 1606 1514 1630 1566
rect 1530 1510 1630 1514
rect 1770 1566 1870 1570
rect 1770 1514 1794 1566
rect 1846 1514 1870 1566
rect 1770 1510 1870 1514
rect 2010 1566 2110 1570
rect 2010 1514 2034 1566
rect 2086 1514 2110 1566
rect 2010 1510 2110 1514
rect 2250 1566 2350 1570
rect 2250 1514 2274 1566
rect 2326 1514 2350 1566
rect 2250 1510 2350 1514
rect 2490 1566 2590 1570
rect 2490 1514 2514 1566
rect 2566 1514 2590 1566
rect 2490 1510 2590 1514
rect 100 1500 180 1510
rect 340 1500 420 1510
rect 580 1500 660 1510
rect 820 1500 900 1510
rect 1060 1500 1140 1510
rect 1300 1500 1380 1510
rect 1540 1500 1620 1510
rect 1780 1500 1860 1510
rect 2020 1500 2100 1510
rect 2260 1500 2340 1510
rect 2500 1500 2580 1510
rect 310 890 390 900
rect 730 890 810 900
rect 1160 890 1240 900
rect 1920 890 2000 900
rect 2310 890 2390 900
rect 300 886 820 890
rect 300 834 324 886
rect 376 834 744 886
rect 796 834 820 886
rect 300 830 820 834
rect 1150 886 2010 890
rect 1150 834 1174 886
rect 1226 834 1934 886
rect 1986 834 2010 886
rect 1150 830 2010 834
rect 2300 886 2400 890
rect 2300 834 2324 886
rect 2376 834 2400 886
rect 2300 830 2400 834
rect 310 820 390 830
rect 730 820 810 830
rect 1160 820 1240 830
rect 1920 820 2000 830
rect 2310 820 2390 830
rect 130 760 210 770
rect 930 760 1010 770
rect 1750 760 1830 770
rect 120 756 1840 760
rect 120 704 144 756
rect 196 704 944 756
rect 996 704 1764 756
rect 1816 704 1840 756
rect 120 700 1840 704
rect 130 690 210 700
rect 930 690 1010 700
rect 1750 690 1830 700
rect 480 630 560 640
rect 1500 630 1580 640
rect 2500 630 2580 640
rect 2660 630 2740 640
rect 470 626 570 630
rect 470 574 494 626
rect 546 574 570 626
rect 470 570 570 574
rect 1490 626 2590 630
rect 1490 574 1514 626
rect 1566 574 2514 626
rect 2566 574 2590 626
rect 1490 570 2590 574
rect 2650 626 2750 630
rect 2650 574 2674 626
rect 2726 574 2750 626
rect 2650 570 2750 574
rect 480 560 560 570
rect 1500 560 1580 570
rect 2500 560 2580 570
rect 2660 560 2740 570
rect 490 500 550 560
rect 2510 550 2570 560
rect 1340 500 1420 510
rect 2020 500 2100 510
rect 490 496 2110 500
rect 490 444 1354 496
rect 1406 444 2034 496
rect 2086 444 2110 496
rect 490 440 2110 444
rect 1340 430 1420 440
rect 2020 430 2100 440
rect 1350 420 1410 430
rect 2030 420 2090 430
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 50 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 50 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 50 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 50 2590 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
rect 1780 40 1860 50
rect 2020 40 2100 50
rect 2260 40 2340 50
rect 2500 40 2580 50
<< labels >>
rlabel metal2 s 100 40 180 120 4 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 100 1500 180 1580 4 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 130 690 210 770 4 A
port 1 nsew signal input
rlabel metal2 s 310 820 390 900 4 B
port 2 nsew signal input
rlabel metal2 s 490 440 550 640 4 CI
port 3 nsew signal input
rlabel metal2 s 2660 560 2740 640 4 CO
port 4 nsew signal output
rlabel metal2 s 2310 820 2390 900 4 S
port 5 nsew signal output
rlabel metal2 s 930 690 1010 770 1 A
port 1 nsew signal input
rlabel metal2 s 1750 690 1830 770 1 A
port 1 nsew signal input
rlabel metal2 s 120 700 1840 760 1 A
port 1 nsew signal input
rlabel metal1 s 120 700 220 760 1 A
port 1 nsew signal input
rlabel metal1 s 920 700 1020 760 1 A
port 1 nsew signal input
rlabel metal1 s 1740 700 1840 760 1 A
port 1 nsew signal input
rlabel metal2 s 730 820 810 900 1 B
port 2 nsew signal input
rlabel metal2 s 300 830 820 890 1 B
port 2 nsew signal input
rlabel metal2 s 1160 820 1240 900 1 B
port 2 nsew signal input
rlabel metal2 s 1920 820 2000 900 1 B
port 2 nsew signal input
rlabel metal2 s 1150 830 2010 890 1 B
port 2 nsew signal input
rlabel metal1 s 300 830 400 890 1 B
port 2 nsew signal input
rlabel metal1 s 720 830 1250 890 1 B
port 2 nsew signal input
rlabel metal1 s 1910 830 2010 890 1 B
port 2 nsew signal input
rlabel metal2 s 480 560 560 640 1 CI
port 3 nsew signal input
rlabel metal2 s 470 570 570 630 1 CI
port 3 nsew signal input
rlabel metal2 s 1350 420 1410 510 1 CI
port 3 nsew signal input
rlabel metal2 s 1340 430 1420 510 1 CI
port 3 nsew signal input
rlabel metal2 s 2030 420 2090 510 1 CI
port 3 nsew signal input
rlabel metal2 s 2020 430 2100 510 1 CI
port 3 nsew signal input
rlabel metal2 s 490 440 2110 500 1 CI
port 3 nsew signal input
rlabel metal1 s 470 570 570 630 1 CI
port 3 nsew signal input
rlabel metal1 s 1330 440 1430 500 1 CI
port 3 nsew signal input
rlabel metal1 s 2010 440 2110 500 1 CI
port 3 nsew signal input
rlabel metal2 s 2650 570 2750 630 1 CO
port 4 nsew signal output
rlabel metal1 s 2640 190 2690 1430 1 CO
port 4 nsew signal output
rlabel metal1 s 2640 560 2720 640 1 CO
port 4 nsew signal output
rlabel metal1 s 2640 570 2750 630 1 CO
port 4 nsew signal output
rlabel metal2 s 2300 830 2400 890 1 S
port 5 nsew signal output
rlabel metal1 s 2320 190 2370 1430 1 S
port 5 nsew signal output
rlabel metal1 s 2320 830 2400 890 1 S
port 5 nsew signal output
rlabel metal2 s 90 1510 190 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 340 1500 420 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 330 1510 430 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 580 1500 660 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 570 1510 670 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 820 1500 900 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 810 1510 910 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1060 1500 1140 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1050 1510 1150 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1300 1500 1380 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1290 1510 1390 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1540 1500 1620 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1530 1510 1630 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1780 1500 1860 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1770 1510 1870 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2020 1500 2100 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2010 1510 2110 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2260 1500 2340 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2250 1510 2350 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2500 1500 2580 1580 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2490 1510 2590 1570 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 280 1090 330 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 960 1090 1010 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 1300 1090 1350 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 2150 1090 2200 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 2470 1090 2520 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 0 1500 2800 1620 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1780 40 1860 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1770 50 1870 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2020 40 2100 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2010 50 2110 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2260 40 2340 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2250 50 2350 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2500 40 2580 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2490 50 2590 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 280 0 330 360 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 960 0 1010 360 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 1300 0 1350 290 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 2150 0 2200 360 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 2470 0 2520 360 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 0 0 2800 120 1 VSS
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2800 1620
string GDS_END 25498
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 136
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
