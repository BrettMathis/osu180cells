magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -63 788 64 828
rect -63 736 -26 788
rect 26 736 64 788
rect -63 570 64 736
rect -63 518 -26 570
rect 26 518 64 570
rect -63 353 64 518
rect -63 301 -26 353
rect 26 301 64 353
rect -63 135 64 301
rect -63 83 -26 135
rect 26 83 64 135
rect -63 -83 64 83
rect -63 -135 -26 -83
rect 26 -135 64 -83
rect -63 -301 64 -135
rect -63 -353 -26 -301
rect 26 -353 64 -301
rect -63 -518 64 -353
rect -63 -570 -26 -518
rect 26 -570 64 -518
rect -63 -736 64 -570
rect -63 -788 -26 -736
rect 26 -788 64 -736
rect -63 -828 64 -788
<< via1 >>
rect -26 736 26 788
rect -26 518 26 570
rect -26 301 26 353
rect -26 83 26 135
rect -26 -135 26 -83
rect -26 -353 26 -301
rect -26 -570 26 -518
rect -26 -788 26 -736
<< metal2 >>
rect -63 788 64 828
rect -63 736 -26 788
rect 26 736 64 788
rect -63 570 64 736
rect -63 518 -26 570
rect 26 518 64 570
rect -63 353 64 518
rect -63 301 -26 353
rect 26 301 64 353
rect -63 135 64 301
rect -63 83 -26 135
rect 26 83 64 135
rect -63 -83 64 83
rect -63 -135 -26 -83
rect 26 -135 64 -83
rect -63 -301 64 -135
rect -63 -353 -26 -301
rect 26 -353 64 -301
rect -63 -518 64 -353
rect -63 -570 -26 -518
rect 26 -570 64 -518
rect -63 -736 64 -570
rect -63 -788 -26 -736
rect 26 -788 64 -736
rect -63 -828 64 -788
<< properties >>
string GDS_END 284024
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 283380
<< end >>
