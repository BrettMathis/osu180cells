magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 6583 57808 9560 58732
rect 13849 58458 15116 58748
rect 13849 58381 15441 58458
rect 10186 57817 10786 57889
rect 13850 57808 15441 58381
rect 6583 57758 8962 57808
rect 16520 57776 21087 58703
<< mvndiff >>
rect 2123 57660 2278 58048
rect 25490 57660 25646 58048
<< mvpsubdiff >>
rect 15782 58582 16254 58639
rect 15782 58536 15837 58582
rect 15883 58536 15995 58582
rect 16041 58536 16153 58582
rect 16199 58536 16254 58582
rect 15782 58479 16254 58536
<< mvnsubdiff >>
rect 13985 58582 14931 58639
rect 13985 58536 14040 58582
rect 14086 58536 14198 58582
rect 14244 58536 14356 58582
rect 14402 58536 14514 58582
rect 14560 58536 14673 58582
rect 14719 58536 14831 58582
rect 14877 58536 14931 58582
rect 13985 58479 14931 58536
<< mvpsubdiffcont >>
rect 15837 58536 15883 58582
rect 15995 58536 16041 58582
rect 16153 58536 16199 58582
<< mvnsubdiffcont >>
rect 14040 58536 14086 58582
rect 14198 58536 14244 58582
rect 14356 58536 14402 58582
rect 14514 58536 14560 58582
rect 14673 58536 14719 58582
rect 14831 58536 14877 58582
<< polysilicon >>
rect 13623 58516 13801 58535
rect 13623 58470 13642 58516
rect 13782 58470 13801 58516
rect 15364 58564 15467 58583
rect 15364 58518 15390 58564
rect 15436 58518 15467 58564
rect 13623 58451 13801 58470
rect 6556 58296 6690 58416
rect 9314 58318 9448 58423
rect 6556 58192 6659 58296
rect 6374 58072 6690 58192
rect 9314 58178 9358 58318
rect 9404 58178 9448 58318
rect 11998 58231 12082 58250
rect 11998 58192 12017 58231
rect 9314 58073 9448 58178
rect 11043 58072 11385 58192
rect 11914 58091 12017 58192
rect 12063 58091 12082 58231
rect 11914 58072 12082 58091
rect 13664 58073 13768 58451
rect 15364 58192 15467 58518
rect 18271 58306 18355 58416
rect 13915 58072 13986 58192
rect 15305 58072 15467 58192
rect 15583 58271 15667 58290
rect 15583 58131 15602 58271
rect 15648 58192 15667 58271
rect 15648 58131 15755 58192
rect 15583 58072 15755 58131
rect 16255 58072 16656 58192
rect 17975 58072 18045 58192
rect 18271 58166 18290 58306
rect 18336 58166 18355 58306
rect 18271 58072 18355 58166
rect 21010 58192 21113 58416
rect 21010 58072 21325 58192
rect 23347 58072 23417 58192
<< polycontact >>
rect 13642 58470 13782 58516
rect 15390 58518 15436 58564
rect 9358 58178 9404 58318
rect 12017 58091 12063 58231
rect 15602 58131 15648 58271
rect 18290 58166 18336 58306
<< metal1 >>
rect 2123 57916 4017 58567
rect 4324 58252 6336 58639
rect 6728 58506 7700 58546
rect 6728 58454 6766 58506
rect 6818 58454 6977 58506
rect 7029 58454 7188 58506
rect 7240 58454 7399 58506
rect 7451 58454 7610 58506
rect 7662 58454 7700 58506
rect 6728 58414 7700 58454
rect 11385 58531 11913 58619
rect 11385 58479 11575 58531
rect 11627 58479 11755 58531
rect 11807 58479 11913 58531
rect 9323 58318 9439 58385
rect 6482 58188 6767 58308
rect 4335 58045 5307 58085
rect 6482 58077 6598 58188
rect 9323 58178 9358 58318
rect 9404 58178 9439 58318
rect 10338 58308 10888 58315
rect 10337 58274 10888 58308
rect 10337 58222 10376 58274
rect 10428 58222 10587 58274
rect 10639 58222 10798 58274
rect 10850 58222 10888 58274
rect 10337 58188 10888 58222
rect 11385 58313 11913 58479
rect 13531 58582 14912 58619
rect 15755 58618 16283 58619
rect 13531 58578 14040 58582
rect 13531 58526 14033 58578
rect 14086 58536 14198 58582
rect 14244 58578 14356 58582
rect 14085 58526 14244 58536
rect 14296 58536 14356 58578
rect 14402 58578 14514 58582
rect 14402 58536 14455 58578
rect 14296 58526 14455 58536
rect 14507 58536 14514 58578
rect 14560 58536 14673 58582
rect 14719 58536 14831 58582
rect 14877 58536 14912 58582
rect 14507 58526 14912 58536
rect 13531 58517 14912 58526
rect 13531 58465 13569 58517
rect 13621 58516 13781 58517
rect 13621 58470 13642 58516
rect 13833 58499 14912 58517
rect 15061 58582 16283 58618
rect 15061 58578 15837 58582
rect 15061 58526 15100 58578
rect 15152 58526 15311 58578
rect 15363 58564 15522 58578
rect 15363 58526 15390 58564
rect 15061 58518 15390 58526
rect 15436 58526 15522 58564
rect 15574 58526 15733 58578
rect 15785 58536 15837 58578
rect 15883 58536 15995 58582
rect 16041 58536 16153 58582
rect 16199 58536 16283 58582
rect 20112 58540 20874 58546
rect 15785 58526 16283 58536
rect 15436 58518 16283 58526
rect 13833 58486 14545 58499
rect 13833 58485 14040 58486
rect 15061 58485 16283 58518
rect 13621 58465 13781 58470
rect 13833 58465 13871 58485
rect 13531 58424 13871 58465
rect 11385 58261 11575 58313
rect 11627 58261 11755 58313
rect 11807 58261 11913 58313
rect 15591 58271 15659 58282
rect 11385 58221 11913 58261
rect 12006 58231 12334 58268
rect 10338 58182 10888 58188
rect 4335 57993 4373 58045
rect 4425 57993 4584 58045
rect 4636 57993 4795 58045
rect 4847 57993 5006 58045
rect 5058 57993 5217 58045
rect 5269 57993 5307 58045
rect 4335 57953 5307 57993
rect 6240 57957 6598 58077
rect 6728 58043 7700 58083
rect 6728 57991 6766 58043
rect 6818 57991 6977 58043
rect 7029 57991 7188 58043
rect 7240 57991 7399 58043
rect 7451 57991 7610 58043
rect 7662 57991 7700 58043
rect 6728 57951 7700 57991
rect 9323 58077 9439 58178
rect 12006 58091 12017 58231
rect 12063 58222 12334 58231
rect 13509 58222 14174 58268
rect 15591 58267 15602 58271
rect 12063 58091 12074 58222
rect 15268 58221 15602 58267
rect 15591 58131 15602 58221
rect 15648 58131 15659 58271
rect 15755 58188 16283 58485
rect 16656 58506 20942 58540
rect 16656 58454 20151 58506
rect 20203 58454 20362 58506
rect 20414 58454 20573 58506
rect 20625 58454 20784 58506
rect 20836 58454 20942 58506
rect 16656 58420 20942 58454
rect 16656 58236 17974 58420
rect 20112 58413 20874 58420
rect 18279 58306 18347 58317
rect 15591 58120 15659 58131
rect 18279 58166 18290 58306
rect 18336 58166 18347 58306
rect 20898 58221 21184 58267
rect 18279 58155 18347 58166
rect 12006 58080 12074 58091
rect 9323 57957 11913 58077
rect 12294 58043 13478 58084
rect 18279 58077 18346 58155
rect 12294 57991 12333 58043
rect 12385 57991 12544 58043
rect 12596 57991 12755 58043
rect 12807 57991 12966 58043
rect 13018 57991 13177 58043
rect 13229 57991 13387 58043
rect 13439 57991 13478 58043
rect 13570 57998 14174 58044
rect 12294 57950 13478 57991
rect 15755 57957 18346 58077
rect 20112 58043 20874 58083
rect 20112 57991 20151 58043
rect 20203 57991 20362 58043
rect 20414 57991 20573 58043
rect 20625 57991 20784 58043
rect 20836 57991 20874 58043
rect 21067 58043 21184 58221
rect 21324 58202 23346 58619
rect 22366 58043 23338 58083
rect 21067 57997 21425 58043
rect 20112 57950 20874 57991
rect 22366 57991 22404 58043
rect 22456 57991 22615 58043
rect 22667 57991 22826 58043
rect 22878 57991 23037 58043
rect 23089 57991 23248 58043
rect 23300 57991 23338 58043
rect 22366 57951 23338 57991
rect 23751 57916 25646 58567
rect 2123 57665 2278 57916
rect 25490 57665 25646 57916
<< via1 >>
rect 6766 58454 6818 58506
rect 6977 58454 7029 58506
rect 7188 58454 7240 58506
rect 7399 58454 7451 58506
rect 7610 58454 7662 58506
rect 11575 58479 11627 58531
rect 11755 58479 11807 58531
rect 10376 58222 10428 58274
rect 10587 58222 10639 58274
rect 10798 58222 10850 58274
rect 14033 58536 14040 58578
rect 14040 58536 14085 58578
rect 14033 58526 14085 58536
rect 14244 58526 14296 58578
rect 14455 58526 14507 58578
rect 13569 58465 13621 58517
rect 13781 58516 13833 58517
rect 13781 58470 13782 58516
rect 13782 58470 13833 58516
rect 15100 58526 15152 58578
rect 15311 58526 15363 58578
rect 15522 58526 15574 58578
rect 15733 58526 15785 58578
rect 13781 58465 13833 58470
rect 11575 58261 11627 58313
rect 11755 58261 11807 58313
rect 4373 57993 4425 58045
rect 4584 57993 4636 58045
rect 4795 57993 4847 58045
rect 5006 57993 5058 58045
rect 5217 57993 5269 58045
rect 6766 57991 6818 58043
rect 6977 57991 7029 58043
rect 7188 57991 7240 58043
rect 7399 57991 7451 58043
rect 7610 57991 7662 58043
rect 20151 58454 20203 58506
rect 20362 58454 20414 58506
rect 20573 58454 20625 58506
rect 20784 58454 20836 58506
rect 12333 57991 12385 58043
rect 12544 57991 12596 58043
rect 12755 57991 12807 58043
rect 12966 57991 13018 58043
rect 13177 57991 13229 58043
rect 13387 57991 13439 58043
rect 20151 57991 20203 58043
rect 20362 57991 20414 58043
rect 20573 57991 20625 58043
rect 20784 57991 20836 58043
rect 22404 57991 22456 58043
rect 22615 57991 22667 58043
rect 22826 57991 22878 58043
rect 23037 57991 23089 58043
rect 23248 57991 23300 58043
<< metal2 >>
rect 2092 57613 4211 58676
rect 5550 58528 6347 58601
rect 5550 58472 5611 58528
rect 5667 58472 5822 58528
rect 5878 58472 6033 58528
rect 6089 58472 6244 58528
rect 6300 58472 6347 58528
rect 4334 58047 5307 58086
rect 4334 57991 4371 58047
rect 4427 57991 4582 58047
rect 4638 57991 4793 58047
rect 4849 57991 5004 58047
rect 5060 57991 5215 58047
rect 5271 57991 5307 58047
rect 4334 57953 5307 57991
rect 5550 57613 6347 58472
rect 6451 58506 7738 58601
rect 6451 58454 6766 58506
rect 6818 58454 6977 58506
rect 7029 58454 7188 58506
rect 7240 58454 7399 58506
rect 7451 58454 7610 58506
rect 7662 58454 7738 58506
rect 6451 58043 7738 58454
rect 6451 57991 6766 58043
rect 6818 57991 6977 58043
rect 7029 57991 7188 58043
rect 7240 57991 7399 58043
rect 7451 57991 7610 58043
rect 7662 57991 7738 58043
rect 6451 57613 7738 57991
rect 8186 58045 9066 58084
rect 8186 57989 8222 58045
rect 8278 57989 8433 58045
rect 8489 57989 8644 58045
rect 8700 57989 8855 58045
rect 8911 57989 9066 58045
rect 8186 57613 9066 57989
rect 9591 57613 10186 58601
rect 10276 58274 10941 58601
rect 10276 58222 10376 58274
rect 10428 58222 10587 58274
rect 10639 58222 10798 58274
rect 10850 58222 10941 58274
rect 10276 57613 10941 58222
rect 11537 58531 11846 58601
rect 13994 58578 14545 58619
rect 11537 58528 11575 58531
rect 11627 58528 11755 58531
rect 11807 58528 11846 58531
rect 11537 58472 11573 58528
rect 11629 58472 11753 58528
rect 11809 58472 11846 58528
rect 11537 58313 11846 58472
rect 13531 58517 13871 58558
rect 13531 58465 13569 58517
rect 13621 58465 13781 58517
rect 13833 58465 13871 58517
rect 13531 58424 13871 58465
rect 13994 58526 14033 58578
rect 14085 58526 14244 58578
rect 14296 58526 14455 58578
rect 14507 58526 14545 58578
rect 11537 58261 11575 58313
rect 11627 58261 11755 58313
rect 11807 58261 11846 58313
rect 11537 57613 11846 58261
rect 12294 58045 13478 58084
rect 12294 57989 12331 58045
rect 12387 57989 12542 58045
rect 12598 57989 12753 58045
rect 12809 57989 12964 58045
rect 13020 57989 13175 58045
rect 13231 57989 13385 58045
rect 13441 57989 13478 58045
rect 12294 57950 13478 57989
rect 13994 58038 14545 58526
rect 13994 57982 14031 58038
rect 14087 57982 14242 58038
rect 14298 57982 14453 58038
rect 14509 57982 14545 58038
rect 13994 57944 14545 57982
rect 15026 58578 15887 58619
rect 15026 58526 15100 58578
rect 15152 58526 15311 58578
rect 15363 58526 15522 58578
rect 15574 58526 15733 58578
rect 15785 58526 15887 58578
rect 12040 57628 12639 57764
rect 12040 57572 12100 57628
rect 12156 57572 12311 57628
rect 12367 57572 12522 57628
rect 12578 57572 12639 57628
rect 15026 57613 15887 58526
rect 20112 58506 21313 58601
rect 20112 58454 20151 58506
rect 20203 58454 20362 58506
rect 20414 58454 20573 58506
rect 20625 58454 20784 58506
rect 20836 58454 21313 58506
rect 20112 58043 21313 58454
rect 20112 57991 20151 58043
rect 20203 57991 20362 58043
rect 20414 57991 20573 58043
rect 20625 57991 20784 58043
rect 20836 57991 21313 58043
rect 20112 57613 21313 57991
rect 21421 58528 22236 58619
rect 21421 58472 21458 58528
rect 21514 58472 21669 58528
rect 21725 58472 21880 58528
rect 21936 58472 22091 58528
rect 22147 58472 22236 58528
rect 21421 57613 22236 58472
rect 22365 58045 23338 58084
rect 22365 57989 22402 58045
rect 22458 57989 22613 58045
rect 22669 57989 22824 58045
rect 22880 57989 23035 58045
rect 23091 57989 23246 58045
rect 23302 57989 23338 58045
rect 22365 57951 23338 57989
rect 23549 57613 25677 58676
rect 12040 57499 12639 57572
rect 8561 -21 8691 112
rect 12841 -164 12971 -31
rect 13219 -164 13348 -31
rect 13597 -164 13726 -31
rect 13974 -164 14104 -31
rect 14352 -164 14481 -31
rect 14730 -164 14859 -31
rect 16882 -164 17011 -31
rect 17260 -164 17389 -31
rect 17637 -164 17767 -31
rect 18015 -164 18144 -31
rect 18393 -164 18522 -31
rect 18770 -164 18900 -31
rect 19148 -164 19277 -31
rect 19526 -164 19655 -31
<< via2 >>
rect 5611 58472 5667 58528
rect 5822 58472 5878 58528
rect 6033 58472 6089 58528
rect 6244 58472 6300 58528
rect 4371 58045 4427 58047
rect 4371 57993 4373 58045
rect 4373 57993 4425 58045
rect 4425 57993 4427 58045
rect 4371 57991 4427 57993
rect 4582 58045 4638 58047
rect 4582 57993 4584 58045
rect 4584 57993 4636 58045
rect 4636 57993 4638 58045
rect 4582 57991 4638 57993
rect 4793 58045 4849 58047
rect 4793 57993 4795 58045
rect 4795 57993 4847 58045
rect 4847 57993 4849 58045
rect 4793 57991 4849 57993
rect 5004 58045 5060 58047
rect 5004 57993 5006 58045
rect 5006 57993 5058 58045
rect 5058 57993 5060 58045
rect 5004 57991 5060 57993
rect 5215 58045 5271 58047
rect 5215 57993 5217 58045
rect 5217 57993 5269 58045
rect 5269 57993 5271 58045
rect 5215 57991 5271 57993
rect 8222 57989 8278 58045
rect 8433 57989 8489 58045
rect 8644 57989 8700 58045
rect 8855 57989 8911 58045
rect 11573 58479 11575 58528
rect 11575 58479 11627 58528
rect 11627 58479 11629 58528
rect 11573 58472 11629 58479
rect 11753 58479 11755 58528
rect 11755 58479 11807 58528
rect 11807 58479 11809 58528
rect 11753 58472 11809 58479
rect 12331 58043 12387 58045
rect 12331 57991 12333 58043
rect 12333 57991 12385 58043
rect 12385 57991 12387 58043
rect 12331 57989 12387 57991
rect 12542 58043 12598 58045
rect 12542 57991 12544 58043
rect 12544 57991 12596 58043
rect 12596 57991 12598 58043
rect 12542 57989 12598 57991
rect 12753 58043 12809 58045
rect 12753 57991 12755 58043
rect 12755 57991 12807 58043
rect 12807 57991 12809 58043
rect 12753 57989 12809 57991
rect 12964 58043 13020 58045
rect 12964 57991 12966 58043
rect 12966 57991 13018 58043
rect 13018 57991 13020 58043
rect 12964 57989 13020 57991
rect 13175 58043 13231 58045
rect 13175 57991 13177 58043
rect 13177 57991 13229 58043
rect 13229 57991 13231 58043
rect 13175 57989 13231 57991
rect 13385 58043 13441 58045
rect 13385 57991 13387 58043
rect 13387 57991 13439 58043
rect 13439 57991 13441 58043
rect 13385 57989 13441 57991
rect 14031 57982 14087 58038
rect 14242 57982 14298 58038
rect 14453 57982 14509 58038
rect 12100 57572 12156 57628
rect 12311 57572 12367 57628
rect 12522 57572 12578 57628
rect 21458 58472 21514 58528
rect 21669 58472 21725 58528
rect 21880 58472 21936 58528
rect 22091 58472 22147 58528
rect 22402 58043 22458 58045
rect 22402 57991 22404 58043
rect 22404 57991 22456 58043
rect 22456 57991 22458 58043
rect 22402 57989 22458 57991
rect 22613 58043 22669 58045
rect 22613 57991 22615 58043
rect 22615 57991 22667 58043
rect 22667 57991 22669 58043
rect 22613 57989 22669 57991
rect 22824 58043 22880 58045
rect 22824 57991 22826 58043
rect 22826 57991 22878 58043
rect 22878 57991 22880 58043
rect 22824 57989 22880 57991
rect 23035 58043 23091 58045
rect 23035 57991 23037 58043
rect 23037 57991 23089 58043
rect 23089 57991 23091 58043
rect 23035 57989 23091 57991
rect 23246 58043 23302 58045
rect 23246 57991 23248 58043
rect 23248 57991 23300 58043
rect 23300 57991 23302 58043
rect 23246 57989 23302 57991
<< metal3 >>
rect 69 58433 199 58567
rect 1725 58528 25945 58601
rect 1725 58472 5611 58528
rect 5667 58472 5822 58528
rect 5878 58472 6033 58528
rect 6089 58472 6244 58528
rect 6300 58472 11573 58528
rect 11629 58472 11753 58528
rect 11809 58472 21458 58528
rect 21514 58472 21669 58528
rect 21725 58472 21880 58528
rect 21936 58472 22091 58528
rect 22147 58472 25945 58528
rect 1725 58399 25945 58472
rect -1 57973 128 58107
rect 1725 58047 5307 58141
rect 1725 57991 4371 58047
rect 4427 57991 4582 58047
rect 4638 57991 4793 58047
rect 4849 57991 5004 58047
rect 5060 57991 5215 58047
rect 5271 57991 5307 58047
rect 1725 57939 5307 57991
rect 8186 58045 13478 58084
rect 8186 57989 8222 58045
rect 8278 57989 8433 58045
rect 8489 57989 8644 58045
rect 8700 57989 8855 58045
rect 8911 57989 12331 58045
rect 12387 57989 12542 58045
rect 12598 57989 12753 58045
rect 12809 57989 12964 58045
rect 13020 57989 13175 58045
rect 13231 57989 13385 58045
rect 13441 57989 13478 58045
rect 13994 58038 14545 58077
rect 13994 58003 14031 58038
rect 8186 57950 13478 57989
rect 13993 57982 14031 58003
rect 14087 57982 14242 58038
rect 14298 57982 14453 58038
rect 14509 57982 14545 58038
rect 13993 57944 14545 57982
rect 22365 58045 25945 58141
rect 22365 57989 22402 58045
rect 22458 57989 22613 58045
rect 22669 57989 22824 58045
rect 22880 57989 23035 58045
rect 23091 57989 23246 58045
rect 23302 57989 25945 58045
rect 69 57533 199 57667
rect 12063 57628 12615 57667
rect 13993 57632 14092 57944
rect 22365 57939 25945 57989
rect 27640 57973 27769 58107
rect 12063 57572 12100 57628
rect 12156 57572 12311 57628
rect 12367 57572 12522 57628
rect 12578 57572 12615 57628
rect 12063 57533 12615 57572
rect -1 57093 128 57227
rect 27640 57093 27769 57227
rect -1 56173 128 56307
rect 27640 56173 27769 56307
rect -1 55293 128 55427
rect 27640 55293 27769 55427
rect -1 54373 128 54507
rect 27640 54373 27769 54507
rect -1 53493 128 53627
rect 27640 53493 27769 53627
rect -1 52573 128 52707
rect 27640 52573 27769 52707
rect -1 51693 128 51827
rect 27640 51693 27769 51827
rect -1 50773 128 50907
rect 27640 50773 27769 50907
rect -1 49893 128 50027
rect 27640 49893 27769 50027
rect -1 48973 128 49107
rect 27640 48973 27769 49107
rect -1 48093 128 48227
rect 27640 48093 27769 48227
rect -1 47173 128 47307
rect 27640 47173 27769 47307
rect -1 46293 128 46427
rect 27640 46293 27769 46427
rect -1 45373 128 45507
rect 27640 45373 27769 45507
rect -1 44493 128 44627
rect 27640 44493 27769 44627
rect -1 43573 128 43707
rect 27640 43573 27769 43707
rect -1 42693 128 42827
rect 27640 42693 27769 42827
rect -1 41773 128 41907
rect 27640 41773 27769 41907
rect -1 40893 128 41027
rect 27640 40893 27769 41027
rect -1 39973 128 40107
rect 27640 39973 27769 40107
rect -1 39093 128 39227
rect 27640 39093 27769 39227
rect -1 38173 128 38307
rect 27640 38173 27769 38307
rect -1 37293 128 37427
rect 27640 37293 27769 37427
rect -1 36373 128 36507
rect 27640 36373 27769 36507
rect -1 35493 128 35627
rect 27640 35493 27769 35627
rect -1 34573 128 34707
rect 27640 34573 27769 34707
rect -1 33693 128 33827
rect 27640 33693 27769 33827
rect -1 32773 128 32907
rect 27640 32773 27769 32907
rect -1 31893 128 32027
rect 27640 31893 27769 32027
rect -1 30973 128 31107
rect 27640 30973 27769 31107
rect -1 30093 128 30227
rect 27640 30093 27769 30227
rect -1 29173 128 29307
rect 27640 29173 27769 29307
rect -1 28273 128 28407
rect 27640 28273 27769 28407
rect -1 27393 128 27527
rect 27640 27393 27769 27527
rect -1 26473 128 26607
rect 27640 26473 27769 26607
rect -1 25593 128 25727
rect 27640 25593 27769 25727
rect -1 24673 128 24807
rect 27640 24673 27769 24807
rect -1 23793 128 23927
rect 27640 23793 27769 23927
rect -1 22873 128 23007
rect 27640 22873 27769 23007
rect -1 21993 128 22127
rect 27640 21993 27769 22127
rect -1 21073 128 21207
rect 27640 21073 27769 21207
rect -1 20193 128 20327
rect 27640 20193 27769 20327
rect -1 19273 128 19407
rect 27640 19273 27769 19407
rect -1 18393 128 18527
rect 27640 18393 27769 18527
rect -1 17473 128 17607
rect 27640 17473 27769 17607
rect -1 16593 128 16727
rect 27640 16593 27769 16727
rect -1 15673 128 15807
rect 27640 15673 27769 15807
rect -1 14793 128 14927
rect 27640 14793 27769 14927
rect -1 13873 128 14007
rect 27640 13873 27769 14007
rect -1 12993 128 13127
rect 27640 12993 27769 13127
rect -1 12073 128 12207
rect 27640 12073 27769 12207
rect -1 11193 128 11327
rect 27640 11193 27769 11327
rect -1 10273 128 10407
rect 27640 10273 27769 10407
rect -1 9393 128 9527
rect 27640 9393 27769 9527
rect -1 8473 128 8607
rect 27640 8473 27769 8607
rect -1 7593 128 7727
rect 27640 7593 27769 7727
rect -1 6673 128 6807
rect 27640 6673 27769 6807
rect -1 5793 128 5927
rect 27640 5793 27769 5927
rect -1 4873 128 5007
rect 27640 4873 27769 5007
rect -1 3993 128 4127
rect 27640 3993 27769 4127
rect -1 3073 128 3207
rect 27640 3073 27769 3207
rect -1 2193 128 2327
rect 27640 2193 27769 2327
rect -1 1273 128 1407
rect 27640 1273 27769 1407
rect -1 393 128 527
rect 27640 393 27769 527
use M1_NACTIVE_02_512x8m81  M1_NACTIVE_02_512x8m81_0
timestamp 1669390400
transform 1 0 14063 0 1 58559
box 0 0 1 1
use M1_NWELL_01_512x8m81  M1_NWELL_01_512x8m81_0
timestamp 1669390400
transform 1 0 2200 0 1 58486
box -221 -717 1960 228
use M1_NWELL_01_512x8m81  M1_NWELL_01_512x8m81_1
timestamp 1669390400
transform -1 0 25568 0 1 58486
box -221 -717 1960 228
use M1_PACTIVE$10_512x8m81  M1_PACTIVE$10_512x8m81_0
timestamp 1669390400
transform 1 0 11463 0 1 58559
box -78 -80 1817 80
use M1_PACTIVE$10_512x8m81  M1_PACTIVE$10_512x8m81_1
timestamp 1669390400
transform 1 0 4390 0 1 58559
box -78 -80 1817 80
use M1_PACTIVE$10_512x8m81  M1_PACTIVE$10_512x8m81_2
timestamp 1669390400
transform 1 0 21475 0 1 58559
box -78 -80 1817 80
use M1_PACTIVE$11_512x8m81  M1_PACTIVE$11_512x8m81_0
timestamp 1669390400
transform 1 0 15860 0 1 58559
box 0 0 1 1
use M1_POLY2$$204150828_512x8m81  M1_POLY2$$204150828_512x8m81_0
timestamp 1669390400
transform 1 0 9381 0 1 58248
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1669390400
transform 1 0 12040 0 1 58161
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1669390400
transform 0 -1 13712 1 0 58493
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1669390400
transform 1 0 15625 0 1 58201
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1669390400
transform 1 0 18313 0 1 58236
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1669390400
transform 1 0 15413 0 1 58541
box 0 0 1 1
use M2_M1$$201262124_512x8m81  M2_M1$$201262124_512x8m81_0
timestamp 1669390400
transform 1 0 13701 0 1 58491
box 0 0 1 1
use M2_M1$$204138540_512x8m81  M2_M1$$204138540_512x8m81_0
timestamp 1669390400
transform 1 0 10402 0 1 58248
box 0 0 1 1
use M2_M1$$204138540_512x8m81  M2_M1$$204138540_512x8m81_1
timestamp 1669390400
transform 1 0 14059 0 1 58552
box 0 0 1 1
use M2_M1$$204139564_512x8m81  M2_M1$$204139564_512x8m81_0
timestamp 1669390400
transform 1 0 11601 0 1 58505
box 0 0 1 1
use M2_M1$$204140588_512x8m81  M2_M1$$204140588_512x8m81_0
timestamp 1669390400
transform 1 0 12359 0 1 58017
box 0 0 1 1
use M2_M1$$204141612_512x8m81  M2_M1$$204141612_512x8m81_0
timestamp 1669390400
transform 1 0 15126 0 1 58552
box 0 0 1 1
use M2_M1$$204141612_512x8m81  M2_M1$$204141612_512x8m81_1
timestamp 1669390400
transform 1 0 20177 0 1 58480
box 0 0 1 1
use M2_M1$$204141612_512x8m81  M2_M1$$204141612_512x8m81_2
timestamp 1669390400
transform 1 0 20177 0 1 58017
box 0 0 1 1
use M2_M1$$204220460_512x8m81  M2_M1$$204220460_512x8m81_0
timestamp 1669390400
transform 1 0 4399 0 1 58019
box 0 0 1 1
use M2_M1$$204220460_512x8m81  M2_M1$$204220460_512x8m81_1
timestamp 1669390400
transform 1 0 6792 0 1 58480
box 0 0 1 1
use M2_M1$$204220460_512x8m81  M2_M1$$204220460_512x8m81_2
timestamp 1669390400
transform 1 0 6792 0 1 58017
box 0 0 1 1
use M2_M1$$204220460_512x8m81  M2_M1$$204220460_512x8m81_3
timestamp 1669390400
transform 1 0 22430 0 1 58017
box 0 0 1 1
use M2_M1$$204221484_512x8m81  M2_M1$$204221484_512x8m81_0
timestamp 1669390400
transform 1 0 2156 0 1 58500
box -65 -502 1751 67
use M2_M1$$204221484_512x8m81  M2_M1$$204221484_512x8m81_1
timestamp 1669390400
transform -1 0 25612 0 1 58500
box -65 -502 1751 67
use M2_M1$$204222508_512x8m81  M2_M1$$204222508_512x8m81_0
timestamp 1669390400
transform 1 0 5639 0 1 58500
box -65 -284 697 67
use M2_M1$$204222508_512x8m81  M2_M1$$204222508_512x8m81_1
timestamp 1669390400
transform 1 0 21486 0 1 58500
box -65 -284 697 67
use M3_M2$$204142636_512x8m81  M3_M2$$204142636_512x8m81_0
timestamp 1669390400
transform 1 0 5639 0 1 58500
box 0 0 1 1
use M3_M2$$204142636_512x8m81  M3_M2$$204142636_512x8m81_1
timestamp 1669390400
transform 1 0 8250 0 1 58017
box 0 0 1 1
use M3_M2$$204142636_512x8m81  M3_M2$$204142636_512x8m81_2
timestamp 1669390400
transform 1 0 21486 0 1 58500
box 0 0 1 1
use M3_M2$$204142636_512x8m81  M3_M2$$204142636_512x8m81_3
timestamp 1669390400
transform 1 0 21486 0 1 58500
box 0 0 1 1
use M3_M2$$204143660_512x8m81  M3_M2$$204143660_512x8m81_0
timestamp 1669390400
transform 1 0 11601 0 1 58500
box 0 0 1 1
use M3_M2$$204144684_512x8m81  M3_M2$$204144684_512x8m81_0
timestamp 1669390400
transform 1 0 4399 0 1 58019
box 0 0 1 1
use M3_M2$$204144684_512x8m81  M3_M2$$204144684_512x8m81_1
timestamp 1669390400
transform 1 0 22430 0 1 58017
box 0 0 1 1
use M3_M2$$204145708_512x8m81  M3_M2$$204145708_512x8m81_0
timestamp 1669390400
transform 1 0 12359 0 1 58017
box 0 0 1 1
use M3_M2$$204146732_512x8m81  M3_M2$$204146732_512x8m81_0
timestamp 1669390400
transform 1 0 14059 0 1 58010
box 0 0 1 1
use M3_M2$$204147756_512x8m81  M3_M2$$204147756_512x8m81_0
timestamp 1669390400
transform 1 0 12339 0 1 57600
box 0 0 1 1
use nmos_1p2_01_R270_512x8m81  nmos_1p2_01_R270_512x8m81_0
timestamp 1669390400
transform 0 -1 13604 -1 0 58162
box -119 -71 177 1389
use nmos_1p2_02_R90_512x8m81  nmos_1p2_02_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 6346 1 0 58103
box -119 -71 177 2091
use nmos_5p04310591302099_512x8m81  nmos_5p04310591302099_512x8m81_0
timestamp 1669390400
transform 0 -1 23346 1 0 58072
box -88 -44 208 2066
use nmos_5p043105913020111_512x8m81  nmos_5p043105913020111_512x8m81_0
timestamp 1669390400
transform 0 -1 11913 1 0 58072
box -88 -44 208 572
use nmos_5p043105913020111_512x8m81  nmos_5p043105913020111_512x8m81_1
timestamp 1669390400
transform 0 -1 16283 1 0 58072
box -88 -44 208 572
use pmos_1p2_01_R90_512x8m81  pmos_1p2_01_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 11004 1 0 58103
box -295 -137 355 1454
use pmos_1p2_02_R90_512x8m81  pmos_1p2_02_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 9245 1 0 58103
box -296 -137 586 2646
use pmos_1p2_02_R90_512x8m81  pmos_1p2_02_R90_512x8m81_1
timestamp 1669390400
transform 0 -1 20950 1 0 58103
box -296 -137 586 2646
use pmos_5p043105913020101_512x8m81  pmos_5p043105913020101_512x8m81_0
timestamp 1669390400
transform 0 -1 17974 1 0 58072
box -208 -120 328 1438
use pmos_5p043105913020101_512x8m81  pmos_5p043105913020101_512x8m81_1
timestamp 1669390400
transform 0 -1 15304 1 0 58072
box -208 -120 328 1438
use pmoscap_L1_W2_R270_512x8m81  pmoscap_L1_W2_R270_512x8m81_0
timestamp 1669390400
transform 0 -1 2203 -1 0 58650
box -60 -407 1259 3251
use pmoscap_L1_W2_R270_512x8m81  pmoscap_L1_W2_R270_512x8m81_1
timestamp 1669390400
transform 0 1 25566 -1 0 58650
box -60 -407 1259 3251
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_0
timestamp 1669390400
transform 0 1 25566 -1 0 16350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_1
timestamp 1669390400
transform 0 1 25566 -1 0 14550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_2
timestamp 1669390400
transform 0 1 25566 -1 0 12750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_3
timestamp 1669390400
transform 0 1 25566 -1 0 10950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_4
timestamp 1669390400
transform 0 1 25566 -1 0 9150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_5
timestamp 1669390400
transform 0 1 25566 -1 0 7350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_6
timestamp 1669390400
transform 0 1 25566 -1 0 5550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_7
timestamp 1669390400
transform 0 1 25566 -1 0 3750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_8
timestamp 1669390400
transform 0 1 25566 -1 0 1950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_9
timestamp 1669390400
transform 0 1 25566 -1 0 28950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_10
timestamp 1669390400
transform 0 1 25566 -1 0 27150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_11
timestamp 1669390400
transform 0 1 25566 -1 0 25350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_12
timestamp 1669390400
transform 0 1 25566 -1 0 23550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_13
timestamp 1669390400
transform 0 1 25566 -1 0 21750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_14
timestamp 1669390400
transform 0 1 25566 -1 0 19950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_15
timestamp 1669390400
transform 0 1 25566 -1 0 18150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_16
timestamp 1669390400
transform 0 -1 2203 -1 0 16350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_17
timestamp 1669390400
transform 0 -1 2203 -1 0 14550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_18
timestamp 1669390400
transform 0 -1 2203 -1 0 12750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_19
timestamp 1669390400
transform 0 -1 2203 -1 0 10950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_20
timestamp 1669390400
transform 0 -1 2203 -1 0 9150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_21
timestamp 1669390400
transform 0 -1 2203 -1 0 7350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_22
timestamp 1669390400
transform 0 -1 2203 -1 0 5550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_23
timestamp 1669390400
transform 0 -1 2203 -1 0 3750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_24
timestamp 1669390400
transform 0 -1 2203 -1 0 1950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_25
timestamp 1669390400
transform 0 -1 2203 -1 0 28950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_26
timestamp 1669390400
transform 0 -1 2203 -1 0 27150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_27
timestamp 1669390400
transform 0 -1 2203 -1 0 25350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_28
timestamp 1669390400
transform 0 -1 2203 -1 0 23550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_29
timestamp 1669390400
transform 0 -1 2203 -1 0 21750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_30
timestamp 1669390400
transform 0 -1 2203 -1 0 19950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_31
timestamp 1669390400
transform 0 -1 2203 -1 0 18150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_32
timestamp 1669390400
transform 0 -1 2203 -1 0 57750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_33
timestamp 1669390400
transform 0 -1 2203 -1 0 55950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_34
timestamp 1669390400
transform 0 -1 2203 -1 0 54150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_35
timestamp 1669390400
transform 0 -1 2203 -1 0 52350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_36
timestamp 1669390400
transform 0 -1 2203 -1 0 50550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_37
timestamp 1669390400
transform 0 -1 2203 -1 0 48750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_38
timestamp 1669390400
transform 0 -1 2203 -1 0 46950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_39
timestamp 1669390400
transform 0 -1 2203 -1 0 45150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_40
timestamp 1669390400
transform 0 -1 2203 -1 0 43350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_41
timestamp 1669390400
transform 0 -1 2203 -1 0 41550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_42
timestamp 1669390400
transform 0 -1 2203 -1 0 39750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_43
timestamp 1669390400
transform 0 -1 2203 -1 0 37950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_44
timestamp 1669390400
transform 0 -1 2203 -1 0 36150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_45
timestamp 1669390400
transform 0 -1 2203 -1 0 34350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_46
timestamp 1669390400
transform 0 -1 2203 -1 0 32550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_47
timestamp 1669390400
transform 0 1 25566 -1 0 57750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_48
timestamp 1669390400
transform 0 1 25566 -1 0 55950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_49
timestamp 1669390400
transform 0 1 25566 -1 0 54150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_50
timestamp 1669390400
transform 0 1 25566 -1 0 52350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_51
timestamp 1669390400
transform 0 1 25566 -1 0 50550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_52
timestamp 1669390400
transform 0 1 25566 -1 0 48750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_53
timestamp 1669390400
transform 0 1 25566 -1 0 46950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_54
timestamp 1669390400
transform 0 1 25566 -1 0 45150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_55
timestamp 1669390400
transform 0 1 25566 -1 0 43350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_56
timestamp 1669390400
transform 0 1 25566 -1 0 41550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_57
timestamp 1669390400
transform 0 1 25566 -1 0 39750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_58
timestamp 1669390400
transform 0 1 25566 -1 0 37950
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_59
timestamp 1669390400
transform 0 1 25566 -1 0 36150
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_60
timestamp 1669390400
transform 0 1 25566 -1 0 34350
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_61
timestamp 1669390400
transform 0 1 25566 -1 0 32550
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_62
timestamp 1669390400
transform 0 -1 2203 -1 0 30750
box -60 -407 2159 5567
use pmoscap_R270_512x8m81  pmoscap_R270_512x8m81_63
timestamp 1669390400
transform 0 1 25566 -1 0 30750
box -60 -407 2159 5567
use xdec32_468_512x8m81  xdec32_468_512x8m81_0
timestamp 1669390400
transform 1 0 1726 0 1 28800
box 0 -228 24219 29028
use xdec32_512x8m81  xdec32_512x8m81_0
timestamp 1669390400
transform 1 0 1726 0 1 0
box 0 -228 24219 29028
<< labels >>
rlabel metal3 s 27705 58040 27705 58040 4 DRWL
port 1 nsew
rlabel metal3 s 27705 30160 27705 30160 4 RWL[33]
port 2 nsew
rlabel metal3 s 27705 31040 27705 31040 4 RWL[34]
port 3 nsew
rlabel metal3 s 27705 31960 27705 31960 4 RWL[35]
port 4 nsew
rlabel metal3 s 27705 32840 27705 32840 4 RWL[36]
port 5 nsew
rlabel metal3 s 27705 33760 27705 33760 4 RWL[37]
port 6 nsew
rlabel metal3 s 27705 34640 27705 34640 4 RWL[38]
port 7 nsew
rlabel metal3 s 27705 35560 27705 35560 4 RWL[39]
port 8 nsew
rlabel metal3 s 27705 36440 27705 36440 4 RWL[40]
port 9 nsew
rlabel metal3 s 27705 37360 27705 37360 4 RWL[41]
port 10 nsew
rlabel metal3 s 27705 38240 27705 38240 4 RWL[42]
port 11 nsew
rlabel metal3 s 27705 39160 27705 39160 4 RWL[43]
port 12 nsew
rlabel metal3 s 27705 40040 27705 40040 4 RWL[44]
port 13 nsew
rlabel metal3 s 27705 40960 27705 40960 4 RWL[45]
port 14 nsew
rlabel metal3 s 27705 41840 27705 41840 4 RWL[46]
port 15 nsew
rlabel metal3 s 27705 42760 27705 42760 4 RWL[47]
port 16 nsew
rlabel metal3 s 27705 43640 27705 43640 4 RWL[48]
port 17 nsew
rlabel metal3 s 27705 44560 27705 44560 4 RWL[49]
port 18 nsew
rlabel metal3 s 27705 45440 27705 45440 4 RWL[50]
port 19 nsew
rlabel metal3 s 27705 46360 27705 46360 4 RWL[51]
port 20 nsew
rlabel metal3 s 27705 47240 27705 47240 4 RWL[52]
port 21 nsew
rlabel metal3 s 27705 48160 27705 48160 4 RWL[53]
port 22 nsew
rlabel metal3 s 27705 49040 27705 49040 4 RWL[54]
port 23 nsew
rlabel metal3 s 27705 49960 27705 49960 4 RWL[55]
port 24 nsew
rlabel metal3 s 27705 50840 27705 50840 4 RWL[56]
port 25 nsew
rlabel metal3 s 27705 51760 27705 51760 4 RWL[57]
port 26 nsew
rlabel metal3 s 27705 52640 27705 52640 4 RWL[58]
port 27 nsew
rlabel metal3 s 27705 53560 27705 53560 4 RWL[59]
port 28 nsew
rlabel metal3 s 27705 54440 27705 54440 4 RWL[60]
port 29 nsew
rlabel metal3 s 27705 55360 27705 55360 4 RWL[61]
port 30 nsew
rlabel metal3 s 27705 56240 27705 56240 4 RWL[62]
port 31 nsew
rlabel metal3 s 27705 57160 27705 57160 4 RWL[63]
port 32 nsew
rlabel metal3 s 64 57160 64 57160 4 LWL[63]
port 33 nsew
rlabel metal3 s 64 56240 64 56240 4 LWL[62]
port 34 nsew
rlabel metal3 s 64 55360 64 55360 4 LWL[61]
port 35 nsew
rlabel metal3 s 64 54440 64 54440 4 LWL[60]
port 36 nsew
rlabel metal3 s 64 53560 64 53560 4 LWL[59]
port 37 nsew
rlabel metal3 s 64 52640 64 52640 4 LWL[58]
port 38 nsew
rlabel metal3 s 64 51760 64 51760 4 LWL[57]
port 39 nsew
rlabel metal3 s 64 50840 64 50840 4 LWL[56]
port 40 nsew
rlabel metal3 s 64 49960 64 49960 4 LWL[55]
port 41 nsew
rlabel metal3 s 64 49040 64 49040 4 LWL[54]
port 42 nsew
rlabel metal3 s 64 48160 64 48160 4 LWL[53]
port 43 nsew
rlabel metal3 s 64 47240 64 47240 4 LWL[52]
port 44 nsew
rlabel metal3 s 64 46360 64 46360 4 LWL[51]
port 45 nsew
rlabel metal3 s 64 45440 64 45440 4 LWL[50]
port 46 nsew
rlabel metal3 s 64 44560 64 44560 4 LWL[49]
port 47 nsew
rlabel metal3 s 64 43640 64 43640 4 LWL[48]
port 48 nsew
rlabel metal3 s 64 42760 64 42760 4 LWL[47]
port 49 nsew
rlabel metal3 s 64 41840 64 41840 4 LWL[46]
port 50 nsew
rlabel metal3 s 64 40960 64 40960 4 LWL[45]
port 51 nsew
rlabel metal3 s 64 40040 64 40040 4 LWL[44]
port 52 nsew
rlabel metal3 s 64 39160 64 39160 4 LWL[43]
port 53 nsew
rlabel metal3 s 64 38240 64 38240 4 LWL[42]
port 54 nsew
rlabel metal3 s 64 37360 64 37360 4 LWL[41]
port 55 nsew
rlabel metal3 s 64 36440 64 36440 4 LWL[40]
port 56 nsew
rlabel metal3 s 64 35560 64 35560 4 LWL[39]
port 57 nsew
rlabel metal3 s 64 34640 64 34640 4 LWL[38]
port 58 nsew
rlabel metal3 s 64 33760 64 33760 4 LWL[37]
port 59 nsew
rlabel metal3 s 64 32840 64 32840 4 LWL[36]
port 60 nsew
rlabel metal3 s 64 31960 64 31960 4 LWL[35]
port 61 nsew
rlabel metal3 s 64 31040 64 31040 4 LWL[34]
port 62 nsew
rlabel metal3 s 64 30160 64 30160 4 LWL[33]
port 63 nsew
rlabel metal3 s 134 58500 134 58500 4 vss
port 64 nsew
rlabel metal3 s 134 57600 134 57600 4 vdd
port 65 nsew
rlabel metal3 s 64 58040 64 58040 4 DLWL
port 66 nsew
rlabel metal3 s 64 28340 64 28340 4 LWL[31]
port 67 nsew
rlabel metal3 s 64 17540 64 17540 4 LWL[19]
port 68 nsew
rlabel metal3 s 64 18460 64 18460 4 LWL[20]
port 69 nsew
rlabel metal3 s 64 19340 64 19340 4 LWL[21]
port 70 nsew
rlabel metal3 s 64 20260 64 20260 4 LWL[22]
port 71 nsew
rlabel metal3 s 64 21140 64 21140 4 LWL[23]
port 72 nsew
rlabel metal3 s 64 22060 64 22060 4 LWL[24]
port 73 nsew
rlabel metal3 s 64 22940 64 22940 4 LWL[25]
port 74 nsew
rlabel metal3 s 64 23860 64 23860 4 LWL[26]
port 75 nsew
rlabel metal3 s 64 24740 64 24740 4 LWL[27]
port 76 nsew
rlabel metal3 s 64 25660 64 25660 4 LWL[28]
port 77 nsew
rlabel metal3 s 64 9460 64 9460 4 LWL[10]
port 78 nsew
rlabel metal3 s 64 10340 64 10340 4 LWL[11]
port 79 nsew
rlabel metal3 s 64 11260 64 11260 4 LWL[12]
port 80 nsew
rlabel metal3 s 64 12140 64 12140 4 LWL[13]
port 81 nsew
rlabel metal3 s 64 13060 64 13060 4 LWL[14]
port 82 nsew
rlabel metal3 s 64 13940 64 13940 4 LWL[15]
port 83 nsew
rlabel metal3 s 64 14860 64 14860 4 LWL[16]
port 84 nsew
rlabel metal3 s 64 15740 64 15740 4 LWL[17]
port 85 nsew
rlabel metal3 s 64 16660 64 16660 4 LWL[18]
port 86 nsew
rlabel metal3 s 64 4940 64 4940 4 LWL[5]
port 87 nsew
rlabel metal3 s 64 4060 64 4060 4 LWL[4]
port 88 nsew
rlabel metal3 s 64 3140 64 3140 4 LWL[3]
port 89 nsew
rlabel metal3 s 64 2260 64 2260 4 LWL[2]
port 90 nsew
rlabel metal3 s 64 1340 64 1340 4 LWL[1]
port 91 nsew
rlabel metal3 s 64 460 64 460 4 LWL[0]
port 92 nsew
rlabel metal3 s 64 7660 64 7660 4 LWL[8]
port 93 nsew
rlabel metal3 s 64 8540 64 8540 4 LWL[9]
port 94 nsew
rlabel metal3 s 64 5860 64 5860 4 LWL[6]
port 95 nsew
rlabel metal3 s 64 29240 64 29240 4 LWL[32]
port 96 nsew
rlabel metal3 s 64 6740 64 6740 4 LWL[7]
port 97 nsew
rlabel metal3 s 64 26540 64 26540 4 LWL[29]
port 98 nsew
rlabel metal3 s 64 27460 64 27460 4 LWL[30]
port 99 nsew
rlabel metal3 s 27705 29240 27705 29240 4 RWL[32]
port 100 nsew
rlabel metal3 s 27705 28340 27705 28340 4 RWL[31]
port 101 nsew
rlabel metal3 s 27705 27460 27705 27460 4 RWL[30]
port 102 nsew
rlabel metal3 s 27705 26540 27705 26540 4 RWL[29]
port 103 nsew
rlabel metal3 s 27705 25660 27705 25660 4 RWL[28]
port 104 nsew
rlabel metal3 s 27705 24740 27705 24740 4 RWL[27]
port 105 nsew
rlabel metal3 s 27705 23860 27705 23860 4 RWL[26]
port 106 nsew
rlabel metal3 s 27705 22940 27705 22940 4 RWL[25]
port 107 nsew
rlabel metal3 s 27705 22060 27705 22060 4 RWL[24]
port 108 nsew
rlabel metal3 s 27705 21140 27705 21140 4 RWL[23]
port 109 nsew
rlabel metal3 s 27705 20260 27705 20260 4 RWL[22]
port 110 nsew
rlabel metal3 s 27705 19340 27705 19340 4 RWL[21]
port 111 nsew
rlabel metal3 s 27705 5860 27705 5860 4 RWL[6]
port 112 nsew
rlabel metal3 s 27705 4060 27705 4060 4 RWL[4]
port 113 nsew
rlabel metal3 s 27705 2260 27705 2260 4 RWL[2]
port 114 nsew
rlabel metal3 s 27705 460 27705 460 4 RWL[0]
port 115 nsew
rlabel metal3 s 27705 1340 27705 1340 4 RWL[1]
port 116 nsew
rlabel metal3 s 27705 3140 27705 3140 4 RWL[3]
port 117 nsew
rlabel metal3 s 27705 4940 27705 4940 4 RWL[5]
port 118 nsew
rlabel metal3 s 27705 6740 27705 6740 4 RWL[7]
port 119 nsew
rlabel metal3 s 27705 7660 27705 7660 4 RWL[8]
port 120 nsew
rlabel metal3 s 27705 8540 27705 8540 4 RWL[9]
port 121 nsew
rlabel metal3 s 27705 9460 27705 9460 4 RWL[10]
port 122 nsew
rlabel metal3 s 27705 10340 27705 10340 4 RWL[11]
port 123 nsew
rlabel metal3 s 27705 11260 27705 11260 4 RWL[12]
port 124 nsew
rlabel metal3 s 27705 12140 27705 12140 4 RWL[13]
port 125 nsew
rlabel metal3 s 27705 13060 27705 13060 4 RWL[14]
port 126 nsew
rlabel metal3 s 27705 13940 27705 13940 4 RWL[15]
port 127 nsew
rlabel metal3 s 27705 14860 27705 14860 4 RWL[16]
port 128 nsew
rlabel metal3 s 27705 15740 27705 15740 4 RWL[17]
port 129 nsew
rlabel metal3 s 27705 16660 27705 16660 4 RWL[18]
port 130 nsew
rlabel metal3 s 27705 17540 27705 17540 4 RWL[19]
port 131 nsew
rlabel metal3 s 27705 18460 27705 18460 4 RWL[20]
port 132 nsew
rlabel metal2 s 14794 -97 14794 -97 4 xb[0]
port 133 nsew
rlabel metal2 s 14417 -97 14417 -97 4 xb[1]
port 134 nsew
rlabel metal2 s 14039 -97 14039 -97 4 xb[2]
port 135 nsew
rlabel metal2 s 13661 -97 13661 -97 4 xb[3]
port 136 nsew
rlabel metal2 s 16947 -97 16947 -97 4 xa[7]
port 137 nsew
rlabel metal2 s 17324 -97 17324 -97 4 xa[6]
port 138 nsew
rlabel metal2 s 17702 -97 17702 -97 4 xa[5]
port 139 nsew
rlabel metal2 s 18080 -97 18080 -97 4 xa[4]
port 140 nsew
rlabel metal2 s 19591 -97 19591 -97 4 xa[0]
port 141 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 142 nsew
rlabel metal2 s 18457 -97 18457 -97 4 xa[3]
port 143 nsew
rlabel metal2 s 18835 -97 18835 -97 4 xa[2]
port 144 nsew
rlabel metal2 s 19213 -97 19213 -97 4 xa[1]
port 145 nsew
rlabel metal2 s 13284 -97 13284 -97 4 xc[0]
port 146 nsew
rlabel metal2 s 12906 -97 12906 -97 4 xc[1]
port 147 nsew
<< properties >>
string GDS_END 2875380
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2848062
<< end >>
