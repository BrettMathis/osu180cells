magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -2594 353 2594 393
rect -2594 301 -2556 353
rect -2504 301 -2345 353
rect -2293 301 -2134 353
rect -2082 301 -1924 353
rect -1872 301 -1713 353
rect -1661 301 -1502 353
rect -1450 301 -1291 353
rect -1239 301 -1080 353
rect -1028 301 -870 353
rect -818 301 -659 353
rect -607 301 -448 353
rect -396 301 -237 353
rect -185 301 -26 353
rect 26 301 185 353
rect 237 301 396 353
rect 448 301 607 353
rect 659 301 818 353
rect 870 301 1028 353
rect 1080 301 1239 353
rect 1291 301 1450 353
rect 1502 301 1661 353
rect 1713 301 1872 353
rect 1924 301 2082 353
rect 2134 301 2293 353
rect 2345 301 2504 353
rect 2556 301 2594 353
rect -2594 135 2594 301
rect -2594 83 -2556 135
rect -2504 83 -2345 135
rect -2293 83 -2134 135
rect -2082 83 -1924 135
rect -1872 83 -1713 135
rect -1661 83 -1502 135
rect -1450 83 -1291 135
rect -1239 83 -1080 135
rect -1028 83 -870 135
rect -818 83 -659 135
rect -607 83 -448 135
rect -396 83 -237 135
rect -185 83 -26 135
rect 26 83 185 135
rect 237 83 396 135
rect 448 83 607 135
rect 659 83 818 135
rect 870 83 1028 135
rect 1080 83 1239 135
rect 1291 83 1450 135
rect 1502 83 1661 135
rect 1713 83 1872 135
rect 1924 83 2082 135
rect 2134 83 2293 135
rect 2345 83 2504 135
rect 2556 83 2594 135
rect -2594 -83 2594 83
rect -2594 -135 -2556 -83
rect -2504 -135 -2345 -83
rect -2293 -135 -2134 -83
rect -2082 -135 -1924 -83
rect -1872 -135 -1713 -83
rect -1661 -135 -1502 -83
rect -1450 -135 -1291 -83
rect -1239 -135 -1080 -83
rect -1028 -135 -870 -83
rect -818 -135 -659 -83
rect -607 -135 -448 -83
rect -396 -135 -237 -83
rect -185 -135 -26 -83
rect 26 -135 185 -83
rect 237 -135 396 -83
rect 448 -135 607 -83
rect 659 -135 818 -83
rect 870 -135 1028 -83
rect 1080 -135 1239 -83
rect 1291 -135 1450 -83
rect 1502 -135 1661 -83
rect 1713 -135 1872 -83
rect 1924 -135 2082 -83
rect 2134 -135 2293 -83
rect 2345 -135 2504 -83
rect 2556 -135 2594 -83
rect -2594 -301 2594 -135
rect -2594 -353 -2556 -301
rect -2504 -353 -2345 -301
rect -2293 -353 -2134 -301
rect -2082 -353 -1924 -301
rect -1872 -353 -1713 -301
rect -1661 -353 -1502 -301
rect -1450 -353 -1291 -301
rect -1239 -353 -1080 -301
rect -1028 -353 -870 -301
rect -818 -353 -659 -301
rect -607 -353 -448 -301
rect -396 -353 -237 -301
rect -185 -353 -26 -301
rect 26 -353 185 -301
rect 237 -353 396 -301
rect 448 -353 607 -301
rect 659 -353 818 -301
rect 870 -353 1028 -301
rect 1080 -353 1239 -301
rect 1291 -353 1450 -301
rect 1502 -353 1661 -301
rect 1713 -353 1872 -301
rect 1924 -353 2082 -301
rect 2134 -353 2293 -301
rect 2345 -353 2504 -301
rect 2556 -353 2594 -301
rect -2594 -393 2594 -353
<< via1 >>
rect -2556 301 -2504 353
rect -2345 301 -2293 353
rect -2134 301 -2082 353
rect -1924 301 -1872 353
rect -1713 301 -1661 353
rect -1502 301 -1450 353
rect -1291 301 -1239 353
rect -1080 301 -1028 353
rect -870 301 -818 353
rect -659 301 -607 353
rect -448 301 -396 353
rect -237 301 -185 353
rect -26 301 26 353
rect 185 301 237 353
rect 396 301 448 353
rect 607 301 659 353
rect 818 301 870 353
rect 1028 301 1080 353
rect 1239 301 1291 353
rect 1450 301 1502 353
rect 1661 301 1713 353
rect 1872 301 1924 353
rect 2082 301 2134 353
rect 2293 301 2345 353
rect 2504 301 2556 353
rect -2556 83 -2504 135
rect -2345 83 -2293 135
rect -2134 83 -2082 135
rect -1924 83 -1872 135
rect -1713 83 -1661 135
rect -1502 83 -1450 135
rect -1291 83 -1239 135
rect -1080 83 -1028 135
rect -870 83 -818 135
rect -659 83 -607 135
rect -448 83 -396 135
rect -237 83 -185 135
rect -26 83 26 135
rect 185 83 237 135
rect 396 83 448 135
rect 607 83 659 135
rect 818 83 870 135
rect 1028 83 1080 135
rect 1239 83 1291 135
rect 1450 83 1502 135
rect 1661 83 1713 135
rect 1872 83 1924 135
rect 2082 83 2134 135
rect 2293 83 2345 135
rect 2504 83 2556 135
rect -2556 -135 -2504 -83
rect -2345 -135 -2293 -83
rect -2134 -135 -2082 -83
rect -1924 -135 -1872 -83
rect -1713 -135 -1661 -83
rect -1502 -135 -1450 -83
rect -1291 -135 -1239 -83
rect -1080 -135 -1028 -83
rect -870 -135 -818 -83
rect -659 -135 -607 -83
rect -448 -135 -396 -83
rect -237 -135 -185 -83
rect -26 -135 26 -83
rect 185 -135 237 -83
rect 396 -135 448 -83
rect 607 -135 659 -83
rect 818 -135 870 -83
rect 1028 -135 1080 -83
rect 1239 -135 1291 -83
rect 1450 -135 1502 -83
rect 1661 -135 1713 -83
rect 1872 -135 1924 -83
rect 2082 -135 2134 -83
rect 2293 -135 2345 -83
rect 2504 -135 2556 -83
rect -2556 -353 -2504 -301
rect -2345 -353 -2293 -301
rect -2134 -353 -2082 -301
rect -1924 -353 -1872 -301
rect -1713 -353 -1661 -301
rect -1502 -353 -1450 -301
rect -1291 -353 -1239 -301
rect -1080 -353 -1028 -301
rect -870 -353 -818 -301
rect -659 -353 -607 -301
rect -448 -353 -396 -301
rect -237 -353 -185 -301
rect -26 -353 26 -301
rect 185 -353 237 -301
rect 396 -353 448 -301
rect 607 -353 659 -301
rect 818 -353 870 -301
rect 1028 -353 1080 -301
rect 1239 -353 1291 -301
rect 1450 -353 1502 -301
rect 1661 -353 1713 -301
rect 1872 -353 1924 -301
rect 2082 -353 2134 -301
rect 2293 -353 2345 -301
rect 2504 -353 2556 -301
<< metal2 >>
rect -2594 353 2594 393
rect -2594 301 -2556 353
rect -2504 301 -2345 353
rect -2293 301 -2134 353
rect -2082 301 -1924 353
rect -1872 301 -1713 353
rect -1661 301 -1502 353
rect -1450 301 -1291 353
rect -1239 301 -1080 353
rect -1028 301 -870 353
rect -818 301 -659 353
rect -607 301 -448 353
rect -396 301 -237 353
rect -185 301 -26 353
rect 26 301 185 353
rect 237 301 396 353
rect 448 301 607 353
rect 659 301 818 353
rect 870 301 1028 353
rect 1080 301 1239 353
rect 1291 301 1450 353
rect 1502 301 1661 353
rect 1713 301 1872 353
rect 1924 301 2082 353
rect 2134 301 2293 353
rect 2345 301 2504 353
rect 2556 301 2594 353
rect -2594 135 2594 301
rect -2594 83 -2556 135
rect -2504 83 -2345 135
rect -2293 83 -2134 135
rect -2082 83 -1924 135
rect -1872 83 -1713 135
rect -1661 83 -1502 135
rect -1450 83 -1291 135
rect -1239 83 -1080 135
rect -1028 83 -870 135
rect -818 83 -659 135
rect -607 83 -448 135
rect -396 83 -237 135
rect -185 83 -26 135
rect 26 83 185 135
rect 237 83 396 135
rect 448 83 607 135
rect 659 83 818 135
rect 870 83 1028 135
rect 1080 83 1239 135
rect 1291 83 1450 135
rect 1502 83 1661 135
rect 1713 83 1872 135
rect 1924 83 2082 135
rect 2134 83 2293 135
rect 2345 83 2504 135
rect 2556 83 2594 135
rect -2594 -83 2594 83
rect -2594 -135 -2556 -83
rect -2504 -135 -2345 -83
rect -2293 -135 -2134 -83
rect -2082 -135 -1924 -83
rect -1872 -135 -1713 -83
rect -1661 -135 -1502 -83
rect -1450 -135 -1291 -83
rect -1239 -135 -1080 -83
rect -1028 -135 -870 -83
rect -818 -135 -659 -83
rect -607 -135 -448 -83
rect -396 -135 -237 -83
rect -185 -135 -26 -83
rect 26 -135 185 -83
rect 237 -135 396 -83
rect 448 -135 607 -83
rect 659 -135 818 -83
rect 870 -135 1028 -83
rect 1080 -135 1239 -83
rect 1291 -135 1450 -83
rect 1502 -135 1661 -83
rect 1713 -135 1872 -83
rect 1924 -135 2082 -83
rect 2134 -135 2293 -83
rect 2345 -135 2504 -83
rect 2556 -135 2594 -83
rect -2594 -301 2594 -135
rect -2594 -353 -2556 -301
rect -2504 -353 -2345 -301
rect -2293 -353 -2134 -301
rect -2082 -353 -1924 -301
rect -1872 -353 -1713 -301
rect -1661 -353 -1502 -301
rect -1450 -353 -1291 -301
rect -1239 -353 -1080 -301
rect -1028 -353 -870 -301
rect -818 -353 -659 -301
rect -607 -353 -448 -301
rect -396 -353 -237 -301
rect -185 -353 -26 -301
rect 26 -353 185 -301
rect 237 -353 396 -301
rect 448 -353 607 -301
rect 659 -353 818 -301
rect 870 -353 1028 -301
rect 1080 -353 1239 -301
rect 1291 -353 1450 -301
rect 1502 -353 1661 -301
rect 1713 -353 1872 -301
rect 1924 -353 2082 -301
rect 2134 -353 2293 -301
rect 2345 -353 2504 -301
rect 2556 -353 2594 -301
rect -2594 -393 2594 -353
<< properties >>
string GDS_END 709854
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 703322
<< end >>
