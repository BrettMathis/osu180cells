magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 272 88 273
rect -31 -73 88 -1
use nmos_5p04310590878157_256x8m81  nmos_5p04310590878157_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 316
<< properties >>
string GDS_END 406604
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 406354
<< end >>
