magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -236 76 236 81
rect -236 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 236 76
rect -236 14 236 48
rect -236 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 236 14
rect -236 -48 236 -14
rect -236 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 236 -48
rect -236 -81 236 -76
<< via2 >>
rect -231 48 -203 76
rect -169 48 -141 76
rect -107 48 -79 76
rect -45 48 -17 76
rect 17 48 45 76
rect 79 48 107 76
rect 141 48 169 76
rect 203 48 231 76
rect -231 -14 -203 14
rect -169 -14 -141 14
rect -107 -14 -79 14
rect -45 -14 -17 14
rect 17 -14 45 14
rect 79 -14 107 14
rect 141 -14 169 14
rect 203 -14 231 14
rect -231 -76 -203 -48
rect -169 -76 -141 -48
rect -107 -76 -79 -48
rect -45 -76 -17 -48
rect 17 -76 45 -48
rect 79 -76 107 -48
rect 141 -76 169 -48
rect 203 -76 231 -48
<< metal3 >>
rect -236 76 236 81
rect -236 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 236 76
rect -236 14 236 48
rect -236 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 236 14
rect -236 -48 236 -14
rect -236 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 236 -48
rect -236 -81 236 -76
<< properties >>
string GDS_END 660286
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 658618
<< end >>
