magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -1962 135 1962 176
rect -1962 83 -1924 135
rect -1872 83 -1713 135
rect -1661 83 -1502 135
rect -1450 83 -1291 135
rect -1239 83 -1080 135
rect -1028 83 -870 135
rect -818 83 -659 135
rect -607 83 -448 135
rect -396 83 -237 135
rect -185 83 -26 135
rect 26 83 185 135
rect 237 83 396 135
rect 448 83 607 135
rect 659 83 818 135
rect 870 83 1028 135
rect 1080 83 1239 135
rect 1291 83 1450 135
rect 1502 83 1661 135
rect 1713 83 1872 135
rect 1924 83 1962 135
rect -1962 -83 1962 83
rect -1962 -135 -1924 -83
rect -1872 -135 -1713 -83
rect -1661 -135 -1502 -83
rect -1450 -135 -1291 -83
rect -1239 -135 -1080 -83
rect -1028 -135 -870 -83
rect -818 -135 -659 -83
rect -607 -135 -448 -83
rect -396 -135 -237 -83
rect -185 -135 -26 -83
rect 26 -135 185 -83
rect 237 -135 396 -83
rect 448 -135 607 -83
rect 659 -135 818 -83
rect 870 -135 1028 -83
rect 1080 -135 1239 -83
rect 1291 -135 1450 -83
rect 1502 -135 1661 -83
rect 1713 -135 1872 -83
rect 1924 -135 1962 -83
rect -1962 -176 1962 -135
<< via1 >>
rect -1924 83 -1872 135
rect -1713 83 -1661 135
rect -1502 83 -1450 135
rect -1291 83 -1239 135
rect -1080 83 -1028 135
rect -870 83 -818 135
rect -659 83 -607 135
rect -448 83 -396 135
rect -237 83 -185 135
rect -26 83 26 135
rect 185 83 237 135
rect 396 83 448 135
rect 607 83 659 135
rect 818 83 870 135
rect 1028 83 1080 135
rect 1239 83 1291 135
rect 1450 83 1502 135
rect 1661 83 1713 135
rect 1872 83 1924 135
rect -1924 -135 -1872 -83
rect -1713 -135 -1661 -83
rect -1502 -135 -1450 -83
rect -1291 -135 -1239 -83
rect -1080 -135 -1028 -83
rect -870 -135 -818 -83
rect -659 -135 -607 -83
rect -448 -135 -396 -83
rect -237 -135 -185 -83
rect -26 -135 26 -83
rect 185 -135 237 -83
rect 396 -135 448 -83
rect 607 -135 659 -83
rect 818 -135 870 -83
rect 1028 -135 1080 -83
rect 1239 -135 1291 -83
rect 1450 -135 1502 -83
rect 1661 -135 1713 -83
rect 1872 -135 1924 -83
<< metal2 >>
rect -1962 135 1962 176
rect -1962 83 -1924 135
rect -1872 83 -1713 135
rect -1661 83 -1502 135
rect -1450 83 -1291 135
rect -1239 83 -1080 135
rect -1028 83 -870 135
rect -818 83 -659 135
rect -607 83 -448 135
rect -396 83 -237 135
rect -185 83 -26 135
rect 26 83 185 135
rect 237 83 396 135
rect 448 83 607 135
rect 659 83 818 135
rect 870 83 1028 135
rect 1080 83 1239 135
rect 1291 83 1450 135
rect 1502 83 1661 135
rect 1713 83 1872 135
rect 1924 83 1962 135
rect -1962 -83 1962 83
rect -1962 -135 -1924 -83
rect -1872 -135 -1713 -83
rect -1661 -135 -1502 -83
rect -1450 -135 -1291 -83
rect -1239 -135 -1080 -83
rect -1028 -135 -870 -83
rect -818 -135 -659 -83
rect -607 -135 -448 -83
rect -396 -135 -237 -83
rect -185 -135 -26 -83
rect 26 -135 185 -83
rect 237 -135 396 -83
rect 448 -135 607 -83
rect 659 -135 818 -83
rect 870 -135 1028 -83
rect 1080 -135 1239 -83
rect 1291 -135 1450 -83
rect 1502 -135 1661 -83
rect 1713 -135 1872 -83
rect 1924 -135 1962 -83
rect -1962 -175 1962 -135
<< properties >>
string GDS_END 945356
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 942792
<< end >>
