magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -9233 -228 9233 228
<< nsubdiff >>
rect -9090 23 9090 80
rect -9090 -23 -9036 23
rect -8990 -23 -8877 23
rect -8831 -23 -8719 23
rect -8673 -23 -8561 23
rect -8515 -23 -8403 23
rect -8357 -23 -8245 23
rect -8199 -23 -8087 23
rect -8041 -23 -7929 23
rect -7883 -23 -7771 23
rect -7725 -23 -7613 23
rect -7567 -23 -7454 23
rect -7408 -23 -7296 23
rect -7250 -23 -7138 23
rect -7092 -23 -6980 23
rect -6934 -23 -6822 23
rect -6776 -23 -6664 23
rect -6618 -23 -6506 23
rect -6460 -23 -6348 23
rect -6302 -23 -6190 23
rect -6144 -23 -6031 23
rect -5985 -23 -5873 23
rect -5827 -23 -5715 23
rect -5669 -23 -5557 23
rect -5511 -23 -5399 23
rect -5353 -23 -5241 23
rect -5195 -23 -5083 23
rect -5037 -23 -4925 23
rect -4879 -23 -4766 23
rect -4720 -23 -4608 23
rect -4562 -23 -4450 23
rect -4404 -23 -4292 23
rect -4246 -23 -4134 23
rect -4088 -23 -3976 23
rect -3930 -23 -3818 23
rect -3772 -23 -3660 23
rect -3614 -23 -3502 23
rect -3456 -23 -3343 23
rect -3297 -23 -3185 23
rect -3139 -23 -3027 23
rect -2981 -23 -2869 23
rect -2823 -23 -2711 23
rect -2665 -23 -2553 23
rect -2507 -23 -2395 23
rect -2349 -23 -2237 23
rect -2191 -23 -2079 23
rect -2033 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 2033 23
rect 2079 -23 2191 23
rect 2237 -23 2349 23
rect 2395 -23 2507 23
rect 2553 -23 2665 23
rect 2711 -23 2823 23
rect 2869 -23 2981 23
rect 3027 -23 3139 23
rect 3185 -23 3297 23
rect 3343 -23 3456 23
rect 3502 -23 3614 23
rect 3660 -23 3772 23
rect 3818 -23 3930 23
rect 3976 -23 4088 23
rect 4134 -23 4246 23
rect 4292 -23 4404 23
rect 4450 -23 4562 23
rect 4608 -23 4720 23
rect 4766 -23 4879 23
rect 4925 -23 5037 23
rect 5083 -23 5195 23
rect 5241 -23 5353 23
rect 5399 -23 5511 23
rect 5557 -23 5669 23
rect 5715 -23 5827 23
rect 5873 -23 5985 23
rect 6031 -23 6144 23
rect 6190 -23 6302 23
rect 6348 -23 6460 23
rect 6506 -23 6618 23
rect 6664 -23 6776 23
rect 6822 -23 6934 23
rect 6980 -23 7092 23
rect 7138 -23 7250 23
rect 7296 -23 7408 23
rect 7454 -23 7567 23
rect 7613 -23 7725 23
rect 7771 -23 7883 23
rect 7929 -23 8041 23
rect 8087 -23 8199 23
rect 8245 -23 8357 23
rect 8403 -23 8515 23
rect 8561 -23 8673 23
rect 8719 -23 8831 23
rect 8877 -23 8990 23
rect 9036 -23 9090 23
rect -9090 -80 9090 -23
<< nsubdiffcont >>
rect -9036 -23 -8990 23
rect -8877 -23 -8831 23
rect -8719 -23 -8673 23
rect -8561 -23 -8515 23
rect -8403 -23 -8357 23
rect -8245 -23 -8199 23
rect -8087 -23 -8041 23
rect -7929 -23 -7883 23
rect -7771 -23 -7725 23
rect -7613 -23 -7567 23
rect -7454 -23 -7408 23
rect -7296 -23 -7250 23
rect -7138 -23 -7092 23
rect -6980 -23 -6934 23
rect -6822 -23 -6776 23
rect -6664 -23 -6618 23
rect -6506 -23 -6460 23
rect -6348 -23 -6302 23
rect -6190 -23 -6144 23
rect -6031 -23 -5985 23
rect -5873 -23 -5827 23
rect -5715 -23 -5669 23
rect -5557 -23 -5511 23
rect -5399 -23 -5353 23
rect -5241 -23 -5195 23
rect -5083 -23 -5037 23
rect -4925 -23 -4879 23
rect -4766 -23 -4720 23
rect -4608 -23 -4562 23
rect -4450 -23 -4404 23
rect -4292 -23 -4246 23
rect -4134 -23 -4088 23
rect -3976 -23 -3930 23
rect -3818 -23 -3772 23
rect -3660 -23 -3614 23
rect -3502 -23 -3456 23
rect -3343 -23 -3297 23
rect -3185 -23 -3139 23
rect -3027 -23 -2981 23
rect -2869 -23 -2823 23
rect -2711 -23 -2665 23
rect -2553 -23 -2507 23
rect -2395 -23 -2349 23
rect -2237 -23 -2191 23
rect -2079 -23 -2033 23
rect -1920 -23 -1874 23
rect -1762 -23 -1716 23
rect -1604 -23 -1558 23
rect -1446 -23 -1400 23
rect -1288 -23 -1242 23
rect -1130 -23 -1084 23
rect -972 -23 -926 23
rect -814 -23 -768 23
rect -656 -23 -610 23
rect -497 -23 -451 23
rect -339 -23 -293 23
rect -181 -23 -135 23
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect 1242 -23 1288 23
rect 1400 -23 1446 23
rect 1558 -23 1604 23
rect 1716 -23 1762 23
rect 1874 -23 1920 23
rect 2033 -23 2079 23
rect 2191 -23 2237 23
rect 2349 -23 2395 23
rect 2507 -23 2553 23
rect 2665 -23 2711 23
rect 2823 -23 2869 23
rect 2981 -23 3027 23
rect 3139 -23 3185 23
rect 3297 -23 3343 23
rect 3456 -23 3502 23
rect 3614 -23 3660 23
rect 3772 -23 3818 23
rect 3930 -23 3976 23
rect 4088 -23 4134 23
rect 4246 -23 4292 23
rect 4404 -23 4450 23
rect 4562 -23 4608 23
rect 4720 -23 4766 23
rect 4879 -23 4925 23
rect 5037 -23 5083 23
rect 5195 -23 5241 23
rect 5353 -23 5399 23
rect 5511 -23 5557 23
rect 5669 -23 5715 23
rect 5827 -23 5873 23
rect 5985 -23 6031 23
rect 6144 -23 6190 23
rect 6302 -23 6348 23
rect 6460 -23 6506 23
rect 6618 -23 6664 23
rect 6776 -23 6822 23
rect 6934 -23 6980 23
rect 7092 -23 7138 23
rect 7250 -23 7296 23
rect 7408 -23 7454 23
rect 7567 -23 7613 23
rect 7725 -23 7771 23
rect 7883 -23 7929 23
rect 8041 -23 8087 23
rect 8199 -23 8245 23
rect 8357 -23 8403 23
rect 8515 -23 8561 23
rect 8673 -23 8719 23
rect 8831 -23 8877 23
rect 8990 -23 9036 23
<< metal1 >>
rect -9070 23 9070 60
rect -9070 -23 -9036 23
rect -8990 -23 -8877 23
rect -8831 -23 -8719 23
rect -8673 -23 -8561 23
rect -8515 -23 -8403 23
rect -8357 -23 -8245 23
rect -8199 -23 -8087 23
rect -8041 -23 -7929 23
rect -7883 -23 -7771 23
rect -7725 -23 -7613 23
rect -7567 -23 -7454 23
rect -7408 -23 -7296 23
rect -7250 -23 -7138 23
rect -7092 -23 -6980 23
rect -6934 -23 -6822 23
rect -6776 -23 -6664 23
rect -6618 -23 -6506 23
rect -6460 -23 -6348 23
rect -6302 -23 -6190 23
rect -6144 -23 -6031 23
rect -5985 -23 -5873 23
rect -5827 -23 -5715 23
rect -5669 -23 -5557 23
rect -5511 -23 -5399 23
rect -5353 -23 -5241 23
rect -5195 -23 -5083 23
rect -5037 -23 -4925 23
rect -4879 -23 -4766 23
rect -4720 -23 -4608 23
rect -4562 -23 -4450 23
rect -4404 -23 -4292 23
rect -4246 -23 -4134 23
rect -4088 -23 -3976 23
rect -3930 -23 -3818 23
rect -3772 -23 -3660 23
rect -3614 -23 -3502 23
rect -3456 -23 -3343 23
rect -3297 -23 -3185 23
rect -3139 -23 -3027 23
rect -2981 -23 -2869 23
rect -2823 -23 -2711 23
rect -2665 -23 -2553 23
rect -2507 -23 -2395 23
rect -2349 -23 -2237 23
rect -2191 -23 -2079 23
rect -2033 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 2033 23
rect 2079 -23 2191 23
rect 2237 -23 2349 23
rect 2395 -23 2507 23
rect 2553 -23 2665 23
rect 2711 -23 2823 23
rect 2869 -23 2981 23
rect 3027 -23 3139 23
rect 3185 -23 3297 23
rect 3343 -23 3456 23
rect 3502 -23 3614 23
rect 3660 -23 3772 23
rect 3818 -23 3930 23
rect 3976 -23 4088 23
rect 4134 -23 4246 23
rect 4292 -23 4404 23
rect 4450 -23 4562 23
rect 4608 -23 4720 23
rect 4766 -23 4879 23
rect 4925 -23 5037 23
rect 5083 -23 5195 23
rect 5241 -23 5353 23
rect 5399 -23 5511 23
rect 5557 -23 5669 23
rect 5715 -23 5827 23
rect 5873 -23 5985 23
rect 6031 -23 6144 23
rect 6190 -23 6302 23
rect 6348 -23 6460 23
rect 6506 -23 6618 23
rect 6664 -23 6776 23
rect 6822 -23 6934 23
rect 6980 -23 7092 23
rect 7138 -23 7250 23
rect 7296 -23 7408 23
rect 7454 -23 7567 23
rect 7613 -23 7725 23
rect 7771 -23 7883 23
rect 7929 -23 8041 23
rect 8087 -23 8199 23
rect 8245 -23 8357 23
rect 8403 -23 8515 23
rect 8561 -23 8673 23
rect 8719 -23 8831 23
rect 8877 -23 8990 23
rect 9036 -23 9070 23
rect -9070 -60 9070 -23
<< properties >>
string GDS_END 820560
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 812940
<< end >>
