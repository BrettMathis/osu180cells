magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect 0 111 64 123
rect 28 70 35 111
rect 47 76 52 104
rect 45 70 55 76
rect 21 57 31 63
rect 28 12 35 36
rect 45 30 55 36
rect 47 19 52 30
rect 0 0 64 12
<< obsm1 >>
rect 11 49 16 104
rect 11 43 44 49
rect 11 19 16 43
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 9 112 19 118
rect 33 112 43 118
rect 10 111 18 112
rect 34 111 42 112
rect 45 69 55 77
rect 22 63 30 64
rect 21 57 31 63
rect 22 56 30 57
rect 47 37 53 69
rect 45 29 55 37
rect 10 11 18 12
rect 34 11 42 12
rect 9 5 19 11
rect 33 5 43 11
rect 10 4 18 5
rect 34 4 42 5
<< labels >>
rlabel metal2 s 22 56 30 64 6 A
port 1 nsew signal input
rlabel metal2 s 21 57 31 63 6 A
port 1 nsew signal input
rlabel metal1 s 21 57 31 63 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 28 70 35 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 64 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 28 0 35 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 64 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 47 29 53 77 6 Y
port 2 nsew signal output
rlabel metal2 s 45 29 55 37 6 Y
port 2 nsew signal output
rlabel metal2 s 45 69 55 77 6 Y
port 2 nsew signal output
rlabel metal1 s 47 70 52 104 6 Y
port 2 nsew signal output
rlabel metal1 s 45 70 55 76 6 Y
port 2 nsew signal output
rlabel metal1 s 47 19 52 36 6 Y
port 2 nsew signal output
rlabel metal1 s 45 30 55 36 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 64 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 118138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 112986
<< end >>
