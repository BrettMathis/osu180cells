magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 459 3110 1094
rect -86 453 86 459
rect 2662 453 3110 459
<< pwell >>
rect 86 453 2662 459
rect -86 -86 3110 453
<< mvnmos >>
rect 387 267 507 339
rect 125 123 245 195
rect 387 123 507 195
rect 819 260 939 332
rect 1187 260 1307 332
rect 819 116 939 188
rect 1187 116 1307 188
rect 1619 260 1739 332
rect 1987 260 2107 332
rect 1619 116 1739 188
rect 1987 116 2107 188
rect 2420 212 2540 284
rect 2420 68 2540 140
rect 2780 68 2900 332
<< mvpmos >>
rect 125 777 225 849
rect 387 777 487 849
rect 387 633 487 705
rect 819 777 919 849
rect 1187 777 1287 849
rect 819 633 919 705
rect 1187 633 1287 705
rect 1619 777 1719 849
rect 1987 777 2087 849
rect 1619 633 1719 705
rect 1987 633 2087 705
rect 2420 777 2520 849
rect 2420 633 2520 705
rect 2780 573 2880 939
<< mvndiff >>
rect 299 326 387 339
rect 299 280 312 326
rect 358 280 387 326
rect 299 267 387 280
rect 507 267 627 339
rect 567 195 627 267
rect 37 182 125 195
rect 37 136 50 182
rect 96 136 125 182
rect 37 123 125 136
rect 245 182 387 195
rect 245 136 274 182
rect 320 136 387 182
rect 245 123 387 136
rect 507 123 627 195
rect 699 260 819 332
rect 939 319 1027 332
rect 939 273 968 319
rect 1014 273 1027 319
rect 939 260 1027 273
rect 1099 319 1187 332
rect 1099 273 1112 319
rect 1158 273 1187 319
rect 1099 260 1187 273
rect 1307 260 1427 332
rect 699 188 759 260
rect 1367 188 1427 260
rect 699 116 819 188
rect 939 175 1187 188
rect 939 129 968 175
rect 1014 129 1187 175
rect 939 116 1187 129
rect 1307 116 1427 188
rect 1499 260 1619 332
rect 1739 319 1827 332
rect 1739 273 1768 319
rect 1814 273 1827 319
rect 1739 260 1827 273
rect 1899 319 1987 332
rect 1899 273 1912 319
rect 1958 273 1987 319
rect 1899 260 1987 273
rect 2107 260 2227 332
rect 1499 188 1559 260
rect 2167 188 2227 260
rect 1499 116 1619 188
rect 1739 175 1987 188
rect 1739 129 1768 175
rect 1814 129 1987 175
rect 1739 116 1987 129
rect 2107 116 2227 188
rect 2300 212 2420 284
rect 2540 271 2628 284
rect 2540 225 2569 271
rect 2615 225 2628 271
rect 2540 212 2628 225
rect 2300 140 2360 212
rect 2700 140 2780 332
rect 2300 68 2420 140
rect 2540 127 2780 140
rect 2540 81 2569 127
rect 2615 81 2780 127
rect 2540 68 2780 81
rect 2900 319 2988 332
rect 2900 179 2929 319
rect 2975 179 2988 319
rect 2900 68 2988 179
<< mvpdiff >>
rect 2700 849 2780 939
rect 37 836 125 849
rect 37 790 50 836
rect 96 790 125 836
rect 37 777 125 790
rect 225 836 387 849
rect 225 790 254 836
rect 300 790 387 836
rect 225 777 387 790
rect 487 777 607 849
rect 547 705 607 777
rect 299 692 387 705
rect 299 646 312 692
rect 358 646 387 692
rect 299 633 387 646
rect 487 633 607 705
rect 699 777 819 849
rect 919 836 1187 849
rect 919 790 948 836
rect 994 790 1187 836
rect 919 777 1187 790
rect 1287 777 1407 849
rect 699 705 759 777
rect 1347 705 1407 777
rect 699 633 819 705
rect 919 692 1007 705
rect 919 646 948 692
rect 994 646 1007 692
rect 919 633 1007 646
rect 1099 692 1187 705
rect 1099 646 1112 692
rect 1158 646 1187 692
rect 1099 633 1187 646
rect 1287 633 1407 705
rect 1499 777 1619 849
rect 1719 836 1987 849
rect 1719 790 1748 836
rect 1794 790 1987 836
rect 1719 777 1987 790
rect 2087 777 2207 849
rect 1499 705 1559 777
rect 2147 705 2207 777
rect 1499 633 1619 705
rect 1719 692 1807 705
rect 1719 646 1748 692
rect 1794 646 1807 692
rect 1719 633 1807 646
rect 1899 692 1987 705
rect 1899 646 1912 692
rect 1958 646 1987 692
rect 1899 633 1987 646
rect 2087 633 2207 705
rect 2300 777 2420 849
rect 2520 836 2780 849
rect 2520 790 2549 836
rect 2595 790 2780 836
rect 2520 777 2780 790
rect 2300 705 2360 777
rect 2300 633 2420 705
rect 2520 692 2608 705
rect 2520 646 2549 692
rect 2595 646 2608 692
rect 2520 633 2608 646
rect 2700 573 2780 777
rect 2880 861 2968 939
rect 2880 721 2909 861
rect 2955 721 2968 861
rect 2880 573 2968 721
<< mvndiffc >>
rect 312 280 358 326
rect 50 136 96 182
rect 274 136 320 182
rect 968 273 1014 319
rect 1112 273 1158 319
rect 968 129 1014 175
rect 1768 273 1814 319
rect 1912 273 1958 319
rect 1768 129 1814 175
rect 2569 225 2615 271
rect 2569 81 2615 127
rect 2929 179 2975 319
<< mvpdiffc >>
rect 50 790 96 836
rect 254 790 300 836
rect 312 646 358 692
rect 948 790 994 836
rect 948 646 994 692
rect 1112 646 1158 692
rect 1748 790 1794 836
rect 1748 646 1794 692
rect 1912 646 1958 692
rect 2549 790 2595 836
rect 2549 646 2595 692
rect 2909 721 2955 861
<< polysilicon >>
rect 2780 939 2880 983
rect 125 849 225 893
rect 387 849 487 893
rect 819 849 919 893
rect 1187 849 1287 893
rect 1619 849 1719 893
rect 1987 849 2087 893
rect 2420 849 2520 893
rect 125 505 225 777
rect 387 705 487 777
rect 819 705 919 777
rect 1187 705 1287 777
rect 1619 705 1719 777
rect 1987 705 2087 777
rect 2420 705 2520 777
rect 125 365 142 505
rect 188 365 225 505
rect 125 239 225 365
rect 387 589 487 633
rect 387 449 400 589
rect 446 449 487 589
rect 387 383 487 449
rect 819 505 919 633
rect 387 339 507 383
rect 819 365 832 505
rect 878 376 919 505
rect 1187 505 1287 633
rect 878 365 939 376
rect 819 332 939 365
rect 1187 365 1200 505
rect 1246 376 1287 505
rect 1619 505 1719 633
rect 1246 365 1307 376
rect 1187 332 1307 365
rect 1619 365 1632 505
rect 1678 376 1719 505
rect 1987 505 2087 633
rect 1678 365 1739 376
rect 1619 332 1739 365
rect 1987 365 2000 505
rect 2046 376 2087 505
rect 2420 505 2520 633
rect 2046 365 2107 376
rect 1987 332 2107 365
rect 2420 365 2433 505
rect 2479 365 2520 505
rect 125 195 245 239
rect 387 195 507 267
rect 819 188 939 260
rect 1187 188 1307 260
rect 125 79 245 123
rect 387 79 507 123
rect 2420 328 2520 365
rect 2780 505 2880 573
rect 2780 365 2793 505
rect 2839 376 2880 505
rect 2839 365 2900 376
rect 2780 332 2900 365
rect 2420 284 2540 328
rect 1619 188 1739 260
rect 1987 188 2107 260
rect 2420 140 2540 212
rect 819 72 939 116
rect 1187 72 1307 116
rect 1619 72 1739 116
rect 1987 72 2107 116
rect 2420 24 2540 68
rect 2780 24 2900 68
<< polycontact >>
rect 142 365 188 505
rect 400 449 446 589
rect 832 365 878 505
rect 1200 365 1246 505
rect 1632 365 1678 505
rect 2000 365 2046 505
rect 2433 365 2479 505
rect 2793 365 2839 505
<< metal1 >>
rect 0 918 3024 1098
rect 39 836 96 847
rect 39 790 50 836
rect 39 608 96 790
rect 254 836 300 918
rect 254 779 300 790
rect 948 836 994 918
rect 948 779 994 790
rect 1748 836 1794 918
rect 1748 779 1794 790
rect 2549 836 2595 918
rect 2549 779 2595 790
rect 2909 861 2994 872
rect 2955 721 2994 861
rect 948 692 994 703
rect 301 646 312 692
rect 358 646 538 692
rect 39 600 275 608
rect 39 589 446 600
rect 39 562 400 589
rect 39 182 85 562
rect 249 554 400 562
rect 142 505 194 516
rect 188 365 194 505
rect 400 438 446 449
rect 142 354 194 365
rect 492 326 538 646
rect 948 516 994 646
rect 1112 692 1158 703
rect 1112 608 1158 646
rect 1748 692 1794 703
rect 1112 562 1338 608
rect 832 505 878 516
rect 832 326 878 365
rect 301 280 312 326
rect 358 280 878 326
rect 948 505 1246 516
rect 948 470 1200 505
rect 948 319 1014 470
rect 1200 354 1246 365
rect 948 273 968 319
rect 948 262 1014 273
rect 1101 273 1112 319
rect 1158 308 1169 319
rect 1292 308 1338 562
rect 1748 516 1794 646
rect 1912 692 1958 703
rect 1912 608 1958 646
rect 2549 692 2595 703
rect 1912 562 2138 608
rect 1632 505 1678 516
rect 1632 308 1678 365
rect 1158 273 1678 308
rect 1101 262 1678 273
rect 1748 505 2046 516
rect 1748 470 2000 505
rect 1748 319 1814 470
rect 2000 354 2046 365
rect 1748 273 1768 319
rect 1748 262 1814 273
rect 1901 273 1912 319
rect 1958 308 1969 319
rect 2092 308 2138 562
rect 2433 505 2479 516
rect 2433 308 2479 365
rect 1958 273 2479 308
rect 1901 262 2479 273
rect 2549 400 2595 646
rect 2793 505 2839 516
rect 2549 365 2793 400
rect 2549 354 2839 365
rect 2549 271 2615 354
rect 2549 225 2569 271
rect 2549 214 2615 225
rect 2909 319 2994 721
rect 274 182 320 193
rect 39 136 50 182
rect 96 136 107 182
rect 274 90 320 136
rect 968 175 1014 186
rect 968 90 1014 129
rect 1768 175 1814 186
rect 2909 179 2929 319
rect 2975 179 2994 319
rect 2909 168 2994 179
rect 1768 90 1814 129
rect 2569 127 2615 138
rect 0 81 2569 90
rect 2615 81 3024 90
rect 0 -90 3024 81
<< labels >>
flabel metal1 s 142 354 194 516 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 3024 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 274 186 320 193 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2909 168 2994 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
rlabel metal1 s 2549 779 2595 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1748 779 1794 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 948 779 994 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 254 779 300 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1768 138 1814 186 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 968 138 1014 186 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 274 138 320 186 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2569 90 2615 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1768 90 1814 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 968 90 1014 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 274 90 320 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3024 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3024 1008
string GDS_END 733646
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 726824
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
