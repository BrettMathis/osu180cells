magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 25 1908 657 2540
rect 1274 1908 1906 2540
rect 25 1008 657 1640
rect 1274 1008 1906 1640
<< mvnsubdiff >>
rect 73 2479 609 2492
rect 73 2433 86 2479
rect 132 2433 202 2479
rect 248 2433 318 2479
rect 364 2433 434 2479
rect 480 2433 550 2479
rect 596 2433 609 2479
rect 73 2420 609 2433
rect 73 2363 145 2420
rect 73 2317 86 2363
rect 132 2317 145 2363
rect 537 2363 609 2420
rect 73 2247 145 2317
rect 73 2201 86 2247
rect 132 2201 145 2247
rect 73 2131 145 2201
rect 73 2085 86 2131
rect 132 2085 145 2131
rect 537 2317 550 2363
rect 596 2317 609 2363
rect 537 2247 609 2317
rect 537 2201 550 2247
rect 596 2201 609 2247
rect 537 2131 609 2201
rect 73 2028 145 2085
rect 537 2085 550 2131
rect 596 2085 609 2131
rect 537 2028 609 2085
rect 73 2015 609 2028
rect 73 1969 86 2015
rect 132 1969 202 2015
rect 248 1969 318 2015
rect 364 1969 434 2015
rect 480 1969 550 2015
rect 596 1969 609 2015
rect 73 1956 609 1969
rect 1322 2479 1858 2492
rect 1322 2433 1335 2479
rect 1381 2433 1451 2479
rect 1497 2433 1567 2479
rect 1613 2433 1683 2479
rect 1729 2433 1799 2479
rect 1845 2433 1858 2479
rect 1322 2420 1858 2433
rect 1322 2363 1394 2420
rect 1322 2317 1335 2363
rect 1381 2317 1394 2363
rect 1786 2363 1858 2420
rect 1322 2247 1394 2317
rect 1322 2201 1335 2247
rect 1381 2201 1394 2247
rect 1322 2131 1394 2201
rect 1322 2085 1335 2131
rect 1381 2085 1394 2131
rect 1786 2317 1799 2363
rect 1845 2317 1858 2363
rect 1786 2247 1858 2317
rect 1786 2201 1799 2247
rect 1845 2201 1858 2247
rect 1786 2131 1858 2201
rect 1322 2028 1394 2085
rect 1786 2085 1799 2131
rect 1845 2085 1858 2131
rect 1786 2028 1858 2085
rect 1322 2015 1858 2028
rect 1322 1969 1335 2015
rect 1381 1969 1451 2015
rect 1497 1969 1567 2015
rect 1613 1969 1683 2015
rect 1729 1969 1799 2015
rect 1845 1969 1858 2015
rect 1322 1956 1858 1969
rect 73 1579 609 1592
rect 73 1533 86 1579
rect 132 1533 202 1579
rect 248 1533 318 1579
rect 364 1533 434 1579
rect 480 1533 550 1579
rect 596 1533 609 1579
rect 73 1520 609 1533
rect 73 1463 145 1520
rect 73 1417 86 1463
rect 132 1417 145 1463
rect 537 1463 609 1520
rect 73 1347 145 1417
rect 73 1301 86 1347
rect 132 1301 145 1347
rect 73 1231 145 1301
rect 73 1185 86 1231
rect 132 1185 145 1231
rect 537 1417 550 1463
rect 596 1417 609 1463
rect 537 1347 609 1417
rect 537 1301 550 1347
rect 596 1301 609 1347
rect 537 1231 609 1301
rect 73 1128 145 1185
rect 537 1185 550 1231
rect 596 1185 609 1231
rect 537 1128 609 1185
rect 73 1115 609 1128
rect 73 1069 86 1115
rect 132 1069 202 1115
rect 248 1069 318 1115
rect 364 1069 434 1115
rect 480 1069 550 1115
rect 596 1069 609 1115
rect 73 1056 609 1069
rect 1322 1579 1858 1592
rect 1322 1533 1335 1579
rect 1381 1533 1451 1579
rect 1497 1533 1567 1579
rect 1613 1533 1683 1579
rect 1729 1533 1799 1579
rect 1845 1533 1858 1579
rect 1322 1520 1858 1533
rect 1322 1463 1394 1520
rect 1322 1417 1335 1463
rect 1381 1417 1394 1463
rect 1786 1463 1858 1520
rect 1322 1347 1394 1417
rect 1322 1301 1335 1347
rect 1381 1301 1394 1347
rect 1322 1231 1394 1301
rect 1322 1185 1335 1231
rect 1381 1185 1394 1231
rect 1786 1417 1799 1463
rect 1845 1417 1858 1463
rect 1786 1347 1858 1417
rect 1786 1301 1799 1347
rect 1845 1301 1858 1347
rect 1786 1231 1858 1301
rect 1322 1128 1394 1185
rect 1786 1185 1799 1231
rect 1845 1185 1858 1231
rect 1786 1128 1858 1185
rect 1322 1115 1858 1128
rect 1322 1069 1335 1115
rect 1381 1069 1451 1115
rect 1497 1069 1567 1115
rect 1613 1069 1683 1115
rect 1729 1069 1799 1115
rect 1845 1069 1858 1115
rect 1322 1056 1858 1069
<< mvnsubdiffcont >>
rect 86 2433 132 2479
rect 202 2433 248 2479
rect 318 2433 364 2479
rect 434 2433 480 2479
rect 550 2433 596 2479
rect 86 2317 132 2363
rect 86 2201 132 2247
rect 86 2085 132 2131
rect 550 2317 596 2363
rect 550 2201 596 2247
rect 550 2085 596 2131
rect 86 1969 132 2015
rect 202 1969 248 2015
rect 318 1969 364 2015
rect 434 1969 480 2015
rect 550 1969 596 2015
rect 1335 2433 1381 2479
rect 1451 2433 1497 2479
rect 1567 2433 1613 2479
rect 1683 2433 1729 2479
rect 1799 2433 1845 2479
rect 1335 2317 1381 2363
rect 1335 2201 1381 2247
rect 1335 2085 1381 2131
rect 1799 2317 1845 2363
rect 1799 2201 1845 2247
rect 1799 2085 1845 2131
rect 1335 1969 1381 2015
rect 1451 1969 1497 2015
rect 1567 1969 1613 2015
rect 1683 1969 1729 2015
rect 1799 1969 1845 2015
rect 86 1533 132 1579
rect 202 1533 248 1579
rect 318 1533 364 1579
rect 434 1533 480 1579
rect 550 1533 596 1579
rect 86 1417 132 1463
rect 86 1301 132 1347
rect 86 1185 132 1231
rect 550 1417 596 1463
rect 550 1301 596 1347
rect 550 1185 596 1231
rect 86 1069 132 1115
rect 202 1069 248 1115
rect 318 1069 364 1115
rect 434 1069 480 1115
rect 550 1069 596 1115
rect 1335 1533 1381 1579
rect 1451 1533 1497 1579
rect 1567 1533 1613 1579
rect 1683 1533 1729 1579
rect 1799 1533 1845 1579
rect 1335 1417 1381 1463
rect 1335 1301 1381 1347
rect 1335 1185 1381 1231
rect 1799 1417 1845 1463
rect 1799 1301 1845 1347
rect 1799 1185 1845 1231
rect 1335 1069 1381 1115
rect 1451 1069 1497 1115
rect 1567 1069 1613 1115
rect 1683 1069 1729 1115
rect 1799 1069 1845 1115
<< mvpdiode >>
rect 241 2311 441 2324
rect 241 2265 254 2311
rect 300 2265 382 2311
rect 428 2265 441 2311
rect 241 2183 441 2265
rect 241 2137 254 2183
rect 300 2137 382 2183
rect 428 2137 441 2183
rect 241 2124 441 2137
rect 1490 2311 1690 2324
rect 1490 2265 1503 2311
rect 1549 2265 1631 2311
rect 1677 2265 1690 2311
rect 1490 2183 1690 2265
rect 1490 2137 1503 2183
rect 1549 2137 1631 2183
rect 1677 2137 1690 2183
rect 1490 2124 1690 2137
rect 241 1411 441 1424
rect 241 1365 254 1411
rect 300 1365 382 1411
rect 428 1365 441 1411
rect 241 1283 441 1365
rect 241 1237 254 1283
rect 300 1237 382 1283
rect 428 1237 441 1283
rect 241 1224 441 1237
rect 1490 1411 1690 1424
rect 1490 1365 1503 1411
rect 1549 1365 1631 1411
rect 1677 1365 1690 1411
rect 1490 1283 1690 1365
rect 1490 1237 1503 1283
rect 1549 1237 1631 1283
rect 1677 1237 1690 1283
rect 1490 1224 1690 1237
<< mvpdiodec >>
rect 254 2265 300 2311
rect 382 2265 428 2311
rect 254 2137 300 2183
rect 382 2137 428 2183
rect 1503 2265 1549 2311
rect 1631 2265 1677 2311
rect 1503 2137 1549 2183
rect 1631 2137 1677 2183
rect 254 1365 300 1411
rect 382 1365 428 1411
rect 254 1237 300 1283
rect 382 1237 428 1283
rect 1503 1365 1549 1411
rect 1631 1365 1677 1411
rect 1503 1237 1549 1283
rect 1631 1237 1677 1283
<< metal1 >>
rect 11094 10853 11274 10865
rect 11094 10801 11106 10853
rect 11262 10801 11274 10853
rect 11094 10789 11274 10801
rect 12354 10691 13432 10703
rect 12354 10602 13368 10691
rect 13356 10535 13368 10602
rect 13420 10535 13432 10691
rect 13356 10523 13432 10535
rect 12164 9812 12240 9824
rect 12164 9656 12176 9812
rect 12228 9656 12240 9812
rect 12164 9644 12240 9656
rect 10095 7859 10347 7871
rect 10095 7703 10107 7859
rect 10159 7703 10347 7859
rect 10095 7691 10347 7703
rect 10275 7369 10351 7381
rect 10275 7213 10287 7369
rect 10339 7213 10351 7369
rect 10275 7201 10351 7213
rect 12136 6514 12316 6526
rect 12136 6462 12148 6514
rect 12304 6462 12316 6514
rect 12136 6450 12316 6462
rect 12736 6381 13432 6393
rect 9570 6301 10171 6313
rect 9570 6249 9582 6301
rect 9738 6249 10003 6301
rect 10159 6249 10171 6301
rect 9570 6237 10171 6249
rect 12736 6225 12748 6381
rect 12800 6306 13368 6381
rect 12800 6225 12812 6306
rect 12736 6213 12812 6225
rect 13356 6225 13368 6306
rect 13420 6225 13432 6381
rect 13356 6213 13432 6225
rect 9726 6165 10351 6177
rect 9726 6113 9738 6165
rect 9894 6113 10183 6165
rect 10339 6113 10351 6165
rect 9726 6101 10351 6113
rect 8310 5571 8815 5639
rect 10027 5362 10103 5374
rect 10027 4894 10039 5362
rect 10091 4894 10103 5362
rect 10027 4882 10103 4894
rect 13168 5362 13452 5374
rect 13168 4894 13388 5362
rect 13440 4894 13452 5362
rect 13168 4882 13452 4894
rect 7991 4446 9118 4522
rect 13356 4458 13432 4470
rect 13356 4439 13368 4458
rect 12910 4326 13368 4439
rect 13356 4302 13368 4326
rect 13420 4302 13432 4458
rect 13356 4290 13432 4302
rect 6820 4270 7000 4278
rect 6733 4266 7000 4270
rect 6733 4214 6832 4266
rect 6988 4214 7000 4266
rect 6733 4202 7000 4214
rect 10027 4176 10103 4188
rect 10027 3708 10039 4176
rect 10091 3708 10103 4176
rect 10027 3696 10103 3708
rect 2969 3347 3149 3359
rect 2969 3295 2981 3347
rect 3137 3295 3149 3347
rect 2969 3283 3149 3295
rect 7841 3169 9118 3245
rect 12136 3225 12316 3237
rect 12136 3173 12148 3225
rect 12304 3173 12316 3225
rect 12136 3161 12316 3173
rect 377 3137 453 3149
rect 377 2981 389 3137
rect 441 3045 453 3137
rect 441 3033 12754 3045
rect 441 2981 12549 3033
rect 12705 2981 12754 3033
rect 377 2969 12754 2981
rect 3171 2896 6287 2908
rect 3171 2844 3183 2896
rect 3339 2844 6119 2896
rect 6275 2844 6287 2896
rect 3171 2832 6287 2844
rect 8058 2897 10072 2909
rect 8058 2845 8070 2897
rect 8226 2845 9904 2897
rect 10060 2845 10072 2897
rect 8058 2833 10072 2845
rect 11457 2782 12859 2794
rect 1784 2761 9490 2773
rect 1784 2709 1796 2761
rect 1952 2709 9426 2761
rect 1784 2697 9426 2709
rect -144 2625 7619 2637
rect -144 2573 -132 2625
rect 24 2573 7451 2625
rect 7607 2573 7619 2625
rect 9414 2605 9426 2697
rect 9478 2605 9490 2761
rect 9726 2761 10142 2773
rect 9414 2593 9490 2605
rect 9570 2729 9646 2741
rect -144 2561 7619 2573
rect 9570 2573 9582 2729
rect 9634 2637 9646 2729
rect 9726 2709 9738 2761
rect 9894 2709 9974 2761
rect 10130 2709 10142 2761
rect 11457 2730 11469 2782
rect 11625 2730 12691 2782
rect 12847 2730 12859 2782
rect 11457 2718 12859 2730
rect 9726 2697 10142 2709
rect 9634 2625 11482 2637
rect 9634 2573 11314 2625
rect 11470 2573 11482 2625
rect 9570 2561 11482 2573
rect 73 2479 609 2492
rect 73 2433 86 2479
rect 132 2433 202 2479
rect 248 2433 318 2479
rect 364 2433 434 2479
rect 480 2433 550 2479
rect 596 2433 609 2479
rect 73 2420 609 2433
rect 73 2363 145 2420
rect 73 2317 86 2363
rect 132 2317 145 2363
rect 537 2363 609 2420
rect 73 2247 145 2317
rect 73 2201 86 2247
rect 132 2201 145 2247
rect 73 2131 145 2201
rect 73 2085 86 2131
rect 132 2085 145 2131
rect 241 2311 441 2324
rect 241 2265 254 2311
rect 300 2265 382 2311
rect 428 2265 441 2311
rect 241 2250 441 2265
rect 241 2198 262 2250
rect 418 2198 441 2250
rect 241 2183 441 2198
rect 241 2137 254 2183
rect 300 2137 382 2183
rect 428 2137 441 2183
rect 241 2124 441 2137
rect 537 2317 550 2363
rect 596 2317 609 2363
rect 537 2247 609 2317
rect 537 2201 550 2247
rect 596 2201 609 2247
rect 537 2131 609 2201
rect 73 2028 145 2085
rect 537 2085 550 2131
rect 596 2085 609 2131
rect 537 2028 609 2085
rect 73 2015 609 2028
rect 73 1969 86 2015
rect 132 1969 202 2015
rect 248 1969 318 2015
rect 364 1969 434 2015
rect 480 1969 550 2015
rect 596 1969 609 2015
rect 73 1956 609 1969
rect 1322 2479 1858 2492
rect 1322 2433 1335 2479
rect 1381 2433 1451 2479
rect 1497 2433 1567 2479
rect 1613 2433 1683 2479
rect 1729 2433 1799 2479
rect 1845 2433 1858 2479
rect 1322 2420 1858 2433
rect 1322 2363 1394 2420
rect 1322 2317 1335 2363
rect 1381 2317 1394 2363
rect 1786 2363 1858 2420
rect 1322 2247 1394 2317
rect 1322 2201 1335 2247
rect 1381 2201 1394 2247
rect 1322 2131 1394 2201
rect 1322 2085 1335 2131
rect 1381 2085 1394 2131
rect 1490 2311 1690 2324
rect 1490 2265 1503 2311
rect 1549 2265 1631 2311
rect 1677 2265 1690 2311
rect 1490 2250 1690 2265
rect 1490 2198 1511 2250
rect 1667 2198 1690 2250
rect 1490 2183 1690 2198
rect 1490 2137 1503 2183
rect 1549 2137 1631 2183
rect 1677 2137 1690 2183
rect 1490 2124 1690 2137
rect 1786 2317 1799 2363
rect 1845 2317 1858 2363
rect 1786 2247 1858 2317
rect 1786 2201 1799 2247
rect 1845 2201 1858 2247
rect 1786 2131 1858 2201
rect 1322 2028 1394 2085
rect 1786 2085 1799 2131
rect 1845 2085 1858 2131
rect 1786 2028 1858 2085
rect 1322 2015 1858 2028
rect 1322 1969 1335 2015
rect 1381 1969 1451 2015
rect 1497 1969 1567 2015
rect 1613 1969 1683 2015
rect 1729 1969 1799 2015
rect 1845 1969 1858 2015
rect 1322 1956 1858 1969
rect 4334 2126 4410 2138
rect 4334 1970 4346 2126
rect 4398 1970 4410 2126
rect 4334 1958 4410 1970
rect 6162 2126 6238 2138
rect 6162 1970 6174 2126
rect 6226 1970 6238 2126
rect 6162 1958 6238 1970
rect 10066 2126 10142 2138
rect 10066 1970 10078 2126
rect 10130 1970 10142 2126
rect 10066 1958 10142 1970
rect 11406 2126 11482 2138
rect 11406 1970 11418 2126
rect 11470 1970 11482 2126
rect 11406 1958 11482 1970
rect 73 1592 1858 1956
rect 73 1579 609 1592
rect 73 1533 86 1579
rect 132 1533 202 1579
rect 248 1533 318 1579
rect 364 1533 434 1579
rect 480 1533 550 1579
rect 596 1533 609 1579
rect 73 1520 609 1533
rect 73 1463 145 1520
rect 73 1417 86 1463
rect 132 1417 145 1463
rect 537 1463 609 1520
rect 73 1347 145 1417
rect 73 1301 86 1347
rect 132 1301 145 1347
rect 73 1231 145 1301
rect 73 1185 86 1231
rect 132 1185 145 1231
rect 241 1411 441 1424
rect 241 1403 254 1411
rect 300 1403 382 1411
rect 241 1247 253 1403
rect 305 1365 382 1403
rect 428 1365 441 1411
rect 305 1283 441 1365
rect 305 1247 382 1283
rect 241 1237 254 1247
rect 300 1237 382 1247
rect 428 1237 441 1283
rect 241 1224 441 1237
rect 537 1417 550 1463
rect 596 1417 609 1463
rect 537 1347 609 1417
rect 537 1301 550 1347
rect 596 1301 609 1347
rect 537 1231 609 1301
rect 73 1128 145 1185
rect 537 1185 550 1231
rect 596 1185 609 1231
rect 537 1128 609 1185
rect 73 1115 609 1128
rect 73 1069 86 1115
rect 132 1069 202 1115
rect 248 1069 318 1115
rect 364 1069 434 1115
rect 480 1069 550 1115
rect 596 1069 609 1115
rect 73 1056 609 1069
rect 1322 1579 1858 1592
rect 1322 1533 1335 1579
rect 1381 1533 1451 1579
rect 1497 1533 1567 1579
rect 1613 1533 1683 1579
rect 1729 1533 1799 1579
rect 1845 1533 1858 1579
rect 1322 1520 1858 1533
rect 1322 1463 1394 1520
rect 1322 1417 1335 1463
rect 1381 1417 1394 1463
rect 1786 1463 1858 1520
rect 1322 1347 1394 1417
rect 1322 1301 1335 1347
rect 1381 1301 1394 1347
rect 1322 1231 1394 1301
rect 1322 1185 1335 1231
rect 1381 1185 1394 1231
rect 1490 1411 1690 1424
rect 1490 1365 1503 1411
rect 1549 1365 1631 1411
rect 1677 1365 1690 1411
rect 1490 1350 1690 1365
rect 1490 1298 1511 1350
rect 1667 1298 1690 1350
rect 1490 1283 1690 1298
rect 1490 1237 1503 1283
rect 1549 1237 1631 1283
rect 1677 1237 1690 1283
rect 1490 1224 1690 1237
rect 1786 1417 1799 1463
rect 1845 1417 1858 1463
rect 1786 1347 1858 1417
rect 1786 1301 1799 1347
rect 1845 1301 1858 1347
rect 2953 1473 3029 1485
rect 2953 1317 2965 1473
rect 3017 1317 3029 1473
rect 2953 1305 3029 1317
rect 7543 1473 7619 1485
rect 7543 1317 7555 1473
rect 7607 1317 7619 1473
rect 7543 1305 7619 1317
rect 8162 1473 8238 1485
rect 8162 1317 8174 1473
rect 8226 1317 8238 1473
rect 8162 1305 8238 1317
rect 12783 1473 12859 1485
rect 12783 1317 12795 1473
rect 12847 1317 12859 1473
rect 12783 1305 12859 1317
rect 1786 1231 1858 1301
rect 1322 1128 1394 1185
rect 1786 1185 1799 1231
rect 1845 1185 1858 1231
rect 1786 1128 1858 1185
rect 1322 1115 1858 1128
rect 1322 1069 1335 1115
rect 1381 1069 1451 1115
rect 1497 1069 1567 1115
rect 1613 1069 1683 1115
rect 1729 1069 1799 1115
rect 1845 1069 1858 1115
rect 1322 1056 1858 1069
rect 73 683 2698 1056
<< via1 >>
rect 11106 10801 11262 10853
rect 13368 10535 13420 10691
rect 12176 9656 12228 9812
rect 10107 7703 10159 7859
rect 10287 7213 10339 7369
rect 12148 6462 12304 6514
rect 9582 6249 9738 6301
rect 10003 6249 10159 6301
rect 12748 6225 12800 6381
rect 13368 6225 13420 6381
rect 9738 6113 9894 6165
rect 10183 6113 10339 6165
rect 10039 4894 10091 5362
rect 13388 4894 13440 5362
rect 13368 4302 13420 4458
rect 6832 4214 6988 4266
rect 10039 3708 10091 4176
rect 2981 3295 3137 3347
rect 12148 3173 12304 3225
rect 389 2981 441 3137
rect 12549 2981 12705 3033
rect 3183 2844 3339 2896
rect 6119 2844 6275 2896
rect 8070 2845 8226 2897
rect 9904 2845 10060 2897
rect 1796 2709 1952 2761
rect -132 2573 24 2625
rect 7451 2573 7607 2625
rect 9426 2605 9478 2761
rect 9582 2573 9634 2729
rect 9738 2709 9894 2761
rect 9974 2709 10130 2761
rect 11469 2730 11625 2782
rect 12691 2730 12847 2782
rect 11314 2573 11470 2625
rect 262 2198 418 2250
rect 1511 2198 1667 2250
rect 4346 1970 4398 2126
rect 6174 1970 6226 2126
rect 10078 1970 10130 2126
rect 11418 1970 11470 2126
rect 253 1365 254 1403
rect 254 1365 300 1403
rect 300 1365 305 1403
rect 253 1283 305 1365
rect 253 1247 254 1283
rect 254 1247 300 1283
rect 300 1247 305 1283
rect 1511 1298 1667 1350
rect 2965 1317 3017 1473
rect 7555 1317 7607 1473
rect 8174 1317 8226 1473
rect 12795 1317 12847 1473
<< metal2 >>
rect 11094 10853 11321 10865
rect 11094 10801 11106 10853
rect 11262 10801 11321 10853
rect 11094 10789 11321 10801
rect 9906 9171 10977 9247
rect 9906 7712 9982 9171
rect 9414 7636 9982 7712
rect 10095 7859 10171 7871
rect 10095 7703 10107 7859
rect 10159 7703 10171 7859
rect 6579 5511 6779 6291
rect 6579 5351 7000 5511
rect 6820 4266 7000 4278
rect 6820 4214 6832 4266
rect 6988 4214 7000 4266
rect 6820 4202 7000 4214
rect 377 3137 453 3149
rect 377 2981 389 3137
rect 441 2981 453 3137
rect 2295 3129 2371 4152
rect 2969 3348 3149 3359
rect 2969 3347 3640 3348
rect 2969 3295 2981 3347
rect 3137 3295 3640 3347
rect 2969 3272 3640 3295
rect 2295 3053 3237 3129
rect -144 2625 36 2637
rect -144 2573 -132 2625
rect 24 2573 36 2625
rect -144 2561 36 2573
rect -144 1415 -68 2561
rect 377 2262 453 2981
rect 3161 2908 3237 3053
rect 3161 2896 3351 2908
rect 3161 2844 3183 2896
rect 3339 2844 3351 2896
rect 3161 2832 3351 2844
rect 1784 2761 1964 2773
rect 1784 2709 1796 2761
rect 1952 2709 1964 2761
rect 1784 2697 1964 2709
rect 1784 2262 1860 2697
rect 250 2250 453 2262
rect 250 2198 262 2250
rect 418 2198 453 2250
rect 250 2186 453 2198
rect 1499 2250 1860 2262
rect 1499 2198 1511 2250
rect 1667 2198 1860 2250
rect 1499 2186 1860 2198
rect -144 1403 317 1415
rect -144 1247 253 1403
rect 305 1247 317 1403
rect -144 1235 317 1247
rect -144 422 -68 1235
rect 377 422 453 2186
rect 3564 1571 3640 3272
rect 6107 2896 6287 2908
rect 6107 2844 6119 2896
rect 6275 2844 6287 2896
rect 6107 2832 6287 2844
rect 8058 2897 8238 2909
rect 8058 2845 8070 2897
rect 8226 2845 8238 2897
rect 8058 2833 8238 2845
rect 4334 2126 4410 2138
rect 4334 1970 4346 2126
rect 4398 1970 4410 2126
rect 4334 1571 4410 1970
rect 6162 2126 6238 2832
rect 7439 2625 7619 2637
rect 7439 2573 7451 2625
rect 7607 2573 7619 2625
rect 7439 2561 7619 2573
rect 6162 1970 6174 2126
rect 6226 1970 6238 2126
rect 6162 1958 6238 1970
rect 3564 1495 4410 1571
rect 2953 1473 3029 1485
rect 2953 1362 2965 1473
rect 1499 1350 2965 1362
rect 1499 1298 1511 1350
rect 1667 1317 2965 1350
rect 3017 1317 3029 1473
rect 1667 1298 3029 1317
rect 7543 1473 7619 2561
rect 7543 1317 7555 1473
rect 7607 1317 7619 1473
rect 7543 1305 7619 1317
rect 8162 1473 8238 2833
rect 9414 2761 9490 7636
rect 10095 6313 10171 7703
rect 9414 2605 9426 2761
rect 9478 2605 9490 2761
rect 9414 2593 9490 2605
rect 9570 6301 9750 6313
rect 9570 6249 9582 6301
rect 9738 6249 9750 6301
rect 9570 6237 9750 6249
rect 9991 6301 10171 6313
rect 9991 6249 10003 6301
rect 10159 6249 10171 6301
rect 9991 6237 10171 6249
rect 10275 7369 10351 7381
rect 10275 7213 10287 7369
rect 10339 7213 10351 7369
rect 9570 2729 9646 6237
rect 10275 6177 10351 7213
rect 9570 2573 9582 2729
rect 9634 2573 9646 2729
rect 9726 6165 9906 6177
rect 9726 6113 9738 6165
rect 9894 6113 9906 6165
rect 9726 6101 9906 6113
rect 10171 6165 10351 6177
rect 10171 6113 10183 6165
rect 10339 6113 10351 6165
rect 10171 6101 10351 6113
rect 9726 2773 9802 6101
rect 11245 5705 11321 10789
rect 13356 10691 13432 10703
rect 13356 10535 13368 10691
rect 13420 10535 13432 10691
rect 12164 9812 12240 9824
rect 12164 9656 12176 9812
rect 12228 9656 12240 9812
rect 12164 7970 12240 9656
rect 9892 5629 11321 5705
rect 11457 7894 12240 7970
rect 9892 2909 9948 5629
rect 10027 5364 10103 5374
rect 10027 4892 10037 5364
rect 10093 4892 10103 5364
rect 10027 4882 10103 4892
rect 10027 4178 10103 4188
rect 10027 3706 10037 4178
rect 10093 3706 10103 4178
rect 10027 3696 10103 3706
rect 9892 2897 10072 2909
rect 9892 2845 9904 2897
rect 10060 2845 10072 2897
rect 9892 2833 10072 2845
rect 11457 2794 11513 7894
rect 12136 6514 12316 6526
rect 12136 6462 12148 6514
rect 12304 6462 12316 6514
rect 12136 3348 12316 6462
rect 12136 3292 12146 3348
rect 12306 3292 12316 3348
rect 12136 3225 12316 3292
rect 12136 3173 12148 3225
rect 12304 3173 12316 3225
rect 12136 3161 12316 3173
rect 12736 6381 12812 6393
rect 12736 6225 12748 6381
rect 12800 6225 12812 6381
rect 12736 3045 12812 6225
rect 13356 6381 13432 10535
rect 13356 6225 13368 6381
rect 13420 6225 13432 6381
rect 13356 6213 13432 6225
rect 13376 5364 13452 5374
rect 13376 4892 13386 5364
rect 13442 4892 13452 5364
rect 13376 4882 13452 4892
rect 13356 4458 13432 4470
rect 13356 4302 13368 4458
rect 13420 4302 13432 4458
rect 13356 4290 13432 4302
rect 12537 3033 12812 3045
rect 12537 2981 12549 3033
rect 12705 2981 12812 3033
rect 12537 2969 12812 2981
rect 11457 2782 11637 2794
rect 9726 2761 9906 2773
rect 9726 2709 9738 2761
rect 9894 2709 9906 2761
rect 9726 2697 9906 2709
rect 9962 2761 10142 2773
rect 9962 2709 9974 2761
rect 10130 2709 10142 2761
rect 11457 2730 11469 2782
rect 11625 2730 11637 2782
rect 11457 2718 11637 2730
rect 12679 2782 12859 2794
rect 12679 2730 12691 2782
rect 12847 2730 12859 2782
rect 12679 2718 12859 2730
rect 9962 2697 10142 2709
rect 9570 2561 9646 2573
rect 10066 2126 10142 2697
rect 11302 2625 11482 2637
rect 11302 2573 11314 2625
rect 11470 2573 11482 2625
rect 11302 2561 11482 2573
rect 10066 1970 10078 2126
rect 10130 1970 10142 2126
rect 10066 1958 10142 1970
rect 11406 2126 11482 2561
rect 11406 1970 11418 2126
rect 11470 1970 11482 2126
rect 11406 1958 11482 1970
rect 8162 1317 8174 1473
rect 8226 1317 8238 1473
rect 8162 1305 8238 1317
rect 12783 1473 12859 2718
rect 12783 1317 12795 1473
rect 12847 1317 12859 1473
rect 12783 1305 12859 1317
rect 1499 1286 3029 1298
<< via2 >>
rect 10037 5362 10093 5364
rect 10037 4894 10039 5362
rect 10039 4894 10091 5362
rect 10091 4894 10093 5362
rect 10037 4892 10093 4894
rect 10037 4176 10093 4178
rect 10037 3708 10039 4176
rect 10039 3708 10091 4176
rect 10091 3708 10093 4176
rect 10037 3706 10093 3708
rect 12146 3292 12306 3348
rect 13386 5362 13442 5364
rect 13386 4894 13388 5362
rect 13388 4894 13440 5362
rect 13440 4894 13442 5362
rect 13386 4892 13442 4894
<< metal3 >>
rect 10027 5364 10103 5374
rect 10027 4892 10037 5364
rect 10093 4892 10103 5364
rect 10027 4882 10103 4892
rect 13376 5364 13452 5374
rect 13376 4892 13386 5364
rect 13442 4892 13452 5364
rect 13376 4882 13452 4892
rect 10027 4178 10103 4188
rect 10027 3706 10037 4178
rect 10093 3706 10103 4178
rect 10027 3696 10103 3706
rect 12136 3348 12316 3358
rect 12136 3292 12146 3348
rect 12306 3292 12316 3348
rect 12136 3282 12316 3292
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_0
timestamp 1669390400
transform 0 1 9452 -1 0 2683
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_1
timestamp 1669390400
transform 0 1 279 -1 0 1325
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_2
timestamp 1669390400
transform 0 -1 415 1 0 3059
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_3
timestamp 1669390400
transform 1 0 1589 0 1 2224
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_4
timestamp 1669390400
transform 1 0 12226 0 1 3199
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_5
timestamp 1669390400
transform 1 0 10261 0 1 6139
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_6
timestamp 1669390400
transform 1 0 6197 0 1 2870
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_7
timestamp 1669390400
transform 1 0 3261 0 1 2870
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_8
timestamp 1669390400
transform 1 0 7529 0 1 2599
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_9
timestamp 1669390400
transform 1 0 1589 0 1 1324
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_10
timestamp 1669390400
transform 1 0 -54 0 1 2599
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_11
timestamp 1669390400
transform 1 0 8148 0 1 2871
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_12
timestamp 1669390400
transform 1 0 12769 0 1 2756
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_13
timestamp 1669390400
transform 1 0 340 0 1 2224
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_14
timestamp 1669390400
transform 1 0 1874 0 1 2735
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_15
timestamp 1669390400
transform 1 0 10052 0 1 2735
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_16
timestamp 1669390400
transform 1 0 11392 0 1 2599
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_17
timestamp 1669390400
transform 1 0 6910 0 1 4240
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_18
timestamp 1669390400
transform 1 0 9982 0 1 2871
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_19
timestamp 1669390400
transform 1 0 11547 0 1 2756
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_20
timestamp 1669390400
transform 1 0 12627 0 1 3007
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_21
timestamp 1669390400
transform 1 0 9816 0 1 6139
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_22
timestamp 1669390400
transform 1 0 9660 0 1 6275
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_23
timestamp 1669390400
transform 1 0 10081 0 1 6275
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_24
timestamp 1669390400
transform 1 0 11184 0 1 10827
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_25
timestamp 1669390400
transform 1 0 12226 0 1 6488
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_26
timestamp 1669390400
transform 1 0 3059 0 1 3321
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1669390400
transform 0 -1 9816 1 0 2735
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1669390400
transform 1 0 10104 0 1 2048
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1669390400
transform 1 0 4372 0 1 2048
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1669390400
transform 1 0 7581 0 1 1395
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1669390400
transform 1 0 2991 0 1 1395
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_5
timestamp 1669390400
transform 1 0 12821 0 1 1395
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_6
timestamp 1669390400
transform 1 0 10313 0 1 7291
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_7
timestamp 1669390400
transform 1 0 10133 0 1 7781
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_8
timestamp 1669390400
transform 1 0 9608 0 1 2651
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_9
timestamp 1669390400
transform 1 0 11444 0 1 2048
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_10
timestamp 1669390400
transform 1 0 6200 0 1 2048
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_11
timestamp 1669390400
transform 1 0 13394 0 1 4380
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_12
timestamp 1669390400
transform 1 0 12774 0 1 6303
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_13
timestamp 1669390400
transform 1 0 8200 0 1 1395
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_14
timestamp 1669390400
transform 1 0 13394 0 1 6303
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_15
timestamp 1669390400
transform 1 0 13394 0 1 10613
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_16
timestamp 1669390400
transform 1 0 12202 0 1 9734
box 0 0 1 1
use M2_M1_CDNS_40661953145312  M2_M1_CDNS_40661953145312_0
timestamp 1669390400
transform 1 0 13414 0 1 5128
box 0 0 1 1
use M2_M1_CDNS_40661953145312  M2_M1_CDNS_40661953145312_1
timestamp 1669390400
transform 1 0 10065 0 1 5128
box 0 0 1 1
use M2_M1_CDNS_40661953145312  M2_M1_CDNS_40661953145312_2
timestamp 1669390400
transform 1 0 10065 0 1 3942
box 0 0 1 1
use M3_M2_CDNS_40661953145313  M3_M2_CDNS_40661953145313_0
timestamp 1669390400
transform 1 0 13414 0 1 5128
box 0 0 1 1
use M3_M2_CDNS_40661953145313  M3_M2_CDNS_40661953145313_1
timestamp 1669390400
transform 1 0 10065 0 1 3942
box 0 0 1 1
use M3_M2_CDNS_40661953145313  M3_M2_CDNS_40661953145313_2
timestamp 1669390400
transform 1 0 10065 0 1 5128
box 0 0 1 1
use M3_M2_CDNS_40661953145314  M3_M2_CDNS_40661953145314_0
timestamp 1669390400
transform 1 0 12226 0 1 3320
box 0 0 1 1
use comp018green_in_cms_smt  comp018green_in_cms_smt_0
timestamp 1669390400
transform 1 0 1532 0 1 3158
box -1402 0 6872 2575
use comp018green_in_drv  comp018green_in_drv_0
timestamp 1669390400
transform 1 0 8900 0 1 3158
box -443 0 4434 2575
use comp018green_in_logic_pupd  comp018green_in_logic_pupd_0
timestamp 1669390400
transform -1 0 13932 0 1 9724
box 428 -3277 3307 2142
use comp018green_in_pupd  comp018green_in_pupd_0
timestamp 1669390400
transform 0 -1 2979 -1 0 14857
box -83 -7722 8992 3035
use comp018green_sigbuf  comp018green_sigbuf_0
timestamp 1669390400
transform 1 0 7863 0 -1 2492
box -83 0 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_1
timestamp 1669390400
transform 1 0 2619 0 -1 2492
box -83 0 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_2
timestamp 1669390400
transform -1 0 13197 0 -1 2492
box -83 0 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_3
timestamp 1669390400
transform -1 0 7953 0 -1 2492
box -83 0 2795 2575
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_0
timestamp 1669390400
transform 1 0 1490 0 1 2124
box 0 0 1 1
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_1
timestamp 1669390400
transform 1 0 241 0 1 1224
box 0 0 1 1
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_2
timestamp 1669390400
transform 1 0 1490 0 1 1224
box 0 0 1 1
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_3
timestamp 1669390400
transform 1 0 241 0 1 2124
box 0 0 1 1
<< labels >>
rlabel metal2 s 6679 6191 6679 6191 4 PAD
port 1 nsew
rlabel metal2 s 2128 1324 2128 1324 4 IE
port 2 nsew
rlabel metal2 s -107 526 -107 526 4 CS
port 3 nsew
rlabel metal2 s 1822 2409 1822 2409 4 PD
port 4 nsew
rlabel metal2 s 414 522 414 522 4 PU
port 5 nsew
rlabel metal1 s 11686 5601 11686 5601 4 VDD
port 6 nsew
<< properties >>
string GDS_END 1654202
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1647262
string path 258.775 153.475 243.150 153.475 
<< end >>
