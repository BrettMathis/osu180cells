magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 153 7068 1633 7462
<< nmos >>
rect 651 486 771 2936
rect 875 486 995 2936
<< ndiff >>
rect 1295 4374 1379 4393
rect 1295 4046 1314 4374
rect 1360 4046 1379 4374
rect 1295 4027 1379 4046
rect 533 2891 651 2936
rect 533 2845 576 2891
rect 622 2845 651 2891
rect 533 2723 651 2845
rect 533 2677 576 2723
rect 622 2677 651 2723
rect 533 2556 651 2677
rect 533 2510 576 2556
rect 622 2510 651 2556
rect 533 2388 651 2510
rect 533 2342 576 2388
rect 622 2342 651 2388
rect 533 2220 651 2342
rect 533 2174 576 2220
rect 622 2174 651 2220
rect 533 2052 651 2174
rect 533 2006 576 2052
rect 622 2006 651 2052
rect 533 1884 651 2006
rect 533 1838 576 1884
rect 622 1838 651 1884
rect 533 1717 651 1838
rect 533 1671 576 1717
rect 622 1671 651 1717
rect 533 1549 651 1671
rect 533 1503 576 1549
rect 622 1503 651 1549
rect 533 1381 651 1503
rect 533 1335 576 1381
rect 622 1335 651 1381
rect 533 1213 651 1335
rect 533 1167 576 1213
rect 622 1167 651 1213
rect 533 1043 651 1167
rect 533 997 576 1043
rect 622 997 651 1043
rect 533 873 651 997
rect 533 827 576 873
rect 622 827 651 873
rect 533 703 651 827
rect 533 657 576 703
rect 622 657 651 703
rect 533 486 651 657
rect 771 486 875 2936
rect 995 2891 1114 2936
rect 995 2845 1025 2891
rect 1071 2845 1114 2891
rect 995 2723 1114 2845
rect 995 2677 1025 2723
rect 1071 2677 1114 2723
rect 995 2556 1114 2677
rect 995 2510 1025 2556
rect 1071 2510 1114 2556
rect 995 2388 1114 2510
rect 995 2342 1025 2388
rect 1071 2342 1114 2388
rect 995 2220 1114 2342
rect 995 2174 1025 2220
rect 1071 2174 1114 2220
rect 995 2052 1114 2174
rect 995 2006 1025 2052
rect 1071 2006 1114 2052
rect 995 1884 1114 2006
rect 995 1838 1025 1884
rect 1071 1838 1114 1884
rect 995 1717 1114 1838
rect 995 1671 1025 1717
rect 1071 1671 1114 1717
rect 995 1549 1114 1671
rect 995 1503 1025 1549
rect 1071 1503 1114 1549
rect 995 1381 1114 1503
rect 995 1335 1025 1381
rect 1071 1335 1114 1381
rect 995 1213 1114 1335
rect 995 1167 1025 1213
rect 1071 1167 1114 1213
rect 995 1043 1114 1167
rect 995 997 1025 1043
rect 1071 997 1114 1043
rect 995 873 1114 997
rect 995 827 1025 873
rect 1071 827 1114 873
rect 995 703 1114 827
rect 995 657 1025 703
rect 1071 657 1114 703
rect 995 486 1114 657
<< ndiffc >>
rect 1314 4046 1360 4374
rect 576 2845 622 2891
rect 576 2677 622 2723
rect 576 2510 622 2556
rect 576 2342 622 2388
rect 576 2174 622 2220
rect 576 2006 622 2052
rect 576 1838 622 1884
rect 576 1671 622 1717
rect 576 1503 622 1549
rect 576 1335 622 1381
rect 576 1167 622 1213
rect 576 997 622 1043
rect 576 827 622 873
rect 576 657 622 703
rect 1025 2845 1071 2891
rect 1025 2677 1071 2723
rect 1025 2510 1071 2556
rect 1025 2342 1071 2388
rect 1025 2174 1071 2220
rect 1025 2006 1071 2052
rect 1025 1838 1071 1884
rect 1025 1671 1071 1717
rect 1025 1503 1071 1549
rect 1025 1335 1071 1381
rect 1025 1167 1071 1213
rect 1025 997 1071 1043
rect 1025 827 1071 873
rect 1025 657 1071 703
<< psubdiff >>
rect 1271 2877 1403 2936
rect 1271 2831 1314 2877
rect 1360 2831 1403 2877
rect 1271 2714 1403 2831
rect 1271 2668 1314 2714
rect 1360 2668 1403 2714
rect 1271 2551 1403 2668
rect 1271 2505 1314 2551
rect 1360 2505 1403 2551
rect 1271 2388 1403 2505
rect 1271 2342 1314 2388
rect 1360 2342 1403 2388
rect 1271 2225 1403 2342
rect 1271 2179 1314 2225
rect 1360 2179 1403 2225
rect 1271 2061 1403 2179
rect 1271 2015 1314 2061
rect 1360 2015 1403 2061
rect 1271 1898 1403 2015
rect 1271 1852 1314 1898
rect 1360 1852 1403 1898
rect 1271 1735 1403 1852
rect 1271 1689 1314 1735
rect 1360 1689 1403 1735
rect 1271 1572 1403 1689
rect 1271 1526 1314 1572
rect 1360 1526 1403 1572
rect 1271 1408 1403 1526
rect 1271 1362 1314 1408
rect 1360 1362 1403 1408
rect 1271 1245 1403 1362
rect 1271 1199 1314 1245
rect 1360 1199 1403 1245
rect 1271 1082 1403 1199
rect 1271 1036 1314 1082
rect 1360 1036 1403 1082
rect 1271 919 1403 1036
rect 1271 873 1314 919
rect 1360 873 1403 919
rect 1271 756 1403 873
rect 1271 710 1314 756
rect 1360 710 1403 756
rect 1271 592 1403 710
rect 1271 546 1314 592
rect 1360 546 1403 592
rect 1271 486 1403 546
rect 440 218 1442 264
rect 440 172 522 218
rect 568 172 680 218
rect 726 172 838 218
rect 884 172 996 218
rect 1042 172 1154 218
rect 1200 172 1442 218
rect 440 126 1442 172
<< nsubdiff >>
rect 295 7239 1490 7296
rect 295 7193 418 7239
rect 464 7193 577 7239
rect 623 7193 1025 7239
rect 1071 7193 1183 7239
rect 1229 7193 1490 7239
rect 295 7136 1490 7193
<< psubdiffcont >>
rect 1314 2831 1360 2877
rect 1314 2668 1360 2714
rect 1314 2505 1360 2551
rect 1314 2342 1360 2388
rect 1314 2179 1360 2225
rect 1314 2015 1360 2061
rect 1314 1852 1360 1898
rect 1314 1689 1360 1735
rect 1314 1526 1360 1572
rect 1314 1362 1360 1408
rect 1314 1199 1360 1245
rect 1314 1036 1360 1082
rect 1314 873 1360 919
rect 1314 710 1360 756
rect 1314 546 1360 592
rect 522 172 568 218
rect 680 172 726 218
rect 838 172 884 218
rect 996 172 1042 218
rect 1154 172 1200 218
<< nsubdiffcont >>
rect 418 7193 464 7239
rect 577 7193 623 7239
rect 1025 7193 1071 7239
rect 1183 7193 1229 7239
<< polysilicon >>
rect 493 10059 613 10100
rect 717 10059 837 10100
rect 941 10059 1061 10100
rect 1165 10059 1285 10100
rect 493 9922 1285 10059
rect 493 9863 613 9922
rect 717 9863 837 9922
rect 941 9863 1061 9922
rect 1165 9863 1285 9922
rect 493 7520 613 7540
rect 717 7520 837 7539
rect 941 7520 1061 7539
rect 1165 7520 1285 7540
rect 493 7473 1285 7520
rect 493 7427 654 7473
rect 1076 7427 1285 7473
rect 493 7383 1285 7427
rect 651 2936 771 3871
rect 875 2936 995 3871
rect 651 414 771 486
rect 875 414 995 486
<< polycontact >>
rect 654 7427 1076 7473
<< metal1 >>
rect 383 11324 515 11392
rect 383 10925 499 11324
rect 831 10925 947 11392
rect 377 10885 505 10925
rect 377 10833 415 10885
rect 467 10833 505 10885
rect 377 10667 505 10833
rect 377 10615 415 10667
rect 467 10615 505 10667
rect 377 10449 505 10615
rect 377 10397 415 10449
rect 467 10397 505 10449
rect 377 10231 505 10397
rect 377 10179 415 10231
rect 467 10179 505 10231
rect 817 10924 947 10925
rect 817 10885 945 10924
rect 817 10833 855 10885
rect 907 10833 945 10885
rect 817 10667 945 10833
rect 817 10615 855 10667
rect 907 10615 945 10667
rect 817 10449 945 10615
rect 817 10397 855 10449
rect 907 10397 945 10449
rect 817 10231 945 10397
rect 377 10139 505 10179
rect 607 10050 723 10180
rect 817 10179 855 10231
rect 907 10179 945 10231
rect 817 10139 945 10179
rect 1049 10885 1177 10925
rect 1279 10924 1395 11392
rect 1049 10833 1087 10885
rect 1139 10833 1177 10885
rect 1049 10667 1177 10833
rect 1049 10615 1087 10667
rect 1139 10615 1177 10667
rect 1049 10449 1177 10615
rect 1049 10397 1087 10449
rect 1139 10397 1177 10449
rect 1049 10231 1177 10397
rect 1049 10179 1087 10231
rect 1139 10179 1177 10231
rect 1049 10139 1177 10179
rect 1055 10050 1171 10139
rect 607 9931 1171 10050
rect 607 9781 723 9931
rect 1055 9781 1171 9931
rect 377 9738 505 9777
rect 377 9686 415 9738
rect 467 9686 505 9738
rect 377 9520 505 9686
rect 377 9468 415 9520
rect 467 9468 505 9520
rect 377 9302 505 9468
rect 377 9250 415 9302
rect 467 9250 505 9302
rect 377 9210 505 9250
rect 825 9738 953 9777
rect 825 9686 863 9738
rect 915 9686 953 9738
rect 825 9520 953 9686
rect 825 9468 863 9520
rect 915 9468 953 9520
rect 825 9302 953 9468
rect 825 9250 863 9302
rect 915 9250 953 9302
rect 825 9210 953 9250
rect 1273 9738 1401 9777
rect 1273 9686 1311 9738
rect 1363 9686 1401 9738
rect 1273 9520 1401 9686
rect 1273 9468 1311 9520
rect 1363 9468 1401 9520
rect 1273 9302 1401 9468
rect 1273 9250 1311 9302
rect 1363 9250 1401 9302
rect 1273 9210 1401 9250
rect 495 7473 1283 7511
rect 495 7427 654 7473
rect 1076 7427 1283 7473
rect 495 7392 1283 7427
rect 765 7391 882 7392
rect 243 7239 657 7275
rect 243 7193 418 7239
rect 464 7193 577 7239
rect 623 7198 657 7239
rect 623 7193 658 7198
rect 243 7156 658 7193
rect 541 6827 658 7156
rect 765 6841 881 7391
rect 989 7239 1490 7275
rect 989 7193 1025 7239
rect 1071 7193 1183 7239
rect 1229 7193 1490 7239
rect 989 7156 1490 7193
rect 989 4374 1395 7156
rect 762 4227 886 4267
rect 762 4175 798 4227
rect 850 4175 886 4227
rect 762 4009 886 4175
rect 762 3957 798 4009
rect 850 3957 886 4009
rect 762 3917 886 3957
rect 989 4046 1314 4374
rect 1360 4046 1395 4374
rect 989 3916 1395 4046
rect 342 3676 1527 3768
rect 342 3474 1527 3567
rect 342 3273 1527 3365
rect 342 3071 1527 3163
rect 540 2891 657 2927
rect 540 2845 576 2891
rect 622 2845 657 2891
rect 540 2723 657 2845
rect 540 2677 576 2723
rect 622 2677 657 2723
rect 540 2556 657 2677
rect 540 2510 576 2556
rect 622 2510 657 2556
rect 540 2388 657 2510
rect 540 2342 576 2388
rect 622 2342 657 2388
rect 540 2220 657 2342
rect 540 2174 576 2220
rect 622 2174 657 2220
rect 540 2052 657 2174
rect 540 2006 576 2052
rect 622 2006 657 2052
rect 540 1884 657 2006
rect 540 1838 576 1884
rect 622 1838 657 1884
rect 540 1717 657 1838
rect 540 1671 576 1717
rect 622 1671 657 1717
rect 540 1549 657 1671
rect 540 1503 576 1549
rect 622 1503 657 1549
rect 540 1381 657 1503
rect 540 1335 576 1381
rect 622 1335 657 1381
rect 540 1270 657 1335
rect 989 2891 1395 2927
rect 989 2845 1025 2891
rect 1071 2877 1395 2891
rect 1071 2845 1314 2877
rect 989 2831 1314 2845
rect 1360 2831 1395 2877
rect 989 2723 1395 2831
rect 989 2677 1025 2723
rect 1071 2714 1395 2723
rect 1071 2677 1314 2714
rect 989 2668 1314 2677
rect 1360 2668 1395 2714
rect 989 2556 1395 2668
rect 989 2510 1025 2556
rect 1071 2551 1395 2556
rect 1071 2510 1314 2551
rect 989 2505 1314 2510
rect 1360 2505 1395 2551
rect 989 2388 1395 2505
rect 989 2342 1025 2388
rect 1071 2342 1314 2388
rect 1360 2342 1395 2388
rect 989 2225 1395 2342
rect 989 2220 1314 2225
rect 989 2174 1025 2220
rect 1071 2179 1314 2220
rect 1360 2179 1395 2225
rect 1071 2174 1395 2179
rect 989 2061 1395 2174
rect 989 2052 1314 2061
rect 989 2006 1025 2052
rect 1071 2015 1314 2052
rect 1360 2015 1395 2061
rect 1071 2006 1395 2015
rect 989 1898 1395 2006
rect 989 1884 1314 1898
rect 989 1838 1025 1884
rect 1071 1852 1314 1884
rect 1360 1852 1395 1898
rect 1071 1838 1395 1852
rect 989 1735 1395 1838
rect 989 1717 1314 1735
rect 989 1671 1025 1717
rect 1071 1689 1314 1717
rect 1360 1689 1395 1735
rect 1071 1671 1395 1689
rect 989 1572 1395 1671
rect 989 1549 1314 1572
rect 989 1503 1025 1549
rect 1071 1526 1314 1549
rect 1360 1526 1395 1572
rect 1071 1503 1395 1526
rect 989 1408 1395 1503
rect 989 1381 1314 1408
rect 989 1335 1025 1381
rect 1071 1362 1314 1381
rect 1360 1362 1395 1408
rect 1071 1335 1395 1362
rect 540 1213 656 1270
rect 540 1167 576 1213
rect 622 1167 656 1213
rect 540 1043 656 1167
rect 540 997 576 1043
rect 622 997 656 1043
rect 540 873 656 997
rect 540 827 576 873
rect 622 827 656 873
rect 540 703 656 827
rect 540 657 576 703
rect 622 657 656 703
rect 540 495 656 657
rect 989 1245 1395 1335
rect 989 1213 1314 1245
rect 989 1167 1025 1213
rect 1071 1199 1314 1213
rect 1360 1199 1395 1245
rect 1071 1167 1395 1199
rect 989 1082 1395 1167
rect 989 1043 1314 1082
rect 989 997 1025 1043
rect 1071 1036 1314 1043
rect 1360 1036 1395 1082
rect 1071 997 1395 1036
rect 989 919 1395 997
rect 989 873 1314 919
rect 1360 873 1395 919
rect 989 827 1025 873
rect 1071 827 1395 873
rect 989 756 1395 827
rect 989 710 1314 756
rect 1360 710 1395 756
rect 989 703 1395 710
rect 989 657 1025 703
rect 1071 657 1395 703
rect 989 592 1395 657
rect 989 546 1314 592
rect 1360 546 1395 592
rect 989 269 1395 546
rect 989 259 1402 269
rect 440 218 1442 259
rect 440 172 522 218
rect 568 172 680 218
rect 726 172 838 218
rect 884 172 996 218
rect 1042 172 1154 218
rect 1200 172 1442 218
rect 440 130 1442 172
<< via1 >>
rect 415 10833 467 10885
rect 415 10615 467 10667
rect 415 10397 467 10449
rect 415 10179 467 10231
rect 855 10833 907 10885
rect 855 10615 907 10667
rect 855 10397 907 10449
rect 855 10179 907 10231
rect 1087 10833 1139 10885
rect 1087 10615 1139 10667
rect 1087 10397 1139 10449
rect 1087 10179 1139 10231
rect 415 9686 467 9738
rect 415 9468 467 9520
rect 415 9250 467 9302
rect 863 9686 915 9738
rect 863 9468 915 9520
rect 863 9250 915 9302
rect 1311 9686 1363 9738
rect 1311 9468 1363 9520
rect 1311 9250 1363 9302
rect 798 4175 850 4227
rect 798 3957 850 4009
<< metal2 >>
rect 377 10887 505 10924
rect 377 10831 413 10887
rect 469 10831 505 10887
rect 377 10669 505 10831
rect 377 10613 413 10669
rect 469 10613 505 10669
rect 377 10451 505 10613
rect 377 10395 413 10451
rect 469 10395 505 10451
rect 377 10233 505 10395
rect 377 10177 413 10233
rect 469 10177 505 10233
rect 377 10139 505 10177
rect 817 10887 945 10924
rect 817 10831 853 10887
rect 909 10831 945 10887
rect 817 10669 945 10831
rect 817 10613 853 10669
rect 909 10613 945 10669
rect 817 10451 945 10613
rect 817 10395 853 10451
rect 909 10395 945 10451
rect 817 10233 945 10395
rect 817 10177 853 10233
rect 909 10177 945 10233
rect 817 10139 945 10177
rect 1049 10885 1270 11157
rect 1049 10833 1087 10885
rect 1139 10833 1270 10885
rect 1049 10667 1270 10833
rect 1049 10615 1087 10667
rect 1139 10615 1270 10667
rect 1049 10449 1270 10615
rect 1049 10397 1087 10449
rect 1139 10397 1270 10449
rect 1049 10231 1270 10397
rect 1049 10179 1087 10231
rect 1139 10179 1270 10231
rect 1049 10139 1270 10179
rect 377 9740 505 9777
rect 377 9684 413 9740
rect 469 9684 505 9740
rect 377 9522 505 9684
rect 377 9466 413 9522
rect 469 9466 505 9522
rect 377 9304 505 9466
rect 377 9248 413 9304
rect 469 9248 505 9304
rect 377 9210 505 9248
rect 825 9740 953 9777
rect 825 9684 861 9740
rect 917 9684 953 9740
rect 825 9522 953 9684
rect 825 9466 861 9522
rect 917 9466 953 9522
rect 825 9304 953 9466
rect 825 9248 861 9304
rect 917 9248 953 9304
rect 825 9210 953 9248
rect 1273 9740 1401 9777
rect 1273 9684 1309 9740
rect 1365 9684 1401 9740
rect 1273 9522 1401 9684
rect 1273 9466 1309 9522
rect 1365 9466 1401 9522
rect 1273 9304 1401 9466
rect 1273 9248 1309 9304
rect 1365 9248 1401 9304
rect 1273 9210 1401 9248
rect 989 5107 1402 7226
rect 535 4227 887 4267
rect 535 4175 798 4227
rect 850 4175 887 4227
rect 535 4009 887 4175
rect 535 3957 798 4009
rect 850 3957 887 4009
rect 535 3916 887 3957
rect 535 2581 663 3916
rect 989 2751 1402 2927
rect 989 2695 1026 2751
rect 1082 2695 1309 2751
rect 1365 2695 1402 2751
rect 989 2533 1402 2695
rect 989 2477 1026 2533
rect 1082 2477 1309 2533
rect 1365 2477 1402 2533
rect 989 2315 1402 2477
rect 989 2259 1026 2315
rect 1082 2259 1309 2315
rect 1365 2259 1402 2315
rect 989 793 1402 2259
rect 989 737 1026 793
rect 1082 737 1309 793
rect 1365 737 1402 793
rect 989 575 1402 737
rect 989 519 1026 575
rect 1082 519 1309 575
rect 1365 519 1402 575
rect 989 357 1402 519
rect 989 301 1026 357
rect 1082 301 1309 357
rect 1365 301 1402 357
rect 989 139 1402 301
rect 989 83 1026 139
rect 1082 83 1309 139
rect 1365 83 1402 139
rect 989 42 1402 83
<< via2 >>
rect 413 10885 469 10887
rect 413 10833 415 10885
rect 415 10833 467 10885
rect 467 10833 469 10885
rect 413 10831 469 10833
rect 413 10667 469 10669
rect 413 10615 415 10667
rect 415 10615 467 10667
rect 467 10615 469 10667
rect 413 10613 469 10615
rect 413 10449 469 10451
rect 413 10397 415 10449
rect 415 10397 467 10449
rect 467 10397 469 10449
rect 413 10395 469 10397
rect 413 10231 469 10233
rect 413 10179 415 10231
rect 415 10179 467 10231
rect 467 10179 469 10231
rect 413 10177 469 10179
rect 853 10885 909 10887
rect 853 10833 855 10885
rect 855 10833 907 10885
rect 907 10833 909 10885
rect 853 10831 909 10833
rect 853 10667 909 10669
rect 853 10615 855 10667
rect 855 10615 907 10667
rect 907 10615 909 10667
rect 853 10613 909 10615
rect 853 10449 909 10451
rect 853 10397 855 10449
rect 855 10397 907 10449
rect 907 10397 909 10449
rect 853 10395 909 10397
rect 853 10231 909 10233
rect 853 10179 855 10231
rect 855 10179 907 10231
rect 907 10179 909 10231
rect 853 10177 909 10179
rect 413 9738 469 9740
rect 413 9686 415 9738
rect 415 9686 467 9738
rect 467 9686 469 9738
rect 413 9684 469 9686
rect 413 9520 469 9522
rect 413 9468 415 9520
rect 415 9468 467 9520
rect 467 9468 469 9520
rect 413 9466 469 9468
rect 413 9302 469 9304
rect 413 9250 415 9302
rect 415 9250 467 9302
rect 467 9250 469 9302
rect 413 9248 469 9250
rect 861 9738 917 9740
rect 861 9686 863 9738
rect 863 9686 915 9738
rect 915 9686 917 9738
rect 861 9684 917 9686
rect 861 9520 917 9522
rect 861 9468 863 9520
rect 863 9468 915 9520
rect 915 9468 917 9520
rect 861 9466 917 9468
rect 861 9302 917 9304
rect 861 9250 863 9302
rect 863 9250 915 9302
rect 915 9250 917 9302
rect 861 9248 917 9250
rect 1309 9738 1365 9740
rect 1309 9686 1311 9738
rect 1311 9686 1363 9738
rect 1363 9686 1365 9738
rect 1309 9684 1365 9686
rect 1309 9520 1365 9522
rect 1309 9468 1311 9520
rect 1311 9468 1363 9520
rect 1363 9468 1365 9520
rect 1309 9466 1365 9468
rect 1309 9302 1365 9304
rect 1309 9250 1311 9302
rect 1311 9250 1363 9302
rect 1363 9250 1365 9302
rect 1309 9248 1365 9250
rect 1026 2695 1082 2751
rect 1309 2695 1365 2751
rect 1026 2477 1082 2533
rect 1309 2477 1365 2533
rect 1026 2259 1082 2315
rect 1309 2259 1365 2315
rect 1026 737 1082 793
rect 1309 737 1365 793
rect 1026 519 1082 575
rect 1309 519 1365 575
rect 1026 301 1082 357
rect 1309 301 1365 357
rect 1026 83 1082 139
rect 1309 83 1365 139
<< metal3 >>
rect 153 10887 1483 10937
rect 153 10831 413 10887
rect 469 10831 853 10887
rect 909 10831 1483 10887
rect 153 10669 1483 10831
rect 153 10613 413 10669
rect 469 10613 853 10669
rect 909 10613 1483 10669
rect 153 10451 1483 10613
rect 153 10395 413 10451
rect 469 10395 853 10451
rect 909 10395 1483 10451
rect 153 10233 1483 10395
rect 153 10177 413 10233
rect 469 10177 853 10233
rect 909 10177 1483 10233
rect 153 9985 1483 10177
rect 153 9740 1483 9873
rect 153 9684 413 9740
rect 469 9684 861 9740
rect 917 9684 1309 9740
rect 1365 9684 1483 9740
rect 153 9522 1483 9684
rect 153 9466 413 9522
rect 469 9466 861 9522
rect 917 9466 1309 9522
rect 1365 9466 1483 9522
rect 153 9304 1483 9466
rect 153 9248 413 9304
rect 469 9248 861 9304
rect 917 9248 1309 9304
rect 1365 9248 1483 9304
rect 153 9160 1483 9248
rect 153 8117 1481 9026
rect 153 5057 1481 7779
rect 855 2751 1483 2882
rect 855 2695 1026 2751
rect 1082 2695 1309 2751
rect 1365 2695 1483 2751
rect 855 2533 1483 2695
rect 855 2477 1026 2533
rect 1082 2477 1309 2533
rect 1365 2477 1483 2533
rect 855 2315 1483 2477
rect 855 2259 1026 2315
rect 1082 2259 1309 2315
rect 1365 2259 1483 2315
rect 855 2200 1483 2259
rect 855 1044 1485 1952
rect 855 793 1488 873
rect 855 737 1026 793
rect 1082 737 1309 793
rect 1365 737 1488 793
rect 855 575 1488 737
rect 855 519 1026 575
rect 1082 519 1309 575
rect 1365 519 1488 575
rect 855 357 1488 519
rect 855 301 1026 357
rect 1082 301 1309 357
rect 1365 301 1488 357
rect 855 139 1488 301
rect 855 83 1026 139
rect 1082 83 1309 139
rect 1365 83 1488 139
rect 855 -35 1488 83
use M1_NACTIVE4310589983229_64x8m81  M1_NACTIVE4310589983229_64x8m81_0
timestamp 1669390400
transform 1 0 1337 0 1 4210
box 0 0 1 1
use M1_POLY24310589983260_64x8m81  M1_POLY24310589983260_64x8m81_0
timestamp 1669390400
transform 1 0 865 0 1 7450
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1669390400
transform -1 0 824 0 1 4092
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_0
timestamp 1669390400
transform -1 0 599 0 1 2099
box -63 -828 64 828
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_0
timestamp 1669390400
transform 1 0 1113 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_1
timestamp 1669390400
transform 1 0 881 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_2
timestamp 1669390400
transform 1 0 441 0 1 10532
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_0
timestamp 1669390400
transform 1 0 441 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_1
timestamp 1669390400
transform 1 0 889 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_2
timestamp 1669390400
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_0
timestamp 1669390400
transform 1 0 1054 0 1 6153
box -64 -1046 64 1046
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_1
timestamp 1669390400
transform 1 0 602 0 1 6153
box -64 -1046 64 1046
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_2
timestamp 1669390400
transform 1 0 1337 0 1 6153
box -64 -1046 64 1046
use M2_M1$$47640620_64x8m81  M2_M1$$47640620_64x8m81_0
timestamp 1669390400
transform 1 0 1337 0 1 1526
box -65 -1264 65 1264
use M2_M1$$47640620_64x8m81  M2_M1$$47640620_64x8m81_1
timestamp 1669390400
transform 1 0 1054 0 1 1526
box -65 -1264 65 1264
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_0
timestamp 1669390400
transform 1 0 1337 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_1
timestamp 1669390400
transform 1 0 1054 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_2
timestamp 1669390400
transform 1 0 441 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_3
timestamp 1669390400
transform 1 0 889 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_4
timestamp 1669390400
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_0
timestamp 1669390400
transform 1 0 1337 0 1 438
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_1
timestamp 1669390400
transform 1 0 1054 0 1 438
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_2
timestamp 1669390400
transform 1 0 881 0 1 10532
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_3
timestamp 1669390400
transform 1 0 441 0 1 10532
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_0
timestamp 1669390400
transform 1 0 1054 0 1 6153
box -65 -1046 65 1046
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_1
timestamp 1669390400
transform 1 0 602 0 1 6153
box -65 -1046 65 1046
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_2
timestamp 1669390400
transform 1 0 1337 0 1 6153
box -65 -1046 65 1046
use nmos_1p2$$47641644_64x8m81  nmos_1p2$$47641644_64x8m81_0
timestamp 1669390400
transform -1 0 1254 0 -1 11038
box -119 -73 177 980
use nmos_1p2$$47641644_64x8m81  nmos_1p2$$47641644_64x8m81_1
timestamp 1669390400
transform -1 0 806 0 -1 11038
box -119 -73 177 980
use nmos_1p2$$47641644_64x8m81  nmos_1p2$$47641644_64x8m81_2
timestamp 1669390400
transform -1 0 582 0 -1 11038
box -119 -73 177 980
use nmos_1p2$$47641644_64x8m81  nmos_1p2$$47641644_64x8m81_3
timestamp 1669390400
transform -1 0 1030 0 -1 11038
box -119 -73 177 980
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_0
timestamp 1669390400
transform -1 0 1030 0 -1 9850
box -286 -141 344 2409
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_1
timestamp 1669390400
transform -1 0 806 0 -1 9850
box -286 -141 344 2409
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_2
timestamp 1669390400
transform -1 0 582 0 -1 9850
box -286 -141 344 2409
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_3
timestamp 1669390400
transform -1 0 1254 0 -1 9850
box -286 -141 344 2409
use pmos_1p2$$47642668_64x8m81  pmos_1p2$$47642668_64x8m81_0
timestamp 1669390400
transform -1 0 964 0 1 3908
box -546 -142 344 3179
use pmos_1p2$$47643692_64x8m81  pmos_1p2$$47643692_64x8m81_0
timestamp 1669390400
transform -1 0 740 0 1 3908
box -286 -142 344 3179
<< properties >>
string GDS_END 430268
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 421950
<< end >>
