magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 3110 870
rect -86 352 1560 377
rect 2713 352 3110 377
<< pwell >>
rect -86 -86 3110 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1736 93 1856 257
rect 1960 93 2080 257
rect 2184 93 2304 257
rect 2408 93 2528 257
rect 2676 68 2796 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 592 497 692 716
rect 796 497 896 716
rect 1020 497 1120 716
rect 1244 497 1344 716
rect 1488 497 1588 716
rect 1756 497 1856 716
rect 1980 497 2080 716
rect 2184 497 2284 716
rect 2408 497 2508 716
rect 2676 497 2776 716
<< mvndiff >>
rect 1648 244 1736 257
rect 1648 232 1661 244
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 127 348 232
rect 244 81 273 127
rect 319 81 348 127
rect 244 68 348 81
rect 468 219 572 232
rect 468 173 497 219
rect 543 173 572 219
rect 468 68 572 173
rect 692 127 796 232
rect 692 81 721 127
rect 767 81 796 127
rect 692 68 796 81
rect 916 219 1020 232
rect 916 173 945 219
rect 991 173 1020 219
rect 916 68 1020 173
rect 1140 127 1244 232
rect 1140 81 1169 127
rect 1215 81 1244 127
rect 1140 68 1244 81
rect 1364 152 1468 232
rect 1364 106 1393 152
rect 1439 106 1468 152
rect 1364 68 1468 106
rect 1588 198 1661 232
rect 1707 198 1736 244
rect 1588 93 1736 198
rect 1856 152 1960 257
rect 1856 106 1885 152
rect 1931 106 1960 152
rect 1856 93 1960 106
rect 2080 244 2184 257
rect 2080 198 2109 244
rect 2155 198 2184 244
rect 2080 93 2184 198
rect 2304 152 2408 257
rect 2304 106 2333 152
rect 2379 106 2408 152
rect 2304 93 2408 106
rect 2528 244 2616 257
rect 2528 198 2557 244
rect 2603 232 2616 244
rect 2603 198 2676 232
rect 2528 93 2676 198
rect 1588 68 1668 93
rect 2596 68 2676 93
rect 2796 152 2884 232
rect 2796 106 2825 152
rect 2871 106 2884 152
rect 2796 68 2884 106
<< mvpdiff >>
rect 56 685 144 716
rect 56 545 69 685
rect 115 545 144 685
rect 56 497 144 545
rect 244 497 368 716
rect 468 497 592 716
rect 692 639 796 716
rect 692 593 721 639
rect 767 593 796 639
rect 692 497 796 593
rect 896 497 1020 716
rect 1120 497 1244 716
rect 1344 703 1488 716
rect 1344 657 1393 703
rect 1439 657 1488 703
rect 1344 497 1488 657
rect 1588 497 1756 716
rect 1856 497 1980 716
rect 2080 639 2184 716
rect 2080 593 2109 639
rect 2155 593 2184 639
rect 2080 497 2184 593
rect 2284 497 2408 716
rect 2508 497 2676 716
rect 2776 685 2864 716
rect 2776 545 2805 685
rect 2851 545 2864 685
rect 2776 497 2864 545
<< mvndiffc >>
rect 49 173 95 219
rect 273 81 319 127
rect 497 173 543 219
rect 721 81 767 127
rect 945 173 991 219
rect 1169 81 1215 127
rect 1393 106 1439 152
rect 1661 198 1707 244
rect 1885 106 1931 152
rect 2109 198 2155 244
rect 2333 106 2379 152
rect 2557 198 2603 244
rect 2825 106 2871 152
<< mvpdiffc >>
rect 69 545 115 685
rect 721 593 767 639
rect 1393 657 1439 703
rect 2109 593 2155 639
rect 2805 545 2851 685
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 592 716 692 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1488 716 1588 760
rect 1756 716 1856 760
rect 1980 716 2080 760
rect 2184 716 2284 760
rect 2408 716 2508 760
rect 2676 716 2776 760
rect 144 416 244 497
rect 144 402 174 416
rect 124 370 174 402
rect 220 370 244 416
rect 368 415 468 497
rect 368 402 395 415
rect 124 232 244 370
rect 348 369 395 402
rect 441 369 468 415
rect 592 415 692 497
rect 592 402 619 415
rect 348 232 468 369
rect 572 369 619 402
rect 665 394 692 415
rect 796 415 896 497
rect 796 394 823 415
rect 665 369 823 394
rect 869 402 896 415
rect 1020 402 1120 497
rect 1244 415 1344 497
rect 869 369 916 402
rect 572 346 916 369
rect 572 232 692 346
rect 796 232 916 346
rect 1020 356 1041 402
rect 1087 356 1140 402
rect 1020 232 1140 356
rect 1244 369 1263 415
rect 1309 402 1344 415
rect 1488 415 1588 497
rect 1488 402 1515 415
rect 1309 369 1364 402
rect 1244 232 1364 369
rect 1468 369 1515 402
rect 1561 369 1588 415
rect 1756 415 1856 497
rect 1756 402 1783 415
rect 1468 232 1588 369
rect 1736 369 1783 402
rect 1829 369 1856 415
rect 1980 402 2080 497
rect 1736 257 1856 369
rect 1960 394 2080 402
rect 2184 402 2284 497
rect 2408 428 2508 497
rect 2184 394 2304 402
rect 1960 346 2304 394
rect 1960 336 2080 346
rect 1960 290 1997 336
rect 2043 290 2080 336
rect 1960 257 2080 290
rect 2184 336 2304 346
rect 2184 290 2221 336
rect 2267 290 2304 336
rect 2184 257 2304 290
rect 2408 382 2435 428
rect 2481 402 2508 428
rect 2676 433 2776 497
rect 2481 382 2528 402
rect 2408 257 2528 382
rect 2676 387 2698 433
rect 2744 402 2776 433
rect 2744 387 2796 402
rect 2676 232 2796 387
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1736 24 1856 93
rect 1960 24 2080 93
rect 2184 24 2304 93
rect 2408 24 2528 93
rect 2676 24 2796 68
<< polycontact >>
rect 174 370 220 416
rect 395 369 441 415
rect 619 369 665 415
rect 823 369 869 415
rect 1041 356 1087 402
rect 1263 369 1309 415
rect 1515 369 1561 415
rect 1783 369 1829 415
rect 1997 290 2043 336
rect 2221 290 2267 336
rect 2435 382 2481 428
rect 2698 387 2744 433
<< metal1 >>
rect 0 724 3024 844
rect 69 685 115 724
rect 1382 703 1450 724
rect 1382 657 1393 703
rect 1439 657 1450 703
rect 2805 685 2851 724
rect 550 639 1332 648
rect 550 593 721 639
rect 767 611 1332 639
rect 1500 639 2243 648
rect 1500 611 2109 639
rect 767 593 2109 611
rect 2155 593 2243 639
rect 550 584 2243 593
rect 1282 565 1550 584
rect 69 526 115 545
rect 165 476 1212 536
rect 165 424 229 476
rect 56 416 229 424
rect 56 370 174 416
rect 220 370 229 416
rect 56 360 229 370
rect 302 415 532 430
rect 302 369 395 415
rect 441 369 532 415
rect 302 354 532 369
rect 578 415 990 424
rect 578 369 619 415
rect 665 369 823 415
rect 869 369 990 415
rect 578 360 990 369
rect 1036 402 1096 430
rect 482 311 532 354
rect 1036 356 1041 402
rect 1087 356 1096 402
rect 1144 424 1212 476
rect 1144 415 1320 424
rect 1144 369 1263 415
rect 1309 369 1320 415
rect 1144 360 1320 369
rect 1036 311 1096 356
rect 482 265 1096 311
rect 1370 244 1430 565
rect 1600 474 2755 536
rect 2805 526 2851 545
rect 1600 428 1646 474
rect 2687 433 2755 474
rect 1488 415 1646 428
rect 1488 369 1515 415
rect 1561 369 1646 415
rect 1488 356 1646 369
rect 1696 415 2435 428
rect 1696 369 1783 415
rect 1829 382 2435 415
rect 2481 382 2508 428
rect 2687 387 2698 433
rect 2744 387 2755 433
rect 2687 382 2755 387
rect 1829 369 1904 382
rect 1696 356 1904 369
rect 2824 336 2888 476
rect 1960 290 1997 336
rect 2043 290 2221 336
rect 2267 290 2888 336
rect 36 173 49 219
rect 95 173 497 219
rect 543 173 945 219
rect 991 173 1322 219
rect 1370 198 1661 244
rect 1707 198 2109 244
rect 2155 198 2557 244
rect 2603 198 2614 244
rect 2676 232 2888 290
rect 1276 152 1322 173
rect 262 81 273 127
rect 319 81 330 127
rect 262 60 330 81
rect 710 81 721 127
rect 767 81 778 127
rect 710 60 778 81
rect 1158 81 1169 127
rect 1215 81 1226 127
rect 1276 106 1393 152
rect 1439 106 1885 152
rect 1931 106 2333 152
rect 2379 106 2825 152
rect 2871 106 2884 152
rect 1158 60 1226 81
rect 0 -60 3024 60
<< labels >>
flabel metal1 s 1600 474 2755 536 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 578 360 990 424 0 FreeSans 400 0 0 0 B1
port 4 nsew default input
flabel metal1 s 1036 354 1096 430 0 FreeSans 400 0 0 0 B2
port 5 nsew default input
flabel metal1 s 165 476 1212 536 0 FreeSans 400 0 0 0 B3
port 6 nsew default input
flabel metal1 s 0 724 3024 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 1158 60 1226 127 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1500 611 2243 648 0 FreeSans 400 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 2824 336 2888 476 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1696 382 2508 428 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
rlabel metal1 s 1960 290 2888 336 1 A1
port 1 nsew default input
rlabel metal1 s 2676 232 2888 290 1 A1
port 1 nsew default input
rlabel metal1 s 1696 356 1904 382 1 A2
port 2 nsew default input
rlabel metal1 s 2687 428 2755 474 1 A3
port 3 nsew default input
rlabel metal1 s 1600 428 1646 474 1 A3
port 3 nsew default input
rlabel metal1 s 2687 382 2755 428 1 A3
port 3 nsew default input
rlabel metal1 s 1488 382 1646 428 1 A3
port 3 nsew default input
rlabel metal1 s 1488 356 1646 382 1 A3
port 3 nsew default input
rlabel metal1 s 302 354 532 430 1 B2
port 5 nsew default input
rlabel metal1 s 1036 311 1096 354 1 B2
port 5 nsew default input
rlabel metal1 s 482 311 532 354 1 B2
port 5 nsew default input
rlabel metal1 s 482 265 1096 311 1 B2
port 5 nsew default input
rlabel metal1 s 1144 424 1212 476 1 B3
port 6 nsew default input
rlabel metal1 s 165 424 229 476 1 B3
port 6 nsew default input
rlabel metal1 s 1144 360 1320 424 1 B3
port 6 nsew default input
rlabel metal1 s 56 360 229 424 1 B3
port 6 nsew default input
rlabel metal1 s 550 611 1332 648 1 ZN
port 7 nsew default output
rlabel metal1 s 550 584 2243 611 1 ZN
port 7 nsew default output
rlabel metal1 s 1282 565 1550 584 1 ZN
port 7 nsew default output
rlabel metal1 s 1370 244 1430 565 1 ZN
port 7 nsew default output
rlabel metal1 s 1370 198 2614 244 1 ZN
port 7 nsew default output
rlabel metal1 s 2805 657 2851 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1382 657 1450 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 69 657 115 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2805 526 2851 657 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 69 526 115 657 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 710 60 778 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3024 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3024 784
string GDS_END 77516
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 71762
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
