magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 1672 560
<< mvpmos >>
rect 0 0 120 440
rect 224 0 344 440
rect 448 0 568 440
rect 672 0 792 440
rect 896 0 1016 440
rect 1120 0 1240 440
rect 1344 0 1464 440
<< mvpdiff >>
rect -88 427 0 440
rect -88 381 -75 427
rect -29 381 0 427
rect -88 305 0 381
rect -88 259 -75 305
rect -29 259 0 305
rect -88 182 0 259
rect -88 136 -75 182
rect -29 136 0 182
rect -88 59 0 136
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 427 224 440
rect 120 381 149 427
rect 195 381 224 427
rect 120 305 224 381
rect 120 259 149 305
rect 195 259 224 305
rect 120 182 224 259
rect 120 136 149 182
rect 195 136 224 182
rect 120 59 224 136
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 427 448 440
rect 344 381 373 427
rect 419 381 448 427
rect 344 305 448 381
rect 344 259 373 305
rect 419 259 448 305
rect 344 182 448 259
rect 344 136 373 182
rect 419 136 448 182
rect 344 59 448 136
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 427 672 440
rect 568 381 597 427
rect 643 381 672 427
rect 568 305 672 381
rect 568 259 597 305
rect 643 259 672 305
rect 568 182 672 259
rect 568 136 597 182
rect 643 136 672 182
rect 568 59 672 136
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 427 896 440
rect 792 381 821 427
rect 867 381 896 427
rect 792 305 896 381
rect 792 259 821 305
rect 867 259 896 305
rect 792 182 896 259
rect 792 136 821 182
rect 867 136 896 182
rect 792 59 896 136
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 427 1120 440
rect 1016 381 1045 427
rect 1091 381 1120 427
rect 1016 305 1120 381
rect 1016 259 1045 305
rect 1091 259 1120 305
rect 1016 182 1120 259
rect 1016 136 1045 182
rect 1091 136 1120 182
rect 1016 59 1120 136
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 427 1344 440
rect 1240 381 1269 427
rect 1315 381 1344 427
rect 1240 305 1344 381
rect 1240 259 1269 305
rect 1315 259 1344 305
rect 1240 182 1344 259
rect 1240 136 1269 182
rect 1315 136 1344 182
rect 1240 59 1344 136
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 427 1552 440
rect 1464 381 1493 427
rect 1539 381 1552 427
rect 1464 305 1552 381
rect 1464 259 1493 305
rect 1539 259 1552 305
rect 1464 182 1552 259
rect 1464 136 1493 182
rect 1539 136 1552 182
rect 1464 59 1552 136
rect 1464 13 1493 59
rect 1539 13 1552 59
rect 1464 0 1552 13
<< mvpdiffc >>
rect -75 381 -29 427
rect -75 259 -29 305
rect -75 136 -29 182
rect -75 13 -29 59
rect 149 381 195 427
rect 149 259 195 305
rect 149 136 195 182
rect 149 13 195 59
rect 373 381 419 427
rect 373 259 419 305
rect 373 136 419 182
rect 373 13 419 59
rect 597 381 643 427
rect 597 259 643 305
rect 597 136 643 182
rect 597 13 643 59
rect 821 381 867 427
rect 821 259 867 305
rect 821 136 867 182
rect 821 13 867 59
rect 1045 381 1091 427
rect 1045 259 1091 305
rect 1045 136 1091 182
rect 1045 13 1091 59
rect 1269 381 1315 427
rect 1269 259 1315 305
rect 1269 136 1315 182
rect 1269 13 1315 59
rect 1493 381 1539 427
rect 1493 259 1539 305
rect 1493 136 1539 182
rect 1493 13 1539 59
<< polysilicon >>
rect 0 440 120 484
rect 224 440 344 484
rect 448 440 568 484
rect 672 440 792 484
rect 896 440 1016 484
rect 1120 440 1240 484
rect 1344 440 1464 484
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
<< metal1 >>
rect -75 427 -29 440
rect -75 305 -29 381
rect -75 182 -29 259
rect -75 59 -29 136
rect -75 0 -29 13
rect 149 427 195 440
rect 149 305 195 381
rect 149 182 195 259
rect 149 59 195 136
rect 149 0 195 13
rect 373 427 419 440
rect 373 305 419 381
rect 373 182 419 259
rect 373 59 419 136
rect 373 0 419 13
rect 597 427 643 440
rect 597 305 643 381
rect 597 182 643 259
rect 597 59 643 136
rect 597 0 643 13
rect 821 427 867 440
rect 821 305 867 381
rect 821 182 867 259
rect 821 59 867 136
rect 821 0 867 13
rect 1045 427 1091 440
rect 1045 305 1091 381
rect 1045 182 1091 259
rect 1045 59 1091 136
rect 1045 0 1091 13
rect 1269 427 1315 440
rect 1269 305 1315 381
rect 1269 182 1315 259
rect 1269 59 1315 136
rect 1269 0 1315 13
rect 1493 427 1539 440
rect 1493 305 1539 381
rect 1493 182 1539 259
rect 1493 59 1539 136
rect 1493 0 1539 13
<< labels >>
flabel metal1 s -52 220 -52 220 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 220 1516 220 0 FreeSans 400 0 0 0 D
flabel metal1 s 172 220 172 220 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 220 396 220 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 220 620 220 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 220 844 220 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 220 1068 220 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 220 1292 220 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 630764
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 625464
<< end >>
