magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 572 89 645
rect 193 572 313 645
rect 417 572 537 645
rect 641 572 761 645
rect 865 572 985 645
rect 1089 572 1209 645
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 641 -74 761 -1
rect 865 -73 985 -1
rect 1089 -74 1209 -1
use nmos_5p04310590878135_256x8m81  nmos_5p04310590878135_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 1328 616
<< properties >>
string GDS_END 240980
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 240090
<< end >>
