magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 776 2120
<< mvpmos >>
rect 0 0 120 2000
rect 224 0 344 2000
rect 448 0 568 2000
<< mvpdiff >>
rect -88 1987 0 2000
rect -88 13 -75 1987
rect -29 13 0 1987
rect -88 0 0 13
rect 120 1987 224 2000
rect 120 13 149 1987
rect 195 13 224 1987
rect 120 0 224 13
rect 344 1987 448 2000
rect 344 13 373 1987
rect 419 13 448 1987
rect 344 0 448 13
rect 568 1987 656 2000
rect 568 13 597 1987
rect 643 13 656 1987
rect 568 0 656 13
<< mvpdiffc >>
rect -75 13 -29 1987
rect 149 13 195 1987
rect 373 13 419 1987
rect 597 13 643 1987
<< polysilicon >>
rect 0 2000 120 2044
rect 224 2000 344 2044
rect 448 2000 568 2044
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
<< metal1 >>
rect -75 1987 -29 2000
rect -75 0 -29 13
rect 149 1987 195 2000
rect 149 0 195 13
rect 373 1987 419 2000
rect 373 0 419 13
rect 597 1987 643 2000
rect 597 0 643 13
<< labels >>
flabel metal1 s -52 1000 -52 1000 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 1000 620 1000 0 FreeSans 400 0 0 0 D
flabel metal1 s 172 1000 172 1000 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 1000 396 1000 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 145604
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 138760
<< end >>
