magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 132
<< mvndiff >>
rect -88 89 0 132
rect -88 43 -75 89
rect -29 43 0 89
rect -88 0 0 43
rect 120 89 208 132
rect 120 43 149 89
rect 195 43 208 89
rect 120 0 208 43
<< mvndiffc >>
rect -75 43 -29 89
rect 149 43 195 89
<< polysilicon >>
rect 0 132 120 176
rect 0 -44 120 0
<< metal1 >>
rect -75 89 -29 132
rect -75 0 -29 43
rect 149 89 195 132
rect 149 0 195 43
<< labels >>
flabel metal1 s -52 66 -52 66 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 66 172 66 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 496018
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 494994
<< end >>
