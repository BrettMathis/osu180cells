magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 1316
<< mvndiff >>
rect -88 1303 0 1316
rect -88 1257 -75 1303
rect -29 1257 0 1303
rect -88 1200 0 1257
rect -88 1154 -75 1200
rect -29 1154 0 1200
rect -88 1097 0 1154
rect -88 1051 -75 1097
rect -29 1051 0 1097
rect -88 994 0 1051
rect -88 948 -75 994
rect -29 948 0 994
rect -88 891 0 948
rect -88 845 -75 891
rect -29 845 0 891
rect -88 787 0 845
rect -88 741 -75 787
rect -29 741 0 787
rect -88 683 0 741
rect -88 637 -75 683
rect -29 637 0 683
rect -88 579 0 637
rect -88 533 -75 579
rect -29 533 0 579
rect -88 475 0 533
rect -88 429 -75 475
rect -29 429 0 475
rect -88 371 0 429
rect -88 325 -75 371
rect -29 325 0 371
rect -88 267 0 325
rect -88 221 -75 267
rect -29 221 0 267
rect -88 163 0 221
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1303 208 1316
rect 120 1257 149 1303
rect 195 1257 208 1303
rect 120 1200 208 1257
rect 120 1154 149 1200
rect 195 1154 208 1200
rect 120 1097 208 1154
rect 120 1051 149 1097
rect 195 1051 208 1097
rect 120 994 208 1051
rect 120 948 149 994
rect 195 948 208 994
rect 120 891 208 948
rect 120 845 149 891
rect 195 845 208 891
rect 120 787 208 845
rect 120 741 149 787
rect 195 741 208 787
rect 120 683 208 741
rect 120 637 149 683
rect 195 637 208 683
rect 120 579 208 637
rect 120 533 149 579
rect 195 533 208 579
rect 120 475 208 533
rect 120 429 149 475
rect 195 429 208 475
rect 120 371 208 429
rect 120 325 149 371
rect 195 325 208 371
rect 120 267 208 325
rect 120 221 149 267
rect 195 221 208 267
rect 120 163 208 221
rect 120 117 149 163
rect 195 117 208 163
rect 120 59 208 117
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 1257 -29 1303
rect -75 1154 -29 1200
rect -75 1051 -29 1097
rect -75 948 -29 994
rect -75 845 -29 891
rect -75 741 -29 787
rect -75 637 -29 683
rect -75 533 -29 579
rect -75 429 -29 475
rect -75 325 -29 371
rect -75 221 -29 267
rect -75 117 -29 163
rect -75 13 -29 59
rect 149 1257 195 1303
rect 149 1154 195 1200
rect 149 1051 195 1097
rect 149 948 195 994
rect 149 845 195 891
rect 149 741 195 787
rect 149 637 195 683
rect 149 533 195 579
rect 149 429 195 475
rect 149 325 195 371
rect 149 221 195 267
rect 149 117 195 163
rect 149 13 195 59
<< polysilicon >>
rect 0 1316 120 1360
rect 0 -44 120 0
<< metal1 >>
rect -75 1303 -29 1316
rect -75 1200 -29 1257
rect -75 1097 -29 1154
rect -75 994 -29 1051
rect -75 891 -29 948
rect -75 787 -29 845
rect -75 683 -29 741
rect -75 579 -29 637
rect -75 475 -29 533
rect -75 371 -29 429
rect -75 267 -29 325
rect -75 163 -29 221
rect -75 59 -29 117
rect -75 0 -29 13
rect 149 1303 195 1316
rect 149 1200 195 1257
rect 149 1097 195 1154
rect 149 994 195 1051
rect 149 891 195 948
rect 149 787 195 845
rect 149 683 195 741
rect 149 579 195 637
rect 149 475 195 533
rect 149 371 195 429
rect 149 267 195 325
rect 149 163 195 221
rect 149 59 195 117
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 658 -52 658 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 658 172 658 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 32490
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 29930
<< end >>
