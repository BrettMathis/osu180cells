magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 4704 844
rect 49 528 95 724
rect 273 611 319 675
rect 466 657 534 724
rect 701 611 747 675
rect 914 657 982 724
rect 1149 611 1195 675
rect 1362 657 1430 724
rect 1597 611 1643 675
rect 1810 657 1878 724
rect 2045 611 2091 675
rect 2258 657 2326 724
rect 2493 611 2539 675
rect 2706 657 2774 724
rect 2941 611 2987 675
rect 3154 657 3222 724
rect 3389 611 3435 675
rect 3602 657 3670 724
rect 3837 611 3883 675
rect 4050 657 4118 724
rect 4285 611 4331 675
rect 273 476 4331 611
rect 4509 528 4555 724
rect 1679 463 2933 476
rect 122 353 1604 430
rect 2206 321 2386 463
rect 2997 353 4475 430
rect 1683 307 2954 321
rect 49 60 95 203
rect 262 173 4351 307
rect 262 146 330 173
rect 721 135 767 173
rect 1169 135 1215 173
rect 1617 135 1663 173
rect 2065 135 2111 173
rect 2513 135 2559 173
rect 2961 135 3007 173
rect 3409 135 3455 173
rect 3857 135 3903 173
rect 4305 135 4351 173
rect 486 60 554 127
rect 934 60 1002 127
rect 1382 60 1450 127
rect 1830 60 1898 127
rect 2278 60 2346 127
rect 2726 60 2794 127
rect 3174 60 3242 127
rect 3622 60 3690 127
rect 4070 60 4138 127
rect 4529 60 4575 203
rect 0 -60 4704 60
<< labels >>
rlabel metal1 s 122 353 1604 430 6 I
port 1 nsew default input
rlabel metal1 s 2997 353 4475 430 6 I
port 1 nsew default input
rlabel metal1 s 4285 611 4331 675 6 ZN
port 2 nsew default output
rlabel metal1 s 3837 611 3883 675 6 ZN
port 2 nsew default output
rlabel metal1 s 3389 611 3435 675 6 ZN
port 2 nsew default output
rlabel metal1 s 2941 611 2987 675 6 ZN
port 2 nsew default output
rlabel metal1 s 2493 611 2539 675 6 ZN
port 2 nsew default output
rlabel metal1 s 2045 611 2091 675 6 ZN
port 2 nsew default output
rlabel metal1 s 1597 611 1643 675 6 ZN
port 2 nsew default output
rlabel metal1 s 1149 611 1195 675 6 ZN
port 2 nsew default output
rlabel metal1 s 701 611 747 675 6 ZN
port 2 nsew default output
rlabel metal1 s 273 611 319 675 6 ZN
port 2 nsew default output
rlabel metal1 s 273 476 4331 611 6 ZN
port 2 nsew default output
rlabel metal1 s 1679 463 2933 476 6 ZN
port 2 nsew default output
rlabel metal1 s 2206 321 2386 463 6 ZN
port 2 nsew default output
rlabel metal1 s 1683 307 2954 321 6 ZN
port 2 nsew default output
rlabel metal1 s 262 173 4351 307 6 ZN
port 2 nsew default output
rlabel metal1 s 4305 146 4351 173 6 ZN
port 2 nsew default output
rlabel metal1 s 3857 146 3903 173 6 ZN
port 2 nsew default output
rlabel metal1 s 3409 146 3455 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2961 146 3007 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2513 146 2559 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2065 146 2111 173 6 ZN
port 2 nsew default output
rlabel metal1 s 1617 146 1663 173 6 ZN
port 2 nsew default output
rlabel metal1 s 1169 146 1215 173 6 ZN
port 2 nsew default output
rlabel metal1 s 721 146 767 173 6 ZN
port 2 nsew default output
rlabel metal1 s 262 146 330 173 6 ZN
port 2 nsew default output
rlabel metal1 s 4305 135 4351 146 6 ZN
port 2 nsew default output
rlabel metal1 s 3857 135 3903 146 6 ZN
port 2 nsew default output
rlabel metal1 s 3409 135 3455 146 6 ZN
port 2 nsew default output
rlabel metal1 s 2961 135 3007 146 6 ZN
port 2 nsew default output
rlabel metal1 s 2513 135 2559 146 6 ZN
port 2 nsew default output
rlabel metal1 s 2065 135 2111 146 6 ZN
port 2 nsew default output
rlabel metal1 s 1617 135 1663 146 6 ZN
port 2 nsew default output
rlabel metal1 s 1169 135 1215 146 6 ZN
port 2 nsew default output
rlabel metal1 s 721 135 767 146 6 ZN
port 2 nsew default output
rlabel metal1 s 0 724 4704 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 657 4555 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4050 657 4118 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3602 657 3670 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3154 657 3222 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2706 657 2774 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2258 657 2326 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1810 657 1878 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1362 657 1430 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 914 657 982 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 466 657 534 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 528 4555 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 528 95 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4529 127 4575 203 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 203 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 60 4575 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4704 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 506656
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 496972
<< end >>
