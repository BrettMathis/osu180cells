magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -143 45 143 50
rect -143 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 143 45
rect -143 -17 143 17
rect -143 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 143 -17
rect -143 -50 143 -45
<< via2 >>
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
<< metal3 >>
rect -143 45 143 50
rect -143 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 143 45
rect -143 -17 143 17
rect -143 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 143 -17
rect -143 -50 143 -45
<< properties >>
string GDS_END 2283700
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2282928
<< end >>
