magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 640 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 520 360
rect 420 252 452 298
rect 498 252 520 298
rect 420 190 520 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 462 1377
rect 508 1143 530 1377
rect 420 1090 530 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 462 1143 508 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
<< psubdiffcont >>
rect 112 52 158 98
<< nsubdiffcont >>
rect 112 1522 158 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 190 990 420 1040
rect 240 800 300 990
rect 210 780 300 800
rect 140 758 300 780
rect 140 712 162 758
rect 208 712 300 758
rect 140 690 300 712
rect 210 680 300 690
rect 240 470 300 680
rect 190 460 300 470
rect 190 400 420 460
rect 190 360 250 400
rect 360 360 420 400
rect 190 140 250 190
rect 360 140 420 190
<< polycontact >>
rect 162 712 208 758
<< metal1 >>
rect 0 1568 640 1620
rect 0 1522 112 1568
rect 158 1566 640 1568
rect 0 1514 114 1522
rect 166 1514 640 1566
rect 0 1470 640 1514
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1060 160 1143
rect 280 1377 330 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 960 330 1143
rect 460 1377 510 1470
rect 460 1143 462 1377
rect 508 1143 510 1377
rect 460 1060 510 1143
rect 280 940 370 960
rect 280 936 400 940
rect 280 884 324 936
rect 376 884 400 936
rect 280 850 400 884
rect 280 820 370 850
rect 130 758 230 760
rect 130 756 162 758
rect 130 704 154 756
rect 208 712 230 758
rect 206 704 230 712
rect 130 670 230 704
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 820
rect 280 252 282 298
rect 328 252 330 298
rect 280 160 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 0 106 640 120
rect 0 98 114 106
rect 0 52 112 98
rect 166 54 640 106
rect 158 52 640 54
rect 0 -30 640 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 114 1514 166 1522
rect 324 884 376 936
rect 154 712 162 756
rect 162 712 206 756
rect 154 704 206 712
rect 114 98 166 106
rect 114 54 158 98
rect 158 54 166 98
<< metal2 >>
rect 100 1570 180 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 100 1470 180 1480
rect 300 936 400 950
rect 300 884 324 936
rect 376 884 400 936
rect 300 840 400 884
rect 130 756 230 770
rect 130 704 154 756
rect 206 704 230 756
rect 130 660 230 704
rect 100 110 180 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 100 10 180 20
<< labels >>
rlabel metal2 s 100 10 180 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 100 1470 180 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 130 660 230 740 4 A
port 1 nsew signal input
rlabel metal2 s 300 840 400 920 4 Y
port 2 nsew signal output
rlabel metal1 s 130 670 230 730 1 A
port 1 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 460 1060 510 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1470 640 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 -30 640 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 820 370 930 1 Y
port 2 nsew signal output
rlabel metal1 s 280 850 400 910 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 640 1590
string GDS_END 174128
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 169808
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
