magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 2800 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
rect 1550 190 1610 360
rect 1720 190 1780 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2230 190 2290 360
rect 2550 190 2610 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 530 700 590 1040
rect 700 700 760 1040
rect 870 700 930 1040
rect 1040 700 1100 1040
rect 1210 700 1270 1040
rect 1380 700 1440 1040
rect 1550 700 1610 1040
rect 1720 700 1780 1040
rect 1890 700 1950 1040
rect 2060 700 2120 1040
rect 2230 700 2290 1040
rect 2550 700 2610 1040
<< ndiff >>
rect 90 258 190 360
rect 90 212 112 258
rect 158 212 190 258
rect 90 190 190 212
rect 250 258 360 360
rect 250 212 282 258
rect 328 212 360 258
rect 250 190 360 212
rect 420 258 530 360
rect 420 212 452 258
rect 498 212 530 258
rect 420 190 530 212
rect 590 258 700 360
rect 590 212 622 258
rect 668 212 700 258
rect 590 190 700 212
rect 760 190 870 360
rect 930 258 1040 360
rect 930 212 962 258
rect 1008 212 1040 258
rect 930 190 1040 212
rect 1100 258 1210 360
rect 1100 212 1132 258
rect 1178 212 1210 258
rect 1100 190 1210 212
rect 1270 258 1380 360
rect 1270 212 1302 258
rect 1348 212 1380 258
rect 1270 190 1380 212
rect 1440 258 1550 360
rect 1440 212 1472 258
rect 1518 212 1550 258
rect 1440 190 1550 212
rect 1610 258 1720 360
rect 1610 212 1642 258
rect 1688 212 1720 258
rect 1610 190 1720 212
rect 1780 190 1890 360
rect 1950 190 2060 360
rect 2120 258 2230 360
rect 2120 212 2152 258
rect 2198 212 2230 258
rect 2120 190 2230 212
rect 2290 258 2390 360
rect 2290 212 2322 258
rect 2368 212 2390 258
rect 2290 190 2390 212
rect 2450 258 2550 360
rect 2450 212 2472 258
rect 2518 212 2550 258
rect 2450 190 2550 212
rect 2610 258 2710 360
rect 2610 212 2642 258
rect 2688 212 2710 258
rect 2610 190 2710 212
<< pdiff >>
rect 90 1013 190 1040
rect 90 967 112 1013
rect 158 967 190 1013
rect 90 700 190 967
rect 250 1013 360 1040
rect 250 967 282 1013
rect 328 967 360 1013
rect 250 700 360 967
rect 420 1013 530 1040
rect 420 967 452 1013
rect 498 967 530 1013
rect 420 700 530 967
rect 590 1018 700 1040
rect 590 972 622 1018
rect 668 972 700 1018
rect 590 700 700 972
rect 760 700 870 1040
rect 930 1013 1040 1040
rect 930 967 962 1013
rect 1008 967 1040 1013
rect 930 700 1040 967
rect 1100 1013 1210 1040
rect 1100 967 1132 1013
rect 1178 967 1210 1013
rect 1100 700 1210 967
rect 1270 1013 1380 1040
rect 1270 967 1302 1013
rect 1348 967 1380 1013
rect 1270 700 1380 967
rect 1440 1013 1550 1040
rect 1440 967 1472 1013
rect 1518 967 1550 1013
rect 1440 700 1550 967
rect 1610 883 1720 1040
rect 1610 837 1642 883
rect 1688 837 1720 883
rect 1610 700 1720 837
rect 1780 700 1890 1040
rect 1950 700 2060 1040
rect 2120 1013 2230 1040
rect 2120 967 2152 1013
rect 2198 967 2230 1013
rect 2120 700 2230 967
rect 2290 1013 2390 1040
rect 2290 967 2322 1013
rect 2368 967 2390 1013
rect 2290 700 2390 967
rect 2450 1013 2550 1040
rect 2450 967 2472 1013
rect 2518 967 2550 1013
rect 2450 700 2550 967
rect 2610 1013 2710 1040
rect 2610 967 2642 1013
rect 2688 967 2710 1013
rect 2610 700 2710 967
<< ndiffc >>
rect 112 212 158 258
rect 282 212 328 258
rect 452 212 498 258
rect 622 212 668 258
rect 962 212 1008 258
rect 1132 212 1178 258
rect 1302 212 1348 258
rect 1472 212 1518 258
rect 1642 212 1688 258
rect 2152 212 2198 258
rect 2322 212 2368 258
rect 2472 212 2518 258
rect 2642 212 2688 258
<< pdiffc >>
rect 112 967 158 1013
rect 282 967 328 1013
rect 452 967 498 1013
rect 622 972 668 1018
rect 962 967 1008 1013
rect 1132 967 1178 1013
rect 1302 967 1348 1013
rect 1472 967 1518 1013
rect 1642 837 1688 883
rect 2152 967 2198 1013
rect 2322 967 2368 1013
rect 2472 967 2518 1013
rect 2642 967 2688 1013
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
rect 1290 1178 1380 1200
rect 1290 1132 1312 1178
rect 1358 1132 1380 1178
rect 1290 1110 1380 1132
rect 1530 1178 1620 1200
rect 1530 1132 1552 1178
rect 1598 1132 1620 1178
rect 1530 1110 1620 1132
rect 1770 1178 1860 1200
rect 1770 1132 1792 1178
rect 1838 1132 1860 1178
rect 1770 1110 1860 1132
rect 2010 1178 2100 1200
rect 2010 1132 2032 1178
rect 2078 1132 2100 1178
rect 2010 1110 2100 1132
rect 2250 1178 2340 1200
rect 2250 1132 2272 1178
rect 2318 1132 2340 1178
rect 2250 1110 2340 1132
rect 2490 1178 2580 1200
rect 2490 1132 2512 1178
rect 2558 1132 2580 1178
rect 2490 1110 2580 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
rect 1312 1132 1358 1178
rect 1552 1132 1598 1178
rect 1792 1132 1838 1178
rect 2032 1132 2078 1178
rect 2272 1132 2318 1178
rect 2512 1132 2558 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 870 1040 930 1090
rect 1040 1040 1100 1090
rect 1210 1040 1270 1090
rect 1380 1040 1440 1090
rect 1550 1040 1610 1090
rect 1720 1040 1780 1090
rect 1890 1040 1950 1090
rect 2060 1040 2120 1090
rect 2230 1040 2290 1090
rect 2550 1040 2610 1090
rect 190 520 250 700
rect 360 650 420 700
rect 300 623 420 650
rect 300 577 327 623
rect 373 577 420 623
rect 300 550 420 577
rect 120 493 250 520
rect 120 447 147 493
rect 193 447 250 493
rect 120 420 250 447
rect 190 360 250 420
rect 360 360 420 550
rect 530 520 590 700
rect 700 680 760 700
rect 870 680 930 700
rect 1040 680 1100 700
rect 1210 680 1270 700
rect 700 653 820 680
rect 700 607 747 653
rect 793 607 820 653
rect 700 580 820 607
rect 870 630 1100 680
rect 1150 653 1270 680
rect 510 493 610 520
rect 510 447 537 493
rect 583 447 610 493
rect 510 420 610 447
rect 530 360 590 420
rect 700 360 760 580
rect 870 550 930 630
rect 1150 607 1177 653
rect 1223 607 1270 653
rect 1150 580 1270 607
rect 870 523 1020 550
rect 870 477 947 523
rect 993 477 1020 523
rect 870 450 1020 477
rect 870 400 1100 450
rect 870 360 930 400
rect 1040 360 1100 400
rect 1210 360 1270 580
rect 1380 550 1440 700
rect 1550 550 1610 700
rect 1720 550 1780 700
rect 1890 680 1950 700
rect 1890 653 2010 680
rect 1890 607 1937 653
rect 1983 607 2010 653
rect 1890 580 2010 607
rect 1380 523 1490 550
rect 1380 477 1417 523
rect 1463 477 1490 523
rect 1380 450 1490 477
rect 1550 523 1660 550
rect 1550 477 1587 523
rect 1633 477 1660 523
rect 1550 450 1660 477
rect 1720 523 1840 550
rect 1720 477 1767 523
rect 1813 477 1840 523
rect 1720 450 1840 477
rect 1380 360 1440 450
rect 1550 360 1610 450
rect 1720 360 1780 450
rect 1890 360 1950 580
rect 2060 530 2120 700
rect 2230 550 2290 700
rect 2550 550 2610 700
rect 2020 503 2120 530
rect 2020 457 2047 503
rect 2093 457 2120 503
rect 2020 430 2120 457
rect 2170 523 2290 550
rect 2170 477 2197 523
rect 2243 477 2290 523
rect 2170 450 2290 477
rect 2490 523 2610 550
rect 2490 477 2517 523
rect 2563 477 2610 523
rect 2490 450 2610 477
rect 2060 360 2120 430
rect 2230 360 2290 450
rect 2550 360 2610 450
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
rect 1550 140 1610 190
rect 1720 140 1780 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2230 140 2290 190
rect 2550 140 2610 190
<< polycontact >>
rect 327 577 373 623
rect 147 447 193 493
rect 747 607 793 653
rect 537 447 583 493
rect 1177 607 1223 653
rect 947 477 993 523
rect 1937 607 1983 653
rect 1417 477 1463 523
rect 1587 477 1633 523
rect 1767 477 1813 523
rect 2047 457 2093 503
rect 2197 477 2243 523
rect 2517 477 2563 523
<< metal1 >>
rect 0 1178 2800 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1312 1178
rect 1358 1176 1552 1178
rect 1598 1176 1792 1178
rect 1838 1176 2032 1178
rect 2078 1176 2272 1178
rect 2318 1176 2512 1178
rect 2558 1176 2800 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 1126 1132 1312 1176
rect 1366 1132 1552 1176
rect 1606 1132 1792 1176
rect 1846 1132 2032 1176
rect 2086 1132 2272 1176
rect 2326 1132 2512 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1314 1132
rect 1366 1124 1554 1132
rect 1606 1124 1794 1132
rect 1846 1124 2034 1132
rect 2086 1124 2274 1132
rect 2326 1124 2514 1132
rect 2566 1124 2800 1176
rect 0 1110 2800 1124
rect 110 1013 160 1040
rect 110 967 112 1013
rect 158 967 160 1013
rect 110 890 160 967
rect 280 1013 330 1110
rect 280 967 282 1013
rect 328 967 330 1013
rect 280 940 330 967
rect 450 1013 500 1040
rect 450 967 452 1013
rect 498 967 500 1013
rect 450 890 500 967
rect 620 1018 680 1040
rect 620 972 622 1018
rect 668 1016 680 1018
rect 620 964 624 972
rect 676 964 680 1016
rect 620 940 680 964
rect 960 1013 1010 1110
rect 960 967 962 1013
rect 1008 967 1010 1013
rect 960 940 1010 967
rect 1130 1013 1180 1040
rect 1130 967 1132 1013
rect 1178 967 1180 1013
rect 110 840 500 890
rect 1130 890 1180 967
rect 1300 1013 1350 1110
rect 1300 967 1302 1013
rect 1348 967 1350 1013
rect 1300 940 1350 967
rect 1470 1013 1520 1040
rect 1470 967 1472 1013
rect 1518 967 1520 1013
rect 1470 890 1520 967
rect 2150 1013 2200 1110
rect 2150 967 2152 1013
rect 2198 967 2200 1013
rect 2150 940 2200 967
rect 2320 1013 2370 1040
rect 2320 967 2322 1013
rect 2368 967 2370 1013
rect 1130 840 1520 890
rect 1620 886 1720 890
rect 1620 883 1644 886
rect 1620 837 1642 883
rect 1620 834 1644 837
rect 1696 834 1720 886
rect 1620 830 1720 834
rect 320 730 800 790
rect 320 626 380 730
rect 320 574 324 626
rect 376 574 380 626
rect 320 550 380 574
rect 430 620 690 680
rect 430 500 480 620
rect 640 530 690 620
rect 740 660 800 730
rect 1170 720 1990 780
rect 1170 660 1230 720
rect 740 653 1230 660
rect 740 607 747 653
rect 793 607 1177 653
rect 1223 607 1230 653
rect 740 600 1230 607
rect 740 580 800 600
rect 1170 580 1230 600
rect 1280 610 1820 670
rect 1280 530 1340 610
rect 640 523 1340 530
rect 120 496 480 500
rect 120 444 144 496
rect 196 444 480 496
rect 120 440 480 444
rect 530 496 590 520
rect 530 444 534 496
rect 586 444 590 496
rect 640 477 947 523
rect 993 477 1340 523
rect 640 470 1340 477
rect 1410 523 1470 550
rect 1760 530 1820 610
rect 1930 653 1990 720
rect 1930 607 1937 653
rect 1983 607 1990 653
rect 1930 580 1990 607
rect 2320 670 2370 967
rect 2470 1013 2520 1110
rect 2470 967 2472 1013
rect 2518 967 2520 1013
rect 2470 940 2520 967
rect 2640 1013 2690 1040
rect 2640 967 2642 1013
rect 2688 967 2690 1013
rect 2640 670 2690 967
rect 2320 660 2380 670
rect 2640 660 2730 670
rect 2320 656 2410 660
rect 2320 604 2334 656
rect 2386 604 2410 656
rect 2320 600 2410 604
rect 2640 656 2750 660
rect 2640 604 2674 656
rect 2726 604 2750 656
rect 2640 600 2750 604
rect 2320 590 2380 600
rect 2640 590 2730 600
rect 1410 477 1417 523
rect 1463 477 1470 523
rect 530 420 590 444
rect 1410 420 1470 477
rect 1560 526 1660 530
rect 1560 474 1584 526
rect 1636 474 1660 526
rect 1560 470 1660 474
rect 1740 523 1840 530
rect 1740 477 1767 523
rect 1813 477 1840 523
rect 2170 526 2270 530
rect 1740 470 1840 477
rect 1950 503 2120 510
rect 1950 457 2047 503
rect 2093 457 2120 503
rect 2170 474 2194 526
rect 2246 474 2270 526
rect 2170 470 2270 474
rect 1950 450 2120 457
rect 1950 420 2010 450
rect 530 360 2010 420
rect 100 266 160 290
rect 100 214 104 266
rect 156 258 160 266
rect 100 212 112 214
rect 158 212 160 258
rect 100 190 160 212
rect 280 258 330 280
rect 280 212 282 258
rect 328 212 330 258
rect 280 120 330 212
rect 440 266 500 290
rect 440 214 444 266
rect 496 258 500 266
rect 440 212 452 214
rect 498 212 500 258
rect 440 190 500 212
rect 620 266 680 290
rect 620 258 624 266
rect 620 212 622 258
rect 676 214 680 266
rect 668 212 680 214
rect 620 190 680 212
rect 960 258 1010 280
rect 960 212 962 258
rect 1008 212 1010 258
rect 960 120 1010 212
rect 1130 266 1190 290
rect 1130 258 1134 266
rect 1130 212 1132 258
rect 1186 214 1190 266
rect 1178 212 1190 214
rect 1130 190 1190 212
rect 1300 258 1350 280
rect 1300 212 1302 258
rect 1348 212 1350 258
rect 1300 120 1350 212
rect 1460 266 1520 290
rect 1460 214 1464 266
rect 1516 258 1520 266
rect 1460 212 1472 214
rect 1518 212 1520 258
rect 1460 190 1520 212
rect 1640 266 1700 290
rect 1640 258 1644 266
rect 1640 212 1642 258
rect 1696 214 1700 266
rect 1688 212 1700 214
rect 1640 190 1700 212
rect 2150 258 2200 280
rect 2150 212 2152 258
rect 2198 212 2200 258
rect 2150 120 2200 212
rect 2320 258 2370 590
rect 2490 526 2590 530
rect 2490 474 2514 526
rect 2566 474 2590 526
rect 2490 470 2590 474
rect 2320 212 2322 258
rect 2368 212 2370 258
rect 2320 190 2370 212
rect 2470 258 2520 280
rect 2470 212 2472 258
rect 2518 212 2520 258
rect 2470 120 2520 212
rect 2640 258 2690 590
rect 2640 212 2642 258
rect 2688 212 2690 258
rect 2640 190 2690 212
rect 0 106 2800 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2800 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2800 54
rect 0 0 2800 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 1314 1132 1358 1176
rect 1358 1132 1366 1176
rect 1554 1132 1598 1176
rect 1598 1132 1606 1176
rect 1794 1132 1838 1176
rect 1838 1132 1846 1176
rect 2034 1132 2078 1176
rect 2078 1132 2086 1176
rect 2274 1132 2318 1176
rect 2318 1132 2326 1176
rect 2514 1132 2558 1176
rect 2558 1132 2566 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 1554 1124 1606 1132
rect 1794 1124 1846 1132
rect 2034 1124 2086 1132
rect 2274 1124 2326 1132
rect 2514 1124 2566 1132
rect 624 972 668 1016
rect 668 972 676 1016
rect 624 964 676 972
rect 1644 883 1696 886
rect 1644 837 1688 883
rect 1688 837 1696 883
rect 1644 834 1696 837
rect 324 623 376 626
rect 324 577 327 623
rect 327 577 373 623
rect 373 577 376 623
rect 324 574 376 577
rect 144 493 196 496
rect 144 447 147 493
rect 147 447 193 493
rect 193 447 196 493
rect 144 444 196 447
rect 534 493 586 496
rect 534 447 537 493
rect 537 447 583 493
rect 583 447 586 493
rect 534 444 586 447
rect 2334 604 2386 656
rect 2674 604 2726 656
rect 1584 523 1636 526
rect 1584 477 1587 523
rect 1587 477 1633 523
rect 1633 477 1636 523
rect 1584 474 1636 477
rect 2194 523 2246 526
rect 2194 477 2197 523
rect 2197 477 2243 523
rect 2243 477 2246 523
rect 2194 474 2246 477
rect 104 258 156 266
rect 104 214 112 258
rect 112 214 156 258
rect 444 258 496 266
rect 444 214 452 258
rect 452 214 496 258
rect 624 258 676 266
rect 624 214 668 258
rect 668 214 676 258
rect 1134 258 1186 266
rect 1134 214 1178 258
rect 1178 214 1186 258
rect 1464 258 1516 266
rect 1464 214 1472 258
rect 1472 214 1516 258
rect 1644 258 1696 266
rect 1644 214 1688 258
rect 1688 214 1696 258
rect 2514 523 2566 526
rect 2514 477 2517 523
rect 2517 477 2563 523
rect 2563 477 2566 523
rect 2514 474 2566 477
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 1540 1180 1620 1190
rect 1780 1180 1860 1190
rect 2020 1180 2100 1190
rect 2260 1180 2340 1190
rect 2500 1180 2580 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 1530 1176 1630 1180
rect 1530 1124 1554 1176
rect 1606 1124 1630 1176
rect 1530 1120 1630 1124
rect 1770 1176 1870 1180
rect 1770 1124 1794 1176
rect 1846 1124 1870 1176
rect 1770 1120 1870 1124
rect 2010 1176 2110 1180
rect 2010 1124 2034 1176
rect 2086 1124 2110 1176
rect 2010 1120 2110 1124
rect 2250 1176 2350 1180
rect 2250 1124 2274 1176
rect 2326 1124 2350 1176
rect 2250 1120 2350 1124
rect 2490 1176 2590 1180
rect 2490 1124 2514 1176
rect 2566 1124 2590 1176
rect 2490 1120 2590 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 1540 1110 1620 1120
rect 1780 1110 1860 1120
rect 2020 1110 2100 1120
rect 2260 1110 2340 1120
rect 2500 1110 2580 1120
rect 620 1030 680 1040
rect 610 1020 690 1030
rect 600 1016 2570 1020
rect 600 964 624 1016
rect 676 964 2570 1016
rect 600 960 2570 964
rect 610 950 690 960
rect 310 630 390 640
rect 300 626 400 630
rect 300 574 324 626
rect 376 574 400 626
rect 300 570 400 574
rect 310 560 390 570
rect 750 530 810 960
rect 1630 890 1710 900
rect 1620 886 2250 890
rect 1620 834 1644 886
rect 1696 834 2250 886
rect 1620 830 2250 834
rect 1630 820 1710 830
rect 1570 530 1650 540
rect 750 526 1660 530
rect 120 496 220 510
rect 520 500 600 510
rect 120 444 144 496
rect 196 444 220 496
rect 120 430 220 444
rect 510 496 610 500
rect 510 444 534 496
rect 586 444 610 496
rect 510 440 610 444
rect 750 474 1584 526
rect 1636 474 1660 526
rect 750 470 1660 474
rect 520 430 600 440
rect 100 280 160 290
rect 440 280 500 290
rect 620 280 680 290
rect 90 270 170 280
rect 430 270 510 280
rect 90 266 510 270
rect 90 214 104 266
rect 156 214 444 266
rect 496 214 510 266
rect 90 210 510 214
rect 90 200 170 210
rect 430 200 510 210
rect 610 270 690 280
rect 750 270 810 470
rect 1570 460 1650 470
rect 1130 280 1190 290
rect 1460 280 1520 290
rect 610 266 810 270
rect 610 214 624 266
rect 676 214 810 266
rect 610 210 810 214
rect 1120 270 1200 280
rect 1450 270 1530 280
rect 1630 270 1710 280
rect 1770 270 1830 830
rect 2190 540 2250 830
rect 2320 660 2400 670
rect 2310 656 2410 660
rect 2310 604 2334 656
rect 2386 604 2410 656
rect 2310 600 2410 604
rect 2320 590 2400 600
rect 2510 540 2570 960
rect 2660 660 2740 670
rect 2650 656 2750 660
rect 2650 604 2674 656
rect 2726 604 2750 656
rect 2650 600 2750 604
rect 2660 590 2740 600
rect 2180 526 2260 540
rect 2500 530 2580 540
rect 2180 474 2194 526
rect 2246 474 2260 526
rect 2180 460 2260 474
rect 2490 526 2590 530
rect 2490 474 2514 526
rect 2566 474 2590 526
rect 2490 470 2590 474
rect 2500 460 2580 470
rect 2190 450 2250 460
rect 2510 450 2570 460
rect 1120 266 1530 270
rect 1120 214 1134 266
rect 1186 214 1464 266
rect 1516 214 1530 266
rect 1120 210 1530 214
rect 1620 266 1830 270
rect 1620 214 1644 266
rect 1696 214 1830 266
rect 1620 210 1830 214
rect 610 200 690 210
rect 1120 200 1200 210
rect 1450 200 1530 210
rect 1630 200 1710 210
rect 100 190 160 200
rect 440 190 500 200
rect 620 190 680 200
rect 1130 190 1190 200
rect 1460 190 1520 200
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 50 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 50 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 50 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 50 2590 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
rect 1780 40 1860 50
rect 2020 40 2100 50
rect 2260 40 2340 50
rect 2500 40 2580 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 120 430 220 510 4 A
port 1 nsew signal input
rlabel metal2 s 310 560 390 640 4 B
port 2 nsew signal input
rlabel metal2 s 520 430 600 510 4 CI
port 3 nsew signal input
rlabel metal2 s 2320 590 2400 670 4 S
port 4 nsew signal output
rlabel metal2 s 2660 590 2740 670 4 CO
port 5 nsew signal output
rlabel metal1 s 120 440 480 500 1 A
port 1 nsew signal input
rlabel metal1 s 430 440 480 680 1 A
port 1 nsew signal input
rlabel metal1 s 640 470 690 680 1 A
port 1 nsew signal input
rlabel metal1 s 430 620 690 680 1 A
port 1 nsew signal input
rlabel metal1 s 640 470 1340 530 1 A
port 1 nsew signal input
rlabel metal1 s 1280 470 1340 670 1 A
port 1 nsew signal input
rlabel metal1 s 1760 470 1820 670 1 A
port 1 nsew signal input
rlabel metal1 s 1280 610 1820 670 1 A
port 1 nsew signal input
rlabel metal1 s 1740 470 1840 530 1 A
port 1 nsew signal input
rlabel metal2 s 300 570 400 630 1 B
port 2 nsew signal input
rlabel metal1 s 320 550 380 790 1 B
port 2 nsew signal input
rlabel metal1 s 740 580 800 790 1 B
port 2 nsew signal input
rlabel metal1 s 320 730 800 790 1 B
port 2 nsew signal input
rlabel metal1 s 740 600 1230 660 1 B
port 2 nsew signal input
rlabel metal1 s 1170 580 1230 780 1 B
port 2 nsew signal input
rlabel metal1 s 1930 580 1990 780 1 B
port 2 nsew signal input
rlabel metal1 s 1170 720 1990 780 1 B
port 2 nsew signal input
rlabel metal2 s 510 440 610 500 1 CI
port 3 nsew signal input
rlabel metal1 s 530 360 590 520 1 CI
port 3 nsew signal input
rlabel metal1 s 1410 360 1470 550 1 CI
port 3 nsew signal input
rlabel metal1 s 530 360 2010 420 1 CI
port 3 nsew signal input
rlabel metal1 s 1950 360 2010 510 1 CI
port 3 nsew signal input
rlabel metal1 s 1950 450 2120 510 1 CI
port 3 nsew signal input
rlabel metal2 s 2650 600 2750 660 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 190 2690 1040 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 590 2730 670 1 CO
port 5 nsew signal output
rlabel metal1 s 2640 600 2750 660 1 CO
port 5 nsew signal output
rlabel metal2 s 2310 600 2410 660 1 S
port 4 nsew signal output
rlabel metal1 s 2320 190 2370 1040 1 S
port 4 nsew signal output
rlabel metal1 s 2320 590 2380 670 1 S
port 4 nsew signal output
rlabel metal1 s 2320 600 2410 660 1 S
port 4 nsew signal output
rlabel metal2 s 90 1120 190 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1540 1110 1620 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1530 1120 1630 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1780 1110 1860 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 1770 1120 1870 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2020 1110 2100 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2010 1120 2110 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2260 1110 2340 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2250 1120 2350 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2500 1110 2580 1190 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 2490 1120 2590 1180 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 280 940 330 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 960 940 1010 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 1300 940 1350 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 2150 940 2200 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 2470 940 2520 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal1 s 0 1110 2800 1230 1 VDD
port 12 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1780 40 1860 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 1770 50 1870 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2020 40 2100 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2010 50 2110 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2260 40 2340 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2250 50 2350 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2500 40 2580 120 1 VSS
port 13 nsew ground bidirectional
rlabel metal2 s 2490 50 2590 110 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 280 0 330 280 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 960 0 1010 280 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 1300 0 1350 280 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 2150 0 2200 280 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 2470 0 2520 280 1 VSS
port 13 nsew ground bidirectional
rlabel metal1 s 0 0 2800 120 1 VSS
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2800 1230
string GDS_END 26072
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 134
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
