magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 111 300 123
rect 11 70 16 111
rect 28 65 33 104
rect 45 70 50 111
rect 62 65 67 104
rect 79 70 84 111
rect 96 65 101 104
rect 113 70 118 111
rect 130 65 135 104
rect 147 70 152 111
rect 164 65 169 104
rect 181 70 186 111
rect 198 65 203 104
rect 215 70 220 111
rect 232 65 237 104
rect 249 70 254 111
rect 266 76 271 104
rect 266 70 277 76
rect 283 70 288 111
rect 266 65 271 70
rect 28 60 271 65
rect 8 44 18 50
rect 28 46 33 60
rect 62 46 67 60
rect 96 46 101 60
rect 130 46 135 60
rect 164 46 169 60
rect 198 46 203 60
rect 232 46 237 60
rect 266 46 271 60
rect 28 41 271 46
rect 11 12 16 36
rect 28 19 33 41
rect 45 12 50 36
rect 62 19 67 41
rect 79 12 84 36
rect 96 19 101 41
rect 113 12 118 36
rect 130 19 135 41
rect 147 12 152 36
rect 164 19 169 41
rect 181 12 186 36
rect 198 19 203 41
rect 215 12 220 36
rect 232 19 237 41
rect 249 12 254 36
rect 266 19 271 41
rect 283 12 288 36
rect 0 0 300 12
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 274 118 282 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 177 112 187 118
rect 201 112 211 118
rect 225 112 235 118
rect 249 112 259 118
rect 273 112 283 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 274 111 282 112
rect 268 76 276 77
rect 267 70 277 76
rect 268 69 276 70
rect 8 43 18 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 274 11 282 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 273 5 283 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
rect 274 4 282 5
<< labels >>
rlabel metal2 s 8 43 18 51 6 A
port 1 nsew signal input
rlabel metal1 s 8 44 18 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 178 111 186 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 177 112 187 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 202 111 210 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 201 112 211 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 226 111 234 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 225 112 235 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 250 111 258 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 249 112 259 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 274 111 282 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 273 112 283 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 45 70 50 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 79 70 84 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 113 70 118 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 147 70 152 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 181 70 186 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 215 70 220 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 249 70 254 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 283 70 288 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 300 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 274 4 282 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 273 5 283 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 0 50 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 79 0 84 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 113 0 118 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 147 0 152 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 181 0 186 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 215 0 220 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 249 0 254 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 283 0 288 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 300 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 268 69 276 77 6 Y
port 2 nsew signal output
rlabel metal2 s 267 70 277 76 6 Y
port 2 nsew signal output
rlabel metal1 s 28 19 33 104 6 Y
port 2 nsew signal output
rlabel metal1 s 62 19 67 104 6 Y
port 2 nsew signal output
rlabel metal1 s 96 19 101 104 6 Y
port 2 nsew signal output
rlabel metal1 s 130 19 135 104 6 Y
port 2 nsew signal output
rlabel metal1 s 164 19 169 104 6 Y
port 2 nsew signal output
rlabel metal1 s 198 19 203 104 6 Y
port 2 nsew signal output
rlabel metal1 s 232 19 237 104 6 Y
port 2 nsew signal output
rlabel metal1 s 28 41 271 46 6 Y
port 2 nsew signal output
rlabel metal1 s 28 60 271 65 6 Y
port 2 nsew signal output
rlabel metal1 s 266 19 271 104 6 Y
port 2 nsew signal output
rlabel metal1 s 266 70 277 76 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 300 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 221814
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 199254
<< end >>
