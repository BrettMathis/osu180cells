magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -221 -1615 221 1615
<< nsubdiff >>
rect -77 1411 77 1467
rect -77 1365 -23 1411
rect 23 1365 77 1411
rect -77 1247 77 1365
rect -77 1201 -23 1247
rect 23 1201 77 1247
rect -77 1084 77 1201
rect -77 1038 -23 1084
rect 23 1038 77 1084
rect -77 921 77 1038
rect -77 875 -23 921
rect 23 875 77 921
rect -77 758 77 875
rect -77 712 -23 758
rect 23 712 77 758
rect -77 595 77 712
rect -77 549 -23 595
rect 23 549 77 595
rect -77 431 77 549
rect -77 385 -23 431
rect 23 385 77 431
rect -77 268 77 385
rect -77 222 -23 268
rect 23 222 77 268
rect -77 105 77 222
rect -77 59 -23 105
rect 23 59 77 105
rect -77 -59 77 59
rect -77 -105 -23 -59
rect 23 -105 77 -59
rect -77 -222 77 -105
rect -77 -268 -23 -222
rect 23 -268 77 -222
rect -77 -385 77 -268
rect -77 -431 -23 -385
rect 23 -431 77 -385
rect -77 -549 77 -431
rect -77 -595 -23 -549
rect 23 -595 77 -549
rect -77 -712 77 -595
rect -77 -758 -23 -712
rect 23 -758 77 -712
rect -77 -875 77 -758
rect -77 -921 -23 -875
rect 23 -921 77 -875
rect -77 -1038 77 -921
rect -77 -1084 -23 -1038
rect 23 -1084 77 -1038
rect -77 -1201 77 -1084
rect -77 -1247 -23 -1201
rect 23 -1247 77 -1201
rect -77 -1365 77 -1247
rect -77 -1411 -23 -1365
rect 23 -1411 77 -1365
rect -77 -1468 77 -1411
<< nsubdiffcont >>
rect -23 1365 23 1411
rect -23 1201 23 1247
rect -23 1038 23 1084
rect -23 875 23 921
rect -23 712 23 758
rect -23 549 23 595
rect -23 385 23 431
rect -23 222 23 268
rect -23 59 23 105
rect -23 -105 23 -59
rect -23 -268 23 -222
rect -23 -431 23 -385
rect -23 -595 23 -549
rect -23 -758 23 -712
rect -23 -921 23 -875
rect -23 -1084 23 -1038
rect -23 -1247 23 -1201
rect -23 -1411 23 -1365
<< metal1 >>
rect -58 1411 58 1447
rect -58 1365 -23 1411
rect 23 1365 58 1411
rect -58 1247 58 1365
rect -58 1201 -23 1247
rect 23 1201 58 1247
rect -58 1084 58 1201
rect -58 1038 -23 1084
rect 23 1038 58 1084
rect -58 921 58 1038
rect -58 875 -23 921
rect 23 875 58 921
rect -58 758 58 875
rect -58 712 -23 758
rect 23 712 58 758
rect -58 595 58 712
rect -58 549 -23 595
rect 23 549 58 595
rect -58 431 58 549
rect -58 385 -23 431
rect 23 385 58 431
rect -58 268 58 385
rect -58 222 -23 268
rect 23 222 58 268
rect -58 105 58 222
rect -58 59 -23 105
rect 23 59 58 105
rect -58 -59 58 59
rect -58 -105 -23 -59
rect 23 -105 58 -59
rect -58 -222 58 -105
rect -58 -268 -23 -222
rect 23 -268 58 -222
rect -58 -385 58 -268
rect -58 -431 -23 -385
rect 23 -431 58 -385
rect -58 -549 58 -431
rect -58 -595 -23 -549
rect 23 -595 58 -549
rect -58 -712 58 -595
rect -58 -758 -23 -712
rect 23 -758 58 -712
rect -58 -875 58 -758
rect -58 -921 -23 -875
rect 23 -921 58 -875
rect -58 -1038 58 -921
rect -58 -1084 -23 -1038
rect 23 -1084 58 -1038
rect -58 -1201 58 -1084
rect -58 -1247 -23 -1201
rect 23 -1247 58 -1201
rect -58 -1365 58 -1247
rect -58 -1411 -23 -1365
rect 23 -1411 58 -1365
rect -58 -1447 58 -1411
<< properties >>
string GDS_END 268830
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 267418
<< end >>
