magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal3 >>
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
<< via3 >>
rect 128 64888 288 64944
rect 128 64776 288 64832
rect 128 64664 288 64720
rect 128 64552 288 64608
rect 128 64440 288 64496
rect 128 64328 288 64384
rect 128 64216 288 64272
rect 128 64104 288 64160
rect 128 63992 288 64048
rect 128 63880 288 63936
rect 128 63768 288 63824
rect 128 63656 288 63712
rect 125 50482 181 50538
rect 237 50482 293 50538
rect 125 50370 181 50426
rect 237 50370 293 50426
rect 125 50258 181 50314
rect 237 50258 293 50314
rect 125 50146 181 50202
rect 237 50146 293 50202
rect 125 50034 181 50090
rect 237 50034 293 50090
rect 125 49922 181 49978
rect 237 49922 293 49978
rect 125 49810 181 49866
rect 237 49810 293 49866
rect 125 49698 181 49754
rect 237 49698 293 49754
rect 125 49586 181 49642
rect 237 49586 293 49642
rect 125 49474 181 49530
rect 237 49474 293 49530
rect 125 49362 181 49418
rect 237 49362 293 49418
rect 125 49250 181 49306
rect 237 49250 293 49306
<< metal4 >>
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
use GF_NI_BRK2_0  GF_NI_BRK2_0_0
timestamp 1669390400
transform 1 0 0 0 1 0
box -32 13097 432 69968
use M4_M3_CDNS_40661954729301  M4_M3_CDNS_40661954729301_0
timestamp 1669390400
transform 1 0 209 0 1 49894
box 0 0 1 1
use M4_M3_CDNS_40661954729302  M4_M3_CDNS_40661954729302_0
timestamp 1669390400
transform 1 0 208 0 1 64300
box 0 0 1 1
<< labels >>
rlabel metal3 s 0 63600 400 65000 4 VSS
port 1 nsew ground bidirectional
rlabel metal4 s 0 63600 400 65000 4 VSS
port 1 nsew ground bidirectional
rlabel metal4 s 0 49200 400 50600 4 VSS
port 1 nsew ground bidirectional
rlabel metal3 s 0 49200 400 50600 4 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 400 70000
string GDS_END 3287678
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3286952
string LEFclass PAD
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
