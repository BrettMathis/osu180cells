magic
tech gf180mcuA
timestamp 1669390400
<< properties >>
string GDS_END 902356
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 901584
<< end >>
