magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -81 447 81 453
rect -81 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 81 447
rect -81 385 81 421
rect -81 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 81 385
rect -81 323 81 359
rect -81 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 81 323
rect -81 261 81 297
rect -81 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 81 261
rect -81 199 81 235
rect -81 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 81 199
rect -81 137 81 173
rect -81 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 81 137
rect -81 75 81 111
rect -81 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 81 75
rect -81 13 81 49
rect -81 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 81 13
rect -81 -49 81 -13
rect -81 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 81 -49
rect -81 -111 81 -75
rect -81 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 81 -111
rect -81 -173 81 -137
rect -81 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 81 -173
rect -81 -235 81 -199
rect -81 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 81 -235
rect -81 -297 81 -261
rect -81 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 81 -297
rect -81 -359 81 -323
rect -81 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 81 -359
rect -81 -421 81 -385
rect -81 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 81 -421
rect -81 -453 81 -447
<< via1 >>
rect -75 421 -49 447
rect -13 421 13 447
rect 49 421 75 447
rect -75 359 -49 385
rect -13 359 13 385
rect 49 359 75 385
rect -75 297 -49 323
rect -13 297 13 323
rect 49 297 75 323
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect -75 -323 -49 -297
rect -13 -323 13 -297
rect 49 -323 75 -297
rect -75 -385 -49 -359
rect -13 -385 13 -359
rect 49 -385 75 -359
rect -75 -447 -49 -421
rect -13 -447 13 -421
rect 49 -447 75 -421
<< metal2 >>
rect -81 447 81 453
rect -81 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 81 447
rect -81 385 81 421
rect -81 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 81 385
rect -81 323 81 359
rect -81 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 81 323
rect -81 261 81 297
rect -81 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 81 261
rect -81 199 81 235
rect -81 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 81 199
rect -81 137 81 173
rect -81 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 81 137
rect -81 75 81 111
rect -81 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 81 75
rect -81 13 81 49
rect -81 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 81 13
rect -81 -49 81 -13
rect -81 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 81 -49
rect -81 -111 81 -75
rect -81 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 81 -111
rect -81 -173 81 -137
rect -81 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 81 -173
rect -81 -235 81 -199
rect -81 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 81 -235
rect -81 -297 81 -261
rect -81 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 81 -297
rect -81 -359 81 -323
rect -81 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 81 -359
rect -81 -421 81 -385
rect -81 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 81 -421
rect -81 -453 81 -447
<< properties >>
string GDS_END 785792
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 782780
<< end >>
