magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 1342 23867 22665 29129
rect 1216 17407 22310 19961
rect 22338 17406 22926 19961
rect 22827 14326 23842 15917
rect 22880 8391 23005 9181
<< mvpmos >>
rect 6089 27950 6209 28632
rect 6314 27950 6434 28632
rect 6780 27950 6900 28632
rect 7005 27950 7125 28632
rect 16889 27950 17009 28632
rect 17114 27950 17234 28632
rect 17580 27950 17700 28632
rect 17805 27950 17925 28632
rect 6089 27175 6209 27857
rect 6314 27175 6434 27857
rect 6780 27175 6900 27857
rect 7005 27175 7125 27857
rect 16889 27175 17009 27857
rect 17114 27175 17234 27857
rect 17580 27175 17700 27857
rect 17805 27175 17925 27857
<< mvpdiff >>
rect 5983 27950 6089 28632
rect 6209 27950 6314 28632
rect 6434 27950 6540 28632
rect 6674 27950 6780 28632
rect 6900 27950 7005 28632
rect 7125 27950 7231 28632
rect 16783 27950 16889 28632
rect 17009 27950 17114 28632
rect 17234 27950 17340 28632
rect 17474 27950 17580 28632
rect 17700 27950 17805 28632
rect 17925 27950 18031 28632
rect 5983 27175 6089 27857
rect 6209 27175 6314 27857
rect 6434 27175 6540 27857
rect 6674 27175 6780 27857
rect 6900 27175 7005 27857
rect 7125 27175 7231 27857
rect 16783 27175 16889 27857
rect 17009 27175 17114 27857
rect 17234 27175 17340 27857
rect 17474 27175 17580 27857
rect 17700 27175 17805 27857
rect 17925 27175 18031 27857
<< metal1 >>
rect 936 29818 1116 29830
rect 936 29766 948 29818
rect 1104 29766 1116 29818
rect 1125 29775 1289 30167
rect 6525 29775 6689 30167
rect 11730 29818 11910 29830
rect 936 29754 1116 29766
rect 11730 29766 11742 29818
rect 11898 29766 11910 29818
rect 11925 29775 12089 30167
rect 17325 29775 17489 30167
rect 22725 29890 22889 30167
rect 22532 29818 24835 29890
rect 11730 29754 11910 29766
rect 22532 29766 22869 29818
rect 23025 29766 24835 29818
rect 22532 29720 24835 29766
rect 22263 27031 22913 27105
rect 23206 18457 23552 19818
rect 23259 4973 23599 5013
rect 23259 4921 23297 4973
rect 23349 4921 23509 4973
rect 23561 4921 23599 4973
rect 23259 4755 23599 4921
rect 23259 4703 23297 4755
rect 23349 4703 23509 4755
rect 23561 4703 23599 4755
rect 23259 4662 23599 4703
<< via1 >>
rect 948 29766 1104 29818
rect 11742 29766 11898 29818
rect 22869 29766 23025 29818
rect 23297 4921 23349 4973
rect 23509 4921 23561 4973
rect 23297 4703 23349 4755
rect 23509 4703 23561 4755
<< metal2 >>
rect 977 29987 1077 31182
rect 977 29931 996 29987
rect 1052 29931 1077 29987
rect 977 29855 1077 29931
rect 977 29830 996 29855
rect 936 29818 996 29830
rect 1052 29830 1077 29855
rect 1052 29818 1116 29830
rect 936 29766 948 29818
rect 1104 29766 1116 29818
rect 936 29754 1116 29766
rect 977 29723 1077 29754
rect 977 29667 996 29723
rect 1052 29667 1077 29723
rect 977 29591 1077 29667
rect 977 29535 996 29591
rect 1052 29535 1077 29591
rect 977 29471 1077 29535
rect 1337 27527 1437 31182
rect 11777 29987 11877 31182
rect 11777 29931 11798 29987
rect 11854 29931 11877 29987
rect 11777 29855 11877 29931
rect 11777 29830 11798 29855
rect 11730 29818 11798 29830
rect 11854 29830 11877 29855
rect 11854 29818 11910 29830
rect 11730 29766 11742 29818
rect 11898 29766 11910 29818
rect 11730 29754 11910 29766
rect 11777 29723 11877 29754
rect 11777 29667 11798 29723
rect 11854 29667 11877 29723
rect 11777 29591 11877 29667
rect 11777 29535 11798 29591
rect 11854 29535 11877 29591
rect 11777 29517 11877 29535
rect 12137 27527 12237 31182
rect 22577 27527 22677 31182
rect 22937 29987 23037 31182
rect 22937 29931 22958 29987
rect 23014 29931 23037 29987
rect 22937 29855 23037 29931
rect 22937 29830 22958 29855
rect 22857 29818 22958 29830
rect 23014 29818 23037 29855
rect 22857 29766 22869 29818
rect 23025 29766 23037 29818
rect 22857 29754 23037 29766
rect 22937 29723 23037 29754
rect 22937 29667 22958 29723
rect 23014 29667 23037 29723
rect 22937 29591 23037 29667
rect 22937 29535 22958 29591
rect 23014 29535 23037 29591
rect 22937 27527 23037 29535
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4757 23599 4919
rect 23259 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 23259 4662 23599 4701
<< via2 >>
rect 996 29931 1052 29987
rect 996 29818 1052 29855
rect 996 29799 1052 29818
rect 996 29667 1052 29723
rect 996 29535 1052 29591
rect 11798 29931 11854 29987
rect 11798 29818 11854 29855
rect 11798 29799 11854 29818
rect 11798 29667 11854 29723
rect 11798 29535 11854 29591
rect 22958 29931 23014 29987
rect 22958 29818 23014 29855
rect 22958 29799 23014 29818
rect 22958 29667 23014 29723
rect 22958 29535 23014 29591
rect 23295 4973 23351 4975
rect 23295 4921 23297 4973
rect 23297 4921 23349 4973
rect 23349 4921 23351 4973
rect 23295 4919 23351 4921
rect 23507 4973 23563 4975
rect 23507 4921 23509 4973
rect 23509 4921 23561 4973
rect 23561 4921 23563 4973
rect 23507 4919 23563 4921
rect 23295 4755 23351 4757
rect 23295 4703 23297 4755
rect 23297 4703 23349 4755
rect 23349 4703 23351 4755
rect 23295 4701 23351 4703
rect 23507 4755 23563 4757
rect 23507 4703 23509 4755
rect 23509 4703 23561 4755
rect 23561 4703 23563 4755
rect 23507 4701 23563 4703
<< metal3 >>
rect -1 89507 23681 89707
rect -1 30537 23681 30897
rect 52 30139 23681 30279
rect -1 29987 24087 29997
rect -1 29931 996 29987
rect 1052 29931 11798 29987
rect 11854 29931 22958 29987
rect 23014 29931 24087 29987
rect -1 29855 24087 29931
rect -1 29799 996 29855
rect 1052 29799 11798 29855
rect 11854 29799 22958 29855
rect 23014 29799 24087 29855
rect -1 29723 24087 29799
rect -1 29667 996 29723
rect 1052 29667 11798 29723
rect 11854 29667 22958 29723
rect 23014 29667 24087 29723
rect -1 29591 24087 29667
rect -1 29535 996 29591
rect 1052 29535 11798 29591
rect 11854 29535 22958 29591
rect 23014 29535 24087 29591
rect -1 29517 24087 29535
rect 800 27296 24087 29105
rect 1314 21089 23252 21304
rect 1314 20767 23252 20983
rect 1314 20446 23252 20661
rect 1314 20124 23252 20339
rect 1314 19432 23252 19648
rect 1314 19110 23252 19326
rect 1314 18789 23252 19004
rect 1314 18467 23252 18682
rect 1314 17918 23252 18361
rect 1314 16807 23252 17263
rect 1314 12996 23252 15720
rect 1314 9308 23252 12711
rect 1262 8442 23710 9158
rect 1262 7016 24488 7827
rect 1314 5154 23971 6474
rect 1165 4923 22567 5011
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4758 23599 4919
rect 1165 4757 23599 4758
rect 1165 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 1165 4662 23599 4701
rect 1314 3133 24166 4495
rect 1314 1961 24276 2576
rect 1314 1286 23252 1855
rect 1314 747 24089 1179
rect 1314 155 24508 610
rect 1277 -959 24602 -504
rect 1277 -1599 23252 -1247
rect 1277 -2041 23252 -1953
rect 1277 -2517 23252 -2165
rect 1277 -3242 23252 -2787
use M2_M1$$43374636_512x8m81  M2_M1$$43374636_512x8m81_0
timestamp 1669390400
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1669390400
transform -1 0 22947 0 -1 29792
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1669390400
transform -1 0 11820 0 -1 29792
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1669390400
transform -1 0 1026 0 -1 29792
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_0
timestamp 1669390400
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_0
timestamp 1669390400
transform 1 0 12186 0 1 28317
box -38 -764 38 764
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_1
timestamp 1669390400
transform 1 0 22626 0 1 28317
box -38 -764 38 764
use M3_M24310591302022_512x8m81  M3_M24310591302022_512x8m81_2
timestamp 1669390400
transform 1 0 1386 0 1 28317
box -38 -764 38 764
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_0
timestamp 1669390400
transform 1 0 1024 0 1 29761
box 0 0 1 1
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_1
timestamp 1669390400
transform 1 0 11826 0 1 29761
box 0 0 1 1
use M3_M24310591302023_512x8m81  M3_M24310591302023_512x8m81_2
timestamp 1669390400
transform 1 0 22986 0 1 29761
box 0 0 1 1
use dcap_103_novia_512x8m81  dcap_103_novia_512x8m81_0
array 0 35 619 0 0 0
timestamp 1669390400
transform 1 0 288 0 1 29009
box -203 -284 822 881
use rarray4_512_512x8m81  rarray4_512_512x8m81_0
timestamp 1669390400
transform 1 0 907 0 1 31107
box -1997 -68 22836 57668
use rdummy_512x4_512x8m81  rdummy_512x4_512x8m81_0
timestamp 1669390400
transform 1 0 307 0 1 30207
box -358 -25410 24098 59488
use saout_R_m2_512x8m81  saout_R_m2_512x8m81_0
timestamp 1669390400
transform -1 0 12194 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_512x8m81  saout_R_m2_512x8m81_1
timestamp 1669390400
transform -1 0 22994 0 1 6
box -269 -3400 7633 31133
use saout_m2_512x8m81  saout_m2_512x8m81_0
timestamp 1669390400
transform 1 0 11820 0 1 -1
box -269 -3393 7633 31140
use saout_m2_512x8m81  saout_m2_512x8m81_1
timestamp 1669390400
transform 1 0 1020 0 1 -1
box -269 -3393 7633 31140
<< labels >>
rlabel metal3 s 1592 60366 1592 60366 4 WL[32]
port 1 nsew
rlabel metal3 s 1592 61266 1592 61266 4 WL[33]
port 2 nsew
rlabel metal3 s 1592 62166 1592 62166 4 WL[34]
port 3 nsew
rlabel metal3 s 1592 63066 1592 63066 4 WL[35]
port 4 nsew
rlabel metal3 s 1592 63966 1592 63966 4 WL[36]
port 5 nsew
rlabel metal3 s 1592 64866 1592 64866 4 WL[37]
port 6 nsew
rlabel metal3 s 1592 69366 1592 69366 4 WL[42]
port 7 nsew
rlabel metal3 s 1592 71166 1592 71166 4 WL[44]
port 8 nsew
rlabel metal3 s 1592 72966 1592 72966 4 WL[46]
port 9 nsew
rlabel metal3 s 1592 74766 1592 74766 4 WL[48]
port 10 nsew
rlabel metal3 s 1592 76566 1592 76566 4 WL[50]
port 11 nsew
rlabel metal3 s 1592 78366 1592 78366 4 WL[52]
port 12 nsew
rlabel metal3 s 1592 80166 1592 80166 4 WL[54]
port 13 nsew
rlabel metal3 s 1592 81966 1592 81966 4 WL[56]
port 14 nsew
rlabel metal3 s 1592 82866 1592 82866 4 WL[57]
port 15 nsew
rlabel metal3 s 1592 84666 1592 84666 4 WL[59]
port 16 nsew
rlabel metal3 s 1592 89157 1592 89157 4 DWL
port 17 nsew
rlabel metal3 s 1777 89717 1777 89717 4 VSS
port 18 nsew
rlabel metal3 s 1592 86465 1592 86465 4 WL[61]
port 19 nsew
rlabel metal3 s 1592 77465 1592 77465 4 WL[51]
port 20 nsew
rlabel metal3 s 1608 57668 1608 57668 4 WL[29]
port 21 nsew
rlabel metal3 s 1608 54068 1608 54068 4 WL[25]
port 22 nsew
rlabel metal3 s 1608 53168 1608 53168 4 WL[24]
port 23 nsew
rlabel metal3 s 1608 52268 1608 52268 4 WL[23]
port 24 nsew
rlabel metal3 s 1608 51368 1608 51368 4 WL[22]
port 25 nsew
rlabel metal3 s 1608 49568 1608 49568 4 WL[20]
port 26 nsew
rlabel metal3 s 1608 55868 1608 55868 4 WL[27]
port 27 nsew
rlabel metal3 s 1608 58568 1608 58568 4 WL[30]
port 28 nsew
rlabel metal3 s 1608 47768 1608 47768 4 WL[18]
port 29 nsew
rlabel metal3 s 1592 68465 1592 68465 4 WL[41]
port 30 nsew
rlabel metal3 s 1608 45068 1608 45068 4 WL[15]
port 31 nsew
rlabel metal3 s 1592 65765 1592 65765 4 WL[38]
port 32 nsew
rlabel metal3 s 1592 72065 1592 72065 4 WL[45]
port 33 nsew
rlabel metal3 s 1592 70265 1592 70265 4 WL[43]
port 34 nsew
rlabel metal3 s 1592 67565 1592 67565 4 WL[40]
port 35 nsew
rlabel metal3 s 1592 66665 1592 66665 4 WL[39]
port 36 nsew
rlabel metal3 s 1608 59468 1608 59468 4 WL[31]
port 37 nsew
rlabel metal3 s 1608 44168 1608 44168 4 WL[14]
port 38 nsew
rlabel metal3 s 1608 45968 1608 45968 4 WL[16]
port 39 nsew
rlabel metal3 s 1608 46868 1608 46868 4 WL[17]
port 40 nsew
rlabel metal3 s 1608 54968 1608 54968 4 WL[26]
port 41 nsew
rlabel metal3 s 1608 48668 1608 48668 4 WL[19]
port 42 nsew
rlabel metal3 s 1592 83765 1592 83765 4 WL[58]
port 43 nsew
rlabel metal3 s 1592 85565 1592 85565 4 WL[60]
port 44 nsew
rlabel metal3 s 1592 87365 1592 87365 4 WL[62]
port 45 nsew
rlabel metal3 s 1608 56768 1608 56768 4 WL[28]
port 46 nsew
rlabel metal3 s 1592 88265 1592 88265 4 WL[63]
port 47 nsew
rlabel metal3 s 1608 50468 1608 50468 4 WL[21]
port 48 nsew
rlabel metal3 s 1592 75665 1592 75665 4 WL[49]
port 49 nsew
rlabel metal3 s 1592 79265 1592 79265 4 WL[53]
port 50 nsew
rlabel metal3 s 1592 73865 1592 73865 4 WL[47]
port 51 nsew
rlabel metal3 s 1592 81065 1592 81065 4 WL[55]
port 52 nsew
rlabel metal3 s 240 30277 240 30277 4 VSS
port 18 nsew
rlabel metal3 s 1777 5806 1777 5806 4 VSS
port 18 nsew
rlabel metal3 s 1608 31568 1608 31568 4 WL[0]
port 53 nsew
rlabel metal3 s 1608 33368 1608 33368 4 WL[2]
port 54 nsew
rlabel metal3 s 1608 42368 1608 42368 4 WL[12]
port 55 nsew
rlabel metal3 s 1608 34268 1608 34268 4 WL[3]
port 56 nsew
rlabel metal3 s 1608 35168 1608 35168 4 WL[4]
port 57 nsew
flabel metal3 s 1659 -781 1659 -781 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
rlabel metal3 s 1608 37868 1608 37868 4 WL[7]
port 59 nsew
rlabel metal3 s 1608 38768 1608 38768 4 WL[8]
port 60 nsew
rlabel metal3 s 1608 39668 1608 39668 4 WL[9]
port 61 nsew
rlabel metal3 s 1608 32468 1608 32468 4 WL[1]
port 62 nsew
rlabel metal3 s 1705 21162 1705 21162 4 ypass[7]
port 63 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 64 nsew
flabel metal3 s 1659 -2347 1659 -2347 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 64 nsew
rlabel metal3 s 1607 36068 1607 36068 4 WL[5]
port 65 nsew
flabel metal3 s 1659 -1446 1659 -1446 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
rlabel metal3 s 1777 1467 1777 1467 4 men
port 64 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 64 nsew
rlabel metal3 s 1704 18591 1704 18591 4 ypass[0]
port 66 nsew
rlabel metal3 s 1608 40568 1608 40568 4 WL[10]
port 67 nsew
rlabel metal3 s 1608 43268 1608 43268 4 WL[13]
port 68 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 64 nsew
rlabel metal3 s 1704 18914 1704 18914 4 ypass[1]
port 69 nsew
rlabel metal3 s 1704 19231 1704 19231 4 ypass[2]
port 70 nsew
rlabel metal3 s 1704 19548 1704 19548 4 ypass[3]
port 71 nsew
rlabel metal3 s 1704 20204 1704 20204 4 ypass[4]
port 72 nsew
rlabel metal3 s 1704 20528 1704 20528 4 ypass[5]
port 73 nsew
rlabel metal3 s 1704 20845 1704 20845 4 ypass[6]
port 74 nsew
rlabel metal3 s 1774 1467 1774 1467 4 men
port 64 nsew
rlabel metal3 s 1607 36968 1607 36968 4 WL[6]
port 75 nsew
rlabel metal3 s 1346 4726 1346 4726 4 tblhl
port 76 nsew
flabel metal3 s 1659 -2004 1659 -2004 0 FreeSans 1000 0 0 0 GWEN
port 77 nsew
flabel metal3 s 1659 -3019 1659 -3019 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
rlabel metal3 s 1346 4983 1346 4983 4 GWE
port 78 nsew
rlabel metal3 s 1777 8832 1777 8832 4 VDD
port 58 nsew
rlabel metal3 s 1608 41468 1608 41468 4 WL[11]
port 79 nsew
flabel metal3 s 1659 390 1659 390 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 3623 1659 3623 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 7598 1659 7598 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 14001 1659 14001 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 18106 1659 18106 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 1659 28191 1659 28191 0 FreeSans 2000 0 0 0 VDD
port 58 nsew
flabel metal3 s 315 29753 315 29753 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 23123 1659 23123 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 16976 1659 16976 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 12236 1659 12236 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 6155 1659 6155 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 2247 1659 2247 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
flabel metal3 s 1659 949 1659 949 0 FreeSans 2000 0 0 0 VSS
port 18 nsew
rlabel metal2 s 1525 104 1525 104 4 din[4]
port 80 nsew
rlabel metal2 s 22492 104 22492 104 4 din[7]
port 81 nsew
rlabel metal2 s 10847 138 10847 138 4 q[5]
port 82 nsew
rlabel metal2 s 13174 104 13174 104 4 q[6]
port 83 nsew
rlabel metal2 s 21634 104 21634 104 4 q[7]
port 84 nsew
rlabel metal2 s 11686 104 11686 104 4 din[5]
port 85 nsew
rlabel metal2 s 12325 104 12325 104 4 din[6]
port 86 nsew
rlabel metal2 s 2371 104 2371 104 4 q[4]
port 87 nsew
rlabel metal1 s 7342 15928 7342 15928 4 pcb[6]
port 88 nsew
rlabel metal1 s 5921 15928 5921 15928 4 pcb[7]
port 89 nsew
rlabel metal1 s 18209 15928 18209 15928 4 pcb[4]
port 90 nsew
rlabel metal1 s 1827 18163 1827 18163 4 vdd
port 91 nsew
flabel metal1 s 22465 -3332 22465 -3332 0 FreeSans 600 0 0 0 WEN[4]
port 92 nsew
flabel metal1 s 1584 -3332 1584 -3332 0 FreeSans 600 0 0 0 WEN[7]
port 93 nsew
rlabel metal1 s 16588 15928 16588 15928 4 pcb[5]
port 94 nsew
flabel metal1 s 12358 -3332 12358 -3332 0 FreeSans 600 0 0 0 WEN[5]
port 95 nsew
flabel metal1 s 11643 -3332 11643 -3332 0 FreeSans 600 0 0 0 WEN[6]
port 96 nsew
<< properties >>
string GDS_END 2831462
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2819088
<< end >>
