magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 343 1502
<< polysilicon >>
rect -31 1361 89 1433
rect -31 -74 89 -1
use pmos_5p0431059087810_256x8m81  pmos_5p0431059087810_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 1482
<< properties >>
string GDS_END 43288
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 42974
<< end >>
