magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 111 134 123
rect 28 76 33 111
rect 64 91 69 104
rect 63 89 69 91
rect 61 83 71 89
rect 100 76 105 111
rect 22 44 32 50
rect 102 46 112 50
rect 47 44 112 46
rect 47 40 109 44
rect 28 12 33 36
rect 63 34 69 35
rect 61 28 71 34
rect 63 26 69 28
rect 64 19 69 26
rect 100 12 105 35
rect 0 0 134 12
<< obsm1 >>
rect 11 65 16 104
rect 54 73 94 78
rect 54 66 60 73
rect 89 68 94 73
rect 117 68 122 104
rect 11 60 47 65
rect 52 61 62 66
rect 11 19 16 60
rect 41 56 47 60
rect 73 56 79 68
rect 89 62 122 68
rect 89 57 95 62
rect 41 51 79 56
rect 87 51 97 57
rect 117 19 122 62
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 63 90 69 91
rect 62 82 70 90
rect 23 50 31 51
rect 22 44 32 50
rect 23 43 31 44
rect 63 35 69 82
rect 103 50 111 51
rect 102 44 112 50
rect 103 43 111 44
rect 61 27 71 35
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
<< labels >>
rlabel metal2 s 23 43 31 51 6 A
port 1 nsew signal input
rlabel metal2 s 22 44 32 50 6 A
port 1 nsew signal input
rlabel metal1 s 22 44 32 50 6 A
port 1 nsew signal input
rlabel metal2 s 103 43 111 51 6 B
port 3 nsew signal input
rlabel metal2 s 102 44 112 50 6 B
port 3 nsew signal input
rlabel metal1 s 47 40 109 46 6 B
port 3 nsew signal input
rlabel metal1 s 102 44 112 50 6 B
port 3 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 28 76 33 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 100 76 105 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 111 134 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 100 0 105 35 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 134 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 63 27 69 91 6 Y
port 2 nsew signal output
rlabel metal2 s 62 82 70 90 6 Y
port 2 nsew signal output
rlabel metal2 s 61 27 71 35 6 Y
port 2 nsew signal output
rlabel metal1 s 63 83 69 91 6 Y
port 2 nsew signal output
rlabel metal1 s 64 83 69 104 6 Y
port 2 nsew signal output
rlabel metal1 s 61 83 71 89 6 Y
port 2 nsew signal output
rlabel metal1 s 64 19 69 35 6 Y
port 2 nsew signal output
rlabel metal1 s 63 26 69 35 6 Y
port 2 nsew signal output
rlabel metal1 s 61 28 71 34 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 134 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 467820
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 456294
<< end >>
