magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -42 51823 342 51842
rect -42 -23 -23 51823
rect 323 -23 342 51823
rect -42 -42 342 -23
<< psubdiffcont >>
rect -23 -23 323 51823
<< metal1 >>
rect -34 51823 334 51834
rect -34 -23 -23 51823
rect 323 -23 334 51823
rect -34 -34 334 -23
<< properties >>
string GDS_END 1463194
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1330134
<< end >>
