magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -208 12637 76 12649
rect -208 11441 -196 12637
rect 64 11441 76 12637
rect -208 11429 76 11441
rect 13388 12637 13672 12649
rect 13388 11441 13400 12637
rect 13660 11441 13672 12637
rect 13388 11429 13672 11441
rect -360 10815 61 10892
rect -360 10763 -293 10815
rect -241 10763 -169 10815
rect -117 10763 -45 10815
rect 7 10763 61 10815
rect -360 10691 61 10763
rect -360 10639 -293 10691
rect -241 10639 -169 10691
rect -117 10639 -45 10691
rect 7 10639 61 10691
rect -360 10567 61 10639
rect -360 10515 -293 10567
rect -241 10515 -169 10567
rect -117 10515 -45 10567
rect 7 10515 61 10567
rect -360 10443 61 10515
rect -360 10391 -293 10443
rect -241 10391 -169 10443
rect -117 10391 -45 10443
rect 7 10391 61 10443
rect -360 10319 61 10391
rect -360 10267 -293 10319
rect -241 10267 -169 10319
rect -117 10267 -45 10319
rect 7 10267 61 10319
rect -360 10195 61 10267
rect -360 10143 -293 10195
rect -241 10143 -169 10195
rect -117 10143 -45 10195
rect 7 10143 61 10195
rect -360 10071 61 10143
rect -360 10019 -293 10071
rect -241 10019 -169 10071
rect -117 10019 -45 10071
rect 7 10019 61 10071
rect 1003 10815 1940 10854
rect 1003 10763 1037 10815
rect 1089 10763 1161 10815
rect 1213 10763 1285 10815
rect 1337 10763 1409 10815
rect 1461 10763 1940 10815
rect 1003 10691 1940 10763
rect 1003 10639 1037 10691
rect 1089 10639 1161 10691
rect 1213 10639 1285 10691
rect 1337 10639 1409 10691
rect 1461 10639 1940 10691
rect 1003 10567 1940 10639
rect 1003 10515 1037 10567
rect 1089 10515 1161 10567
rect 1213 10515 1285 10567
rect 1337 10515 1409 10567
rect 1461 10515 1940 10567
rect 1003 10443 1940 10515
rect 1003 10391 1037 10443
rect 1089 10391 1161 10443
rect 1213 10391 1285 10443
rect 1337 10391 1409 10443
rect 1461 10391 1940 10443
rect 1003 10319 1940 10391
rect 1003 10267 1037 10319
rect 1089 10267 1161 10319
rect 1213 10267 1285 10319
rect 1337 10267 1409 10319
rect 1461 10267 1940 10319
rect 1003 10195 1940 10267
rect 1003 10143 1037 10195
rect 1089 10143 1161 10195
rect 1213 10143 1285 10195
rect 1337 10143 1409 10195
rect 1461 10143 1940 10195
rect 1003 10071 1940 10143
rect 1003 10058 1037 10071
rect -360 9947 61 10019
rect -360 9895 -293 9947
rect -241 9895 -169 9947
rect -117 9895 -45 9947
rect 7 9895 61 9947
rect -360 9823 61 9895
rect -360 9771 -293 9823
rect -241 9771 -169 9823
rect -117 9771 -45 9823
rect 7 9771 61 9823
rect -360 8855 61 9771
rect 1025 10019 1037 10058
rect 1089 10019 1161 10071
rect 1213 10019 1285 10071
rect 1337 10019 1409 10071
rect 1461 10058 1940 10071
rect 11505 10815 12426 10854
rect 11505 10763 11968 10815
rect 12020 10763 12092 10815
rect 12144 10763 12216 10815
rect 12268 10763 12340 10815
rect 12392 10763 12426 10815
rect 11505 10691 12426 10763
rect 11505 10639 11968 10691
rect 12020 10639 12092 10691
rect 12144 10639 12216 10691
rect 12268 10639 12340 10691
rect 12392 10639 12426 10691
rect 11505 10567 12426 10639
rect 11505 10515 11968 10567
rect 12020 10515 12092 10567
rect 12144 10515 12216 10567
rect 12268 10515 12340 10567
rect 12392 10515 12426 10567
rect 11505 10443 12426 10515
rect 11505 10391 11968 10443
rect 12020 10391 12092 10443
rect 12144 10391 12216 10443
rect 12268 10391 12340 10443
rect 12392 10391 12426 10443
rect 11505 10319 12426 10391
rect 11505 10267 11968 10319
rect 12020 10267 12092 10319
rect 12144 10267 12216 10319
rect 12268 10267 12340 10319
rect 12392 10267 12426 10319
rect 11505 10195 12426 10267
rect 11505 10143 11968 10195
rect 12020 10143 12092 10195
rect 12144 10143 12216 10195
rect 12268 10143 12340 10195
rect 12392 10143 12426 10195
rect 11505 10071 12426 10143
rect 11505 10058 11968 10071
rect 1461 10019 1473 10058
rect 1025 9947 1473 10019
rect 1025 9895 1037 9947
rect 1089 9895 1161 9947
rect 1213 9895 1285 9947
rect 1337 9895 1409 9947
rect 1461 9895 1473 9947
rect 1025 9823 1473 9895
rect 1025 9771 1037 9823
rect 1089 9771 1161 9823
rect 1213 9771 1285 9823
rect 1337 9771 1409 9823
rect 1461 9771 1473 9823
rect 1025 9759 1473 9771
rect 11956 10019 11968 10058
rect 12020 10019 12092 10071
rect 12144 10019 12216 10071
rect 12268 10019 12340 10071
rect 12392 10058 12426 10071
rect 13364 10815 13785 10892
rect 13364 10763 13418 10815
rect 13470 10763 13542 10815
rect 13594 10763 13666 10815
rect 13718 10763 13785 10815
rect 13364 10691 13785 10763
rect 13364 10639 13418 10691
rect 13470 10639 13542 10691
rect 13594 10639 13666 10691
rect 13718 10639 13785 10691
rect 13364 10567 13785 10639
rect 13364 10515 13418 10567
rect 13470 10515 13542 10567
rect 13594 10515 13666 10567
rect 13718 10515 13785 10567
rect 13364 10443 13785 10515
rect 13364 10391 13418 10443
rect 13470 10391 13542 10443
rect 13594 10391 13666 10443
rect 13718 10391 13785 10443
rect 13364 10319 13785 10391
rect 13364 10267 13418 10319
rect 13470 10267 13542 10319
rect 13594 10267 13666 10319
rect 13718 10267 13785 10319
rect 13364 10195 13785 10267
rect 13364 10143 13418 10195
rect 13470 10143 13542 10195
rect 13594 10143 13666 10195
rect 13718 10143 13785 10195
rect 13364 10071 13785 10143
rect 12392 10019 12404 10058
rect 11956 9947 12404 10019
rect 11956 9895 11968 9947
rect 12020 9895 12092 9947
rect 12144 9895 12216 9947
rect 12268 9895 12340 9947
rect 12392 9895 12404 9947
rect 11956 9823 12404 9895
rect 11956 9771 11968 9823
rect 12020 9771 12092 9823
rect 12144 9771 12216 9823
rect 12268 9771 12340 9823
rect 12392 9771 12404 9823
rect 11956 9759 12404 9771
rect 13364 10019 13418 10071
rect 13470 10019 13542 10071
rect 13594 10019 13666 10071
rect 13718 10019 13785 10071
rect 13364 9947 13785 10019
rect 13364 9895 13418 9947
rect 13470 9895 13542 9947
rect 13594 9895 13666 9947
rect 13718 9895 13785 9947
rect 13364 9823 13785 9895
rect 13364 9771 13418 9823
rect 13470 9771 13542 9823
rect 13594 9771 13666 9823
rect 13718 9771 13785 9823
rect 1417 9510 1597 9522
rect 1417 9458 1429 9510
rect 1585 9458 1597 9510
rect 1417 9446 1597 9458
rect 11881 9510 12061 9522
rect 11881 9458 11893 9510
rect 12049 9458 12061 9510
rect 11881 9446 12061 9458
rect 1417 9342 1597 9354
rect 1417 9290 1429 9342
rect 1585 9290 1597 9342
rect 1417 9278 1597 9290
rect 11881 9342 12061 9354
rect 11881 9290 11893 9342
rect 12049 9290 12061 9342
rect 11881 9278 12061 9290
rect 1417 9182 1597 9194
rect 1417 9130 1429 9182
rect 1585 9130 1597 9182
rect 1417 9118 1597 9130
rect 11881 9182 12061 9194
rect 11881 9130 11893 9182
rect 12049 9130 12061 9182
rect 11881 9118 12061 9130
rect 1417 9016 1597 9028
rect 1417 8964 1429 9016
rect 1585 8964 1597 9016
rect 1417 8952 1597 8964
rect 11881 9016 12061 9028
rect 11881 8964 11893 9016
rect 12049 8964 12061 9016
rect 11881 8952 12061 8964
rect 13364 8877 13785 9771
rect -360 8482 971 8855
rect 2014 8824 2090 8836
rect 2014 6588 2026 8824
rect 2078 6588 2090 8824
rect 2014 6576 2090 6588
rect 11339 8824 11415 8836
rect 11339 6588 11351 8824
rect 11403 6588 11415 8824
rect 12360 8482 13785 8877
rect 11339 6576 11415 6588
rect 2014 6263 2090 6275
rect 2014 3403 2026 6263
rect 2078 3403 2090 6263
rect 2014 3391 2090 3403
rect 11339 6263 11415 6275
rect 11339 3403 11351 6263
rect 11403 3403 11415 6263
rect 11339 3391 11415 3403
rect 2014 3067 2090 3079
rect 2014 519 2026 3067
rect 2078 519 2090 3067
rect 2014 507 2090 519
rect 11339 3067 11415 3079
rect 11339 519 11351 3067
rect 11403 519 11415 3067
rect 11339 507 11415 519
<< via1 >>
rect -196 11441 64 12637
rect 13400 11441 13660 12637
rect -293 10763 -241 10815
rect -169 10763 -117 10815
rect -45 10763 7 10815
rect -293 10639 -241 10691
rect -169 10639 -117 10691
rect -45 10639 7 10691
rect -293 10515 -241 10567
rect -169 10515 -117 10567
rect -45 10515 7 10567
rect -293 10391 -241 10443
rect -169 10391 -117 10443
rect -45 10391 7 10443
rect -293 10267 -241 10319
rect -169 10267 -117 10319
rect -45 10267 7 10319
rect -293 10143 -241 10195
rect -169 10143 -117 10195
rect -45 10143 7 10195
rect -293 10019 -241 10071
rect -169 10019 -117 10071
rect -45 10019 7 10071
rect 1037 10763 1089 10815
rect 1161 10763 1213 10815
rect 1285 10763 1337 10815
rect 1409 10763 1461 10815
rect 1037 10639 1089 10691
rect 1161 10639 1213 10691
rect 1285 10639 1337 10691
rect 1409 10639 1461 10691
rect 1037 10515 1089 10567
rect 1161 10515 1213 10567
rect 1285 10515 1337 10567
rect 1409 10515 1461 10567
rect 1037 10391 1089 10443
rect 1161 10391 1213 10443
rect 1285 10391 1337 10443
rect 1409 10391 1461 10443
rect 1037 10267 1089 10319
rect 1161 10267 1213 10319
rect 1285 10267 1337 10319
rect 1409 10267 1461 10319
rect 1037 10143 1089 10195
rect 1161 10143 1213 10195
rect 1285 10143 1337 10195
rect 1409 10143 1461 10195
rect -293 9895 -241 9947
rect -169 9895 -117 9947
rect -45 9895 7 9947
rect -293 9771 -241 9823
rect -169 9771 -117 9823
rect -45 9771 7 9823
rect 1037 10019 1089 10071
rect 1161 10019 1213 10071
rect 1285 10019 1337 10071
rect 1409 10019 1461 10071
rect 11968 10763 12020 10815
rect 12092 10763 12144 10815
rect 12216 10763 12268 10815
rect 12340 10763 12392 10815
rect 11968 10639 12020 10691
rect 12092 10639 12144 10691
rect 12216 10639 12268 10691
rect 12340 10639 12392 10691
rect 11968 10515 12020 10567
rect 12092 10515 12144 10567
rect 12216 10515 12268 10567
rect 12340 10515 12392 10567
rect 11968 10391 12020 10443
rect 12092 10391 12144 10443
rect 12216 10391 12268 10443
rect 12340 10391 12392 10443
rect 11968 10267 12020 10319
rect 12092 10267 12144 10319
rect 12216 10267 12268 10319
rect 12340 10267 12392 10319
rect 11968 10143 12020 10195
rect 12092 10143 12144 10195
rect 12216 10143 12268 10195
rect 12340 10143 12392 10195
rect 1037 9895 1089 9947
rect 1161 9895 1213 9947
rect 1285 9895 1337 9947
rect 1409 9895 1461 9947
rect 1037 9771 1089 9823
rect 1161 9771 1213 9823
rect 1285 9771 1337 9823
rect 1409 9771 1461 9823
rect 11968 10019 12020 10071
rect 12092 10019 12144 10071
rect 12216 10019 12268 10071
rect 12340 10019 12392 10071
rect 13418 10763 13470 10815
rect 13542 10763 13594 10815
rect 13666 10763 13718 10815
rect 13418 10639 13470 10691
rect 13542 10639 13594 10691
rect 13666 10639 13718 10691
rect 13418 10515 13470 10567
rect 13542 10515 13594 10567
rect 13666 10515 13718 10567
rect 13418 10391 13470 10443
rect 13542 10391 13594 10443
rect 13666 10391 13718 10443
rect 13418 10267 13470 10319
rect 13542 10267 13594 10319
rect 13666 10267 13718 10319
rect 13418 10143 13470 10195
rect 13542 10143 13594 10195
rect 13666 10143 13718 10195
rect 11968 9895 12020 9947
rect 12092 9895 12144 9947
rect 12216 9895 12268 9947
rect 12340 9895 12392 9947
rect 11968 9771 12020 9823
rect 12092 9771 12144 9823
rect 12216 9771 12268 9823
rect 12340 9771 12392 9823
rect 13418 10019 13470 10071
rect 13542 10019 13594 10071
rect 13666 10019 13718 10071
rect 13418 9895 13470 9947
rect 13542 9895 13594 9947
rect 13666 9895 13718 9947
rect 13418 9771 13470 9823
rect 13542 9771 13594 9823
rect 13666 9771 13718 9823
rect 1429 9458 1585 9510
rect 11893 9458 12049 9510
rect 1429 9290 1585 9342
rect 11893 9290 12049 9342
rect 1429 9130 1585 9182
rect 11893 9130 12049 9182
rect 1429 8964 1585 9016
rect 11893 8964 12049 9016
rect 2026 6588 2078 8824
rect 11351 6588 11403 8824
rect 2026 3403 2078 6263
rect 11351 3403 11403 6263
rect 2026 519 2078 3067
rect 11351 519 11403 3067
<< metal2 >>
rect -208 12637 76 12649
rect -208 11441 -196 12637
rect 64 11441 76 12637
rect -208 11429 76 11441
rect -310 10818 50 10828
rect -310 10762 -300 10818
rect -244 10815 -158 10818
rect -102 10815 -16 10818
rect -241 10763 -169 10815
rect -102 10763 -45 10815
rect -244 10762 -158 10763
rect -102 10762 -16 10763
rect 40 10762 50 10818
rect -310 10691 50 10762
rect -310 10676 -293 10691
rect -310 10620 -300 10676
rect -241 10639 -169 10691
rect -117 10676 -45 10691
rect 7 10676 50 10691
rect -102 10639 -45 10676
rect -244 10620 -158 10639
rect -102 10620 -16 10639
rect 40 10620 50 10676
rect -310 10567 50 10620
rect -310 10534 -293 10567
rect -310 10478 -300 10534
rect -241 10515 -169 10567
rect -117 10534 -45 10567
rect 7 10534 50 10567
rect -102 10515 -45 10534
rect -244 10478 -158 10515
rect -102 10478 -16 10515
rect 40 10478 50 10534
rect -310 10443 50 10478
rect -310 10392 -293 10443
rect -310 10336 -300 10392
rect -241 10391 -169 10443
rect -117 10392 -45 10443
rect 7 10392 50 10443
rect -102 10391 -45 10392
rect -244 10336 -158 10391
rect -102 10336 -16 10391
rect 40 10336 50 10392
rect -310 10319 50 10336
rect -310 10267 -293 10319
rect -241 10267 -169 10319
rect -117 10267 -45 10319
rect 7 10267 50 10319
rect -310 10250 50 10267
rect -310 10194 -300 10250
rect -244 10195 -158 10250
rect -102 10195 -16 10250
rect -310 10143 -293 10194
rect -241 10143 -169 10195
rect -102 10194 -45 10195
rect 40 10194 50 10250
rect -117 10143 -45 10194
rect 7 10143 50 10194
rect -310 10108 50 10143
rect -310 10052 -300 10108
rect -244 10071 -158 10108
rect -102 10071 -16 10108
rect -310 10019 -293 10052
rect -241 10019 -169 10071
rect -102 10052 -45 10071
rect 40 10052 50 10108
rect -117 10019 -45 10052
rect 7 10019 50 10052
rect -310 9966 50 10019
rect -310 9910 -300 9966
rect -244 9947 -158 9966
rect -102 9947 -16 9966
rect -310 9895 -293 9910
rect -241 9895 -169 9947
rect -102 9910 -45 9947
rect 40 9910 50 9966
rect -117 9895 -45 9910
rect 7 9895 50 9910
rect -310 9824 50 9895
rect -310 9768 -300 9824
rect -244 9823 -158 9824
rect -102 9823 -16 9824
rect -241 9771 -169 9823
rect -102 9771 -45 9823
rect -244 9768 -158 9771
rect -102 9768 -16 9771
rect 40 9768 50 9824
rect -310 9758 50 9768
rect 213 9051 313 26936
rect 393 9211 493 26936
rect 573 9371 673 26936
rect 753 9539 861 26936
rect 1697 26000 11785 26600
rect 1697 24843 2941 26000
rect 3465 24843 4709 26000
rect 5233 24843 6477 26000
rect 7001 24843 8245 26000
rect 8769 24843 10013 26000
rect 10537 24843 11781 26000
rect 1697 12658 2941 12843
rect 3465 12658 4709 12843
rect 5233 12658 6477 12843
rect 7001 12658 8245 12843
rect 8769 12658 10013 12843
rect 10537 12658 11781 12843
rect 1025 10818 1473 10828
rect 1025 10815 1079 10818
rect 1135 10815 1221 10818
rect 1025 10763 1037 10815
rect 1135 10763 1161 10815
rect 1213 10763 1221 10815
rect 1025 10762 1079 10763
rect 1135 10762 1221 10763
rect 1277 10815 1363 10818
rect 1419 10815 1473 10818
rect 1277 10763 1285 10815
rect 1337 10763 1363 10815
rect 1461 10763 1473 10815
rect 1277 10762 1363 10763
rect 1419 10762 1473 10763
rect 1025 10691 1473 10762
rect 1025 10639 1037 10691
rect 1089 10676 1161 10691
rect 1135 10639 1161 10676
rect 1213 10676 1285 10691
rect 1213 10639 1221 10676
rect 1025 10620 1079 10639
rect 1135 10620 1221 10639
rect 1277 10639 1285 10676
rect 1337 10676 1409 10691
rect 1337 10639 1363 10676
rect 1461 10639 1473 10691
rect 1277 10620 1363 10639
rect 1419 10620 1473 10639
rect 1025 10567 1473 10620
rect 1025 10515 1037 10567
rect 1089 10534 1161 10567
rect 1135 10515 1161 10534
rect 1213 10534 1285 10567
rect 1213 10515 1221 10534
rect 1025 10478 1079 10515
rect 1135 10478 1221 10515
rect 1277 10515 1285 10534
rect 1337 10534 1409 10567
rect 1337 10515 1363 10534
rect 1461 10515 1473 10567
rect 1277 10478 1363 10515
rect 1419 10478 1473 10515
rect 1025 10443 1473 10478
rect 1025 10391 1037 10443
rect 1089 10392 1161 10443
rect 1135 10391 1161 10392
rect 1213 10392 1285 10443
rect 1213 10391 1221 10392
rect 1025 10336 1079 10391
rect 1135 10336 1221 10391
rect 1277 10391 1285 10392
rect 1337 10392 1409 10443
rect 1337 10391 1363 10392
rect 1461 10391 1473 10443
rect 1277 10336 1363 10391
rect 1419 10336 1473 10391
rect 1025 10319 1473 10336
rect 1025 10267 1037 10319
rect 1089 10267 1161 10319
rect 1213 10267 1285 10319
rect 1337 10267 1409 10319
rect 1461 10267 1473 10319
rect 1025 10250 1473 10267
rect 1025 10195 1079 10250
rect 1135 10195 1221 10250
rect 1025 10143 1037 10195
rect 1135 10194 1161 10195
rect 1089 10143 1161 10194
rect 1213 10194 1221 10195
rect 1277 10195 1363 10250
rect 1419 10195 1473 10250
rect 1277 10194 1285 10195
rect 1213 10143 1285 10194
rect 1337 10194 1363 10195
rect 1337 10143 1409 10194
rect 1461 10143 1473 10195
rect 1025 10108 1473 10143
rect 1025 10071 1079 10108
rect 1135 10071 1221 10108
rect 1025 10019 1037 10071
rect 1135 10052 1161 10071
rect 1089 10019 1161 10052
rect 1213 10052 1221 10071
rect 1277 10071 1363 10108
rect 1419 10071 1473 10108
rect 1277 10052 1285 10071
rect 1213 10019 1285 10052
rect 1337 10052 1363 10071
rect 1337 10019 1409 10052
rect 1461 10019 1473 10071
rect 1025 9966 1473 10019
rect 1025 9947 1079 9966
rect 1135 9947 1221 9966
rect 1025 9895 1037 9947
rect 1135 9910 1161 9947
rect 1089 9895 1161 9910
rect 1213 9910 1221 9947
rect 1277 9947 1363 9966
rect 1419 9947 1473 9966
rect 1277 9910 1285 9947
rect 1213 9895 1285 9910
rect 1337 9910 1363 9947
rect 1337 9895 1409 9910
rect 1461 9895 1473 9947
rect 1025 9824 1473 9895
rect 1025 9823 1079 9824
rect 1135 9823 1221 9824
rect 1025 9771 1037 9823
rect 1135 9771 1161 9823
rect 1213 9771 1221 9823
rect 1025 9768 1079 9771
rect 1135 9768 1221 9771
rect 1277 9823 1363 9824
rect 1419 9823 1473 9824
rect 1277 9771 1285 9823
rect 1337 9771 1363 9823
rect 1461 9771 1473 9823
rect 1277 9768 1363 9771
rect 1419 9768 1473 9771
rect 1025 9758 1473 9768
rect 753 9510 1597 9539
rect 753 9458 1429 9510
rect 1585 9458 1597 9510
rect 753 9431 1597 9458
rect 573 9342 1597 9371
rect 573 9290 1429 9342
rect 1585 9290 1597 9342
rect 573 9271 1597 9290
rect 393 9182 1597 9211
rect 393 9130 1429 9182
rect 1585 9130 1597 9182
rect 393 9111 1597 9130
rect 213 9016 1597 9051
rect 213 8964 1429 9016
rect 1585 8964 1597 9016
rect 213 8951 1597 8964
rect 1697 8943 11781 12658
rect 11956 10818 12404 10828
rect 11956 10815 12010 10818
rect 12066 10815 12152 10818
rect 11956 10763 11968 10815
rect 12066 10763 12092 10815
rect 12144 10763 12152 10815
rect 11956 10762 12010 10763
rect 12066 10762 12152 10763
rect 12208 10815 12294 10818
rect 12350 10815 12404 10818
rect 12208 10763 12216 10815
rect 12268 10763 12294 10815
rect 12392 10763 12404 10815
rect 12208 10762 12294 10763
rect 12350 10762 12404 10763
rect 11956 10691 12404 10762
rect 11956 10639 11968 10691
rect 12020 10676 12092 10691
rect 12066 10639 12092 10676
rect 12144 10676 12216 10691
rect 12144 10639 12152 10676
rect 11956 10620 12010 10639
rect 12066 10620 12152 10639
rect 12208 10639 12216 10676
rect 12268 10676 12340 10691
rect 12268 10639 12294 10676
rect 12392 10639 12404 10691
rect 12208 10620 12294 10639
rect 12350 10620 12404 10639
rect 11956 10567 12404 10620
rect 11956 10515 11968 10567
rect 12020 10534 12092 10567
rect 12066 10515 12092 10534
rect 12144 10534 12216 10567
rect 12144 10515 12152 10534
rect 11956 10478 12010 10515
rect 12066 10478 12152 10515
rect 12208 10515 12216 10534
rect 12268 10534 12340 10567
rect 12268 10515 12294 10534
rect 12392 10515 12404 10567
rect 12208 10478 12294 10515
rect 12350 10478 12404 10515
rect 11956 10443 12404 10478
rect 11956 10391 11968 10443
rect 12020 10392 12092 10443
rect 12066 10391 12092 10392
rect 12144 10392 12216 10443
rect 12144 10391 12152 10392
rect 11956 10336 12010 10391
rect 12066 10336 12152 10391
rect 12208 10391 12216 10392
rect 12268 10392 12340 10443
rect 12268 10391 12294 10392
rect 12392 10391 12404 10443
rect 12208 10336 12294 10391
rect 12350 10336 12404 10391
rect 11956 10319 12404 10336
rect 11956 10267 11968 10319
rect 12020 10267 12092 10319
rect 12144 10267 12216 10319
rect 12268 10267 12340 10319
rect 12392 10267 12404 10319
rect 11956 10250 12404 10267
rect 11956 10195 12010 10250
rect 12066 10195 12152 10250
rect 11956 10143 11968 10195
rect 12066 10194 12092 10195
rect 12020 10143 12092 10194
rect 12144 10194 12152 10195
rect 12208 10195 12294 10250
rect 12350 10195 12404 10250
rect 12208 10194 12216 10195
rect 12144 10143 12216 10194
rect 12268 10194 12294 10195
rect 12268 10143 12340 10194
rect 12392 10143 12404 10195
rect 11956 10108 12404 10143
rect 11956 10071 12010 10108
rect 12066 10071 12152 10108
rect 11956 10019 11968 10071
rect 12066 10052 12092 10071
rect 12020 10019 12092 10052
rect 12144 10052 12152 10071
rect 12208 10071 12294 10108
rect 12350 10071 12404 10108
rect 12208 10052 12216 10071
rect 12144 10019 12216 10052
rect 12268 10052 12294 10071
rect 12268 10019 12340 10052
rect 12392 10019 12404 10071
rect 11956 9966 12404 10019
rect 11956 9947 12010 9966
rect 12066 9947 12152 9966
rect 11956 9895 11968 9947
rect 12066 9910 12092 9947
rect 12020 9895 12092 9910
rect 12144 9910 12152 9947
rect 12208 9947 12294 9966
rect 12350 9947 12404 9966
rect 12208 9910 12216 9947
rect 12144 9895 12216 9910
rect 12268 9910 12294 9947
rect 12268 9895 12340 9910
rect 12392 9895 12404 9947
rect 11956 9824 12404 9895
rect 11956 9823 12010 9824
rect 12066 9823 12152 9824
rect 11956 9771 11968 9823
rect 12066 9771 12092 9823
rect 12144 9771 12152 9823
rect 11956 9768 12010 9771
rect 12066 9768 12152 9771
rect 12208 9823 12294 9824
rect 12350 9823 12404 9824
rect 12208 9771 12216 9823
rect 12268 9771 12294 9823
rect 12392 9771 12404 9823
rect 12208 9768 12294 9771
rect 12350 9768 12404 9771
rect 11956 9758 12404 9768
rect 12617 9539 12725 26936
rect 11881 9510 12725 9539
rect 11881 9458 11893 9510
rect 12049 9458 12725 9510
rect 11881 9431 12725 9458
rect 12805 9371 12905 26936
rect 11881 9342 12905 9371
rect 11881 9290 11893 9342
rect 12049 9290 12905 9342
rect 11881 9271 12905 9290
rect 12985 9211 13085 26936
rect 11881 9182 13085 9211
rect 11881 9130 11893 9182
rect 12049 9130 13085 9182
rect 11881 9111 13085 9130
rect 13165 9051 13265 26936
rect 13388 12637 13672 12649
rect 13388 11441 13400 12637
rect 13660 11441 13672 12637
rect 13388 11429 13672 11441
rect 13375 10818 13735 10828
rect 13375 10762 13385 10818
rect 13441 10815 13527 10818
rect 13583 10815 13669 10818
rect 13470 10763 13527 10815
rect 13594 10763 13666 10815
rect 13441 10762 13527 10763
rect 13583 10762 13669 10763
rect 13725 10762 13735 10818
rect 13375 10691 13735 10762
rect 13375 10676 13418 10691
rect 13470 10676 13542 10691
rect 13375 10620 13385 10676
rect 13470 10639 13527 10676
rect 13594 10639 13666 10691
rect 13718 10676 13735 10691
rect 13441 10620 13527 10639
rect 13583 10620 13669 10639
rect 13725 10620 13735 10676
rect 13375 10567 13735 10620
rect 13375 10534 13418 10567
rect 13470 10534 13542 10567
rect 13375 10478 13385 10534
rect 13470 10515 13527 10534
rect 13594 10515 13666 10567
rect 13718 10534 13735 10567
rect 13441 10478 13527 10515
rect 13583 10478 13669 10515
rect 13725 10478 13735 10534
rect 13375 10443 13735 10478
rect 13375 10392 13418 10443
rect 13470 10392 13542 10443
rect 13375 10336 13385 10392
rect 13470 10391 13527 10392
rect 13594 10391 13666 10443
rect 13718 10392 13735 10443
rect 13441 10336 13527 10391
rect 13583 10336 13669 10391
rect 13725 10336 13735 10392
rect 13375 10319 13735 10336
rect 13375 10267 13418 10319
rect 13470 10267 13542 10319
rect 13594 10267 13666 10319
rect 13718 10267 13735 10319
rect 13375 10250 13735 10267
rect 13375 10194 13385 10250
rect 13441 10195 13527 10250
rect 13583 10195 13669 10250
rect 13470 10194 13527 10195
rect 13375 10143 13418 10194
rect 13470 10143 13542 10194
rect 13594 10143 13666 10195
rect 13725 10194 13735 10250
rect 13718 10143 13735 10194
rect 13375 10108 13735 10143
rect 13375 10052 13385 10108
rect 13441 10071 13527 10108
rect 13583 10071 13669 10108
rect 13470 10052 13527 10071
rect 13375 10019 13418 10052
rect 13470 10019 13542 10052
rect 13594 10019 13666 10071
rect 13725 10052 13735 10108
rect 13718 10019 13735 10052
rect 13375 9966 13735 10019
rect 13375 9910 13385 9966
rect 13441 9947 13527 9966
rect 13583 9947 13669 9966
rect 13470 9910 13527 9947
rect 13375 9895 13418 9910
rect 13470 9895 13542 9910
rect 13594 9895 13666 9947
rect 13725 9910 13735 9966
rect 13718 9895 13735 9910
rect 13375 9824 13735 9895
rect 13375 9768 13385 9824
rect 13441 9823 13527 9824
rect 13583 9823 13669 9824
rect 13470 9771 13527 9823
rect 13594 9771 13666 9823
rect 13441 9768 13527 9771
rect 13583 9768 13669 9771
rect 13725 9768 13735 9824
rect 13375 9758 13735 9768
rect 11881 9016 13265 9051
rect 11881 8964 11893 9016
rect 12049 8964 13265 9016
rect 11881 8951 13265 8964
rect 1698 -1081 1896 8943
rect 2014 8824 2168 8843
rect 2014 8799 2026 8824
rect 2078 8799 2168 8824
rect 2014 8743 2024 8799
rect 2080 8743 2168 8799
rect 2014 8657 2026 8743
rect 2078 8657 2168 8743
rect 2014 8601 2024 8657
rect 2080 8601 2168 8657
rect 2014 8515 2026 8601
rect 2078 8515 2168 8601
rect 2014 8459 2024 8515
rect 2080 8459 2168 8515
rect 2014 8373 2026 8459
rect 2078 8373 2168 8459
rect 2014 8317 2024 8373
rect 2080 8317 2168 8373
rect 2014 8231 2026 8317
rect 2078 8231 2168 8317
rect 2014 8175 2024 8231
rect 2080 8175 2168 8231
rect 2014 8089 2026 8175
rect 2078 8089 2168 8175
rect 2014 8033 2024 8089
rect 2080 8033 2168 8089
rect 2014 7947 2026 8033
rect 2078 7947 2168 8033
rect 2014 7891 2024 7947
rect 2080 7891 2168 7947
rect 2014 7805 2026 7891
rect 2078 7805 2168 7891
rect 2014 7749 2024 7805
rect 2080 7749 2168 7805
rect 2014 7663 2026 7749
rect 2078 7663 2168 7749
rect 2014 7607 2024 7663
rect 2080 7607 2168 7663
rect 2014 7521 2026 7607
rect 2078 7521 2168 7607
rect 2014 7465 2024 7521
rect 2080 7465 2168 7521
rect 2014 7379 2026 7465
rect 2078 7379 2168 7465
rect 2014 7323 2024 7379
rect 2080 7323 2168 7379
rect 2014 7237 2026 7323
rect 2078 7237 2168 7323
rect 2014 7181 2024 7237
rect 2080 7181 2168 7237
rect 2014 7095 2026 7181
rect 2078 7095 2168 7181
rect 2014 7039 2024 7095
rect 2080 7039 2168 7095
rect 2014 6953 2026 7039
rect 2078 6953 2168 7039
rect 2014 6897 2024 6953
rect 2080 6897 2168 6953
rect 2014 6811 2026 6897
rect 2078 6811 2168 6897
rect 2014 6755 2024 6811
rect 2080 6755 2168 6811
rect 2014 6669 2026 6755
rect 2078 6669 2168 6755
rect 2014 6613 2024 6669
rect 2080 6613 2168 6669
rect 2014 6588 2026 6613
rect 2078 6588 2168 6613
rect 2014 6263 2168 6588
rect 2014 6217 2026 6263
rect 2078 6217 2168 6263
rect 2014 6161 2024 6217
rect 2080 6161 2168 6217
rect 2014 6075 2026 6161
rect 2078 6075 2168 6161
rect 2014 6019 2024 6075
rect 2080 6019 2168 6075
rect 2014 5933 2026 6019
rect 2078 5933 2168 6019
rect 2014 5877 2024 5933
rect 2080 5877 2168 5933
rect 2014 5791 2026 5877
rect 2078 5791 2168 5877
rect 2014 5735 2024 5791
rect 2080 5735 2168 5791
rect 2014 5649 2026 5735
rect 2078 5649 2168 5735
rect 2014 5593 2024 5649
rect 2080 5593 2168 5649
rect 2014 5507 2026 5593
rect 2078 5507 2168 5593
rect 2014 5451 2024 5507
rect 2080 5451 2168 5507
rect 2014 5365 2026 5451
rect 2078 5365 2168 5451
rect 2014 5309 2024 5365
rect 2080 5309 2168 5365
rect 2014 5223 2026 5309
rect 2078 5223 2168 5309
rect 2014 5167 2024 5223
rect 2080 5167 2168 5223
rect 2014 5081 2026 5167
rect 2078 5081 2168 5167
rect 2014 5025 2024 5081
rect 2080 5025 2168 5081
rect 2014 4939 2026 5025
rect 2078 4939 2168 5025
rect 2014 4883 2024 4939
rect 2080 4883 2168 4939
rect 2014 4797 2026 4883
rect 2078 4797 2168 4883
rect 2014 4741 2024 4797
rect 2080 4741 2168 4797
rect 2014 4655 2026 4741
rect 2078 4655 2168 4741
rect 2014 4599 2024 4655
rect 2080 4599 2168 4655
rect 2014 4513 2026 4599
rect 2078 4513 2168 4599
rect 2014 4457 2024 4513
rect 2080 4457 2168 4513
rect 2014 4371 2026 4457
rect 2078 4371 2168 4457
rect 2014 4315 2024 4371
rect 2080 4315 2168 4371
rect 2014 4229 2026 4315
rect 2078 4229 2168 4315
rect 2014 4173 2024 4229
rect 2080 4173 2168 4229
rect 2014 4087 2026 4173
rect 2078 4087 2168 4173
rect 2014 4031 2024 4087
rect 2080 4031 2168 4087
rect 2014 3945 2026 4031
rect 2078 3945 2168 4031
rect 2014 3889 2024 3945
rect 2080 3889 2168 3945
rect 2014 3803 2026 3889
rect 2078 3803 2168 3889
rect 2014 3747 2024 3803
rect 2080 3747 2168 3803
rect 2014 3661 2026 3747
rect 2078 3661 2168 3747
rect 2014 3605 2024 3661
rect 2080 3605 2168 3661
rect 2014 3519 2026 3605
rect 2078 3519 2168 3605
rect 2014 3463 2024 3519
rect 2080 3463 2168 3519
rect 2014 3403 2026 3463
rect 2078 3403 2168 3463
rect 2014 3090 2168 3403
rect 2014 3034 2024 3090
rect 2080 3034 2168 3090
rect 2014 2948 2026 3034
rect 2078 2948 2168 3034
rect 2014 2892 2024 2948
rect 2080 2892 2168 2948
rect 2014 2806 2026 2892
rect 2078 2806 2168 2892
rect 2014 2750 2024 2806
rect 2080 2750 2168 2806
rect 2014 2664 2026 2750
rect 2078 2664 2168 2750
rect 2014 2608 2024 2664
rect 2080 2608 2168 2664
rect 2014 2522 2026 2608
rect 2078 2522 2168 2608
rect 2014 2466 2024 2522
rect 2080 2466 2168 2522
rect 2014 2380 2026 2466
rect 2078 2380 2168 2466
rect 2014 2324 2024 2380
rect 2080 2324 2168 2380
rect 2014 2238 2026 2324
rect 2078 2238 2168 2324
rect 2014 2182 2024 2238
rect 2080 2182 2168 2238
rect 2014 2096 2026 2182
rect 2078 2096 2168 2182
rect 2014 2040 2024 2096
rect 2080 2040 2168 2096
rect 2014 1954 2026 2040
rect 2078 1954 2168 2040
rect 2014 1898 2024 1954
rect 2080 1898 2168 1954
rect 2014 1812 2026 1898
rect 2078 1812 2168 1898
rect 2014 1756 2024 1812
rect 2080 1756 2168 1812
rect 2014 1670 2026 1756
rect 2078 1670 2168 1756
rect 2014 1614 2024 1670
rect 2080 1614 2168 1670
rect 2014 1528 2026 1614
rect 2078 1528 2168 1614
rect 2014 1472 2024 1528
rect 2080 1472 2168 1528
rect 2014 1386 2026 1472
rect 2078 1386 2168 1472
rect 2014 1330 2024 1386
rect 2080 1330 2168 1386
rect 2014 1244 2026 1330
rect 2078 1244 2168 1330
rect 2014 1188 2024 1244
rect 2080 1188 2168 1244
rect 2014 1102 2026 1188
rect 2078 1102 2168 1188
rect 2014 1046 2024 1102
rect 2080 1046 2168 1102
rect 2014 960 2026 1046
rect 2078 960 2168 1046
rect 2014 904 2024 960
rect 2080 904 2168 960
rect 2014 818 2026 904
rect 2078 843 2168 904
rect 2078 818 2090 843
rect 2014 762 2024 818
rect 2080 762 2090 818
rect 2014 676 2026 762
rect 2078 676 2090 762
rect 2014 620 2024 676
rect 2080 620 2090 676
rect 2014 519 2026 620
rect 2078 519 2090 620
rect 2014 507 2090 519
rect 2572 -1095 4216 8943
rect 4780 -1095 6424 8943
rect 6988 -1095 8632 8943
rect 9196 -1095 10840 8943
rect 11244 8836 11341 8843
rect 11244 8824 11415 8836
rect 11244 8799 11351 8824
rect 11403 8799 11415 8824
rect 11244 8743 11349 8799
rect 11405 8743 11415 8799
rect 11244 8657 11351 8743
rect 11403 8657 11415 8743
rect 11244 8601 11349 8657
rect 11405 8601 11415 8657
rect 11244 8515 11351 8601
rect 11403 8515 11415 8601
rect 11244 8459 11349 8515
rect 11405 8459 11415 8515
rect 11244 8373 11351 8459
rect 11403 8373 11415 8459
rect 11244 8317 11349 8373
rect 11405 8317 11415 8373
rect 11244 8231 11351 8317
rect 11403 8231 11415 8317
rect 11244 8175 11349 8231
rect 11405 8175 11415 8231
rect 11244 8089 11351 8175
rect 11403 8089 11415 8175
rect 11244 8033 11349 8089
rect 11405 8033 11415 8089
rect 11244 7947 11351 8033
rect 11403 7947 11415 8033
rect 11244 7891 11349 7947
rect 11405 7891 11415 7947
rect 11244 7805 11351 7891
rect 11403 7805 11415 7891
rect 11244 7749 11349 7805
rect 11405 7749 11415 7805
rect 11244 7663 11351 7749
rect 11403 7663 11415 7749
rect 11244 7607 11349 7663
rect 11405 7607 11415 7663
rect 11244 7521 11351 7607
rect 11403 7521 11415 7607
rect 11244 7465 11349 7521
rect 11405 7465 11415 7521
rect 11244 7379 11351 7465
rect 11403 7379 11415 7465
rect 11244 7323 11349 7379
rect 11405 7323 11415 7379
rect 11244 7237 11351 7323
rect 11403 7237 11415 7323
rect 11244 7181 11349 7237
rect 11405 7181 11415 7237
rect 11244 7095 11351 7181
rect 11403 7095 11415 7181
rect 11244 7039 11349 7095
rect 11405 7039 11415 7095
rect 11244 6953 11351 7039
rect 11403 6953 11415 7039
rect 11244 6897 11349 6953
rect 11405 6897 11415 6953
rect 11244 6811 11351 6897
rect 11403 6811 11415 6897
rect 11244 6755 11349 6811
rect 11405 6755 11415 6811
rect 11244 6669 11351 6755
rect 11403 6669 11415 6755
rect 11244 6613 11349 6669
rect 11405 6613 11415 6669
rect 11244 6588 11351 6613
rect 11403 6588 11415 6613
rect 11244 6576 11415 6588
rect 11244 6275 11341 6576
rect 11244 6263 11415 6275
rect 11244 6217 11351 6263
rect 11403 6217 11415 6263
rect 11244 6161 11349 6217
rect 11405 6161 11415 6217
rect 11244 6075 11351 6161
rect 11403 6075 11415 6161
rect 11244 6019 11349 6075
rect 11405 6019 11415 6075
rect 11244 5933 11351 6019
rect 11403 5933 11415 6019
rect 11244 5877 11349 5933
rect 11405 5877 11415 5933
rect 11244 5791 11351 5877
rect 11403 5791 11415 5877
rect 11244 5735 11349 5791
rect 11405 5735 11415 5791
rect 11244 5649 11351 5735
rect 11403 5649 11415 5735
rect 11244 5593 11349 5649
rect 11405 5593 11415 5649
rect 11244 5507 11351 5593
rect 11403 5507 11415 5593
rect 11244 5451 11349 5507
rect 11405 5451 11415 5507
rect 11244 5365 11351 5451
rect 11403 5365 11415 5451
rect 11244 5309 11349 5365
rect 11405 5309 11415 5365
rect 11244 5223 11351 5309
rect 11403 5223 11415 5309
rect 11244 5167 11349 5223
rect 11405 5167 11415 5223
rect 11244 5081 11351 5167
rect 11403 5081 11415 5167
rect 11244 5025 11349 5081
rect 11405 5025 11415 5081
rect 11244 4939 11351 5025
rect 11403 4939 11415 5025
rect 11244 4883 11349 4939
rect 11405 4883 11415 4939
rect 11244 4797 11351 4883
rect 11403 4797 11415 4883
rect 11244 4741 11349 4797
rect 11405 4741 11415 4797
rect 11244 4655 11351 4741
rect 11403 4655 11415 4741
rect 11244 4599 11349 4655
rect 11405 4599 11415 4655
rect 11244 4513 11351 4599
rect 11403 4513 11415 4599
rect 11244 4457 11349 4513
rect 11405 4457 11415 4513
rect 11244 4371 11351 4457
rect 11403 4371 11415 4457
rect 11244 4315 11349 4371
rect 11405 4315 11415 4371
rect 11244 4229 11351 4315
rect 11403 4229 11415 4315
rect 11244 4173 11349 4229
rect 11405 4173 11415 4229
rect 11244 4087 11351 4173
rect 11403 4087 11415 4173
rect 11244 4031 11349 4087
rect 11405 4031 11415 4087
rect 11244 3945 11351 4031
rect 11403 3945 11415 4031
rect 11244 3889 11349 3945
rect 11405 3889 11415 3945
rect 11244 3803 11351 3889
rect 11403 3803 11415 3889
rect 11244 3747 11349 3803
rect 11405 3747 11415 3803
rect 11244 3661 11351 3747
rect 11403 3661 11415 3747
rect 11244 3605 11349 3661
rect 11405 3605 11415 3661
rect 11244 3519 11351 3605
rect 11403 3519 11415 3605
rect 11244 3463 11349 3519
rect 11405 3463 11415 3519
rect 11244 3403 11351 3463
rect 11403 3403 11415 3463
rect 11244 3391 11415 3403
rect 11244 3100 11341 3391
rect 11244 3090 11415 3100
rect 11244 3034 11349 3090
rect 11405 3034 11415 3090
rect 11244 2948 11351 3034
rect 11403 2948 11415 3034
rect 11244 2892 11349 2948
rect 11405 2892 11415 2948
rect 11244 2806 11351 2892
rect 11403 2806 11415 2892
rect 11244 2750 11349 2806
rect 11405 2750 11415 2806
rect 11244 2664 11351 2750
rect 11403 2664 11415 2750
rect 11244 2608 11349 2664
rect 11405 2608 11415 2664
rect 11244 2522 11351 2608
rect 11403 2522 11415 2608
rect 11244 2466 11349 2522
rect 11405 2466 11415 2522
rect 11244 2380 11351 2466
rect 11403 2380 11415 2466
rect 11244 2324 11349 2380
rect 11405 2324 11415 2380
rect 11244 2238 11351 2324
rect 11403 2238 11415 2324
rect 11244 2182 11349 2238
rect 11405 2182 11415 2238
rect 11244 2096 11351 2182
rect 11403 2096 11415 2182
rect 11244 2040 11349 2096
rect 11405 2040 11415 2096
rect 11244 1954 11351 2040
rect 11403 1954 11415 2040
rect 11244 1898 11349 1954
rect 11405 1898 11415 1954
rect 11244 1812 11351 1898
rect 11403 1812 11415 1898
rect 11244 1756 11349 1812
rect 11405 1756 11415 1812
rect 11244 1670 11351 1756
rect 11403 1670 11415 1756
rect 11244 1614 11349 1670
rect 11405 1614 11415 1670
rect 11244 1528 11351 1614
rect 11403 1528 11415 1614
rect 11244 1472 11349 1528
rect 11405 1472 11415 1528
rect 11244 1386 11351 1472
rect 11403 1386 11415 1472
rect 11244 1330 11349 1386
rect 11405 1330 11415 1386
rect 11244 1244 11351 1330
rect 11403 1244 11415 1330
rect 11244 1188 11349 1244
rect 11405 1188 11415 1244
rect 11244 1102 11351 1188
rect 11403 1102 11415 1188
rect 11244 1046 11349 1102
rect 11405 1046 11415 1102
rect 11244 960 11351 1046
rect 11403 960 11415 1046
rect 11244 904 11349 960
rect 11405 904 11415 960
rect 11244 843 11351 904
rect 11339 818 11351 843
rect 11403 818 11415 904
rect 11339 762 11349 818
rect 11405 762 11415 818
rect 11339 676 11351 762
rect 11403 676 11415 762
rect 11339 620 11349 676
rect 11405 620 11415 676
rect 11339 519 11351 620
rect 11403 519 11415 620
rect 11339 507 11415 519
rect 11541 -1081 11781 8943
<< via2 >>
rect -165 12508 -109 12564
rect -23 12508 33 12564
rect -165 12366 -109 12422
rect -23 12366 33 12422
rect -165 12224 -109 12280
rect -23 12224 33 12280
rect -165 12082 -109 12138
rect -23 12082 33 12138
rect -165 11940 -109 11996
rect -23 11940 33 11996
rect -165 11798 -109 11854
rect -23 11798 33 11854
rect -165 11656 -109 11712
rect -23 11656 33 11712
rect -165 11514 -109 11570
rect -23 11514 33 11570
rect -300 10815 -244 10818
rect -158 10815 -102 10818
rect -16 10815 40 10818
rect -300 10763 -293 10815
rect -293 10763 -244 10815
rect -158 10763 -117 10815
rect -117 10763 -102 10815
rect -16 10763 7 10815
rect 7 10763 40 10815
rect -300 10762 -244 10763
rect -158 10762 -102 10763
rect -16 10762 40 10763
rect -300 10639 -293 10676
rect -293 10639 -244 10676
rect -158 10639 -117 10676
rect -117 10639 -102 10676
rect -16 10639 7 10676
rect 7 10639 40 10676
rect -300 10620 -244 10639
rect -158 10620 -102 10639
rect -16 10620 40 10639
rect -300 10515 -293 10534
rect -293 10515 -244 10534
rect -158 10515 -117 10534
rect -117 10515 -102 10534
rect -16 10515 7 10534
rect 7 10515 40 10534
rect -300 10478 -244 10515
rect -158 10478 -102 10515
rect -16 10478 40 10515
rect -300 10391 -293 10392
rect -293 10391 -244 10392
rect -158 10391 -117 10392
rect -117 10391 -102 10392
rect -16 10391 7 10392
rect 7 10391 40 10392
rect -300 10336 -244 10391
rect -158 10336 -102 10391
rect -16 10336 40 10391
rect -300 10195 -244 10250
rect -158 10195 -102 10250
rect -16 10195 40 10250
rect -300 10194 -293 10195
rect -293 10194 -244 10195
rect -158 10194 -117 10195
rect -117 10194 -102 10195
rect -16 10194 7 10195
rect 7 10194 40 10195
rect -300 10071 -244 10108
rect -158 10071 -102 10108
rect -16 10071 40 10108
rect -300 10052 -293 10071
rect -293 10052 -244 10071
rect -158 10052 -117 10071
rect -117 10052 -102 10071
rect -16 10052 7 10071
rect 7 10052 40 10071
rect -300 9947 -244 9966
rect -158 9947 -102 9966
rect -16 9947 40 9966
rect -300 9910 -293 9947
rect -293 9910 -244 9947
rect -158 9910 -117 9947
rect -117 9910 -102 9947
rect -16 9910 7 9947
rect 7 9910 40 9947
rect -300 9823 -244 9824
rect -158 9823 -102 9824
rect -16 9823 40 9824
rect -300 9771 -293 9823
rect -293 9771 -244 9823
rect -158 9771 -117 9823
rect -117 9771 -102 9823
rect -16 9771 7 9823
rect 7 9771 40 9823
rect -300 9768 -244 9771
rect -158 9768 -102 9771
rect -16 9768 40 9771
rect 1079 10815 1135 10818
rect 1079 10763 1089 10815
rect 1089 10763 1135 10815
rect 1079 10762 1135 10763
rect 1221 10762 1277 10818
rect 1363 10815 1419 10818
rect 1363 10763 1409 10815
rect 1409 10763 1419 10815
rect 1363 10762 1419 10763
rect 1079 10639 1089 10676
rect 1089 10639 1135 10676
rect 1079 10620 1135 10639
rect 1221 10620 1277 10676
rect 1363 10639 1409 10676
rect 1409 10639 1419 10676
rect 1363 10620 1419 10639
rect 1079 10515 1089 10534
rect 1089 10515 1135 10534
rect 1079 10478 1135 10515
rect 1221 10478 1277 10534
rect 1363 10515 1409 10534
rect 1409 10515 1419 10534
rect 1363 10478 1419 10515
rect 1079 10391 1089 10392
rect 1089 10391 1135 10392
rect 1079 10336 1135 10391
rect 1221 10336 1277 10392
rect 1363 10391 1409 10392
rect 1409 10391 1419 10392
rect 1363 10336 1419 10391
rect 1079 10195 1135 10250
rect 1079 10194 1089 10195
rect 1089 10194 1135 10195
rect 1221 10194 1277 10250
rect 1363 10195 1419 10250
rect 1363 10194 1409 10195
rect 1409 10194 1419 10195
rect 1079 10071 1135 10108
rect 1079 10052 1089 10071
rect 1089 10052 1135 10071
rect 1221 10052 1277 10108
rect 1363 10071 1419 10108
rect 1363 10052 1409 10071
rect 1409 10052 1419 10071
rect 1079 9947 1135 9966
rect 1079 9910 1089 9947
rect 1089 9910 1135 9947
rect 1221 9910 1277 9966
rect 1363 9947 1419 9966
rect 1363 9910 1409 9947
rect 1409 9910 1419 9947
rect 1079 9823 1135 9824
rect 1079 9771 1089 9823
rect 1089 9771 1135 9823
rect 1079 9768 1135 9771
rect 1221 9768 1277 9824
rect 1363 9823 1419 9824
rect 1363 9771 1409 9823
rect 1409 9771 1419 9823
rect 1363 9768 1419 9771
rect 12010 10815 12066 10818
rect 12010 10763 12020 10815
rect 12020 10763 12066 10815
rect 12010 10762 12066 10763
rect 12152 10762 12208 10818
rect 12294 10815 12350 10818
rect 12294 10763 12340 10815
rect 12340 10763 12350 10815
rect 12294 10762 12350 10763
rect 12010 10639 12020 10676
rect 12020 10639 12066 10676
rect 12010 10620 12066 10639
rect 12152 10620 12208 10676
rect 12294 10639 12340 10676
rect 12340 10639 12350 10676
rect 12294 10620 12350 10639
rect 12010 10515 12020 10534
rect 12020 10515 12066 10534
rect 12010 10478 12066 10515
rect 12152 10478 12208 10534
rect 12294 10515 12340 10534
rect 12340 10515 12350 10534
rect 12294 10478 12350 10515
rect 12010 10391 12020 10392
rect 12020 10391 12066 10392
rect 12010 10336 12066 10391
rect 12152 10336 12208 10392
rect 12294 10391 12340 10392
rect 12340 10391 12350 10392
rect 12294 10336 12350 10391
rect 12010 10195 12066 10250
rect 12010 10194 12020 10195
rect 12020 10194 12066 10195
rect 12152 10194 12208 10250
rect 12294 10195 12350 10250
rect 12294 10194 12340 10195
rect 12340 10194 12350 10195
rect 12010 10071 12066 10108
rect 12010 10052 12020 10071
rect 12020 10052 12066 10071
rect 12152 10052 12208 10108
rect 12294 10071 12350 10108
rect 12294 10052 12340 10071
rect 12340 10052 12350 10071
rect 12010 9947 12066 9966
rect 12010 9910 12020 9947
rect 12020 9910 12066 9947
rect 12152 9910 12208 9966
rect 12294 9947 12350 9966
rect 12294 9910 12340 9947
rect 12340 9910 12350 9947
rect 12010 9823 12066 9824
rect 12010 9771 12020 9823
rect 12020 9771 12066 9823
rect 12010 9768 12066 9771
rect 12152 9768 12208 9824
rect 12294 9823 12350 9824
rect 12294 9771 12340 9823
rect 12340 9771 12350 9823
rect 12294 9768 12350 9771
rect 13431 12508 13487 12564
rect 13573 12508 13629 12564
rect 13431 12366 13487 12422
rect 13573 12366 13629 12422
rect 13431 12224 13487 12280
rect 13573 12224 13629 12280
rect 13431 12082 13487 12138
rect 13573 12082 13629 12138
rect 13431 11940 13487 11996
rect 13573 11940 13629 11996
rect 13431 11798 13487 11854
rect 13573 11798 13629 11854
rect 13431 11656 13487 11712
rect 13573 11656 13629 11712
rect 13431 11514 13487 11570
rect 13573 11514 13629 11570
rect 13385 10815 13441 10818
rect 13527 10815 13583 10818
rect 13669 10815 13725 10818
rect 13385 10763 13418 10815
rect 13418 10763 13441 10815
rect 13527 10763 13542 10815
rect 13542 10763 13583 10815
rect 13669 10763 13718 10815
rect 13718 10763 13725 10815
rect 13385 10762 13441 10763
rect 13527 10762 13583 10763
rect 13669 10762 13725 10763
rect 13385 10639 13418 10676
rect 13418 10639 13441 10676
rect 13527 10639 13542 10676
rect 13542 10639 13583 10676
rect 13669 10639 13718 10676
rect 13718 10639 13725 10676
rect 13385 10620 13441 10639
rect 13527 10620 13583 10639
rect 13669 10620 13725 10639
rect 13385 10515 13418 10534
rect 13418 10515 13441 10534
rect 13527 10515 13542 10534
rect 13542 10515 13583 10534
rect 13669 10515 13718 10534
rect 13718 10515 13725 10534
rect 13385 10478 13441 10515
rect 13527 10478 13583 10515
rect 13669 10478 13725 10515
rect 13385 10391 13418 10392
rect 13418 10391 13441 10392
rect 13527 10391 13542 10392
rect 13542 10391 13583 10392
rect 13669 10391 13718 10392
rect 13718 10391 13725 10392
rect 13385 10336 13441 10391
rect 13527 10336 13583 10391
rect 13669 10336 13725 10391
rect 13385 10195 13441 10250
rect 13527 10195 13583 10250
rect 13669 10195 13725 10250
rect 13385 10194 13418 10195
rect 13418 10194 13441 10195
rect 13527 10194 13542 10195
rect 13542 10194 13583 10195
rect 13669 10194 13718 10195
rect 13718 10194 13725 10195
rect 13385 10071 13441 10108
rect 13527 10071 13583 10108
rect 13669 10071 13725 10108
rect 13385 10052 13418 10071
rect 13418 10052 13441 10071
rect 13527 10052 13542 10071
rect 13542 10052 13583 10071
rect 13669 10052 13718 10071
rect 13718 10052 13725 10071
rect 13385 9947 13441 9966
rect 13527 9947 13583 9966
rect 13669 9947 13725 9966
rect 13385 9910 13418 9947
rect 13418 9910 13441 9947
rect 13527 9910 13542 9947
rect 13542 9910 13583 9947
rect 13669 9910 13718 9947
rect 13718 9910 13725 9947
rect 13385 9823 13441 9824
rect 13527 9823 13583 9824
rect 13669 9823 13725 9824
rect 13385 9771 13418 9823
rect 13418 9771 13441 9823
rect 13527 9771 13542 9823
rect 13542 9771 13583 9823
rect 13669 9771 13718 9823
rect 13718 9771 13725 9823
rect 13385 9768 13441 9771
rect 13527 9768 13583 9771
rect 13669 9768 13725 9771
rect 2024 8743 2026 8799
rect 2026 8743 2078 8799
rect 2078 8743 2080 8799
rect 2024 8601 2026 8657
rect 2026 8601 2078 8657
rect 2078 8601 2080 8657
rect 2024 8459 2026 8515
rect 2026 8459 2078 8515
rect 2078 8459 2080 8515
rect 2024 8317 2026 8373
rect 2026 8317 2078 8373
rect 2078 8317 2080 8373
rect 2024 8175 2026 8231
rect 2026 8175 2078 8231
rect 2078 8175 2080 8231
rect 2024 8033 2026 8089
rect 2026 8033 2078 8089
rect 2078 8033 2080 8089
rect 2024 7891 2026 7947
rect 2026 7891 2078 7947
rect 2078 7891 2080 7947
rect 2024 7749 2026 7805
rect 2026 7749 2078 7805
rect 2078 7749 2080 7805
rect 2024 7607 2026 7663
rect 2026 7607 2078 7663
rect 2078 7607 2080 7663
rect 2024 7465 2026 7521
rect 2026 7465 2078 7521
rect 2078 7465 2080 7521
rect 2024 7323 2026 7379
rect 2026 7323 2078 7379
rect 2078 7323 2080 7379
rect 2024 7181 2026 7237
rect 2026 7181 2078 7237
rect 2078 7181 2080 7237
rect 2024 7039 2026 7095
rect 2026 7039 2078 7095
rect 2078 7039 2080 7095
rect 2024 6897 2026 6953
rect 2026 6897 2078 6953
rect 2078 6897 2080 6953
rect 2024 6755 2026 6811
rect 2026 6755 2078 6811
rect 2078 6755 2080 6811
rect 2024 6613 2026 6669
rect 2026 6613 2078 6669
rect 2078 6613 2080 6669
rect 2024 6161 2026 6217
rect 2026 6161 2078 6217
rect 2078 6161 2080 6217
rect 2024 6019 2026 6075
rect 2026 6019 2078 6075
rect 2078 6019 2080 6075
rect 2024 5877 2026 5933
rect 2026 5877 2078 5933
rect 2078 5877 2080 5933
rect 2024 5735 2026 5791
rect 2026 5735 2078 5791
rect 2078 5735 2080 5791
rect 2024 5593 2026 5649
rect 2026 5593 2078 5649
rect 2078 5593 2080 5649
rect 2024 5451 2026 5507
rect 2026 5451 2078 5507
rect 2078 5451 2080 5507
rect 2024 5309 2026 5365
rect 2026 5309 2078 5365
rect 2078 5309 2080 5365
rect 2024 5167 2026 5223
rect 2026 5167 2078 5223
rect 2078 5167 2080 5223
rect 2024 5025 2026 5081
rect 2026 5025 2078 5081
rect 2078 5025 2080 5081
rect 2024 4883 2026 4939
rect 2026 4883 2078 4939
rect 2078 4883 2080 4939
rect 2024 4741 2026 4797
rect 2026 4741 2078 4797
rect 2078 4741 2080 4797
rect 2024 4599 2026 4655
rect 2026 4599 2078 4655
rect 2078 4599 2080 4655
rect 2024 4457 2026 4513
rect 2026 4457 2078 4513
rect 2078 4457 2080 4513
rect 2024 4315 2026 4371
rect 2026 4315 2078 4371
rect 2078 4315 2080 4371
rect 2024 4173 2026 4229
rect 2026 4173 2078 4229
rect 2078 4173 2080 4229
rect 2024 4031 2026 4087
rect 2026 4031 2078 4087
rect 2078 4031 2080 4087
rect 2024 3889 2026 3945
rect 2026 3889 2078 3945
rect 2078 3889 2080 3945
rect 2024 3747 2026 3803
rect 2026 3747 2078 3803
rect 2078 3747 2080 3803
rect 2024 3605 2026 3661
rect 2026 3605 2078 3661
rect 2078 3605 2080 3661
rect 2024 3463 2026 3519
rect 2026 3463 2078 3519
rect 2078 3463 2080 3519
rect 2024 3067 2080 3090
rect 2024 3034 2026 3067
rect 2026 3034 2078 3067
rect 2078 3034 2080 3067
rect 2024 2892 2026 2948
rect 2026 2892 2078 2948
rect 2078 2892 2080 2948
rect 2024 2750 2026 2806
rect 2026 2750 2078 2806
rect 2078 2750 2080 2806
rect 2024 2608 2026 2664
rect 2026 2608 2078 2664
rect 2078 2608 2080 2664
rect 2024 2466 2026 2522
rect 2026 2466 2078 2522
rect 2078 2466 2080 2522
rect 2024 2324 2026 2380
rect 2026 2324 2078 2380
rect 2078 2324 2080 2380
rect 2024 2182 2026 2238
rect 2026 2182 2078 2238
rect 2078 2182 2080 2238
rect 2024 2040 2026 2096
rect 2026 2040 2078 2096
rect 2078 2040 2080 2096
rect 2024 1898 2026 1954
rect 2026 1898 2078 1954
rect 2078 1898 2080 1954
rect 2024 1756 2026 1812
rect 2026 1756 2078 1812
rect 2078 1756 2080 1812
rect 2024 1614 2026 1670
rect 2026 1614 2078 1670
rect 2078 1614 2080 1670
rect 2024 1472 2026 1528
rect 2026 1472 2078 1528
rect 2078 1472 2080 1528
rect 2024 1330 2026 1386
rect 2026 1330 2078 1386
rect 2078 1330 2080 1386
rect 2024 1188 2026 1244
rect 2026 1188 2078 1244
rect 2078 1188 2080 1244
rect 2024 1046 2026 1102
rect 2026 1046 2078 1102
rect 2078 1046 2080 1102
rect 2024 904 2026 960
rect 2026 904 2078 960
rect 2078 904 2080 960
rect 2024 762 2026 818
rect 2026 762 2078 818
rect 2078 762 2080 818
rect 2024 620 2026 676
rect 2026 620 2078 676
rect 2078 620 2080 676
rect 11349 8743 11351 8799
rect 11351 8743 11403 8799
rect 11403 8743 11405 8799
rect 11349 8601 11351 8657
rect 11351 8601 11403 8657
rect 11403 8601 11405 8657
rect 11349 8459 11351 8515
rect 11351 8459 11403 8515
rect 11403 8459 11405 8515
rect 11349 8317 11351 8373
rect 11351 8317 11403 8373
rect 11403 8317 11405 8373
rect 11349 8175 11351 8231
rect 11351 8175 11403 8231
rect 11403 8175 11405 8231
rect 11349 8033 11351 8089
rect 11351 8033 11403 8089
rect 11403 8033 11405 8089
rect 11349 7891 11351 7947
rect 11351 7891 11403 7947
rect 11403 7891 11405 7947
rect 11349 7749 11351 7805
rect 11351 7749 11403 7805
rect 11403 7749 11405 7805
rect 11349 7607 11351 7663
rect 11351 7607 11403 7663
rect 11403 7607 11405 7663
rect 11349 7465 11351 7521
rect 11351 7465 11403 7521
rect 11403 7465 11405 7521
rect 11349 7323 11351 7379
rect 11351 7323 11403 7379
rect 11403 7323 11405 7379
rect 11349 7181 11351 7237
rect 11351 7181 11403 7237
rect 11403 7181 11405 7237
rect 11349 7039 11351 7095
rect 11351 7039 11403 7095
rect 11403 7039 11405 7095
rect 11349 6897 11351 6953
rect 11351 6897 11403 6953
rect 11403 6897 11405 6953
rect 11349 6755 11351 6811
rect 11351 6755 11403 6811
rect 11403 6755 11405 6811
rect 11349 6613 11351 6669
rect 11351 6613 11403 6669
rect 11403 6613 11405 6669
rect 11349 6161 11351 6217
rect 11351 6161 11403 6217
rect 11403 6161 11405 6217
rect 11349 6019 11351 6075
rect 11351 6019 11403 6075
rect 11403 6019 11405 6075
rect 11349 5877 11351 5933
rect 11351 5877 11403 5933
rect 11403 5877 11405 5933
rect 11349 5735 11351 5791
rect 11351 5735 11403 5791
rect 11403 5735 11405 5791
rect 11349 5593 11351 5649
rect 11351 5593 11403 5649
rect 11403 5593 11405 5649
rect 11349 5451 11351 5507
rect 11351 5451 11403 5507
rect 11403 5451 11405 5507
rect 11349 5309 11351 5365
rect 11351 5309 11403 5365
rect 11403 5309 11405 5365
rect 11349 5167 11351 5223
rect 11351 5167 11403 5223
rect 11403 5167 11405 5223
rect 11349 5025 11351 5081
rect 11351 5025 11403 5081
rect 11403 5025 11405 5081
rect 11349 4883 11351 4939
rect 11351 4883 11403 4939
rect 11403 4883 11405 4939
rect 11349 4741 11351 4797
rect 11351 4741 11403 4797
rect 11403 4741 11405 4797
rect 11349 4599 11351 4655
rect 11351 4599 11403 4655
rect 11403 4599 11405 4655
rect 11349 4457 11351 4513
rect 11351 4457 11403 4513
rect 11403 4457 11405 4513
rect 11349 4315 11351 4371
rect 11351 4315 11403 4371
rect 11403 4315 11405 4371
rect 11349 4173 11351 4229
rect 11351 4173 11403 4229
rect 11403 4173 11405 4229
rect 11349 4031 11351 4087
rect 11351 4031 11403 4087
rect 11403 4031 11405 4087
rect 11349 3889 11351 3945
rect 11351 3889 11403 3945
rect 11403 3889 11405 3945
rect 11349 3747 11351 3803
rect 11351 3747 11403 3803
rect 11403 3747 11405 3803
rect 11349 3605 11351 3661
rect 11351 3605 11403 3661
rect 11403 3605 11405 3661
rect 11349 3463 11351 3519
rect 11351 3463 11403 3519
rect 11403 3463 11405 3519
rect 11349 3067 11405 3090
rect 11349 3034 11351 3067
rect 11351 3034 11403 3067
rect 11403 3034 11405 3067
rect 11349 2892 11351 2948
rect 11351 2892 11403 2948
rect 11403 2892 11405 2948
rect 11349 2750 11351 2806
rect 11351 2750 11403 2806
rect 11403 2750 11405 2806
rect 11349 2608 11351 2664
rect 11351 2608 11403 2664
rect 11403 2608 11405 2664
rect 11349 2466 11351 2522
rect 11351 2466 11403 2522
rect 11403 2466 11405 2522
rect 11349 2324 11351 2380
rect 11351 2324 11403 2380
rect 11403 2324 11405 2380
rect 11349 2182 11351 2238
rect 11351 2182 11403 2238
rect 11403 2182 11405 2238
rect 11349 2040 11351 2096
rect 11351 2040 11403 2096
rect 11403 2040 11405 2096
rect 11349 1898 11351 1954
rect 11351 1898 11403 1954
rect 11403 1898 11405 1954
rect 11349 1756 11351 1812
rect 11351 1756 11403 1812
rect 11403 1756 11405 1812
rect 11349 1614 11351 1670
rect 11351 1614 11403 1670
rect 11403 1614 11405 1670
rect 11349 1472 11351 1528
rect 11351 1472 11403 1528
rect 11403 1472 11405 1528
rect 11349 1330 11351 1386
rect 11351 1330 11403 1386
rect 11403 1330 11405 1386
rect 11349 1188 11351 1244
rect 11351 1188 11403 1244
rect 11403 1188 11405 1244
rect 11349 1046 11351 1102
rect 11351 1046 11403 1102
rect 11403 1046 11405 1102
rect 11349 904 11351 960
rect 11351 904 11403 960
rect 11403 904 11405 960
rect 11349 762 11351 818
rect 11351 762 11403 818
rect 11403 762 11405 818
rect 11349 620 11351 676
rect 11351 620 11403 676
rect 11403 620 11405 676
<< metal3 >>
rect -175 12564 43 12574
rect -175 12508 -165 12564
rect -109 12508 -23 12564
rect 33 12508 43 12564
rect -175 12422 43 12508
rect -175 12366 -165 12422
rect -109 12366 -23 12422
rect 33 12366 43 12422
rect -175 12280 43 12366
rect -175 12224 -165 12280
rect -109 12224 -23 12280
rect 33 12224 43 12280
rect -175 12138 43 12224
rect -175 12082 -165 12138
rect -109 12082 -23 12138
rect 33 12082 43 12138
rect -175 11996 43 12082
rect -175 11940 -165 11996
rect -109 11940 -23 11996
rect 33 11940 43 11996
rect -175 11854 43 11940
rect -175 11798 -165 11854
rect -109 11798 -23 11854
rect 33 11798 43 11854
rect -175 11712 43 11798
rect -175 11656 -165 11712
rect -109 11656 -23 11712
rect 33 11656 43 11712
rect -175 11570 43 11656
rect -175 11514 -165 11570
rect -109 11514 -23 11570
rect 33 11514 43 11570
rect -175 11504 43 11514
rect 13421 12564 13639 12574
rect 13421 12508 13431 12564
rect 13487 12508 13573 12564
rect 13629 12508 13639 12564
rect 13421 12422 13639 12508
rect 13421 12366 13431 12422
rect 13487 12366 13573 12422
rect 13629 12366 13639 12422
rect 13421 12280 13639 12366
rect 13421 12224 13431 12280
rect 13487 12224 13573 12280
rect 13629 12224 13639 12280
rect 13421 12138 13639 12224
rect 13421 12082 13431 12138
rect 13487 12082 13573 12138
rect 13629 12082 13639 12138
rect 13421 11996 13639 12082
rect 13421 11940 13431 11996
rect 13487 11940 13573 11996
rect 13629 11940 13639 11996
rect 13421 11854 13639 11940
rect 13421 11798 13431 11854
rect 13487 11798 13573 11854
rect 13629 11798 13639 11854
rect 13421 11712 13639 11798
rect 13421 11656 13431 11712
rect 13487 11656 13573 11712
rect 13629 11656 13639 11712
rect 13421 11570 13639 11656
rect 13421 11514 13431 11570
rect 13487 11514 13573 11570
rect 13629 11514 13639 11570
rect 13421 11504 13639 11514
rect -310 10818 50 10828
rect -310 10762 -300 10818
rect -244 10762 -158 10818
rect -102 10762 -16 10818
rect 40 10762 50 10818
rect -310 10676 50 10762
rect -310 10620 -300 10676
rect -244 10620 -158 10676
rect -102 10620 -16 10676
rect 40 10620 50 10676
rect -310 10534 50 10620
rect -310 10478 -300 10534
rect -244 10478 -158 10534
rect -102 10478 -16 10534
rect 40 10478 50 10534
rect -310 10392 50 10478
rect -310 10336 -300 10392
rect -244 10336 -158 10392
rect -102 10336 -16 10392
rect 40 10336 50 10392
rect -310 10250 50 10336
rect -310 10194 -300 10250
rect -244 10194 -158 10250
rect -102 10194 -16 10250
rect 40 10194 50 10250
rect -310 10108 50 10194
rect -310 10052 -300 10108
rect -244 10052 -158 10108
rect -102 10052 -16 10108
rect 40 10052 50 10108
rect -310 9966 50 10052
rect -310 9910 -300 9966
rect -244 9910 -158 9966
rect -102 9910 -16 9966
rect 40 9910 50 9966
rect -310 9824 50 9910
rect -310 9768 -300 9824
rect -244 9768 -158 9824
rect -102 9768 -16 9824
rect 40 9768 50 9824
rect -310 9758 50 9768
rect 1069 10818 1429 10828
rect 1069 10762 1079 10818
rect 1135 10762 1221 10818
rect 1277 10762 1363 10818
rect 1419 10762 1429 10818
rect 1069 10676 1429 10762
rect 1069 10620 1079 10676
rect 1135 10620 1221 10676
rect 1277 10620 1363 10676
rect 1419 10620 1429 10676
rect 1069 10534 1429 10620
rect 1069 10478 1079 10534
rect 1135 10478 1221 10534
rect 1277 10478 1363 10534
rect 1419 10478 1429 10534
rect 1069 10392 1429 10478
rect 1069 10336 1079 10392
rect 1135 10336 1221 10392
rect 1277 10336 1363 10392
rect 1419 10336 1429 10392
rect 1069 10250 1429 10336
rect 1069 10194 1079 10250
rect 1135 10194 1221 10250
rect 1277 10194 1363 10250
rect 1419 10194 1429 10250
rect 1069 10108 1429 10194
rect 1069 10052 1079 10108
rect 1135 10052 1221 10108
rect 1277 10052 1363 10108
rect 1419 10052 1429 10108
rect 1069 9966 1429 10052
rect 1069 9910 1079 9966
rect 1135 9910 1221 9966
rect 1277 9910 1363 9966
rect 1419 9910 1429 9966
rect 1069 9824 1429 9910
rect 1069 9768 1079 9824
rect 1135 9768 1221 9824
rect 1277 9768 1363 9824
rect 1419 9768 1429 9824
rect 1069 9758 1429 9768
rect 12000 10818 12360 10828
rect 12000 10762 12010 10818
rect 12066 10762 12152 10818
rect 12208 10762 12294 10818
rect 12350 10762 12360 10818
rect 12000 10676 12360 10762
rect 12000 10620 12010 10676
rect 12066 10620 12152 10676
rect 12208 10620 12294 10676
rect 12350 10620 12360 10676
rect 12000 10534 12360 10620
rect 12000 10478 12010 10534
rect 12066 10478 12152 10534
rect 12208 10478 12294 10534
rect 12350 10478 12360 10534
rect 12000 10392 12360 10478
rect 12000 10336 12010 10392
rect 12066 10336 12152 10392
rect 12208 10336 12294 10392
rect 12350 10336 12360 10392
rect 12000 10250 12360 10336
rect 12000 10194 12010 10250
rect 12066 10194 12152 10250
rect 12208 10194 12294 10250
rect 12350 10194 12360 10250
rect 12000 10108 12360 10194
rect 12000 10052 12010 10108
rect 12066 10052 12152 10108
rect 12208 10052 12294 10108
rect 12350 10052 12360 10108
rect 12000 9966 12360 10052
rect 12000 9910 12010 9966
rect 12066 9910 12152 9966
rect 12208 9910 12294 9966
rect 12350 9910 12360 9966
rect 12000 9824 12360 9910
rect 12000 9768 12010 9824
rect 12066 9768 12152 9824
rect 12208 9768 12294 9824
rect 12350 9768 12360 9824
rect 12000 9758 12360 9768
rect 13375 10818 13735 10828
rect 13375 10762 13385 10818
rect 13441 10762 13527 10818
rect 13583 10762 13669 10818
rect 13725 10762 13735 10818
rect 13375 10676 13735 10762
rect 13375 10620 13385 10676
rect 13441 10620 13527 10676
rect 13583 10620 13669 10676
rect 13725 10620 13735 10676
rect 13375 10534 13735 10620
rect 13375 10478 13385 10534
rect 13441 10478 13527 10534
rect 13583 10478 13669 10534
rect 13725 10478 13735 10534
rect 13375 10392 13735 10478
rect 13375 10336 13385 10392
rect 13441 10336 13527 10392
rect 13583 10336 13669 10392
rect 13725 10336 13735 10392
rect 13375 10250 13735 10336
rect 13375 10194 13385 10250
rect 13441 10194 13527 10250
rect 13583 10194 13669 10250
rect 13725 10194 13735 10250
rect 13375 10108 13735 10194
rect 13375 10052 13385 10108
rect 13441 10052 13527 10108
rect 13583 10052 13669 10108
rect 13725 10052 13735 10108
rect 13375 9966 13735 10052
rect 13375 9910 13385 9966
rect 13441 9910 13527 9966
rect 13583 9910 13669 9966
rect 13725 9910 13735 9966
rect 13375 9824 13735 9910
rect 13375 9768 13385 9824
rect 13441 9768 13527 9824
rect 13583 9768 13669 9824
rect 13725 9768 13735 9824
rect 13375 9758 13735 9768
rect 2014 8799 2090 8809
rect 2014 8743 2024 8799
rect 2080 8743 2090 8799
rect 2014 8657 2090 8743
rect 2014 8601 2024 8657
rect 2080 8601 2090 8657
rect 2014 8515 2090 8601
rect 2014 8459 2024 8515
rect 2080 8459 2090 8515
rect 2014 8373 2090 8459
rect 2014 8317 2024 8373
rect 2080 8317 2090 8373
rect 2014 8231 2090 8317
rect 2014 8175 2024 8231
rect 2080 8175 2090 8231
rect 2014 8089 2090 8175
rect 2014 8033 2024 8089
rect 2080 8033 2090 8089
rect 2014 7947 2090 8033
rect 2014 7891 2024 7947
rect 2080 7891 2090 7947
rect 2014 7805 2090 7891
rect 2014 7749 2024 7805
rect 2080 7749 2090 7805
rect 2014 7663 2090 7749
rect 2014 7607 2024 7663
rect 2080 7607 2090 7663
rect 2014 7521 2090 7607
rect 2014 7465 2024 7521
rect 2080 7465 2090 7521
rect 2014 7379 2090 7465
rect 2014 7323 2024 7379
rect 2080 7323 2090 7379
rect 2014 7237 2090 7323
rect 2014 7181 2024 7237
rect 2080 7181 2090 7237
rect 2014 7095 2090 7181
rect 2014 7039 2024 7095
rect 2080 7039 2090 7095
rect 2014 6953 2090 7039
rect 2014 6897 2024 6953
rect 2080 6897 2090 6953
rect 2014 6811 2090 6897
rect 2014 6755 2024 6811
rect 2080 6755 2090 6811
rect 2014 6669 2090 6755
rect 2014 6613 2024 6669
rect 2080 6613 2090 6669
rect 2014 6603 2090 6613
rect 11339 8799 11415 8809
rect 11339 8743 11349 8799
rect 11405 8743 11415 8799
rect 11339 8657 11415 8743
rect 11339 8601 11349 8657
rect 11405 8601 11415 8657
rect 11339 8515 11415 8601
rect 11339 8459 11349 8515
rect 11405 8459 11415 8515
rect 11339 8373 11415 8459
rect 11339 8317 11349 8373
rect 11405 8317 11415 8373
rect 11339 8231 11415 8317
rect 11339 8175 11349 8231
rect 11405 8175 11415 8231
rect 11339 8089 11415 8175
rect 11339 8033 11349 8089
rect 11405 8033 11415 8089
rect 11339 7947 11415 8033
rect 11339 7891 11349 7947
rect 11405 7891 11415 7947
rect 11339 7805 11415 7891
rect 11339 7749 11349 7805
rect 11405 7749 11415 7805
rect 11339 7663 11415 7749
rect 11339 7607 11349 7663
rect 11405 7607 11415 7663
rect 11339 7521 11415 7607
rect 11339 7465 11349 7521
rect 11405 7465 11415 7521
rect 11339 7379 11415 7465
rect 11339 7323 11349 7379
rect 11405 7323 11415 7379
rect 11339 7237 11415 7323
rect 11339 7181 11349 7237
rect 11405 7181 11415 7237
rect 11339 7095 11415 7181
rect 11339 7039 11349 7095
rect 11405 7039 11415 7095
rect 11339 6953 11415 7039
rect 11339 6897 11349 6953
rect 11405 6897 11415 6953
rect 11339 6811 11415 6897
rect 11339 6755 11349 6811
rect 11405 6755 11415 6811
rect 11339 6669 11415 6755
rect 11339 6613 11349 6669
rect 11405 6613 11415 6669
rect 11339 6603 11415 6613
rect 2014 6217 2090 6227
rect 2014 6161 2024 6217
rect 2080 6161 2090 6217
rect 2014 6075 2090 6161
rect 2014 6019 2024 6075
rect 2080 6019 2090 6075
rect 2014 5933 2090 6019
rect 2014 5877 2024 5933
rect 2080 5877 2090 5933
rect 2014 5791 2090 5877
rect 2014 5735 2024 5791
rect 2080 5735 2090 5791
rect 2014 5649 2090 5735
rect 2014 5593 2024 5649
rect 2080 5593 2090 5649
rect 2014 5507 2090 5593
rect 2014 5451 2024 5507
rect 2080 5451 2090 5507
rect 2014 5365 2090 5451
rect 2014 5309 2024 5365
rect 2080 5309 2090 5365
rect 2014 5223 2090 5309
rect 2014 5167 2024 5223
rect 2080 5167 2090 5223
rect 2014 5081 2090 5167
rect 2014 5025 2024 5081
rect 2080 5025 2090 5081
rect 2014 4939 2090 5025
rect 2014 4883 2024 4939
rect 2080 4883 2090 4939
rect 2014 4797 2090 4883
rect 2014 4741 2024 4797
rect 2080 4741 2090 4797
rect 2014 4655 2090 4741
rect 2014 4599 2024 4655
rect 2080 4599 2090 4655
rect 2014 4513 2090 4599
rect 2014 4457 2024 4513
rect 2080 4457 2090 4513
rect 2014 4371 2090 4457
rect 2014 4315 2024 4371
rect 2080 4315 2090 4371
rect 2014 4229 2090 4315
rect 2014 4173 2024 4229
rect 2080 4173 2090 4229
rect 2014 4087 2090 4173
rect 2014 4031 2024 4087
rect 2080 4031 2090 4087
rect 2014 3945 2090 4031
rect 2014 3889 2024 3945
rect 2080 3889 2090 3945
rect 2014 3803 2090 3889
rect 2014 3747 2024 3803
rect 2080 3747 2090 3803
rect 2014 3661 2090 3747
rect 2014 3605 2024 3661
rect 2080 3605 2090 3661
rect 2014 3519 2090 3605
rect 2014 3463 2024 3519
rect 2080 3463 2090 3519
rect 2014 3453 2090 3463
rect 11339 6217 11415 6227
rect 11339 6161 11349 6217
rect 11405 6161 11415 6217
rect 11339 6075 11415 6161
rect 11339 6019 11349 6075
rect 11405 6019 11415 6075
rect 11339 5933 11415 6019
rect 11339 5877 11349 5933
rect 11405 5877 11415 5933
rect 11339 5791 11415 5877
rect 11339 5735 11349 5791
rect 11405 5735 11415 5791
rect 11339 5649 11415 5735
rect 11339 5593 11349 5649
rect 11405 5593 11415 5649
rect 11339 5507 11415 5593
rect 11339 5451 11349 5507
rect 11405 5451 11415 5507
rect 11339 5365 11415 5451
rect 11339 5309 11349 5365
rect 11405 5309 11415 5365
rect 11339 5223 11415 5309
rect 11339 5167 11349 5223
rect 11405 5167 11415 5223
rect 11339 5081 11415 5167
rect 11339 5025 11349 5081
rect 11405 5025 11415 5081
rect 11339 4939 11415 5025
rect 11339 4883 11349 4939
rect 11405 4883 11415 4939
rect 11339 4797 11415 4883
rect 11339 4741 11349 4797
rect 11405 4741 11415 4797
rect 11339 4655 11415 4741
rect 11339 4599 11349 4655
rect 11405 4599 11415 4655
rect 11339 4513 11415 4599
rect 11339 4457 11349 4513
rect 11405 4457 11415 4513
rect 11339 4371 11415 4457
rect 11339 4315 11349 4371
rect 11405 4315 11415 4371
rect 11339 4229 11415 4315
rect 11339 4173 11349 4229
rect 11405 4173 11415 4229
rect 11339 4087 11415 4173
rect 11339 4031 11349 4087
rect 11405 4031 11415 4087
rect 11339 3945 11415 4031
rect 11339 3889 11349 3945
rect 11405 3889 11415 3945
rect 11339 3803 11415 3889
rect 11339 3747 11349 3803
rect 11405 3747 11415 3803
rect 11339 3661 11415 3747
rect 11339 3605 11349 3661
rect 11405 3605 11415 3661
rect 11339 3519 11415 3605
rect 11339 3463 11349 3519
rect 11405 3463 11415 3519
rect 11339 3453 11415 3463
rect 2014 3090 2090 3100
rect 2014 3034 2024 3090
rect 2080 3034 2090 3090
rect 2014 2948 2090 3034
rect 2014 2892 2024 2948
rect 2080 2892 2090 2948
rect 2014 2806 2090 2892
rect 2014 2750 2024 2806
rect 2080 2750 2090 2806
rect 2014 2664 2090 2750
rect 2014 2608 2024 2664
rect 2080 2608 2090 2664
rect 2014 2522 2090 2608
rect 2014 2466 2024 2522
rect 2080 2466 2090 2522
rect 2014 2380 2090 2466
rect 2014 2324 2024 2380
rect 2080 2324 2090 2380
rect 2014 2238 2090 2324
rect 2014 2182 2024 2238
rect 2080 2182 2090 2238
rect 2014 2096 2090 2182
rect 2014 2040 2024 2096
rect 2080 2040 2090 2096
rect 2014 1954 2090 2040
rect 2014 1898 2024 1954
rect 2080 1898 2090 1954
rect 2014 1812 2090 1898
rect 2014 1756 2024 1812
rect 2080 1756 2090 1812
rect 2014 1670 2090 1756
rect 2014 1614 2024 1670
rect 2080 1614 2090 1670
rect 2014 1528 2090 1614
rect 2014 1472 2024 1528
rect 2080 1472 2090 1528
rect 2014 1386 2090 1472
rect 2014 1330 2024 1386
rect 2080 1330 2090 1386
rect 2014 1244 2090 1330
rect 2014 1188 2024 1244
rect 2080 1188 2090 1244
rect 2014 1102 2090 1188
rect 2014 1046 2024 1102
rect 2080 1046 2090 1102
rect 2014 960 2090 1046
rect 2014 904 2024 960
rect 2080 904 2090 960
rect 2014 818 2090 904
rect 2014 762 2024 818
rect 2080 762 2090 818
rect 2014 676 2090 762
rect 2014 620 2024 676
rect 2080 620 2090 676
rect 2014 610 2090 620
rect 11339 3090 11415 3100
rect 11339 3034 11349 3090
rect 11405 3034 11415 3090
rect 11339 2948 11415 3034
rect 11339 2892 11349 2948
rect 11405 2892 11415 2948
rect 11339 2806 11415 2892
rect 11339 2750 11349 2806
rect 11405 2750 11415 2806
rect 11339 2664 11415 2750
rect 11339 2608 11349 2664
rect 11405 2608 11415 2664
rect 11339 2522 11415 2608
rect 11339 2466 11349 2522
rect 11405 2466 11415 2522
rect 11339 2380 11415 2466
rect 11339 2324 11349 2380
rect 11405 2324 11415 2380
rect 11339 2238 11415 2324
rect 11339 2182 11349 2238
rect 11405 2182 11415 2238
rect 11339 2096 11415 2182
rect 11339 2040 11349 2096
rect 11405 2040 11415 2096
rect 11339 1954 11415 2040
rect 11339 1898 11349 1954
rect 11405 1898 11415 1954
rect 11339 1812 11415 1898
rect 11339 1756 11349 1812
rect 11405 1756 11415 1812
rect 11339 1670 11415 1756
rect 11339 1614 11349 1670
rect 11405 1614 11415 1670
rect 11339 1528 11415 1614
rect 11339 1472 11349 1528
rect 11405 1472 11415 1528
rect 11339 1386 11415 1472
rect 11339 1330 11349 1386
rect 11405 1330 11415 1386
rect 11339 1244 11415 1330
rect 11339 1188 11349 1244
rect 11405 1188 11415 1244
rect 11339 1102 11415 1188
rect 11339 1046 11349 1102
rect 11405 1046 11415 1102
rect 11339 960 11415 1046
rect 11339 904 11349 960
rect 11405 904 11415 960
rect 11339 818 11415 904
rect 11339 762 11349 818
rect 11405 762 11415 818
rect 11339 676 11415 762
rect 11339 620 11349 676
rect 11405 620 11415 676
rect 11339 610 11415 620
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1669390400
transform 0 1 11971 1 0 8990
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1669390400
transform 0 1 11971 1 0 9156
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1669390400
transform 0 1 11971 1 0 9316
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1669390400
transform 0 1 11971 1 0 9484
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1669390400
transform 0 -1 1507 1 0 9484
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_5
timestamp 1669390400
transform 0 -1 1507 1 0 8990
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_6
timestamp 1669390400
transform 0 -1 1507 1 0 9156
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_7
timestamp 1669390400
transform 0 -1 1507 1 0 9316
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_0
timestamp 1669390400
transform 1 0 2052 0 1 7706
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_1
timestamp 1669390400
transform 1 0 11377 0 1 7706
box 0 0 1 1
use M2_M1_CDNS_40661953145276  M2_M1_CDNS_40661953145276_0
timestamp 1669390400
transform 1 0 -66 0 1 12039
box 0 0 1 1
use M2_M1_CDNS_40661953145276  M2_M1_CDNS_40661953145276_1
timestamp 1669390400
transform 1 0 13530 0 1 12039
box 0 0 1 1
use M2_M1_CDNS_40661953145279  M2_M1_CDNS_40661953145279_0
timestamp 1669390400
transform 1 0 2052 0 1 4833
box 0 0 1 1
use M2_M1_CDNS_40661953145279  M2_M1_CDNS_40661953145279_1
timestamp 1669390400
transform 1 0 11377 0 1 4833
box 0 0 1 1
use M2_M1_CDNS_40661953145280  M2_M1_CDNS_40661953145280_0
timestamp 1669390400
transform 1 0 2052 0 1 1793
box 0 0 1 1
use M2_M1_CDNS_40661953145280  M2_M1_CDNS_40661953145280_1
timestamp 1669390400
transform 1 0 11377 0 1 1793
box 0 0 1 1
use M2_M1_CDNS_40661953145281  M2_M1_CDNS_40661953145281_0
timestamp 1669390400
transform 1 0 1249 0 1 10293
box 0 0 1 1
use M2_M1_CDNS_40661953145281  M2_M1_CDNS_40661953145281_1
timestamp 1669390400
transform 1 0 12180 0 1 10293
box 0 0 1 1
use M2_M1_CDNS_40661953145282  M2_M1_CDNS_40661953145282_0
timestamp 1669390400
transform -1 0 13568 0 1 10293
box 0 0 1 1
use M2_M1_CDNS_40661953145282  M2_M1_CDNS_40661953145282_1
timestamp 1669390400
transform 1 0 -143 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145199  M3_M2_CDNS_40661953145199_0
timestamp 1669390400
transform 1 0 11377 0 1 1855
box 0 0 1 1
use M3_M2_CDNS_40661953145199  M3_M2_CDNS_40661953145199_1
timestamp 1669390400
transform 1 0 2052 0 1 1855
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_0
timestamp 1669390400
transform 1 0 11377 0 1 7706
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_1
timestamp 1669390400
transform 1 0 2052 0 1 7706
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_0
timestamp 1669390400
transform -1 0 13555 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_1
timestamp 1669390400
transform 1 0 12180 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_2
timestamp 1669390400
transform 1 0 1249 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145263  M3_M2_CDNS_40661953145263_3
timestamp 1669390400
transform 1 0 -130 0 1 10293
box 0 0 1 1
use M3_M2_CDNS_40661953145277  M3_M2_CDNS_40661953145277_0
timestamp 1669390400
transform 1 0 2052 0 1 4840
box 0 0 1 1
use M3_M2_CDNS_40661953145277  M3_M2_CDNS_40661953145277_1
timestamp 1669390400
transform 1 0 11377 0 1 4840
box 0 0 1 1
use M3_M2_CDNS_40661953145278  M3_M2_CDNS_40661953145278_0
timestamp 1669390400
transform 1 0 -66 0 1 12039
box 0 0 1 1
use M3_M2_CDNS_40661953145278  M3_M2_CDNS_40661953145278_1
timestamp 1669390400
transform 1 0 13530 0 1 12039
box 0 0 1 1
use comp018green_out_paddrv_6T_NMOS_GROUP  comp018green_out_paddrv_6T_NMOS_GROUP_0
timestamp 1669390400
transform 1 0 1609 0 1 31
box -1426 -398 11585 10917
use comp018green_out_paddrv_6T_PMOS_GROUP  comp018green_out_paddrv_6T_PMOS_GROUP_0
timestamp 1669390400
transform 1 0 548 0 1 12347
box -975 -1312 13355 15294
<< properties >>
string GDS_END 2695084
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2689506
string path 42.425 657.500 294.625 657.500 
<< end >>
