magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 1990 870
rect -86 352 678 377
rect 1051 352 1990 377
<< pwell >>
rect 678 352 1051 377
rect -86 -86 1990 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 572 93 692 165
rect 1037 68 1157 232
rect 1405 93 1525 165
rect 1660 93 1780 165
<< mvpmos >>
rect 124 560 224 684
rect 328 560 428 684
rect 532 560 632 684
rect 994 497 1094 716
rect 1425 592 1525 716
rect 1660 592 1760 716
<< mvndiff >>
rect 752 244 824 257
rect 752 198 765 244
rect 811 198 824 244
rect 752 165 824 198
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 572 165
rect 468 106 497 152
rect 543 106 572 152
rect 468 93 572 106
rect 692 93 824 165
rect 904 244 977 257
rect 904 198 917 244
rect 963 232 977 244
rect 963 198 1037 232
rect 904 68 1037 198
rect 1157 142 1245 232
rect 1157 96 1186 142
rect 1232 96 1245 142
rect 1157 68 1245 96
rect 1317 152 1405 165
rect 1317 106 1330 152
rect 1376 106 1405 152
rect 1317 93 1405 106
rect 1525 152 1660 165
rect 1525 106 1554 152
rect 1600 106 1660 152
rect 1525 93 1660 106
rect 1780 152 1868 165
rect 1780 106 1809 152
rect 1855 106 1868 152
rect 1780 93 1868 106
<< mvpdiff >>
rect 36 645 124 684
rect 36 599 49 645
rect 95 599 124 645
rect 36 560 124 599
rect 224 645 328 684
rect 224 599 253 645
rect 299 599 328 645
rect 224 560 328 599
rect 428 645 532 684
rect 428 599 457 645
rect 503 599 532 645
rect 428 560 532 599
rect 632 581 764 684
rect 632 560 705 581
rect 692 535 705 560
rect 751 535 764 581
rect 692 522 764 535
rect 906 567 994 716
rect 906 521 919 567
rect 965 521 994 567
rect 906 497 994 521
rect 1094 687 1182 716
rect 1094 641 1123 687
rect 1169 641 1182 687
rect 1094 497 1182 641
rect 1337 662 1425 716
rect 1337 616 1350 662
rect 1396 616 1425 662
rect 1337 592 1425 616
rect 1525 680 1660 716
rect 1525 634 1554 680
rect 1600 634 1660 680
rect 1525 592 1660 634
rect 1760 662 1848 716
rect 1760 616 1789 662
rect 1835 616 1848 662
rect 1760 592 1848 616
<< mvndiffc >>
rect 765 198 811 244
rect 49 106 95 152
rect 273 106 319 152
rect 497 106 543 152
rect 917 198 963 244
rect 1186 96 1232 142
rect 1330 106 1376 152
rect 1554 106 1600 152
rect 1809 106 1855 152
<< mvpdiffc >>
rect 49 599 95 645
rect 253 599 299 645
rect 457 599 503 645
rect 705 535 751 581
rect 919 521 965 567
rect 1123 641 1169 687
rect 1350 616 1396 662
rect 1554 634 1600 680
rect 1789 616 1835 662
<< polysilicon >>
rect 124 684 224 728
rect 328 684 428 728
rect 532 684 632 728
rect 994 716 1094 760
rect 1425 716 1525 760
rect 1660 716 1760 760
rect 124 412 224 560
rect 328 412 428 560
rect 532 527 632 560
rect 532 481 545 527
rect 591 481 632 527
rect 1425 557 1525 592
rect 532 468 632 481
rect 994 439 1094 497
rect 124 399 692 412
rect 124 353 137 399
rect 465 353 692 399
rect 994 393 1030 439
rect 1076 393 1094 439
rect 994 380 1094 393
rect 124 340 692 353
rect 124 165 244 340
rect 348 245 468 258
rect 348 199 385 245
rect 431 199 468 245
rect 348 165 468 199
rect 572 165 692 340
rect 1037 311 1157 324
rect 1037 265 1069 311
rect 1115 265 1157 311
rect 1425 287 1452 557
rect 1037 232 1157 265
rect 124 24 244 93
rect 348 24 468 93
rect 572 24 692 93
rect 1405 229 1452 287
rect 1498 229 1525 557
rect 1405 165 1525 229
rect 1660 463 1760 592
rect 1660 323 1688 463
rect 1734 323 1760 463
rect 1660 287 1760 323
rect 1660 165 1780 287
rect 1037 24 1157 68
rect 1405 49 1525 93
rect 1660 49 1780 93
<< polycontact >>
rect 545 481 591 527
rect 137 353 465 399
rect 1030 393 1076 439
rect 385 199 431 245
rect 1069 265 1115 311
rect 1452 229 1498 557
rect 1688 323 1734 463
<< metal1 >>
rect 0 724 1904 844
rect 49 645 95 678
rect 49 527 95 599
rect 253 645 299 724
rect 1123 687 1169 724
rect 253 573 299 599
rect 457 645 1077 678
rect 503 632 1077 645
rect 457 573 503 599
rect 648 581 764 582
rect 648 535 705 581
rect 751 535 764 581
rect 49 481 545 527
rect 591 481 602 527
rect 82 399 485 424
rect 82 353 137 399
rect 465 353 485 399
rect 82 340 485 353
rect 542 245 602 481
rect 36 199 385 245
rect 431 199 602 245
rect 648 522 764 535
rect 36 152 108 199
rect 648 152 694 522
rect 810 476 856 632
rect 754 430 856 476
rect 906 567 984 586
rect 906 521 919 567
rect 965 521 984 567
rect 754 244 822 430
rect 754 198 765 244
rect 811 198 822 244
rect 906 244 984 521
rect 1030 554 1077 632
rect 1554 680 1600 724
rect 1123 600 1169 641
rect 1350 662 1396 675
rect 1554 623 1600 634
rect 1789 662 1835 675
rect 1350 554 1396 616
rect 1789 577 1835 616
rect 1030 507 1396 554
rect 1452 557 1835 577
rect 1030 439 1076 507
rect 1030 380 1076 393
rect 906 198 917 244
rect 963 198 984 244
rect 1069 311 1115 324
rect 1115 265 1387 273
rect 1069 227 1387 265
rect 1069 152 1115 227
rect 36 106 49 152
rect 95 106 108 152
rect 262 106 273 152
rect 319 106 330 152
rect 480 106 497 152
rect 543 106 1115 152
rect 1186 142 1232 181
rect 262 60 330 106
rect 1317 152 1387 227
rect 1498 530 1835 557
rect 1548 463 1880 475
rect 1548 323 1688 463
rect 1734 323 1880 463
rect 1548 312 1880 323
rect 1498 229 1692 255
rect 1452 209 1692 229
rect 1317 106 1330 152
rect 1376 106 1387 152
rect 1554 152 1600 163
rect 1646 152 1692 209
rect 1646 106 1809 152
rect 1855 106 1868 152
rect 1186 60 1232 96
rect 1554 60 1600 106
rect 0 -60 1904 60
<< labels >>
flabel metal1 s 0 724 1904 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1186 163 1232 181 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 906 198 984 586 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 82 340 485 424 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1548 312 1880 475 0 FreeSans 400 0 0 0 I
port 2 nsew default input
rlabel metal1 s 1554 623 1600 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1123 623 1169 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 623 299 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1123 600 1169 623 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 600 299 623 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 573 299 600 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1554 152 1600 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1186 152 1232 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1554 60 1600 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1186 60 1232 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1904 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 784
string GDS_END 512146
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 506720
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
