magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 3334 870
rect -86 352 2159 377
rect 2379 352 3334 377
<< pwell >>
rect 2159 352 2379 377
rect -86 -86 3334 352
<< mvnmos >>
rect 157 93 277 165
rect 381 93 501 165
rect 605 93 725 165
rect 829 93 949 165
rect 1013 93 1133 165
rect 1385 93 1505 165
rect 1569 93 1689 165
rect 1829 68 1949 232
rect 2053 68 2173 232
rect 2365 68 2485 232
rect 2733 68 2853 232
rect 2957 68 3077 232
<< mvpmos >>
rect 177 534 277 606
rect 391 534 491 606
rect 631 494 731 606
rect 835 494 935 606
rect 1039 494 1139 606
rect 1391 497 1491 609
rect 1595 497 1695 609
rect 1843 497 1943 716
rect 2053 497 2153 716
rect 2267 497 2367 716
rect 2733 472 2833 716
rect 2957 472 3057 716
<< mvndiff >>
rect 2233 244 2305 257
rect 2233 232 2246 244
rect 1749 165 1829 232
rect 69 152 157 165
rect 69 106 82 152
rect 128 106 157 152
rect 69 93 157 106
rect 277 152 381 165
rect 277 106 306 152
rect 352 106 381 152
rect 277 93 381 106
rect 501 152 605 165
rect 501 106 530 152
rect 576 106 605 152
rect 501 93 605 106
rect 725 152 829 165
rect 725 106 754 152
rect 800 106 829 152
rect 725 93 829 106
rect 949 93 1013 165
rect 1133 152 1221 165
rect 1133 106 1162 152
rect 1208 106 1221 152
rect 1133 93 1221 106
rect 1297 152 1385 165
rect 1297 106 1310 152
rect 1356 106 1385 152
rect 1297 93 1385 106
rect 1505 93 1569 165
rect 1689 152 1829 165
rect 1689 106 1718 152
rect 1764 106 1829 152
rect 1689 93 1829 106
rect 1749 68 1829 93
rect 1949 152 2053 232
rect 1949 106 1978 152
rect 2024 106 2053 152
rect 1949 68 2053 106
rect 2173 198 2246 232
rect 2292 232 2305 244
rect 2292 198 2365 232
rect 2173 68 2365 198
rect 2485 152 2573 232
rect 2485 106 2514 152
rect 2560 106 2573 152
rect 2485 68 2573 106
rect 2645 204 2733 232
rect 2645 158 2658 204
rect 2704 158 2733 204
rect 2645 68 2733 158
rect 2853 142 2957 232
rect 2853 96 2882 142
rect 2928 96 2957 142
rect 2853 68 2957 96
rect 3077 204 3165 232
rect 3077 158 3106 204
rect 3152 158 3165 204
rect 3077 68 3165 158
<< mvpdiff >>
rect 1755 701 1843 716
rect 1755 609 1768 701
rect 89 593 177 606
rect 89 547 102 593
rect 148 547 177 593
rect 89 534 177 547
rect 277 534 391 606
rect 491 593 631 606
rect 491 547 556 593
rect 602 547 631 593
rect 491 534 631 547
rect 551 494 631 534
rect 731 593 835 606
rect 731 547 760 593
rect 806 547 835 593
rect 731 494 835 547
rect 935 567 1039 606
rect 935 521 964 567
rect 1010 521 1039 567
rect 935 494 1039 521
rect 1139 593 1227 606
rect 1139 547 1168 593
rect 1214 547 1227 593
rect 1139 494 1227 547
rect 1303 593 1391 609
rect 1303 547 1316 593
rect 1362 547 1391 593
rect 1303 497 1391 547
rect 1491 556 1595 609
rect 1491 510 1520 556
rect 1566 510 1595 556
rect 1491 497 1595 510
rect 1695 561 1768 609
rect 1814 561 1843 701
rect 1695 497 1843 561
rect 1943 610 2053 716
rect 1943 564 1972 610
rect 2018 564 2053 610
rect 1943 497 2053 564
rect 2153 497 2267 716
rect 2367 703 2471 716
rect 2367 657 2411 703
rect 2457 657 2471 703
rect 2367 497 2471 657
rect 2645 653 2733 716
rect 2645 513 2658 653
rect 2704 513 2733 653
rect 2645 472 2733 513
rect 2833 689 2957 716
rect 2833 643 2862 689
rect 2908 643 2957 689
rect 2833 472 2957 643
rect 3057 653 3145 716
rect 3057 513 3086 653
rect 3132 513 3145 653
rect 3057 472 3145 513
<< mvndiffc >>
rect 82 106 128 152
rect 306 106 352 152
rect 530 106 576 152
rect 754 106 800 152
rect 1162 106 1208 152
rect 1310 106 1356 152
rect 1718 106 1764 152
rect 1978 106 2024 152
rect 2246 198 2292 244
rect 2514 106 2560 152
rect 2658 158 2704 204
rect 2882 96 2928 142
rect 3106 158 3152 204
<< mvpdiffc >>
rect 102 547 148 593
rect 556 547 602 593
rect 760 547 806 593
rect 964 521 1010 567
rect 1168 547 1214 593
rect 1316 547 1362 593
rect 1520 510 1566 556
rect 1768 561 1814 701
rect 1972 564 2018 610
rect 2411 657 2457 703
rect 2658 513 2704 653
rect 2862 643 2908 689
rect 3086 513 3132 653
<< polysilicon >>
rect 1843 716 1943 760
rect 2053 716 2153 760
rect 2267 716 2367 760
rect 2733 716 2833 760
rect 2957 716 3057 760
rect 177 606 277 651
rect 391 606 491 651
rect 631 606 731 651
rect 835 606 935 651
rect 1039 606 1139 651
rect 1391 609 1491 653
rect 1595 609 1695 653
rect 177 472 277 534
rect 177 332 215 472
rect 261 332 277 472
rect 177 209 277 332
rect 391 303 491 534
rect 391 257 429 303
rect 475 257 491 303
rect 391 209 491 257
rect 631 399 731 494
rect 631 353 650 399
rect 696 353 731 399
rect 631 225 731 353
rect 835 303 935 494
rect 835 257 849 303
rect 895 257 935 303
rect 631 209 725 225
rect 835 209 935 257
rect 1039 344 1139 494
rect 1391 362 1491 497
rect 1039 298 1068 344
rect 1114 298 1139 344
rect 1039 225 1139 298
rect 1385 347 1491 362
rect 1385 301 1405 347
rect 1451 301 1491 347
rect 1039 209 1133 225
rect 157 165 277 209
rect 381 165 501 209
rect 605 165 725 209
rect 829 165 949 209
rect 1013 165 1133 209
rect 1385 209 1491 301
rect 1595 415 1695 497
rect 1595 369 1634 415
rect 1680 369 1695 415
rect 1595 354 1695 369
rect 1595 209 1689 354
rect 1843 311 1943 497
rect 1843 276 1865 311
rect 1829 265 1865 276
rect 1911 276 1943 311
rect 2053 415 2153 497
rect 2053 369 2080 415
rect 2126 369 2153 415
rect 2053 276 2153 369
rect 2267 395 2367 497
rect 2733 415 2833 472
rect 2267 380 2485 395
rect 2267 334 2294 380
rect 2340 334 2485 380
rect 2267 319 2485 334
rect 1911 265 1949 276
rect 1829 232 1949 265
rect 2053 232 2173 276
rect 1385 165 1505 209
rect 1569 165 1689 209
rect 157 49 277 93
rect 381 49 501 93
rect 605 49 725 93
rect 829 49 949 93
rect 1013 49 1133 93
rect 1385 49 1505 93
rect 1569 49 1689 93
rect 2365 232 2485 319
rect 2733 369 2754 415
rect 2800 369 2833 415
rect 2733 357 2833 369
rect 2957 415 3057 472
rect 2957 369 2978 415
rect 3024 369 3057 415
rect 2957 357 3057 369
rect 2733 311 3057 357
rect 2733 232 2853 311
rect 2957 288 3057 311
rect 2957 232 3077 288
rect 1829 24 1949 68
rect 2053 24 2173 68
rect 2365 24 2485 68
rect 2733 24 2853 68
rect 2957 24 3077 68
<< polycontact >>
rect 215 332 261 472
rect 429 257 475 303
rect 650 353 696 399
rect 849 257 895 303
rect 1068 298 1114 344
rect 1405 301 1451 347
rect 1634 369 1680 415
rect 1865 265 1911 311
rect 2080 369 2126 415
rect 2294 334 2340 380
rect 2754 369 2800 415
rect 2978 369 3024 415
<< metal1 >>
rect 0 724 3248 844
rect 102 593 148 606
rect 545 593 613 724
rect 545 547 556 593
rect 602 547 613 593
rect 747 632 1214 678
rect 747 593 819 632
rect 747 547 760 593
rect 806 547 819 593
rect 1157 593 1214 632
rect 102 244 148 547
rect 215 491 455 532
rect 944 521 964 567
rect 1010 521 1111 567
rect 1157 547 1168 593
rect 1157 536 1214 547
rect 1305 593 1362 724
rect 1755 701 1827 724
rect 1305 547 1316 593
rect 1305 536 1362 547
rect 1408 602 1689 648
rect 215 472 813 491
rect 261 445 813 472
rect 767 419 813 445
rect 1065 444 1111 521
rect 1408 444 1454 602
rect 215 298 261 332
rect 307 353 650 399
rect 696 353 712 399
rect 767 353 1019 419
rect 1065 398 1454 444
rect 307 244 363 353
rect 960 344 1019 353
rect 1402 347 1454 398
rect 410 303 907 307
rect 410 257 429 303
rect 475 257 849 303
rect 895 257 907 303
rect 960 298 1068 344
rect 1114 298 1139 344
rect 960 297 1139 298
rect 1402 301 1405 347
rect 1451 301 1454 347
rect 410 253 907 257
rect 1402 244 1454 301
rect 102 198 363 244
rect 295 152 363 198
rect 1048 198 1454 244
rect 1509 510 1520 556
rect 1566 510 1577 556
rect 1509 244 1577 510
rect 1632 513 1689 602
rect 1755 561 1768 701
rect 1814 561 1827 701
rect 2398 703 2471 724
rect 2398 657 2411 703
rect 2457 657 2471 703
rect 2862 689 2908 724
rect 2398 656 2471 657
rect 2658 653 2704 672
rect 1950 564 1972 610
rect 2018 564 2471 610
rect 1950 563 2471 564
rect 1755 559 1827 561
rect 1632 466 2267 513
rect 1623 415 2142 419
rect 1623 369 1634 415
rect 1680 369 2080 415
rect 2126 369 2142 415
rect 1623 365 2142 369
rect 2221 380 2267 466
rect 2425 419 2471 563
rect 2862 603 2908 643
rect 3048 653 3152 672
rect 3048 536 3086 653
rect 2704 513 3086 536
rect 3132 513 3152 653
rect 2658 472 3152 513
rect 2425 415 3042 419
rect 2221 334 2294 380
rect 2340 334 2352 380
rect 2425 369 2754 415
rect 2800 369 2978 415
rect 3024 369 3042 415
rect 2425 365 3042 369
rect 1854 265 1865 311
rect 1911 265 1922 311
rect 1854 244 1922 265
rect 2425 244 2471 365
rect 3092 312 3152 472
rect 1509 198 1922 244
rect 2234 198 2246 244
rect 2292 198 2471 244
rect 2658 248 3152 312
rect 2658 204 2704 248
rect 71 106 82 152
rect 128 106 139 152
rect 295 106 306 152
rect 352 106 363 152
rect 519 152 587 155
rect 1048 152 1094 198
rect 1509 152 1577 198
rect 3106 204 3152 248
rect 519 106 530 152
rect 576 106 587 152
rect 725 106 754 152
rect 800 106 1094 152
rect 1151 106 1162 152
rect 1208 106 1219 152
rect 1297 106 1310 152
rect 1356 106 1577 152
rect 1707 106 1718 152
rect 1764 106 1776 152
rect 1959 106 1978 152
rect 2024 106 2514 152
rect 2560 106 2573 152
rect 2658 131 2704 158
rect 2882 142 2928 181
rect 71 60 139 106
rect 519 60 587 106
rect 1151 60 1219 106
rect 1707 60 1776 106
rect 3106 131 3152 158
rect 2882 60 2928 96
rect 0 -60 3248 60
<< labels >>
flabel metal1 s 1623 365 2142 419 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 3248 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2882 155 2928 181 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 3048 536 3152 672 0 FreeSans 400 0 0 0 Z
port 4 nsew default output
flabel metal1 s 410 253 907 307 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 215 491 455 532 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
rlabel metal1 s 215 445 813 491 1 A2
port 2 nsew default input
rlabel metal1 s 767 419 813 445 1 A2
port 2 nsew default input
rlabel metal1 s 215 419 261 445 1 A2
port 2 nsew default input
rlabel metal1 s 767 353 1019 419 1 A2
port 2 nsew default input
rlabel metal1 s 215 353 261 419 1 A2
port 2 nsew default input
rlabel metal1 s 960 344 1019 353 1 A2
port 2 nsew default input
rlabel metal1 s 215 344 261 353 1 A2
port 2 nsew default input
rlabel metal1 s 960 298 1139 344 1 A2
port 2 nsew default input
rlabel metal1 s 215 298 261 344 1 A2
port 2 nsew default input
rlabel metal1 s 960 297 1139 298 1 A2
port 2 nsew default input
rlabel metal1 s 2658 536 2704 672 1 Z
port 4 nsew default output
rlabel metal1 s 2658 472 3152 536 1 Z
port 4 nsew default output
rlabel metal1 s 3092 312 3152 472 1 Z
port 4 nsew default output
rlabel metal1 s 2658 248 3152 312 1 Z
port 4 nsew default output
rlabel metal1 s 3106 131 3152 248 1 Z
port 4 nsew default output
rlabel metal1 s 2658 131 2704 248 1 Z
port 4 nsew default output
rlabel metal1 s 2862 656 2908 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2398 656 2471 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1755 656 1827 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1305 656 1362 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 545 656 613 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2862 603 2908 656 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1755 603 1827 656 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1305 603 1362 656 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 545 603 613 656 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1755 559 1827 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1305 559 1362 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 545 559 613 603 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1305 547 1362 559 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 545 547 613 559 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1305 536 1362 547 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2882 152 2928 155 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 519 152 587 155 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2882 60 2928 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1707 60 1776 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1151 60 1219 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 519 60 587 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 71 60 139 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3248 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3248 784
string GDS_END 377010
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 369794
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
