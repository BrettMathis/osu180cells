magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4230 1094
<< pwell >>
rect -86 -86 4230 453
<< mvnmos >>
rect 128 175 248 333
rect 352 175 472 333
rect 732 215 852 333
rect 956 215 1076 333
rect 1180 215 1300 333
rect 1348 215 1468 333
rect 1568 215 1688 333
rect 1792 215 1912 333
rect 1960 215 2080 333
rect 2184 215 2304 333
rect 2408 215 2528 333
rect 2955 175 3075 333
rect 3123 175 3243 333
rect 3347 175 3467 333
rect 3515 175 3635 333
rect 3900 69 4020 333
<< mvpmos >>
rect 124 586 224 862
rect 328 586 428 862
rect 676 582 776 782
rect 880 582 980 782
rect 1084 582 1184 782
rect 1288 582 1388 782
rect 1568 690 1668 890
rect 1916 690 2016 890
rect 2196 573 2296 773
rect 2400 573 2500 773
rect 2604 573 2704 773
rect 2952 584 3052 860
rect 3156 584 3256 860
rect 3360 584 3460 860
rect 3564 584 3664 860
rect 3912 573 4012 939
<< mvndiff >>
rect 40 320 128 333
rect 40 274 53 320
rect 99 274 128 320
rect 40 175 128 274
rect 248 234 352 333
rect 248 188 277 234
rect 323 188 352 234
rect 248 175 352 188
rect 472 320 560 333
rect 472 274 501 320
rect 547 274 560 320
rect 472 175 560 274
rect 644 274 732 333
rect 644 228 657 274
rect 703 228 732 274
rect 644 215 732 228
rect 852 320 956 333
rect 852 274 881 320
rect 927 274 956 320
rect 852 215 956 274
rect 1076 320 1180 333
rect 1076 274 1105 320
rect 1151 274 1180 320
rect 1076 215 1180 274
rect 1300 215 1348 333
rect 1468 215 1568 333
rect 1688 274 1792 333
rect 1688 228 1717 274
rect 1763 228 1792 274
rect 1688 215 1792 228
rect 1912 215 1960 333
rect 2080 320 2184 333
rect 2080 274 2109 320
rect 2155 274 2184 320
rect 2080 215 2184 274
rect 2304 320 2408 333
rect 2304 274 2333 320
rect 2379 274 2408 320
rect 2304 215 2408 274
rect 2528 320 2616 333
rect 2528 274 2557 320
rect 2603 274 2616 320
rect 2528 215 2616 274
rect 2867 320 2955 333
rect 2867 274 2880 320
rect 2926 274 2955 320
rect 2867 175 2955 274
rect 3075 175 3123 333
rect 3243 234 3347 333
rect 3243 188 3272 234
rect 3318 188 3347 234
rect 3243 175 3347 188
rect 3467 175 3515 333
rect 3635 320 3723 333
rect 3635 274 3664 320
rect 3710 274 3723 320
rect 3635 175 3723 274
rect 3812 320 3900 333
rect 3812 180 3825 320
rect 3871 180 3900 320
rect 3812 69 3900 180
rect 4020 222 4108 333
rect 4020 82 4049 222
rect 4095 82 4108 222
rect 4020 69 4108 82
<< mvpdiff >>
rect 36 735 124 862
rect 36 689 49 735
rect 95 689 124 735
rect 36 586 124 689
rect 224 849 328 862
rect 224 803 253 849
rect 299 803 328 849
rect 224 586 328 803
rect 428 739 516 862
rect 1436 955 1508 968
rect 1436 909 1449 955
rect 1495 909 1508 955
rect 2076 955 2148 968
rect 1436 896 1508 909
rect 1448 890 1508 896
rect 2076 909 2089 955
rect 2135 909 2148 955
rect 2076 896 2148 909
rect 2076 890 2136 896
rect 1448 782 1568 890
rect 428 599 457 739
rect 503 599 516 739
rect 428 586 516 599
rect 588 769 676 782
rect 588 723 601 769
rect 647 723 676 769
rect 588 582 676 723
rect 776 735 880 782
rect 776 595 805 735
rect 851 595 880 735
rect 776 582 880 595
rect 980 735 1084 782
rect 980 595 1009 735
rect 1055 595 1084 735
rect 980 582 1084 595
rect 1184 727 1288 782
rect 1184 681 1213 727
rect 1259 681 1288 727
rect 1184 582 1288 681
rect 1388 690 1568 782
rect 1668 749 1756 890
rect 1668 703 1697 749
rect 1743 703 1756 749
rect 1668 690 1756 703
rect 1828 749 1916 890
rect 1828 703 1841 749
rect 1887 703 1916 749
rect 1828 690 1916 703
rect 2016 773 2136 890
rect 2864 847 2952 860
rect 2864 801 2877 847
rect 2923 801 2952 847
rect 2016 690 2196 773
rect 1388 582 1468 690
rect 2116 573 2196 690
rect 2296 726 2400 773
rect 2296 586 2325 726
rect 2371 586 2400 726
rect 2296 573 2400 586
rect 2500 744 2604 773
rect 2500 604 2529 744
rect 2575 604 2604 744
rect 2500 573 2604 604
rect 2704 632 2792 773
rect 2704 586 2733 632
rect 2779 586 2792 632
rect 2704 573 2792 586
rect 2864 584 2952 801
rect 3052 643 3156 860
rect 3052 597 3081 643
rect 3127 597 3156 643
rect 3052 584 3156 597
rect 3256 847 3360 860
rect 3256 801 3285 847
rect 3331 801 3360 847
rect 3256 584 3360 801
rect 3460 643 3564 860
rect 3460 597 3489 643
rect 3535 597 3564 643
rect 3460 584 3564 597
rect 3664 847 3752 860
rect 3664 707 3693 847
rect 3739 707 3752 847
rect 3664 584 3752 707
rect 3824 726 3912 939
rect 3824 586 3837 726
rect 3883 586 3912 726
rect 3824 573 3912 586
rect 4012 926 4100 939
rect 4012 786 4041 926
rect 4087 786 4100 926
rect 4012 573 4100 786
<< mvndiffc >>
rect 53 274 99 320
rect 277 188 323 234
rect 501 274 547 320
rect 657 228 703 274
rect 881 274 927 320
rect 1105 274 1151 320
rect 1717 228 1763 274
rect 2109 274 2155 320
rect 2333 274 2379 320
rect 2557 274 2603 320
rect 2880 274 2926 320
rect 3272 188 3318 234
rect 3664 274 3710 320
rect 3825 180 3871 320
rect 4049 82 4095 222
<< mvpdiffc >>
rect 49 689 95 735
rect 253 803 299 849
rect 1449 909 1495 955
rect 2089 909 2135 955
rect 457 599 503 739
rect 601 723 647 769
rect 805 595 851 735
rect 1009 595 1055 735
rect 1213 681 1259 727
rect 1697 703 1743 749
rect 1841 703 1887 749
rect 2877 801 2923 847
rect 2325 586 2371 726
rect 2529 604 2575 744
rect 2733 586 2779 632
rect 3081 597 3127 643
rect 3285 801 3331 847
rect 3489 597 3535 643
rect 3693 707 3739 847
rect 3837 586 3883 726
rect 4041 786 4087 926
<< polysilicon >>
rect 328 922 1184 962
rect 124 862 224 906
rect 328 862 428 922
rect 880 861 980 874
rect 676 782 776 826
rect 880 815 921 861
rect 967 815 980 861
rect 880 782 980 815
rect 1084 861 1184 922
rect 1084 815 1125 861
rect 1171 815 1184 861
rect 1568 890 1668 934
rect 1916 890 2016 934
rect 2208 920 3052 960
rect 3912 939 4012 983
rect 1084 782 1184 815
rect 1288 782 1388 826
rect 124 553 224 586
rect 124 542 142 553
rect 128 507 142 542
rect 188 507 224 553
rect 328 542 428 586
rect 2208 847 2296 920
rect 2196 773 2296 847
rect 2400 852 2500 865
rect 2952 860 3052 920
rect 3156 860 3256 904
rect 3360 860 3460 904
rect 3564 860 3664 904
rect 2400 806 2441 852
rect 2487 806 2500 852
rect 2400 773 2500 806
rect 2604 773 2704 817
rect 128 377 224 507
rect 352 412 428 542
rect 676 538 776 582
rect 880 538 980 582
rect 1084 538 1184 582
rect 1288 538 1388 582
rect 128 333 248 377
rect 352 366 365 412
rect 411 377 428 412
rect 732 522 776 538
rect 732 509 804 522
rect 732 463 745 509
rect 791 463 804 509
rect 732 377 804 463
rect 940 465 980 538
rect 1348 493 1388 538
rect 1348 480 1468 493
rect 940 425 1300 465
rect 1180 412 1300 425
rect 411 366 472 377
rect 352 333 472 366
rect 732 333 852 377
rect 956 333 1076 377
rect 1180 366 1197 412
rect 1243 366 1300 412
rect 1180 333 1300 366
rect 1348 434 1361 480
rect 1407 434 1468 480
rect 1348 333 1468 434
rect 1568 377 1668 690
rect 1916 585 2016 690
rect 1792 572 2016 585
rect 1792 526 1853 572
rect 1899 545 2016 572
rect 1899 526 1912 545
rect 1568 333 1688 377
rect 1792 333 1912 526
rect 2196 465 2296 573
rect 2400 529 2500 573
rect 1960 425 2296 465
rect 1960 333 2080 425
rect 2408 377 2500 529
rect 2604 457 2704 573
rect 2952 551 3052 584
rect 2952 505 2965 551
rect 3011 505 3052 551
rect 2952 497 3052 505
rect 2604 444 2718 457
rect 2604 398 2659 444
rect 2705 398 2718 444
rect 2604 393 2718 398
rect 2646 385 2718 393
rect 2955 377 3052 497
rect 3156 540 3256 584
rect 3360 551 3460 584
rect 3156 412 3243 540
rect 3156 377 3184 412
rect 2184 333 2304 377
rect 2408 333 2528 377
rect 2955 333 3075 377
rect 3123 366 3184 377
rect 3230 366 3243 412
rect 3360 505 3390 551
rect 3436 505 3460 551
rect 3360 377 3460 505
rect 3564 551 3664 584
rect 3564 505 3581 551
rect 3627 505 3664 551
rect 3564 492 3664 505
rect 3564 377 3634 492
rect 3912 465 4012 573
rect 3720 452 4012 465
rect 3720 406 3733 452
rect 3779 406 4012 452
rect 3720 393 4012 406
rect 3900 377 4012 393
rect 3123 333 3243 366
rect 3347 333 3467 377
rect 3515 333 3635 377
rect 3900 333 4020 377
rect 128 131 248 175
rect 352 115 472 175
rect 732 171 852 215
rect 956 115 1076 215
rect 1180 171 1300 215
rect 1348 171 1468 215
rect 352 75 1076 115
rect 1568 75 1688 215
rect 1792 171 1912 215
rect 1960 171 2080 215
rect 2184 182 2304 215
rect 2184 136 2197 182
rect 2243 136 2304 182
rect 2408 171 2528 215
rect 2184 123 2304 136
rect 2955 131 3075 175
rect 3123 131 3243 175
rect 3347 75 3467 175
rect 3515 131 3635 175
rect 1568 35 3467 75
rect 3900 25 4020 69
<< polycontact >>
rect 921 815 967 861
rect 1125 815 1171 861
rect 142 507 188 553
rect 2441 806 2487 852
rect 365 366 411 412
rect 745 463 791 509
rect 1197 366 1243 412
rect 1361 434 1407 480
rect 1853 526 1899 572
rect 2965 505 3011 551
rect 2659 398 2705 444
rect 3184 366 3230 412
rect 3390 505 3436 551
rect 3581 505 3627 551
rect 3733 406 3779 452
rect 2197 136 2243 182
<< metal1 >>
rect 0 955 4144 1098
rect 0 918 1449 955
rect 253 849 299 918
rect 253 792 299 803
rect 601 769 647 918
rect 1495 918 2089 955
rect 1449 898 1495 909
rect 2135 926 4144 955
rect 2135 918 4041 926
rect 2089 898 2135 909
rect 49 735 411 746
rect 95 700 411 735
rect 49 678 95 689
rect 142 553 316 654
rect 188 507 316 553
rect 142 496 316 507
rect 365 412 411 700
rect 365 348 411 366
rect 53 320 411 348
rect 99 302 411 320
rect 457 739 503 750
rect 601 712 647 723
rect 693 861 967 872
rect 693 815 921 861
rect 693 804 967 815
rect 1114 815 1125 861
rect 1171 852 1182 861
rect 1171 815 2441 852
rect 1114 806 2441 815
rect 2487 806 2498 852
rect 2866 847 2934 918
rect 693 666 739 804
rect 2866 801 2877 847
rect 2923 801 2934 847
rect 3274 847 3342 918
rect 3274 801 3285 847
rect 3331 801 3342 847
rect 3693 847 3739 918
rect 1213 749 1743 760
rect 503 620 739 666
rect 805 735 851 746
rect 503 599 547 620
rect 457 320 547 599
rect 1009 735 1055 746
rect 851 595 927 601
rect 805 555 927 595
rect 593 509 754 542
rect 593 463 745 509
rect 791 463 802 509
rect 53 263 99 274
rect 457 274 501 320
rect 881 320 927 555
rect 1213 727 1697 749
rect 1259 703 1697 727
rect 1259 681 1743 703
rect 1841 749 2371 760
rect 1887 726 2371 749
rect 1887 714 2325 726
rect 1887 703 1991 714
rect 1841 692 1991 703
rect 1213 670 1743 681
rect 1009 583 1055 595
rect 1009 572 1899 583
rect 1009 537 1853 572
rect 457 263 547 274
rect 657 274 703 285
rect 277 234 323 245
rect 277 90 323 188
rect 881 263 927 274
rect 1105 320 1151 537
rect 1853 515 1899 526
rect 1361 480 1407 491
rect 1945 469 1991 692
rect 2529 744 3627 755
rect 2325 575 2371 586
rect 2417 604 2529 639
rect 2575 709 3627 744
rect 2417 593 2575 604
rect 2733 632 2779 643
rect 2417 529 2463 593
rect 2733 547 2779 586
rect 2942 578 3011 654
rect 2965 551 3011 578
rect 2333 483 2463 529
rect 2557 501 2899 547
rect 1407 434 2155 469
rect 1361 423 2155 434
rect 1197 412 1243 423
rect 1243 366 2063 377
rect 1197 331 2063 366
rect 1105 263 1151 274
rect 1717 274 1763 285
rect 657 90 703 228
rect 1717 90 1763 228
rect 2017 182 2063 331
rect 2109 320 2155 423
rect 2109 263 2155 274
rect 2333 320 2379 483
rect 2333 263 2379 274
rect 2557 320 2603 501
rect 2557 263 2603 274
rect 2659 444 2705 455
rect 2659 182 2705 398
rect 2853 448 2899 501
rect 2965 494 3011 505
rect 3081 643 3127 654
rect 3081 448 3127 597
rect 3489 643 3535 654
rect 3260 551 3442 578
rect 3260 505 3390 551
rect 3436 505 3442 551
rect 3260 466 3442 505
rect 2853 402 3127 448
rect 3489 412 3535 597
rect 3581 551 3627 709
rect 4087 918 4144 926
rect 4041 775 4087 786
rect 3693 696 3739 707
rect 3825 726 3890 737
rect 3581 494 3627 505
rect 3825 586 3837 726
rect 3883 586 3890 726
rect 3664 452 3779 463
rect 3664 412 3733 452
rect 2853 320 2926 402
rect 3173 366 3184 412
rect 3230 406 3733 412
rect 3230 395 3779 406
rect 3230 366 3710 395
rect 2853 274 2880 320
rect 2853 263 2926 274
rect 3664 320 3710 366
rect 3664 263 3710 274
rect 3825 320 3890 586
rect 2017 136 2197 182
rect 2243 136 2705 182
rect 3272 234 3318 245
rect 3272 90 3318 188
rect 3871 180 3890 320
rect 3825 169 3890 180
rect 4049 222 4095 233
rect 0 82 4049 90
rect 4095 82 4144 90
rect 0 -90 4144 82
<< labels >>
flabel metal1 s 142 496 316 654 0 FreeSans 200 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 593 509 754 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3825 169 3890 737 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3260 466 3442 578 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 2942 578 3011 654 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 4144 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1717 245 1763 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 593 463 802 509 1 D
port 1 nsew default input
rlabel metal1 s 2965 494 3011 578 1 SETN
port 3 nsew default input
rlabel metal1 s 4041 898 4087 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 898 3739 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3274 898 3342 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2866 898 2934 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2089 898 2135 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1449 898 1495 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 898 647 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 898 299 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4041 801 4087 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 801 3739 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3274 801 3342 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2866 801 2934 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 801 647 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 801 299 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4041 792 4087 801 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 792 3739 801 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 792 647 801 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 792 299 801 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4041 775 4087 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 775 3739 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 775 647 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 712 3739 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 712 647 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3693 696 3739 712 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 657 245 703 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3272 233 3318 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1717 233 1763 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 657 233 703 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 277 233 323 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4049 90 4095 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3272 90 3318 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1717 90 1763 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 657 90 703 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 277 90 323 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4144 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4144 1008
string GDS_END 630974
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 621210
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
