magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 498
<< mvpmos >>
rect 0 0 120 378
<< mvpdiff >>
rect -88 365 0 378
rect -88 13 -75 365
rect -29 13 0 365
rect -88 0 0 13
rect 120 365 208 378
rect 120 13 149 365
rect 195 13 208 365
rect 120 0 208 13
<< mvpdiffc >>
rect -75 13 -29 365
rect 149 13 195 365
<< polysilicon >>
rect 0 378 120 422
rect 0 -44 120 0
<< metal1 >>
rect -75 365 -29 378
rect -75 0 -29 13
rect 149 365 195 378
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 189 -52 189 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 189 172 189 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 801958
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 800486
<< end >>
