magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 111 181 123
rect 28 70 33 111
rect 45 65 50 104
rect 62 70 67 111
rect 79 65 84 104
rect 96 70 101 111
rect 113 65 118 104
rect 130 70 135 111
rect 147 76 152 104
rect 145 70 155 76
rect 164 70 169 111
rect 147 65 152 70
rect 45 59 152 65
rect 21 44 31 50
rect 45 47 50 59
rect 79 47 84 59
rect 113 47 118 59
rect 147 47 152 59
rect 45 41 152 47
rect 28 12 33 36
rect 45 19 50 41
rect 62 12 67 36
rect 79 19 84 41
rect 96 12 101 36
rect 113 19 118 41
rect 130 12 135 36
rect 147 19 152 41
rect 164 12 169 36
rect 0 0 181 12
<< obsm1 >>
rect 11 65 16 104
rect 11 59 40 65
rect 11 19 16 59
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 145 69 155 77
rect 22 50 30 51
rect 21 44 31 50
rect 22 43 30 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
<< labels >>
rlabel metal2 s 22 43 30 51 6 A
port 1 nsew signal input
rlabel metal2 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal1 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 28 70 33 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 62 70 67 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 96 70 101 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 130 70 135 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 164 70 169 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 181 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 62 0 67 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 96 0 101 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 130 0 135 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 164 0 169 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 181 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 145 69 155 77 6 Y
port 2 nsew signal output
rlabel metal1 s 45 19 50 104 6 Y
port 2 nsew signal output
rlabel metal1 s 79 19 84 104 6 Y
port 2 nsew signal output
rlabel metal1 s 113 19 118 104 6 Y
port 2 nsew signal output
rlabel metal1 s 45 41 152 47 6 Y
port 2 nsew signal output
rlabel metal1 s 45 59 152 65 6 Y
port 2 nsew signal output
rlabel metal1 s 147 19 152 104 6 Y
port 2 nsew signal output
rlabel metal1 s 145 70 155 76 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 181 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 147790
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 133870
<< end >>
