magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 960 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 530 700 590 1040
rect 700 700 760 1040
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 860 360
rect 760 252 792 298
rect 838 252 860 298
rect 760 190 860 252
<< pdiff >>
rect 90 987 190 1040
rect 90 753 112 987
rect 158 753 190 987
rect 90 700 190 753
rect 250 987 360 1040
rect 250 753 282 987
rect 328 753 360 987
rect 250 700 360 753
rect 420 987 530 1040
rect 420 753 452 987
rect 498 753 530 987
rect 420 700 530 753
rect 590 987 700 1040
rect 590 753 622 987
rect 668 753 700 987
rect 590 700 700 753
rect 760 987 870 1040
rect 760 753 802 987
rect 848 753 870 987
rect 760 700 870 753
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
<< pdiffc >>
rect 112 753 158 987
rect 282 753 328 987
rect 452 753 498 987
rect 622 753 668 987
rect 802 753 848 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 190 650 250 700
rect 360 650 420 700
rect 530 650 590 700
rect 700 650 760 700
rect 190 600 760 650
rect 190 520 250 600
rect 90 498 250 520
rect 90 452 112 498
rect 158 460 250 498
rect 158 452 760 460
rect 90 430 760 452
rect 190 400 760 430
rect 190 360 250 400
rect 360 360 420 400
rect 530 360 590 400
rect 700 360 760 400
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
<< polycontact >>
rect 112 452 158 498
<< metal1 >>
rect 0 1178 960 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 960 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 960 1176
rect 0 1110 960 1124
rect 110 987 160 1110
rect 110 753 112 987
rect 158 753 160 987
rect 110 700 160 753
rect 280 987 330 1040
rect 280 753 282 987
rect 328 753 330 987
rect 280 650 330 753
rect 450 987 500 1110
rect 450 753 452 987
rect 498 753 500 987
rect 450 700 500 753
rect 620 987 670 1040
rect 620 753 622 987
rect 668 760 670 987
rect 800 987 850 1110
rect 668 756 750 760
rect 668 753 674 756
rect 620 704 674 753
rect 726 704 750 756
rect 620 700 750 704
rect 800 753 802 987
rect 848 753 850 987
rect 800 700 850 753
rect 620 650 670 700
rect 280 600 670 650
rect 80 498 180 500
rect 80 496 112 498
rect 80 444 104 496
rect 158 452 180 498
rect 156 444 180 452
rect 80 440 180 444
rect 280 460 330 600
rect 620 460 670 600
rect 280 410 670 460
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 410
rect 280 252 282 298
rect 328 252 330 298
rect 280 190 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 410
rect 620 252 622 298
rect 668 252 670 298
rect 620 190 670 252
rect 790 298 840 360
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 0 106 960 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 960 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 960 54
rect 0 0 960 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 674 704 726 756
rect 104 452 112 496
rect 112 452 156 496
rect 104 444 156 452
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 660 760 740 770
rect 650 756 750 760
rect 650 704 674 756
rect 726 704 750 756
rect 650 700 750 704
rect 660 690 740 700
rect 80 496 180 510
rect 80 444 104 496
rect 156 444 180 496
rect 80 430 180 444
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 80 430 180 510 4 A
port 1 nsew signal input
rlabel metal2 s 660 690 740 770 4 Y
port 2 nsew signal output
rlabel metal1 s 80 440 180 500 1 A
port 1 nsew signal input
rlabel metal2 s 90 1120 190 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 700 160 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 700 500 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 800 700 850 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1110 960 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 0 160 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 0 500 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 0 840 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 960 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 650 700 750 760 1 Y
port 2 nsew signal output
rlabel metal1 s 280 190 330 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 280 410 670 460 1 Y
port 2 nsew signal output
rlabel metal1 s 280 600 670 650 1 Y
port 2 nsew signal output
rlabel metal1 s 620 190 670 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 620 700 750 760 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 960 1230
string GDS_END 369802
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 362410
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
