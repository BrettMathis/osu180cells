magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 4902 870
rect -86 352 2765 377
rect 4596 352 4902 377
<< pwell >>
rect -86 -86 4902 352
<< mvnmos >>
rect 165 68 285 232
rect 389 68 509 232
rect 613 68 733 232
rect 837 68 957 232
rect 1061 68 1181 232
rect 1285 68 1405 232
rect 1509 68 1629 232
rect 1733 68 1853 232
rect 1957 68 2077 232
rect 2181 68 2301 232
rect 2405 68 2525 232
rect 2629 68 2749 232
rect 2957 93 3077 257
rect 3181 93 3301 257
rect 3405 93 3525 257
rect 3629 93 3749 257
rect 3853 93 3973 257
rect 4077 93 4197 257
rect 4301 93 4421 257
rect 4569 68 4689 232
<< mvpmos >>
rect 185 497 285 716
rect 409 497 509 716
rect 613 497 713 716
rect 857 497 957 716
rect 1061 497 1161 716
rect 1305 497 1405 716
rect 1509 497 1609 716
rect 1753 497 1853 716
rect 1977 497 2077 716
rect 2181 497 2281 716
rect 2425 497 2525 716
rect 2629 497 2729 716
rect 2977 497 3077 716
rect 3201 497 3301 716
rect 3405 497 3505 716
rect 3649 497 3749 716
rect 3853 497 3953 716
rect 4097 497 4197 716
rect 4301 497 4401 716
rect 4569 497 4669 716
<< mvndiff >>
rect 2857 232 2957 257
rect 77 219 165 232
rect 77 173 90 219
rect 136 173 165 219
rect 77 68 165 173
rect 285 127 389 232
rect 285 81 314 127
rect 360 81 389 127
rect 285 68 389 81
rect 509 219 613 232
rect 509 173 538 219
rect 584 173 613 219
rect 509 68 613 173
rect 733 127 837 232
rect 733 81 762 127
rect 808 81 837 127
rect 733 68 837 81
rect 957 219 1061 232
rect 957 173 986 219
rect 1032 173 1061 219
rect 957 68 1061 173
rect 1181 127 1285 232
rect 1181 81 1210 127
rect 1256 81 1285 127
rect 1181 68 1285 81
rect 1405 219 1509 232
rect 1405 173 1434 219
rect 1480 173 1509 219
rect 1405 68 1509 173
rect 1629 127 1733 232
rect 1629 81 1658 127
rect 1704 81 1733 127
rect 1629 68 1733 81
rect 1853 219 1957 232
rect 1853 173 1882 219
rect 1928 173 1957 219
rect 1853 68 1957 173
rect 2077 127 2181 232
rect 2077 81 2106 127
rect 2152 81 2181 127
rect 2077 68 2181 81
rect 2301 219 2405 232
rect 2301 173 2330 219
rect 2376 173 2405 219
rect 2301 68 2405 173
rect 2525 127 2629 232
rect 2525 81 2554 127
rect 2600 81 2629 127
rect 2525 68 2629 81
rect 2749 152 2957 232
rect 2749 106 2778 152
rect 2824 106 2957 152
rect 2749 93 2957 106
rect 3077 244 3181 257
rect 3077 198 3106 244
rect 3152 198 3181 244
rect 3077 93 3181 198
rect 3301 152 3405 257
rect 3301 106 3330 152
rect 3376 106 3405 152
rect 3301 93 3405 106
rect 3525 244 3629 257
rect 3525 198 3554 244
rect 3600 198 3629 244
rect 3525 93 3629 198
rect 3749 152 3853 257
rect 3749 106 3778 152
rect 3824 106 3853 152
rect 3749 93 3853 106
rect 3973 244 4077 257
rect 3973 198 4002 244
rect 4048 198 4077 244
rect 3973 93 4077 198
rect 4197 152 4301 257
rect 4197 106 4226 152
rect 4272 106 4301 152
rect 4197 93 4301 106
rect 4421 244 4509 257
rect 4421 198 4450 244
rect 4496 232 4509 244
rect 4496 198 4569 232
rect 4421 93 4569 198
rect 2749 68 2877 93
rect 4489 68 4569 93
rect 4689 152 4777 232
rect 4689 106 4718 152
rect 4764 106 4777 152
rect 4689 68 4777 106
<< mvpdiff >>
rect 87 665 185 716
rect 87 525 100 665
rect 146 525 185 665
rect 87 497 185 525
rect 285 497 409 716
rect 509 703 613 716
rect 509 657 538 703
rect 584 657 613 703
rect 509 497 613 657
rect 713 497 857 716
rect 957 634 1061 716
rect 957 588 986 634
rect 1032 588 1061 634
rect 957 497 1061 588
rect 1161 497 1305 716
rect 1405 703 1509 716
rect 1405 657 1434 703
rect 1480 657 1509 703
rect 1405 497 1509 657
rect 1609 497 1753 716
rect 1853 497 1977 716
rect 2077 562 2181 716
rect 2077 516 2106 562
rect 2152 516 2181 562
rect 2077 497 2181 516
rect 2281 674 2425 716
rect 2281 628 2330 674
rect 2376 628 2425 674
rect 2281 497 2425 628
rect 2525 562 2629 716
rect 2525 516 2554 562
rect 2600 516 2629 562
rect 2525 497 2629 516
rect 2729 674 2817 716
rect 2729 628 2758 674
rect 2804 628 2817 674
rect 2729 497 2817 628
rect 2889 703 2977 716
rect 2889 657 2902 703
rect 2948 657 2977 703
rect 2889 497 2977 657
rect 3077 497 3201 716
rect 3301 639 3405 716
rect 3301 593 3330 639
rect 3376 593 3405 639
rect 3301 497 3405 593
rect 3505 497 3649 716
rect 3749 703 3853 716
rect 3749 657 3778 703
rect 3824 657 3853 703
rect 3749 497 3853 657
rect 3953 497 4097 716
rect 4197 639 4301 716
rect 4197 593 4226 639
rect 4272 593 4301 639
rect 4197 497 4301 593
rect 4401 497 4569 716
rect 4669 665 4759 716
rect 4669 525 4700 665
rect 4746 525 4759 665
rect 4669 497 4759 525
<< mvndiffc >>
rect 90 173 136 219
rect 314 81 360 127
rect 538 173 584 219
rect 762 81 808 127
rect 986 173 1032 219
rect 1210 81 1256 127
rect 1434 173 1480 219
rect 1658 81 1704 127
rect 1882 173 1928 219
rect 2106 81 2152 127
rect 2330 173 2376 219
rect 2554 81 2600 127
rect 2778 106 2824 152
rect 3106 198 3152 244
rect 3330 106 3376 152
rect 3554 198 3600 244
rect 3778 106 3824 152
rect 4002 198 4048 244
rect 4226 106 4272 152
rect 4450 198 4496 244
rect 4718 106 4764 152
<< mvpdiffc >>
rect 100 525 146 665
rect 538 657 584 703
rect 986 588 1032 634
rect 1434 657 1480 703
rect 2106 516 2152 562
rect 2330 628 2376 674
rect 2554 516 2600 562
rect 2758 628 2804 674
rect 2902 657 2948 703
rect 3330 593 3376 639
rect 3778 657 3824 703
rect 4226 593 4272 639
rect 4700 525 4746 665
<< polysilicon >>
rect 185 716 285 760
rect 409 716 509 760
rect 613 716 713 760
rect 857 716 957 760
rect 1061 716 1161 760
rect 1305 716 1405 760
rect 1509 716 1609 760
rect 1753 716 1853 760
rect 1977 716 2077 760
rect 2181 716 2281 760
rect 2425 716 2525 760
rect 2629 716 2729 760
rect 2977 716 3077 760
rect 3201 716 3301 760
rect 3405 716 3505 760
rect 3649 716 3749 760
rect 3853 716 3953 760
rect 4097 716 4197 760
rect 4301 716 4401 760
rect 4569 716 4669 760
rect 185 415 285 497
rect 185 402 212 415
rect 165 369 212 402
rect 258 369 285 415
rect 409 415 509 497
rect 409 402 436 415
rect 165 232 285 369
rect 389 369 436 402
rect 482 394 509 415
rect 613 415 713 497
rect 613 394 640 415
rect 482 369 640 394
rect 686 402 713 415
rect 857 415 957 497
rect 857 402 884 415
rect 686 369 733 402
rect 389 348 733 369
rect 389 232 509 348
rect 613 232 733 348
rect 837 369 884 402
rect 930 394 957 415
rect 1061 415 1161 497
rect 1061 394 1088 415
rect 930 369 1088 394
rect 1134 402 1161 415
rect 1305 415 1405 497
rect 1305 402 1332 415
rect 1134 369 1181 402
rect 837 348 1181 369
rect 837 232 957 348
rect 1061 232 1181 348
rect 1285 369 1332 402
rect 1378 394 1405 415
rect 1509 415 1609 497
rect 1509 394 1536 415
rect 1378 369 1536 394
rect 1582 402 1609 415
rect 1753 415 1853 497
rect 1753 402 1780 415
rect 1582 369 1629 402
rect 1285 348 1629 369
rect 1285 232 1405 348
rect 1509 232 1629 348
rect 1733 369 1780 402
rect 1826 369 1853 415
rect 1977 415 2077 497
rect 1977 402 2004 415
rect 1733 232 1853 369
rect 1957 369 2004 402
rect 2050 402 2077 415
rect 2181 415 2281 497
rect 2181 402 2208 415
rect 2050 369 2208 402
rect 2254 402 2281 415
rect 2425 415 2525 497
rect 2425 402 2452 415
rect 2254 369 2452 402
rect 2498 402 2525 415
rect 2629 415 2729 497
rect 2629 402 2656 415
rect 2498 369 2656 402
rect 2702 402 2729 415
rect 2977 415 3077 497
rect 2977 402 3004 415
rect 2702 369 2749 402
rect 1957 348 2749 369
rect 1957 232 2077 348
rect 2181 232 2301 348
rect 2405 232 2525 348
rect 2629 232 2749 348
rect 2957 369 3004 402
rect 3050 369 3077 415
rect 3201 415 3301 497
rect 3201 402 3228 415
rect 2957 257 3077 369
rect 3181 369 3228 402
rect 3274 394 3301 415
rect 3405 415 3505 497
rect 3405 394 3432 415
rect 3274 369 3432 394
rect 3478 402 3505 415
rect 3649 433 3749 497
rect 3649 402 3676 433
rect 3478 369 3525 402
rect 3181 348 3525 369
rect 3181 257 3301 348
rect 3405 257 3525 348
rect 3629 387 3676 402
rect 3722 394 3749 433
rect 3853 433 3953 497
rect 3853 394 3880 433
rect 3722 387 3880 394
rect 3926 402 3953 433
rect 4097 415 4197 497
rect 4097 402 4124 415
rect 3926 387 3973 402
rect 3629 348 3973 387
rect 3629 257 3749 348
rect 3853 257 3973 348
rect 4077 369 4124 402
rect 4170 394 4197 415
rect 4301 415 4401 497
rect 4301 394 4328 415
rect 4170 369 4328 394
rect 4374 402 4401 415
rect 4569 415 4669 497
rect 4374 369 4421 402
rect 4077 348 4421 369
rect 4077 257 4197 348
rect 4301 257 4421 348
rect 4569 369 4596 415
rect 4642 402 4669 415
rect 4642 369 4689 402
rect 4569 232 4689 369
rect 165 24 285 68
rect 389 24 509 68
rect 613 24 733 68
rect 837 24 957 68
rect 1061 24 1181 68
rect 1285 24 1405 68
rect 1509 24 1629 68
rect 1733 24 1853 68
rect 1957 24 2077 68
rect 2181 24 2301 68
rect 2405 24 2525 68
rect 2629 24 2749 68
rect 2957 24 3077 93
rect 3181 24 3301 93
rect 3405 24 3525 93
rect 3629 24 3749 93
rect 3853 24 3973 93
rect 4077 24 4197 93
rect 4301 24 4421 93
rect 4569 24 4689 68
<< polycontact >>
rect 212 369 258 415
rect 436 369 482 415
rect 640 369 686 415
rect 884 369 930 415
rect 1088 369 1134 415
rect 1332 369 1378 415
rect 1536 369 1582 415
rect 1780 369 1826 415
rect 2004 369 2050 415
rect 2208 369 2254 415
rect 2452 369 2498 415
rect 2656 369 2702 415
rect 3004 369 3050 415
rect 3228 369 3274 415
rect 3432 369 3478 415
rect 3676 387 3722 433
rect 3880 387 3926 433
rect 4124 369 4170 415
rect 4328 369 4374 415
rect 4596 369 4642 415
<< metal1 >>
rect 0 724 4816 844
rect 527 703 595 724
rect 100 665 146 676
rect 527 657 538 703
rect 584 657 595 703
rect 1423 703 1491 724
rect 1423 657 1434 703
rect 1480 657 1491 703
rect 2891 703 2959 724
rect 646 611 986 634
rect 146 588 986 611
rect 1032 611 1373 634
rect 1638 628 2330 674
rect 2376 628 2758 674
rect 2804 628 2817 674
rect 2891 657 2902 703
rect 2948 657 2959 703
rect 3767 703 3835 724
rect 3767 657 3778 703
rect 3824 657 3835 703
rect 4700 665 4746 724
rect 3009 639 3717 648
rect 1638 611 1684 628
rect 1032 588 1684 611
rect 146 565 696 588
rect 1323 565 1684 588
rect 3009 593 3330 639
rect 3376 611 3717 639
rect 3885 639 4362 648
rect 3885 611 4226 639
rect 3376 593 4226 611
rect 4272 593 4362 639
rect 3009 584 4362 593
rect 3009 563 3059 584
rect 3667 565 3931 584
rect 1914 562 3059 563
rect 100 506 146 525
rect 746 516 1273 538
rect 1914 516 2106 562
rect 2152 516 2554 562
rect 2600 516 3059 562
rect 211 470 1827 516
rect 1914 472 3059 516
rect 3109 519 3610 536
rect 3989 519 4645 536
rect 3109 472 4645 519
rect 4700 506 4746 525
rect 211 415 259 470
rect 211 369 212 415
rect 258 369 259 415
rect 211 352 259 369
rect 346 415 774 424
rect 346 369 436 415
rect 482 369 640 415
rect 686 369 774 415
rect 346 360 774 369
rect 873 415 1145 470
rect 873 369 884 415
rect 930 369 1088 415
rect 1134 369 1145 415
rect 873 365 1145 369
rect 1242 415 1670 424
rect 1242 369 1332 415
rect 1378 369 1536 415
rect 1582 369 1670 415
rect 728 315 774 360
rect 1242 360 1670 369
rect 1779 415 1827 470
rect 1779 369 1780 415
rect 1826 369 1827 415
rect 1242 315 1288 360
rect 1779 352 1827 369
rect 1914 415 2776 424
rect 1914 369 2004 415
rect 2050 369 2208 415
rect 2254 369 2452 415
rect 2498 369 2656 415
rect 2702 369 2776 415
rect 1914 360 2776 369
rect 728 269 1288 315
rect 2824 244 2884 472
rect 3109 424 3155 472
rect 3665 433 3937 472
rect 2930 415 3155 424
rect 2930 369 3004 415
rect 3050 369 3155 415
rect 2930 360 3155 369
rect 3201 415 3574 424
rect 3201 369 3228 415
rect 3274 369 3432 415
rect 3478 369 3574 415
rect 3665 387 3676 433
rect 3722 387 3880 433
rect 3926 387 3937 433
rect 3665 382 3937 387
rect 4042 415 4470 424
rect 3201 360 3574 369
rect 3528 336 3574 360
rect 4042 369 4124 415
rect 4170 369 4328 415
rect 4374 369 4470 415
rect 4042 360 4470 369
rect 4593 415 4645 472
rect 4593 369 4596 415
rect 4642 369 4645 415
rect 4042 336 4088 360
rect 4593 352 4645 369
rect 3528 290 4088 336
rect 77 173 90 219
rect 136 173 538 219
rect 584 173 986 219
rect 1032 173 1434 219
rect 1480 173 1882 219
rect 1928 173 2330 219
rect 2376 173 2727 219
rect 2824 198 3106 244
rect 3152 198 3554 244
rect 3600 198 4002 244
rect 4048 198 4450 244
rect 4496 198 4507 244
rect 2681 152 2727 173
rect 303 81 314 127
rect 360 81 371 127
rect 303 60 371 81
rect 751 81 762 127
rect 808 81 819 127
rect 751 60 819 81
rect 1199 81 1210 127
rect 1256 81 1267 127
rect 1199 60 1267 81
rect 1647 81 1658 127
rect 1704 81 1715 127
rect 1647 60 1715 81
rect 2095 81 2106 127
rect 2152 81 2163 127
rect 2095 60 2163 81
rect 2543 81 2554 127
rect 2600 81 2611 127
rect 2681 106 2778 152
rect 2824 106 3330 152
rect 3376 106 3778 152
rect 3824 106 4226 152
rect 4272 106 4718 152
rect 4764 106 4777 152
rect 2543 60 2611 81
rect 0 -60 4816 60
<< labels >>
flabel metal1 s 1242 360 1670 424 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 4042 360 4470 424 0 FreeSans 400 0 0 0 B1
port 4 nsew default input
flabel metal1 s 3989 519 4645 536 0 FreeSans 400 0 0 0 B2
port 5 nsew default input
flabel metal1 s 0 724 4816 844 0 FreeSans 400 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 2543 60 2611 127 0 FreeSans 400 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 3885 611 4362 648 0 FreeSans 400 0 0 0 ZN
port 6 nsew default output
flabel metal1 s 1914 360 2776 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 746 516 1273 538 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
rlabel metal1 s 211 470 1827 516 1 A2
port 2 nsew default input
rlabel metal1 s 1779 365 1827 470 1 A2
port 2 nsew default input
rlabel metal1 s 873 365 1145 470 1 A2
port 2 nsew default input
rlabel metal1 s 211 365 259 470 1 A2
port 2 nsew default input
rlabel metal1 s 1779 352 1827 365 1 A2
port 2 nsew default input
rlabel metal1 s 211 352 259 365 1 A2
port 2 nsew default input
rlabel metal1 s 346 360 774 424 1 A3
port 3 nsew default input
rlabel metal1 s 1242 315 1288 360 1 A3
port 3 nsew default input
rlabel metal1 s 728 315 774 360 1 A3
port 3 nsew default input
rlabel metal1 s 728 269 1288 315 1 A3
port 3 nsew default input
rlabel metal1 s 3201 360 3574 424 1 B1
port 4 nsew default input
rlabel metal1 s 4042 336 4088 360 1 B1
port 4 nsew default input
rlabel metal1 s 3528 336 3574 360 1 B1
port 4 nsew default input
rlabel metal1 s 3528 290 4088 336 1 B1
port 4 nsew default input
rlabel metal1 s 3109 519 3610 536 1 B2
port 5 nsew default input
rlabel metal1 s 3109 472 4645 519 1 B2
port 5 nsew default input
rlabel metal1 s 4593 424 4645 472 1 B2
port 5 nsew default input
rlabel metal1 s 3665 424 3937 472 1 B2
port 5 nsew default input
rlabel metal1 s 3109 424 3155 472 1 B2
port 5 nsew default input
rlabel metal1 s 4593 382 4645 424 1 B2
port 5 nsew default input
rlabel metal1 s 3665 382 3937 424 1 B2
port 5 nsew default input
rlabel metal1 s 2930 382 3155 424 1 B2
port 5 nsew default input
rlabel metal1 s 4593 360 4645 382 1 B2
port 5 nsew default input
rlabel metal1 s 2930 360 3155 382 1 B2
port 5 nsew default input
rlabel metal1 s 4593 352 4645 360 1 B2
port 5 nsew default input
rlabel metal1 s 3009 611 3717 648 1 ZN
port 6 nsew default output
rlabel metal1 s 3009 584 4362 611 1 ZN
port 6 nsew default output
rlabel metal1 s 3667 565 3931 584 1 ZN
port 6 nsew default output
rlabel metal1 s 3009 565 3059 584 1 ZN
port 6 nsew default output
rlabel metal1 s 3009 563 3059 565 1 ZN
port 6 nsew default output
rlabel metal1 s 1914 472 3059 563 1 ZN
port 6 nsew default output
rlabel metal1 s 2824 244 2884 472 1 ZN
port 6 nsew default output
rlabel metal1 s 2824 198 4507 244 1 ZN
port 6 nsew default output
rlabel metal1 s 4700 657 4746 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3767 657 3835 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2891 657 2959 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1423 657 1491 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 527 657 595 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4700 506 4746 657 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2095 60 2163 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1647 60 1715 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1199 60 1267 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 751 60 819 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 303 60 371 127 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4816 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 784
string GDS_END 67528
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 59180
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
