magic
tech gf180mcuB
timestamp 1669390400
<< properties >>
string GDS_END 1306198
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1305746
<< end >>
