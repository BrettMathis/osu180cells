magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 3386
<< mvpmos >>
rect 0 0 120 3266
<< mvpdiff >>
rect -88 3253 0 3266
rect -88 3207 -75 3253
rect -29 3207 0 3253
rect -88 3150 0 3207
rect -88 3104 -75 3150
rect -29 3104 0 3150
rect -88 3047 0 3104
rect -88 3001 -75 3047
rect -29 3001 0 3047
rect -88 2944 0 3001
rect -88 2898 -75 2944
rect -29 2898 0 2944
rect -88 2841 0 2898
rect -88 2795 -75 2841
rect -29 2795 0 2841
rect -88 2738 0 2795
rect -88 2692 -75 2738
rect -29 2692 0 2738
rect -88 2635 0 2692
rect -88 2589 -75 2635
rect -29 2589 0 2635
rect -88 2532 0 2589
rect -88 2486 -75 2532
rect -29 2486 0 2532
rect -88 2429 0 2486
rect -88 2383 -75 2429
rect -29 2383 0 2429
rect -88 2326 0 2383
rect -88 2280 -75 2326
rect -29 2280 0 2326
rect -88 2223 0 2280
rect -88 2177 -75 2223
rect -29 2177 0 2223
rect -88 2120 0 2177
rect -88 2074 -75 2120
rect -29 2074 0 2120
rect -88 2017 0 2074
rect -88 1971 -75 2017
rect -29 1971 0 2017
rect -88 1914 0 1971
rect -88 1868 -75 1914
rect -29 1868 0 1914
rect -88 1811 0 1868
rect -88 1765 -75 1811
rect -29 1765 0 1811
rect -88 1708 0 1765
rect -88 1662 -75 1708
rect -29 1662 0 1708
rect -88 1605 0 1662
rect -88 1559 -75 1605
rect -29 1559 0 1605
rect -88 1502 0 1559
rect -88 1456 -75 1502
rect -29 1456 0 1502
rect -88 1399 0 1456
rect -88 1353 -75 1399
rect -29 1353 0 1399
rect -88 1296 0 1353
rect -88 1250 -75 1296
rect -29 1250 0 1296
rect -88 1193 0 1250
rect -88 1147 -75 1193
rect -29 1147 0 1193
rect -88 1090 0 1147
rect -88 1044 -75 1090
rect -29 1044 0 1090
rect -88 987 0 1044
rect -88 941 -75 987
rect -29 941 0 987
rect -88 884 0 941
rect -88 838 -75 884
rect -29 838 0 884
rect -88 781 0 838
rect -88 735 -75 781
rect -29 735 0 781
rect -88 678 0 735
rect -88 632 -75 678
rect -29 632 0 678
rect -88 575 0 632
rect -88 529 -75 575
rect -29 529 0 575
rect -88 472 0 529
rect -88 426 -75 472
rect -29 426 0 472
rect -88 369 0 426
rect -88 323 -75 369
rect -29 323 0 369
rect -88 266 0 323
rect -88 220 -75 266
rect -29 220 0 266
rect -88 163 0 220
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 3253 208 3266
rect 120 3207 149 3253
rect 195 3207 208 3253
rect 120 3150 208 3207
rect 120 3104 149 3150
rect 195 3104 208 3150
rect 120 3047 208 3104
rect 120 3001 149 3047
rect 195 3001 208 3047
rect 120 2944 208 3001
rect 120 2898 149 2944
rect 195 2898 208 2944
rect 120 2841 208 2898
rect 120 2795 149 2841
rect 195 2795 208 2841
rect 120 2738 208 2795
rect 120 2692 149 2738
rect 195 2692 208 2738
rect 120 2635 208 2692
rect 120 2589 149 2635
rect 195 2589 208 2635
rect 120 2532 208 2589
rect 120 2486 149 2532
rect 195 2486 208 2532
rect 120 2429 208 2486
rect 120 2383 149 2429
rect 195 2383 208 2429
rect 120 2326 208 2383
rect 120 2280 149 2326
rect 195 2280 208 2326
rect 120 2223 208 2280
rect 120 2177 149 2223
rect 195 2177 208 2223
rect 120 2120 208 2177
rect 120 2074 149 2120
rect 195 2074 208 2120
rect 120 2017 208 2074
rect 120 1971 149 2017
rect 195 1971 208 2017
rect 120 1914 208 1971
rect 120 1868 149 1914
rect 195 1868 208 1914
rect 120 1811 208 1868
rect 120 1765 149 1811
rect 195 1765 208 1811
rect 120 1708 208 1765
rect 120 1662 149 1708
rect 195 1662 208 1708
rect 120 1605 208 1662
rect 120 1559 149 1605
rect 195 1559 208 1605
rect 120 1502 208 1559
rect 120 1456 149 1502
rect 195 1456 208 1502
rect 120 1399 208 1456
rect 120 1353 149 1399
rect 195 1353 208 1399
rect 120 1296 208 1353
rect 120 1250 149 1296
rect 195 1250 208 1296
rect 120 1193 208 1250
rect 120 1147 149 1193
rect 195 1147 208 1193
rect 120 1090 208 1147
rect 120 1044 149 1090
rect 195 1044 208 1090
rect 120 987 208 1044
rect 120 941 149 987
rect 195 941 208 987
rect 120 884 208 941
rect 120 838 149 884
rect 195 838 208 884
rect 120 781 208 838
rect 120 735 149 781
rect 195 735 208 781
rect 120 678 208 735
rect 120 632 149 678
rect 195 632 208 678
rect 120 575 208 632
rect 120 529 149 575
rect 195 529 208 575
rect 120 472 208 529
rect 120 426 149 472
rect 195 426 208 472
rect 120 369 208 426
rect 120 323 149 369
rect 195 323 208 369
rect 120 266 208 323
rect 120 220 149 266
rect 195 220 208 266
rect 120 163 208 220
rect 120 117 149 163
rect 195 117 208 163
rect 120 59 208 117
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 3207 -29 3253
rect -75 3104 -29 3150
rect -75 3001 -29 3047
rect -75 2898 -29 2944
rect -75 2795 -29 2841
rect -75 2692 -29 2738
rect -75 2589 -29 2635
rect -75 2486 -29 2532
rect -75 2383 -29 2429
rect -75 2280 -29 2326
rect -75 2177 -29 2223
rect -75 2074 -29 2120
rect -75 1971 -29 2017
rect -75 1868 -29 1914
rect -75 1765 -29 1811
rect -75 1662 -29 1708
rect -75 1559 -29 1605
rect -75 1456 -29 1502
rect -75 1353 -29 1399
rect -75 1250 -29 1296
rect -75 1147 -29 1193
rect -75 1044 -29 1090
rect -75 941 -29 987
rect -75 838 -29 884
rect -75 735 -29 781
rect -75 632 -29 678
rect -75 529 -29 575
rect -75 426 -29 472
rect -75 323 -29 369
rect -75 220 -29 266
rect -75 117 -29 163
rect -75 13 -29 59
rect 149 3207 195 3253
rect 149 3104 195 3150
rect 149 3001 195 3047
rect 149 2898 195 2944
rect 149 2795 195 2841
rect 149 2692 195 2738
rect 149 2589 195 2635
rect 149 2486 195 2532
rect 149 2383 195 2429
rect 149 2280 195 2326
rect 149 2177 195 2223
rect 149 2074 195 2120
rect 149 1971 195 2017
rect 149 1868 195 1914
rect 149 1765 195 1811
rect 149 1662 195 1708
rect 149 1559 195 1605
rect 149 1456 195 1502
rect 149 1353 195 1399
rect 149 1250 195 1296
rect 149 1147 195 1193
rect 149 1044 195 1090
rect 149 941 195 987
rect 149 838 195 884
rect 149 735 195 781
rect 149 632 195 678
rect 149 529 195 575
rect 149 426 195 472
rect 149 323 195 369
rect 149 220 195 266
rect 149 117 195 163
rect 149 13 195 59
<< polysilicon >>
rect 0 3266 120 3310
rect 0 -44 120 0
<< metal1 >>
rect -75 3253 -29 3266
rect -75 3150 -29 3207
rect -75 3047 -29 3104
rect -75 2944 -29 3001
rect -75 2841 -29 2898
rect -75 2738 -29 2795
rect -75 2635 -29 2692
rect -75 2532 -29 2589
rect -75 2429 -29 2486
rect -75 2326 -29 2383
rect -75 2223 -29 2280
rect -75 2120 -29 2177
rect -75 2017 -29 2074
rect -75 1914 -29 1971
rect -75 1811 -29 1868
rect -75 1708 -29 1765
rect -75 1605 -29 1662
rect -75 1502 -29 1559
rect -75 1399 -29 1456
rect -75 1296 -29 1353
rect -75 1193 -29 1250
rect -75 1090 -29 1147
rect -75 987 -29 1044
rect -75 884 -29 941
rect -75 781 -29 838
rect -75 678 -29 735
rect -75 575 -29 632
rect -75 472 -29 529
rect -75 369 -29 426
rect -75 266 -29 323
rect -75 163 -29 220
rect -75 59 -29 117
rect -75 0 -29 13
rect 149 3253 195 3266
rect 149 3150 195 3207
rect 149 3047 195 3104
rect 149 2944 195 3001
rect 149 2841 195 2898
rect 149 2738 195 2795
rect 149 2635 195 2692
rect 149 2532 195 2589
rect 149 2429 195 2486
rect 149 2326 195 2383
rect 149 2223 195 2280
rect 149 2120 195 2177
rect 149 2017 195 2074
rect 149 1914 195 1971
rect 149 1811 195 1868
rect 149 1708 195 1765
rect 149 1605 195 1662
rect 149 1502 195 1559
rect 149 1399 195 1456
rect 149 1296 195 1353
rect 149 1193 195 1250
rect 149 1090 195 1147
rect 149 987 195 1044
rect 149 884 195 941
rect 149 781 195 838
rect 149 678 195 735
rect 149 575 195 632
rect 149 472 195 529
rect 149 369 195 426
rect 149 266 195 323
rect 149 163 195 220
rect 149 59 195 117
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1633 -52 1633 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1633 172 1633 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 126684
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 121628
<< end >>
