magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 4020
<< mvpmos >>
rect 0 0 120 3900
<< mvpdiff >>
rect -88 3887 0 3900
rect -88 13 -75 3887
rect -29 13 0 3887
rect -88 0 0 13
rect 120 3887 208 3900
rect 120 13 149 3887
rect 195 13 208 3887
rect 120 0 208 13
<< mvpdiffc >>
rect -75 13 -29 3887
rect 149 13 195 3887
<< polysilicon >>
rect 0 3900 120 3944
rect 0 -44 120 0
<< metal1 >>
rect -75 3887 -29 3900
rect -75 0 -29 13
rect 149 3887 195 3900
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1950 -52 1950 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1950 172 1950 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 409418
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 403466
<< end >>
