magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -141 344 4041
<< polysilicon >>
rect -31 3900 88 3973
rect -31 -74 88 0
use pmos_5p04310589983294_64x8m81  pmos_5p04310589983294_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 4020
<< properties >>
string GDS_END 862794
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 862480
<< end >>
