magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 5488 844
rect 262 601 330 724
rect 610 600 678 724
rect 1517 633 1586 724
rect 56 354 318 430
rect 578 354 810 430
rect 262 60 330 210
rect 654 60 722 215
rect 2690 607 2736 724
rect 2116 60 2184 183
rect 3541 588 3609 724
rect 3490 354 3708 430
rect 3645 264 3708 354
rect 3949 588 4017 724
rect 3876 354 4126 430
rect 4368 483 4414 724
rect 4516 514 4562 724
rect 4709 466 4777 676
rect 4924 514 4970 724
rect 5117 466 5246 676
rect 5332 514 5378 724
rect 4709 420 5246 466
rect 3949 60 4017 215
rect 5170 234 5246 420
rect 4720 188 5246 234
rect 4496 60 4542 153
rect 4720 110 4766 188
rect 4933 60 5001 142
rect 5168 110 5246 188
rect 5392 60 5438 153
rect 0 -60 5488 60
<< obsm1 >>
rect 69 534 115 660
rect 477 554 523 660
rect 757 621 1419 667
rect 757 554 803 621
rect 1373 587 1419 621
rect 1656 632 2644 678
rect 1656 587 1702 632
rect 69 487 411 534
rect 365 302 411 487
rect 49 256 411 302
rect 477 508 803 554
rect 49 162 95 256
rect 477 230 523 508
rect 477 162 543 230
rect 858 169 946 566
rect 1062 403 1130 566
rect 1281 495 1327 574
rect 1373 541 1702 587
rect 2102 563 2170 575
rect 1748 517 2170 563
rect 2358 529 2552 575
rect 1748 495 1794 517
rect 1281 449 1794 495
rect 2506 469 2552 529
rect 2598 561 2644 632
rect 2835 632 3096 678
rect 2835 561 2881 632
rect 2598 515 2881 561
rect 2927 469 2995 575
rect 1840 414 2460 460
rect 2506 425 2995 469
rect 2506 423 2950 425
rect 1840 403 1886 414
rect 1062 357 1886 403
rect 1113 158 1159 357
rect 1932 321 2368 367
rect 1932 311 1978 321
rect 1227 204 1295 311
rect 1406 265 1978 311
rect 2024 229 2276 275
rect 2024 204 2070 229
rect 1227 158 2070 204
rect 2230 152 2276 229
rect 2322 263 2368 321
rect 2414 355 2460 414
rect 2414 309 2494 355
rect 2893 263 2950 423
rect 3050 414 3096 632
rect 3142 632 3495 678
rect 3142 263 3188 632
rect 3335 274 3403 579
rect 3449 542 3495 632
rect 3655 617 3894 664
rect 3655 542 3701 617
rect 3449 495 3701 542
rect 2322 217 2950 263
rect 2996 217 3188 263
rect 3234 263 3403 274
rect 3234 217 3592 263
rect 3234 206 3291 217
rect 3535 215 3592 217
rect 3756 215 3802 571
rect 3848 542 3894 617
rect 4063 617 4322 664
rect 4063 542 4109 617
rect 3848 496 4109 542
rect 4164 503 4230 571
rect 4184 312 4230 503
rect 4276 382 4322 617
rect 4593 312 5078 364
rect 4184 308 5078 312
rect 3861 295 5078 308
rect 3861 266 4661 295
rect 3861 262 4398 266
rect 2886 152 2954 171
rect 3355 152 3423 171
rect 3535 158 3802 215
rect 2230 106 3423 152
rect 4352 158 4398 262
<< labels >>
rlabel metal1 s 578 354 810 430 6 D
port 1 nsew default input
rlabel metal1 s 3876 354 4126 430 6 RN
port 2 nsew default input
rlabel metal1 s 3490 354 3708 430 6 SETN
port 3 nsew default input
rlabel metal1 s 3645 264 3708 354 6 SETN
port 3 nsew default input
rlabel metal1 s 56 354 318 430 6 CLKN
port 4 nsew clock input
rlabel metal1 s 5117 466 5246 676 6 Q
port 5 nsew default output
rlabel metal1 s 4709 466 4777 676 6 Q
port 5 nsew default output
rlabel metal1 s 4709 420 5246 466 6 Q
port 5 nsew default output
rlabel metal1 s 5170 234 5246 420 6 Q
port 5 nsew default output
rlabel metal1 s 4720 188 5246 234 6 Q
port 5 nsew default output
rlabel metal1 s 5168 110 5246 188 6 Q
port 5 nsew default output
rlabel metal1 s 4720 110 4766 188 6 Q
port 5 nsew default output
rlabel metal1 s 0 724 5488 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 633 5378 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 633 4970 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 633 4562 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 633 4414 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 633 4017 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 633 3609 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2690 633 2736 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1517 633 1586 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 633 678 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 633 330 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 607 5378 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 607 4970 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 607 4562 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 607 4414 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 607 4017 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 607 3609 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2690 607 2736 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 607 678 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 607 330 633 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 601 5378 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 601 4970 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 601 4562 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 601 4414 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 601 4017 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 601 3609 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 601 678 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 601 330 607 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 600 5378 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 600 4970 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 600 4562 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 600 4414 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 600 4017 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 600 3609 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 600 678 601 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 588 5378 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 588 4970 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 588 4562 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 588 4414 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 588 4017 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 588 3609 600 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 514 5378 588 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 514 4970 588 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 514 4562 588 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 514 4414 588 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 483 4414 514 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 210 4017 215 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 210 722 215 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 183 4017 210 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 183 722 210 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 183 330 210 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 153 4017 183 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 153 2184 183 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 153 722 183 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 153 330 183 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5392 142 5438 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4496 142 4542 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 142 4017 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 142 2184 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 142 722 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 142 330 153 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5392 60 5438 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4933 60 5001 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4496 60 4542 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 60 4017 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 60 2184 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 60 722 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 142 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5488 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5488 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 922820
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 911874
<< end >>
