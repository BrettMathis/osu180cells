magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 1240 595
<< polysilicon >>
rect -31 454 88 527
rect 193 454 312 527
rect 417 454 536 527
rect 641 454 760 527
rect 865 454 984 527
rect -31 -74 88 -1
rect 193 -74 312 -1
rect 417 -74 536 -1
rect 641 -74 760 -1
rect 865 -74 984 -1
use pmos_5p04310590878137_256x8m81  pmos_5p04310590878137_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 1224 574
<< properties >>
string GDS_END 309054
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 308228
<< end >>
