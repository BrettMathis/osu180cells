magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -300 635 81 636
rect -300 -636 300 635
<< nsubdiff >>
rect -156 431 157 488
rect -156 385 -102 431
rect -56 385 56 431
rect 102 385 157 431
rect -156 268 157 385
rect -156 222 -102 268
rect -56 222 56 268
rect 102 222 157 268
rect -156 105 157 222
rect -156 59 -102 105
rect -56 59 56 105
rect 102 59 157 105
rect -156 -59 157 59
rect -156 -105 -102 -59
rect -56 -105 56 -59
rect 102 -105 157 -59
rect -156 -222 157 -105
rect -156 -268 -102 -222
rect -56 -268 56 -222
rect 102 -268 157 -222
rect -156 -385 157 -268
rect -156 -431 -102 -385
rect -56 -431 56 -385
rect 102 -431 157 -385
rect -156 -488 157 -431
<< nsubdiffcont >>
rect -102 385 -56 431
rect 56 385 102 431
rect -102 222 -56 268
rect 56 222 102 268
rect -102 59 -56 105
rect 56 59 102 105
rect -102 -105 -56 -59
rect 56 -105 102 -59
rect -102 -268 -56 -222
rect 56 -268 102 -222
rect -102 -431 -56 -385
rect 56 -431 102 -385
<< metal1 >>
rect -137 431 137 468
rect -137 385 -102 431
rect -56 385 56 431
rect 102 385 137 431
rect -137 268 137 385
rect -137 222 -102 268
rect -56 222 56 268
rect 102 222 137 268
rect -137 105 137 222
rect -137 59 -102 105
rect -56 59 56 105
rect 102 59 137 105
rect -137 -59 137 59
rect -137 -105 -102 -59
rect -56 -105 56 -59
rect 102 -105 137 -59
rect -137 -222 137 -105
rect -137 -268 -102 -222
rect -56 -268 56 -222
rect 102 -268 137 -222
rect -137 -385 137 -268
rect -137 -431 -102 -385
rect -56 -431 56 -385
rect 102 -431 137 -385
rect -137 -468 137 -431
<< properties >>
string GDS_END 377326
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 376282
<< end >>
