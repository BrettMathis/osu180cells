magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 2721 89 2794
rect -31 -74 89 -1
use nmos_5p0431059054877_128x8m81  nmos_5p0431059054877_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 2766
<< properties >>
string GDS_END 313002
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 312752
<< end >>
