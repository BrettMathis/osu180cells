magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 918 448 1098
rect 353 710 399 918
rect 49 90 95 298
rect 0 -90 448 90
<< obsm1 >>
rect 49 412 95 872
rect 254 494 399 540
rect 49 366 194 412
rect 353 136 399 494
<< labels >>
rlabel metal1 s 0 918 448 1098 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 710 399 918 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 49 90 95 298 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 448 90 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 1008
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 760750
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 758596
<< end >>
