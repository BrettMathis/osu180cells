magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -71 222 71 227
rect -71 -222 -66 222
rect 66 -222 71 222
rect -71 -227 71 -222
<< via2 >>
rect -66 -222 66 222
<< metal3 >>
rect -71 222 71 227
rect -71 -222 -66 222
rect 66 -222 71 222
rect -71 -227 71 -222
<< properties >>
string GDS_END 1822708
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1820848
<< end >>
