magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -19 449 19 454
rect -19 421 -14 449
rect 14 421 19 449
rect -19 391 19 421
rect -19 363 -14 391
rect 14 363 19 391
rect -19 333 19 363
rect -19 305 -14 333
rect 14 305 19 333
rect -19 275 19 305
rect -19 247 -14 275
rect 14 247 19 275
rect -19 217 19 247
rect -19 189 -14 217
rect 14 189 19 217
rect -19 159 19 189
rect -19 131 -14 159
rect 14 131 19 159
rect -19 101 19 131
rect -19 73 -14 101
rect 14 73 19 101
rect -19 43 19 73
rect -19 15 -14 43
rect 14 15 19 43
rect -19 -15 19 15
rect -19 -43 -14 -15
rect 14 -43 19 -15
rect -19 -73 19 -43
rect -19 -101 -14 -73
rect 14 -101 19 -73
rect -19 -131 19 -101
rect -19 -159 -14 -131
rect 14 -159 19 -131
rect -19 -189 19 -159
rect -19 -217 -14 -189
rect 14 -217 19 -189
rect -19 -247 19 -217
rect -19 -275 -14 -247
rect 14 -275 19 -247
rect -19 -305 19 -275
rect -19 -333 -14 -305
rect 14 -333 19 -305
rect -19 -363 19 -333
rect -19 -391 -14 -363
rect 14 -391 19 -363
rect -19 -421 19 -391
rect -19 -449 -14 -421
rect 14 -449 19 -421
rect -19 -454 19 -449
<< via2 >>
rect -14 421 14 449
rect -14 363 14 391
rect -14 305 14 333
rect -14 247 14 275
rect -14 189 14 217
rect -14 131 14 159
rect -14 73 14 101
rect -14 15 14 43
rect -14 -43 14 -15
rect -14 -101 14 -73
rect -14 -159 14 -131
rect -14 -217 14 -189
rect -14 -275 14 -247
rect -14 -333 14 -305
rect -14 -391 14 -363
rect -14 -449 14 -421
<< metal3 >>
rect -19 449 19 454
rect -19 421 -14 449
rect 14 421 19 449
rect -19 391 19 421
rect -19 363 -14 391
rect 14 363 19 391
rect -19 333 19 363
rect -19 305 -14 333
rect 14 305 19 333
rect -19 275 19 305
rect -19 247 -14 275
rect 14 247 19 275
rect -19 217 19 247
rect -19 189 -14 217
rect 14 189 19 217
rect -19 159 19 189
rect -19 131 -14 159
rect 14 131 19 159
rect -19 101 19 131
rect -19 73 -14 101
rect 14 73 19 101
rect -19 43 19 73
rect -19 15 -14 43
rect 14 15 19 43
rect -19 -15 19 15
rect -19 -43 -14 -15
rect 14 -43 19 -15
rect -19 -73 19 -43
rect -19 -101 -14 -73
rect 14 -101 19 -73
rect -19 -131 19 -101
rect -19 -159 -14 -131
rect 14 -159 19 -131
rect -19 -189 19 -159
rect -19 -217 -14 -189
rect 14 -217 19 -189
rect -19 -247 19 -217
rect -19 -275 -14 -247
rect 14 -275 19 -247
rect -19 -305 19 -275
rect -19 -333 -14 -305
rect 14 -333 19 -305
rect -19 -363 19 -333
rect -19 -391 -14 -363
rect 14 -391 19 -363
rect -19 -421 19 -391
rect -19 -449 -14 -421
rect 14 -449 19 -421
rect -19 -454 19 -449
<< properties >>
string GDS_END 1312768
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1311612
<< end >>
