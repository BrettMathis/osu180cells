magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -256 -141 344 595
<< polysilicon >>
rect -31 454 88 527
rect -31 -74 88 0
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 574
<< properties >>
string GDS_END 218762
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 218448
<< end >>
