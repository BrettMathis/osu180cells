magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
use nmos_5p04310590548788_128x8m81  nmos_5p04310590548788_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 4464 1518
<< properties >>
string GDS_END 846222
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 846100
<< end >>
