magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1456 844
rect 266 608 312 724
rect 530 472 1191 540
rect 116 360 456 425
rect 530 220 594 472
rect 658 360 1345 424
rect 658 280 726 360
rect 800 248 1345 312
rect 194 174 665 220
rect 62 60 108 153
rect 194 112 449 174
rect 619 161 665 174
rect 499 60 567 128
rect 619 115 995 161
rect 1330 60 1376 153
rect 0 -60 1456 60
<< obsm1 >>
rect 62 552 108 676
rect 360 619 1376 665
rect 360 552 407 619
rect 62 506 407 552
rect 1330 487 1376 619
<< labels >>
rlabel metal1 s 800 248 1345 312 6 A1
port 1 nsew default input
rlabel metal1 s 658 360 1345 424 6 A2
port 2 nsew default input
rlabel metal1 s 658 280 726 360 6 A2
port 2 nsew default input
rlabel metal1 s 116 360 456 425 6 B
port 3 nsew default input
rlabel metal1 s 530 472 1191 540 6 ZN
port 4 nsew default output
rlabel metal1 s 530 220 594 472 6 ZN
port 4 nsew default output
rlabel metal1 s 194 174 665 220 6 ZN
port 4 nsew default output
rlabel metal1 s 619 161 665 174 6 ZN
port 4 nsew default output
rlabel metal1 s 194 161 449 174 6 ZN
port 4 nsew default output
rlabel metal1 s 619 115 995 161 6 ZN
port 4 nsew default output
rlabel metal1 s 194 115 449 161 6 ZN
port 4 nsew default output
rlabel metal1 s 194 112 449 115 6 ZN
port 4 nsew default output
rlabel metal1 s 0 724 1456 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 266 608 312 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1330 128 1376 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 62 128 108 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1330 60 1376 128 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 499 60 567 128 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 62 60 108 128 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1456 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1230370
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1226642
<< end >>
