magic
tech gf180mcuC
magscale 1 10
timestamp 1669650257
<< checkpaint >>
rect 34400 34400 73000 73000
<< metal4 >>
rect 36400 55421 39400 71000
tri 39400 55421 40644 56665 sw
tri 36400 53376 38445 55421 ne
rect 38445 53376 40644 55421
tri 40644 53376 42689 55421 sw
tri 38445 49132 42689 53376 ne
tri 42689 49132 46933 53376 sw
tri 42689 44888 46933 49132 ne
tri 46933 44888 51177 49132 sw
tri 46933 40644 51177 44888 ne
tri 51177 40644 55421 44888 sw
tri 51177 36400 55421 40644 ne
tri 55421 39400 56665 40644 sw
rect 55421 36400 71000 39400
<< end >>
