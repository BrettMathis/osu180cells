magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -30 907 88 980
rect -30 -73 88 0
use nmos_5p04310591302057_512x8m81  nmos_5p04310591302057_512x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 952
<< properties >>
string GDS_END 312302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 312052
<< end >>
