magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 1900 1230
<< nmos >>
rect 200 190 260 360
rect 400 190 460 360
rect 540 190 600 360
rect 710 190 770 360
rect 950 190 1010 360
rect 1150 190 1210 360
rect 1470 190 1530 360
rect 1640 190 1700 360
<< pmos >>
rect 200 700 260 1040
rect 370 700 430 1040
rect 540 700 600 1040
rect 710 700 770 1040
rect 980 700 1040 1040
rect 1150 700 1210 1040
rect 1470 700 1530 1040
rect 1640 700 1700 1040
<< ndiff >>
rect 100 298 200 360
rect 100 252 122 298
rect 168 252 200 298
rect 100 190 200 252
rect 260 268 400 360
rect 260 222 307 268
rect 353 222 400 268
rect 260 190 400 222
rect 460 190 540 360
rect 600 273 710 360
rect 600 227 632 273
rect 678 227 710 273
rect 600 190 710 227
rect 770 190 950 360
rect 1010 263 1150 360
rect 1010 217 1057 263
rect 1103 217 1150 263
rect 1010 190 1150 217
rect 1210 298 1310 360
rect 1210 252 1242 298
rect 1288 252 1310 298
rect 1210 190 1310 252
rect 1370 298 1470 360
rect 1370 252 1392 298
rect 1438 252 1470 298
rect 1370 190 1470 252
rect 1530 263 1640 360
rect 1530 217 1562 263
rect 1608 217 1640 263
rect 1530 190 1640 217
rect 1700 298 1800 360
rect 1700 252 1732 298
rect 1778 252 1800 298
rect 1700 190 1800 252
<< pdiff >>
rect 100 987 200 1040
rect 100 753 122 987
rect 168 753 200 987
rect 100 700 200 753
rect 260 1020 370 1040
rect 260 880 292 1020
rect 338 880 370 1020
rect 260 700 370 880
rect 430 700 540 1040
rect 600 1017 710 1040
rect 600 783 632 1017
rect 678 783 710 1017
rect 600 700 710 783
rect 770 700 980 1040
rect 1040 1012 1150 1040
rect 1040 778 1072 1012
rect 1118 778 1150 1012
rect 1040 700 1150 778
rect 1210 1017 1310 1040
rect 1210 783 1242 1017
rect 1288 783 1310 1017
rect 1210 700 1310 783
rect 1370 992 1470 1040
rect 1370 758 1392 992
rect 1438 758 1470 992
rect 1370 700 1470 758
rect 1530 1010 1640 1040
rect 1530 870 1562 1010
rect 1608 870 1640 1010
rect 1530 700 1640 870
rect 1700 987 1800 1040
rect 1700 753 1732 987
rect 1778 753 1800 987
rect 1700 700 1800 753
<< ndiffc >>
rect 122 252 168 298
rect 307 222 353 268
rect 632 227 678 273
rect 1057 217 1103 263
rect 1242 252 1288 298
rect 1392 252 1438 298
rect 1562 217 1608 263
rect 1732 252 1778 298
<< pdiffc >>
rect 122 753 168 987
rect 292 880 338 1020
rect 632 783 678 1017
rect 1072 778 1118 1012
rect 1242 783 1288 1017
rect 1392 758 1438 992
rect 1562 870 1608 1010
rect 1732 753 1778 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 340 98 430 120
rect 340 52 362 98
rect 408 52 430 98
rect 340 30 430 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1060 98 1150 120
rect 1060 52 1082 98
rect 1128 52 1150 98
rect 1060 30 1150 52
rect 1290 98 1390 120
rect 1290 52 1312 98
rect 1358 52 1390 98
rect 1290 30 1390 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 340 1178 430 1200
rect 340 1132 362 1178
rect 408 1132 430 1178
rect 340 1110 430 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1060 1178 1150 1200
rect 1060 1132 1082 1178
rect 1128 1132 1150 1178
rect 1060 1110 1150 1132
rect 1300 1178 1390 1200
rect 1300 1132 1322 1178
rect 1368 1132 1390 1178
rect 1300 1110 1390 1132
rect 1540 1178 1630 1200
rect 1540 1132 1562 1178
rect 1608 1132 1630 1178
rect 1540 1110 1630 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 362 52 408 98
rect 592 52 638 98
rect 832 52 878 98
rect 1082 52 1128 98
rect 1312 52 1358 98
rect 1552 52 1598 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 362 1132 408 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1082 1132 1128 1178
rect 1322 1132 1368 1178
rect 1562 1132 1608 1178
<< polysilicon >>
rect 200 1040 260 1090
rect 370 1040 430 1090
rect 540 1040 600 1090
rect 710 1040 770 1090
rect 980 1040 1040 1090
rect 1150 1040 1210 1090
rect 1470 1040 1530 1090
rect 1640 1040 1700 1090
rect 200 680 260 700
rect 200 653 320 680
rect 200 607 237 653
rect 283 607 320 653
rect 200 580 320 607
rect 370 650 430 700
rect 540 680 600 700
rect 710 680 770 700
rect 520 653 620 680
rect 370 623 470 650
rect 200 360 260 580
rect 370 577 397 623
rect 443 577 470 623
rect 520 607 547 653
rect 593 607 620 653
rect 520 580 620 607
rect 680 653 780 680
rect 680 607 707 653
rect 753 607 780 653
rect 680 580 780 607
rect 370 550 470 577
rect 370 420 430 550
rect 710 530 770 580
rect 540 490 770 530
rect 830 543 930 570
rect 830 497 857 543
rect 903 497 930 543
rect 370 380 460 420
rect 400 360 460 380
rect 540 360 600 490
rect 830 470 930 497
rect 980 550 1040 700
rect 1150 680 1210 700
rect 1140 653 1240 680
rect 1140 607 1167 653
rect 1213 607 1240 653
rect 1140 580 1240 607
rect 980 523 1100 550
rect 980 477 1027 523
rect 1073 477 1100 523
rect 830 440 900 470
rect 710 400 900 440
rect 980 450 1100 477
rect 980 420 1040 450
rect 710 360 770 400
rect 950 380 1040 420
rect 950 360 1010 380
rect 1150 360 1210 580
rect 1470 550 1530 700
rect 1640 550 1700 700
rect 1440 528 1530 550
rect 1440 482 1462 528
rect 1508 482 1530 528
rect 1440 460 1530 482
rect 1470 360 1530 460
rect 1580 523 1700 550
rect 1580 477 1607 523
rect 1653 477 1700 523
rect 1580 450 1700 477
rect 1640 360 1700 450
rect 200 140 260 190
rect 400 140 460 190
rect 540 140 600 190
rect 710 140 770 190
rect 950 140 1010 190
rect 1150 140 1210 190
rect 1470 140 1530 190
rect 1640 140 1700 190
<< polycontact >>
rect 237 607 283 653
rect 397 577 443 623
rect 547 607 593 653
rect 707 607 753 653
rect 857 497 903 543
rect 1167 607 1213 653
rect 1027 477 1073 523
rect 1462 482 1508 528
rect 1607 477 1653 523
<< metal1 >>
rect 0 1178 1900 1230
rect 0 1132 112 1178
rect 158 1176 362 1178
rect 0 1124 114 1132
rect 166 1124 354 1176
rect 408 1132 592 1178
rect 638 1176 832 1178
rect 878 1176 1082 1178
rect 1128 1176 1322 1178
rect 1368 1176 1562 1178
rect 646 1132 832 1176
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1176
rect 1128 1132 1314 1176
rect 1368 1132 1554 1176
rect 1608 1132 1900 1178
rect 1126 1124 1314 1132
rect 1366 1124 1554 1132
rect 1606 1124 1900 1132
rect 0 1110 1900 1124
rect 120 987 170 1040
rect 120 753 122 987
rect 168 753 170 987
rect 290 1020 340 1110
rect 290 880 292 1020
rect 338 880 340 1020
rect 290 860 340 880
rect 630 1017 680 1040
rect 630 810 632 1017
rect 120 510 170 753
rect 230 783 632 810
rect 678 783 680 1017
rect 230 760 680 783
rect 1070 1012 1120 1110
rect 1070 778 1072 1012
rect 1118 778 1120 1012
rect 230 660 280 760
rect 1070 750 1120 778
rect 1240 1017 1290 1040
rect 1240 783 1242 1017
rect 1288 783 1290 1017
rect 1240 780 1290 783
rect 1390 992 1440 1040
rect 1240 730 1340 780
rect 220 653 310 660
rect 220 607 237 653
rect 283 607 310 653
rect 520 653 620 660
rect 220 600 310 607
rect 370 626 470 630
rect 100 500 170 510
rect 70 496 170 500
rect 70 444 94 496
rect 146 444 170 496
rect 70 440 170 444
rect 90 430 170 440
rect 120 298 170 430
rect 230 430 280 600
rect 370 574 394 626
rect 446 574 470 626
rect 520 607 547 653
rect 593 607 620 653
rect 520 600 620 607
rect 680 653 780 660
rect 680 626 707 653
rect 753 626 780 653
rect 370 570 470 574
rect 540 520 600 600
rect 680 574 704 626
rect 756 574 780 626
rect 1140 656 1240 660
rect 1140 604 1164 656
rect 1216 604 1240 656
rect 1140 600 1240 604
rect 680 570 780 574
rect 830 543 930 550
rect 830 520 857 543
rect 540 497 857 520
rect 903 497 930 543
rect 540 490 930 497
rect 1000 526 1100 530
rect 540 470 910 490
rect 1000 474 1024 526
rect 1076 474 1100 526
rect 1000 470 1100 474
rect 540 460 900 470
rect 230 380 480 430
rect 120 252 122 298
rect 168 252 170 298
rect 120 190 170 252
rect 290 268 370 300
rect 290 222 307 268
rect 353 222 370 268
rect 430 290 480 380
rect 840 390 900 460
rect 1290 450 1340 730
rect 1390 758 1392 992
rect 1438 758 1440 992
rect 1560 1010 1610 1110
rect 1560 870 1562 1010
rect 1608 870 1610 1010
rect 1560 840 1610 870
rect 1730 987 1780 1040
rect 1390 720 1440 758
rect 1730 753 1732 987
rect 1778 753 1780 987
rect 1390 670 1660 720
rect 1440 528 1540 530
rect 1440 482 1462 528
rect 1508 526 1540 528
rect 1440 474 1464 482
rect 1516 474 1540 526
rect 1440 470 1540 474
rect 1600 523 1660 670
rect 1600 477 1607 523
rect 1653 477 1660 523
rect 1240 400 1340 450
rect 1600 420 1660 477
rect 1240 390 1290 400
rect 840 340 1290 390
rect 630 290 680 310
rect 1240 298 1290 340
rect 430 273 680 290
rect 430 240 632 273
rect 290 120 370 222
rect 630 227 632 240
rect 678 227 680 273
rect 630 190 680 227
rect 1040 263 1120 290
rect 1040 217 1057 263
rect 1103 217 1120 263
rect 1040 120 1120 217
rect 1240 252 1242 298
rect 1288 252 1290 298
rect 1240 190 1290 252
rect 1390 370 1660 420
rect 1730 640 1780 753
rect 1730 630 1810 640
rect 1730 626 1830 630
rect 1730 574 1754 626
rect 1806 574 1830 626
rect 1730 570 1830 574
rect 1730 560 1810 570
rect 1390 298 1440 370
rect 1390 252 1392 298
rect 1438 252 1440 298
rect 1730 298 1780 560
rect 1390 190 1440 252
rect 1560 263 1610 290
rect 1560 217 1562 263
rect 1608 217 1610 263
rect 1560 120 1610 217
rect 1730 252 1732 298
rect 1778 252 1780 298
rect 1730 190 1780 252
rect 0 106 1900 120
rect 0 98 114 106
rect 0 52 112 98
rect 166 54 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 158 52 362 54
rect 408 52 592 98
rect 646 54 832 98
rect 886 54 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 638 52 832 54
rect 878 52 1082 54
rect 1128 52 1312 98
rect 1366 54 1552 98
rect 1606 54 1900 106
rect 1358 52 1552 54
rect 1598 52 1900 54
rect 0 0 1900 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 114 1124 166 1132
rect 354 1132 362 1176
rect 362 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1132 1082 1176
rect 1082 1132 1126 1176
rect 1314 1132 1322 1176
rect 1322 1132 1366 1176
rect 1554 1132 1562 1176
rect 1562 1132 1606 1176
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 1554 1124 1606 1132
rect 94 444 146 496
rect 394 623 446 626
rect 394 577 397 623
rect 397 577 443 623
rect 443 577 446 623
rect 394 574 446 577
rect 704 607 707 626
rect 707 607 753 626
rect 753 607 756 626
rect 704 574 756 607
rect 1164 653 1216 656
rect 1164 607 1167 653
rect 1167 607 1213 653
rect 1213 607 1216 653
rect 1164 604 1216 607
rect 1024 523 1076 526
rect 1024 477 1027 523
rect 1027 477 1073 523
rect 1073 477 1076 523
rect 1024 474 1076 477
rect 1464 482 1508 526
rect 1508 482 1516 526
rect 1464 474 1516 482
rect 1754 574 1806 626
rect 114 98 166 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 354 54 362 98
rect 362 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1074 54 1082 98
rect 1082 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 1540 1180 1620 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 1530 1176 1630 1180
rect 1530 1124 1554 1176
rect 1606 1124 1630 1176
rect 1530 1120 1630 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 1540 1110 1620 1120
rect 1140 660 1240 670
rect 700 656 1240 660
rect 700 640 1164 656
rect 370 626 470 640
rect 690 630 1164 640
rect 370 574 394 626
rect 446 574 470 626
rect 370 560 470 574
rect 680 626 1164 630
rect 680 574 704 626
rect 756 604 1164 626
rect 1216 604 1240 656
rect 1740 630 1820 640
rect 756 600 1240 604
rect 756 574 780 600
rect 1140 590 1240 600
rect 1730 626 1830 630
rect 680 570 780 574
rect 1730 574 1754 626
rect 1806 574 1830 626
rect 1730 570 1830 574
rect 690 560 770 570
rect 1740 560 1820 570
rect 1010 530 1090 540
rect 1440 530 1540 540
rect 920 526 1540 530
rect 70 500 170 510
rect 920 500 1024 526
rect 70 496 1024 500
rect 70 444 94 496
rect 146 474 1024 496
rect 1076 474 1464 526
rect 1516 474 1540 526
rect 146 470 1540 474
rect 146 460 1090 470
rect 1440 460 1540 470
rect 146 444 980 460
rect 70 440 980 444
rect 70 430 170 440
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 370 560 470 640 4 D
port 1 nsew signal input
rlabel metal2 s 1740 560 1820 640 4 Q
port 2 nsew signal output
rlabel metal2 s 690 560 770 640 4 CLK
port 3 nsew clock input
rlabel metal2 s 680 570 780 630 1 CLK
port 3 nsew clock input
rlabel metal2 s 700 600 1240 660 1 CLK
port 3 nsew clock input
rlabel metal2 s 1140 590 1240 670 1 CLK
port 3 nsew clock input
rlabel metal1 s 680 570 780 660 1 CLK
port 3 nsew clock input
rlabel metal1 s 1140 600 1240 660 1 CLK
port 3 nsew clock input
rlabel metal1 s 370 570 470 630 1 D
port 1 nsew signal input
rlabel metal2 s 1730 570 1830 630 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 190 1780 1040 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 560 1810 640 1 Q
port 2 nsew signal output
rlabel metal1 s 1730 570 1830 630 1 Q
port 2 nsew signal output
rlabel metal2 s 90 1120 190 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1540 1110 1620 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1530 1120 1630 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 290 860 340 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1070 750 1120 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1560 840 1610 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1110 1900 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 290 0 370 300 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 1040 0 1120 290 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 1560 0 1610 290 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 0 1900 120 1 VSS
port 9 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1900 1230
string GDS_END 334522
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 316786
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
