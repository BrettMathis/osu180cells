magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4790 1094
<< pwell >>
rect -86 -86 4790 453
<< mvnmos >>
rect 124 156 244 274
rect 348 156 468 274
rect 516 156 636 274
rect 740 156 860 274
rect 908 156 1028 274
rect 1317 166 1437 324
rect 1541 166 1661 324
rect 1913 195 2033 313
rect 2137 195 2257 313
rect 2305 195 2425 313
rect 2477 195 2597 313
rect 2701 195 2821 313
rect 2925 195 3045 313
rect 3153 195 3273 313
rect 3421 195 3541 313
rect 3681 124 3801 324
rect 3849 124 3969 324
rect 4236 68 4356 332
rect 4460 68 4580 332
<< mvpmos >>
rect 144 652 244 852
rect 348 652 448 852
rect 496 652 596 852
rect 740 652 840 852
rect 888 652 988 852
rect 1317 580 1417 856
rect 1521 580 1621 856
rect 1869 652 1969 852
rect 2073 652 2173 852
rect 2277 652 2377 852
rect 2481 652 2581 852
rect 2829 652 2929 852
rect 3033 652 3133 852
rect 3237 652 3337 852
rect 3441 652 3541 852
rect 3733 663 3833 939
rect 3937 663 4037 939
rect 4246 573 4346 939
rect 4454 573 4554 939
<< mvndiff >>
rect 1229 311 1317 324
rect 36 217 124 274
rect 36 171 49 217
rect 95 171 124 217
rect 36 156 124 171
rect 244 217 348 274
rect 244 171 273 217
rect 319 171 348 217
rect 244 156 348 171
rect 468 156 516 274
rect 636 217 740 274
rect 636 171 665 217
rect 711 171 740 217
rect 636 156 740 171
rect 860 156 908 274
rect 1028 156 1152 274
rect 1229 265 1242 311
rect 1288 265 1317 311
rect 1229 166 1317 265
rect 1437 225 1541 324
rect 1437 179 1466 225
rect 1512 179 1541 225
rect 1437 166 1541 179
rect 1661 300 1749 324
rect 3601 313 3681 324
rect 1661 254 1690 300
rect 1736 254 1749 300
rect 1661 166 1749 254
rect 1825 254 1913 313
rect 1825 208 1838 254
rect 1884 208 1913 254
rect 1825 195 1913 208
rect 2033 254 2137 313
rect 2033 208 2062 254
rect 2108 208 2137 254
rect 2033 195 2137 208
rect 2257 195 2305 313
rect 2425 195 2477 313
rect 2597 254 2701 313
rect 2597 208 2626 254
rect 2672 208 2701 254
rect 2597 195 2701 208
rect 2821 300 2925 313
rect 2821 254 2850 300
rect 2896 254 2925 300
rect 2821 195 2925 254
rect 3045 300 3153 313
rect 3045 254 3078 300
rect 3124 254 3153 300
rect 3045 195 3153 254
rect 3273 300 3421 313
rect 3273 254 3346 300
rect 3392 254 3421 300
rect 3273 195 3421 254
rect 3541 254 3681 313
rect 3541 208 3570 254
rect 3616 208 3681 254
rect 3541 195 3681 208
rect 1088 122 1152 156
rect 1088 110 1160 122
rect 1088 64 1101 110
rect 1147 64 1160 110
rect 1088 51 1160 64
rect 3601 124 3681 195
rect 3801 124 3849 324
rect 3969 311 4057 324
rect 3969 171 3998 311
rect 4044 171 4057 311
rect 3969 124 4057 171
rect 4148 221 4236 332
rect 4148 81 4161 221
rect 4207 81 4236 221
rect 4148 68 4236 81
rect 4356 319 4460 332
rect 4356 179 4385 319
rect 4431 179 4460 319
rect 4356 68 4460 179
rect 4580 221 4668 332
rect 4580 81 4609 221
rect 4655 81 4668 221
rect 4580 68 4668 81
<< mvpdiff >>
rect 56 839 144 852
rect 56 699 69 839
rect 115 699 144 839
rect 56 652 144 699
rect 244 839 348 852
rect 244 699 273 839
rect 319 699 348 839
rect 244 652 348 699
rect 448 652 496 852
rect 596 839 740 852
rect 596 699 625 839
rect 671 699 740 839
rect 596 652 740 699
rect 840 652 888 852
rect 988 839 1076 852
rect 988 699 1017 839
rect 1063 699 1076 839
rect 988 652 1076 699
rect 1229 639 1317 856
rect 1229 593 1242 639
rect 1288 593 1317 639
rect 1229 580 1317 593
rect 1417 834 1521 856
rect 1417 788 1446 834
rect 1492 788 1521 834
rect 1417 580 1521 788
rect 1621 639 1709 856
rect 3601 953 3673 966
rect 3601 907 3614 953
rect 3660 939 3673 953
rect 3660 907 3733 939
rect 3601 852 3733 907
rect 1781 839 1869 852
rect 1781 699 1794 839
rect 1840 699 1869 839
rect 1781 652 1869 699
rect 1969 839 2073 852
rect 1969 699 1998 839
rect 2044 699 2073 839
rect 1969 652 2073 699
rect 2173 839 2277 852
rect 2173 699 2202 839
rect 2248 699 2277 839
rect 2173 652 2277 699
rect 2377 745 2481 852
rect 2377 699 2406 745
rect 2452 699 2481 745
rect 2377 652 2481 699
rect 2581 839 2669 852
rect 2581 699 2610 839
rect 2656 699 2669 839
rect 2581 652 2669 699
rect 2741 839 2829 852
rect 2741 699 2754 839
rect 2800 699 2829 839
rect 2741 652 2829 699
rect 2929 839 3033 852
rect 2929 699 2958 839
rect 3004 699 3033 839
rect 2929 652 3033 699
rect 3133 839 3237 852
rect 3133 699 3162 839
rect 3208 699 3237 839
rect 3133 652 3237 699
rect 3337 745 3441 852
rect 3337 699 3366 745
rect 3412 699 3441 745
rect 3337 652 3441 699
rect 3541 663 3733 852
rect 3833 745 3937 939
rect 3833 699 3862 745
rect 3908 699 3937 745
rect 3833 663 3937 699
rect 4037 839 4246 939
rect 4037 699 4066 839
rect 4112 699 4246 839
rect 4037 663 4246 699
rect 3541 652 3621 663
rect 1621 593 1650 639
rect 1696 593 1709 639
rect 1621 580 1709 593
rect 4166 573 4246 663
rect 4346 839 4454 939
rect 4346 699 4379 839
rect 4425 699 4454 839
rect 4346 573 4454 699
rect 4554 839 4642 939
rect 4554 699 4583 839
rect 4629 699 4642 839
rect 4554 573 4642 699
<< mvndiffc >>
rect 49 171 95 217
rect 273 171 319 217
rect 665 171 711 217
rect 1242 265 1288 311
rect 1466 179 1512 225
rect 1690 254 1736 300
rect 1838 208 1884 254
rect 2062 208 2108 254
rect 2626 208 2672 254
rect 2850 254 2896 300
rect 3078 254 3124 300
rect 3346 254 3392 300
rect 3570 208 3616 254
rect 1101 64 1147 110
rect 3998 171 4044 311
rect 4161 81 4207 221
rect 4385 179 4431 319
rect 4609 81 4655 221
<< mvpdiffc >>
rect 69 699 115 839
rect 273 699 319 839
rect 625 699 671 839
rect 1017 699 1063 839
rect 1242 593 1288 639
rect 1446 788 1492 834
rect 3614 907 3660 953
rect 1794 699 1840 839
rect 1998 699 2044 839
rect 2202 699 2248 839
rect 2406 699 2452 745
rect 2610 699 2656 839
rect 2754 699 2800 839
rect 2958 699 3004 839
rect 3162 699 3208 839
rect 3366 699 3412 745
rect 3862 699 3908 745
rect 4066 699 4112 839
rect 1650 593 1696 639
rect 4379 699 4425 839
rect 4583 699 4629 839
<< polysilicon >>
rect 144 944 988 984
rect 144 852 244 944
rect 348 852 448 896
rect 496 852 596 896
rect 740 852 840 896
rect 888 852 988 944
rect 1521 944 3133 984
rect 1317 856 1417 900
rect 1521 856 1621 944
rect 144 547 244 652
rect 144 501 157 547
rect 203 501 244 547
rect 144 318 244 501
rect 124 274 244 318
rect 348 539 448 652
rect 348 493 361 539
rect 407 493 448 539
rect 348 318 448 493
rect 496 547 596 652
rect 496 501 509 547
rect 555 501 596 547
rect 496 488 596 501
rect 740 547 840 652
rect 888 608 988 652
rect 1869 852 1969 896
rect 2073 852 2173 944
rect 2277 852 2377 896
rect 2481 852 2581 896
rect 2829 852 2929 896
rect 3033 852 3133 944
rect 3733 939 3833 983
rect 3937 939 4037 983
rect 4246 939 4346 983
rect 4454 939 4554 983
rect 3237 852 3337 896
rect 3441 852 3541 896
rect 740 501 753 547
rect 799 501 840 547
rect 740 318 840 501
rect 908 547 1028 560
rect 908 501 941 547
rect 987 501 1028 547
rect 348 274 468 318
rect 516 274 636 318
rect 740 274 860 318
rect 908 274 1028 501
rect 1317 547 1417 580
rect 1317 501 1330 547
rect 1376 501 1417 547
rect 1317 368 1417 501
rect 1521 547 1621 580
rect 1521 501 1534 547
rect 1580 501 1621 547
rect 1521 488 1621 501
rect 1541 368 1621 488
rect 1869 550 1969 652
rect 2073 608 2173 652
rect 2277 608 2377 652
rect 1869 547 2257 550
rect 1869 501 1882 547
rect 1928 501 2257 547
rect 1869 478 2257 501
rect 2137 392 2257 478
rect 1317 324 1437 368
rect 1541 324 1661 368
rect 1913 313 2033 357
rect 2137 346 2178 392
rect 2224 346 2257 392
rect 2137 313 2257 346
rect 2305 455 2377 608
rect 2305 409 2318 455
rect 2364 409 2377 455
rect 2305 357 2377 409
rect 2481 357 2581 652
rect 2829 608 2929 652
rect 3033 608 3133 652
rect 2829 560 2869 608
rect 2701 547 2869 560
rect 2701 501 2734 547
rect 2780 501 2869 547
rect 2701 488 2869 501
rect 2925 547 3045 560
rect 2925 501 2958 547
rect 3004 501 3045 547
rect 2305 313 2425 357
rect 2477 313 2597 357
rect 2701 313 2821 488
rect 2925 313 3045 501
rect 3093 468 3133 608
rect 3237 547 3337 652
rect 3237 501 3254 547
rect 3300 501 3337 547
rect 3237 488 3337 501
rect 3441 547 3541 652
rect 3733 619 3833 663
rect 3733 560 3801 619
rect 3937 568 4037 663
rect 3441 501 3482 547
rect 3528 501 3541 547
rect 3093 396 3193 468
rect 3153 357 3193 396
rect 3441 357 3541 501
rect 3153 313 3273 357
rect 3421 313 3541 357
rect 3681 547 3801 560
rect 3681 501 3722 547
rect 3768 501 3801 547
rect 3681 324 3801 501
rect 3849 562 4037 568
rect 3849 516 3954 562
rect 4000 516 4037 562
rect 3849 503 4037 516
rect 3849 324 3969 503
rect 4246 464 4346 573
rect 4454 464 4554 573
rect 4246 456 4554 464
rect 4047 443 4554 456
rect 4047 397 4060 443
rect 4106 397 4554 443
rect 4047 392 4554 397
rect 4047 384 4118 392
rect 4236 332 4356 392
rect 4460 376 4554 392
rect 4460 332 4580 376
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1317 122 1437 166
rect 124 24 636 64
rect 1541 96 1661 166
rect 1913 96 2033 195
rect 2137 151 2257 195
rect 2305 151 2425 195
rect 1541 24 2033 96
rect 2477 64 2597 195
rect 2701 151 2821 195
rect 2925 151 3045 195
rect 3153 151 3273 195
rect 3421 151 3541 195
rect 3681 64 3801 124
rect 3849 80 3969 124
rect 2477 24 3801 64
rect 4236 24 4356 68
rect 4460 24 4580 68
<< polycontact >>
rect 157 501 203 547
rect 361 493 407 539
rect 509 501 555 547
rect 753 501 799 547
rect 941 501 987 547
rect 1330 501 1376 547
rect 1534 501 1580 547
rect 1882 501 1928 547
rect 2178 346 2224 392
rect 2318 409 2364 455
rect 2734 501 2780 547
rect 2958 501 3004 547
rect 3254 501 3300 547
rect 3482 501 3528 547
rect 3722 501 3768 547
rect 3954 516 4000 562
rect 4060 397 4106 443
<< metal1 >>
rect 0 953 4704 1098
rect 0 918 3614 953
rect 69 839 115 850
rect 69 642 115 699
rect 273 839 319 918
rect 273 688 319 699
rect 625 839 971 850
rect 671 804 971 839
rect 625 688 671 699
rect 69 596 555 642
rect 142 501 157 547
rect 203 501 306 547
rect 142 466 306 501
rect 354 539 430 550
rect 354 493 361 539
rect 407 493 430 539
rect 354 366 430 493
rect 509 547 555 596
rect 509 320 555 501
rect 702 547 799 654
rect 925 642 971 804
rect 1017 839 1063 918
rect 1435 834 1503 918
rect 1435 788 1446 834
rect 1492 788 1503 834
rect 1794 839 1840 850
rect 1017 688 1063 699
rect 1109 699 1794 742
rect 1109 696 1840 699
rect 1109 642 1155 696
rect 1794 688 1840 696
rect 1998 839 2044 850
rect 925 596 1155 642
rect 1650 639 1707 650
rect 1231 593 1242 639
rect 1288 593 1518 639
rect 1472 547 1518 593
rect 1696 593 1707 639
rect 1650 547 1707 593
rect 1998 583 2044 699
rect 2202 839 2248 850
rect 2202 642 2248 699
rect 2406 745 2452 918
rect 2406 688 2452 699
rect 2610 839 2656 850
rect 2610 642 2656 699
rect 2754 839 2800 918
rect 3660 918 4704 953
rect 3614 896 3660 907
rect 2754 688 2800 699
rect 2958 839 3004 850
rect 2958 650 3004 699
rect 2202 596 2656 642
rect 2850 604 3004 650
rect 3162 839 4000 850
rect 3208 804 4000 839
rect 1998 547 2107 583
rect 702 501 753 547
rect 702 466 799 501
rect 930 501 941 547
rect 987 501 998 547
rect 930 320 998 501
rect 1262 501 1330 547
rect 1376 501 1426 547
rect 1262 466 1426 501
rect 1472 501 1534 547
rect 1580 501 1591 547
rect 1650 504 1882 547
rect 1690 501 1882 504
rect 1928 501 1939 547
rect 1998 537 2734 547
rect 2062 501 2734 537
rect 2780 501 2791 547
rect 1472 420 1518 501
rect 49 274 998 320
rect 1242 374 1518 420
rect 1242 311 1288 374
rect 49 217 95 274
rect 1242 254 1288 265
rect 1334 282 1644 328
rect 49 160 95 171
rect 273 217 319 228
rect 273 90 319 171
rect 654 171 665 217
rect 711 213 722 217
rect 711 208 1221 213
rect 1334 208 1380 282
rect 711 171 1380 208
rect 654 167 1380 171
rect 1200 162 1380 167
rect 1466 225 1512 236
rect 1101 110 1147 121
rect 0 64 1101 90
rect 1466 90 1512 179
rect 1598 197 1644 282
rect 1690 300 1736 501
rect 1690 243 1736 254
rect 1838 254 1884 265
rect 1838 197 1884 208
rect 2062 254 2108 501
rect 2850 455 2896 604
rect 2307 409 2318 455
rect 2364 409 2896 455
rect 2167 346 2178 392
rect 2224 363 2235 392
rect 2224 346 2804 363
rect 2167 317 2804 346
rect 2062 197 2108 208
rect 2626 254 2672 265
rect 1598 151 1884 197
rect 2626 90 2672 208
rect 2758 197 2804 317
rect 2850 300 2896 409
rect 2850 243 2896 254
rect 2958 547 3004 558
rect 2958 197 3004 501
rect 3162 311 3208 699
rect 3346 745 3412 756
rect 3346 699 3366 745
rect 3078 300 3208 311
rect 3124 254 3208 300
rect 3078 243 3208 254
rect 3254 547 3300 558
rect 3254 197 3300 501
rect 3346 300 3412 699
rect 3482 745 3908 756
rect 3482 710 3862 745
rect 3482 547 3528 710
rect 3614 578 3778 654
rect 3482 490 3528 501
rect 3722 547 3778 578
rect 3768 501 3778 547
rect 3722 354 3778 501
rect 3862 443 3908 699
rect 3954 562 4000 804
rect 4066 839 4112 918
rect 4066 688 4112 699
rect 4379 839 4450 850
rect 4425 699 4450 839
rect 3954 505 4000 516
rect 3862 397 4060 443
rect 4106 397 4117 443
rect 3392 254 3412 300
rect 3998 311 4044 397
rect 3346 243 3412 254
rect 3570 254 3616 265
rect 2758 151 3300 197
rect 3570 90 3616 208
rect 4379 319 4450 699
rect 4583 839 4629 918
rect 4583 688 4629 699
rect 3998 160 4044 171
rect 4161 221 4207 232
rect 1147 81 4161 90
rect 4379 179 4385 319
rect 4431 179 4450 319
rect 4379 168 4450 179
rect 4609 221 4655 232
rect 4207 81 4609 90
rect 4655 81 4704 90
rect 1147 64 4704 81
rect 0 -90 4704 64
<< labels >>
flabel metal1 s 1262 466 1426 547 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 702 466 799 654 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4379 168 4450 850 0 FreeSans 200 0 0 0 Q
port 6 nsew default output
flabel metal1 s 3614 578 3778 654 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 142 466 306 547 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 354 366 430 550 0 FreeSans 200 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 918 4704 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 3570 236 3616 265 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 3722 354 3778 578 1 RN
port 2 nsew default input
rlabel metal1 s 4583 896 4629 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4066 896 4112 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3614 896 3660 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2754 896 2800 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2406 896 2452 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1435 896 1503 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 896 1063 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 273 896 319 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4583 788 4629 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4066 788 4112 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2754 788 2800 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2406 788 2452 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1435 788 1503 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 788 1063 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 273 788 319 896 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4583 688 4629 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4066 688 4112 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2754 688 2800 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2406 688 2452 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1017 688 1063 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 273 688 319 788 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2626 236 2672 265 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3570 232 3616 236 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2626 232 2672 236 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1466 232 1512 236 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4609 228 4655 232 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4161 228 4207 232 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3570 228 3616 232 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2626 228 2672 232 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1466 228 1512 232 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4609 121 4655 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4161 121 4207 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3570 121 3616 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2626 121 2672 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1466 121 1512 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 121 319 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4609 90 4655 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4161 90 4207 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3570 90 3616 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2626 90 2672 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1466 90 1512 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1101 90 1147 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 121 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4704 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 1008
string GDS_END 347706
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 336698
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
