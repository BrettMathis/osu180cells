magic
tech gf180mcuC
magscale 1 5
timestamp 1675314274
<< obsm1 >>
rect 120 2430 89880 57225
<< metal2 >>
rect 5768 59600 5824 60000
rect 16968 59600 17024 60000
rect 28168 59600 28224 60000
rect 39368 59600 39424 60000
rect 50568 59600 50624 60000
rect 61768 59600 61824 60000
rect 72968 59600 73024 60000
rect 84168 59600 84224 60000
rect 5768 0 5824 400
rect 16968 0 17024 400
rect 28168 0 28224 400
rect 39368 0 39424 400
rect 50568 0 50624 400
rect 61768 0 61824 400
rect 72968 0 73024 400
rect 84168 0 84224 400
<< obsm2 >>
rect 1686 59570 5738 59600
rect 5854 59570 16938 59600
rect 17054 59570 28138 59600
rect 28254 59570 39338 59600
rect 39454 59570 50538 59600
rect 50654 59570 61738 59600
rect 61854 59570 72938 59600
rect 73054 59570 84138 59600
rect 84254 59570 89810 59600
rect 1686 430 89810 59570
rect 1686 350 5738 430
rect 5854 350 16938 430
rect 17054 350 28138 430
rect 28254 350 39338 430
rect 39454 350 50538 430
rect 50654 350 61738 430
rect 61854 350 72938 430
rect 73054 350 84138 430
rect 84254 350 89810 430
<< metal3 >>
rect 89600 56000 90000 56056
rect 89600 48552 90000 48608
rect 89600 41104 90000 41160
rect 89600 33656 90000 33712
rect 89600 26208 90000 26264
rect 89600 18760 90000 18816
rect 89600 11312 90000 11368
rect 89600 3864 90000 3920
<< obsm3 >>
rect 1681 56086 89815 57209
rect 1681 55970 89570 56086
rect 1681 48638 89815 55970
rect 1681 48522 89570 48638
rect 1681 41190 89815 48522
rect 1681 41074 89570 41190
rect 1681 33742 89815 41074
rect 1681 33626 89570 33742
rect 1681 26294 89815 33626
rect 1681 26178 89570 26294
rect 1681 18846 89815 26178
rect 1681 18730 89570 18846
rect 1681 11398 89815 18730
rect 1681 11282 89570 11398
rect 1681 3950 89815 11282
rect 1681 3834 89570 3950
rect 1681 2446 89815 3834
<< metal4 >>
rect 1672 2430 1832 57225
rect 9352 2430 9512 57225
rect 17032 2430 17192 57225
rect 24712 2430 24872 57225
rect 32392 2430 32552 57225
rect 40072 2430 40232 57225
rect 47752 2430 47912 57225
rect 55432 2430 55592 57225
rect 63112 2430 63272 57225
rect 70792 2430 70952 57225
rect 78472 2430 78632 57225
rect 86152 2430 86312 57225
<< obsm4 >>
rect 39158 24201 39410 25611
<< labels >>
rlabel metal2 s 5768 0 5824 400 6 a_in[0]
port 1 nsew signal input
rlabel metal2 s 16968 0 17024 400 6 a_in[1]
port 2 nsew signal input
rlabel metal2 s 28168 0 28224 400 6 a_in[2]
port 3 nsew signal input
rlabel metal2 s 39368 0 39424 400 6 a_in[3]
port 4 nsew signal input
rlabel metal2 s 50568 0 50624 400 6 a_in[4]
port 5 nsew signal input
rlabel metal2 s 61768 0 61824 400 6 a_in[5]
port 6 nsew signal input
rlabel metal2 s 72968 0 73024 400 6 a_in[6]
port 7 nsew signal input
rlabel metal2 s 84168 0 84224 400 6 a_in[7]
port 8 nsew signal input
rlabel metal3 s 89600 3864 90000 3920 6 b_in[0]
port 9 nsew signal input
rlabel metal3 s 89600 11312 90000 11368 6 b_in[1]
port 10 nsew signal input
rlabel metal3 s 89600 18760 90000 18816 6 b_in[2]
port 11 nsew signal input
rlabel metal3 s 89600 26208 90000 26264 6 b_in[3]
port 12 nsew signal input
rlabel metal3 s 89600 33656 90000 33712 6 b_in[4]
port 13 nsew signal input
rlabel metal3 s 89600 41104 90000 41160 6 b_in[5]
port 14 nsew signal input
rlabel metal3 s 89600 48552 90000 48608 6 b_in[6]
port 15 nsew signal input
rlabel metal3 s 89600 56000 90000 56056 6 b_in[7]
port 16 nsew signal input
rlabel metal2 s 5768 59600 5824 60000 6 sum[0]
port 17 nsew signal output
rlabel metal2 s 16968 59600 17024 60000 6 sum[1]
port 18 nsew signal output
rlabel metal2 s 28168 59600 28224 60000 6 sum[2]
port 19 nsew signal output
rlabel metal2 s 39368 59600 39424 60000 6 sum[3]
port 20 nsew signal output
rlabel metal2 s 50568 59600 50624 60000 6 sum[4]
port 21 nsew signal output
rlabel metal2 s 61768 59600 61824 60000 6 sum[5]
port 22 nsew signal output
rlabel metal2 s 72968 59600 73024 60000 6 sum[6]
port 23 nsew signal output
rlabel metal2 s 84168 59600 84224 60000 6 sum[7]
port 24 nsew signal output
rlabel metal4 s 1672 2430 1832 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 17032 2430 17192 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 32392 2430 32552 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 47752 2430 47912 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 63112 2430 63272 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 78472 2430 78632 57225 6 vdd
port 25 nsew power bidirectional
rlabel metal4 s 9352 2430 9512 57225 6 vss
port 26 nsew ground bidirectional
rlabel metal4 s 24712 2430 24872 57225 6 vss
port 26 nsew ground bidirectional
rlabel metal4 s 40072 2430 40232 57225 6 vss
port 26 nsew ground bidirectional
rlabel metal4 s 55432 2430 55592 57225 6 vss
port 26 nsew ground bidirectional
rlabel metal4 s 70792 2430 70952 57225 6 vss
port 26 nsew ground bidirectional
rlabel metal4 s 86152 2430 86312 57225 6 vss
port 26 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4796970
string GDS_FILE /home/brettcm/caravel/main/osu180cells/openlane/adder/runs/23_02_01_23_03/results/signoff/adder.magic.gds
string GDS_START 64376
<< end >>

