magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 111 164 123
rect 11 70 16 111
rect 28 65 33 104
rect 45 70 50 111
rect 62 65 67 104
rect 79 70 84 111
rect 96 65 101 104
rect 113 70 118 111
rect 130 76 135 104
rect 130 70 143 76
rect 148 70 153 111
rect 130 65 135 70
rect 28 60 135 65
rect 8 44 18 50
rect 28 46 33 60
rect 62 46 67 60
rect 96 46 101 60
rect 130 46 135 60
rect 28 41 135 46
rect 11 12 16 36
rect 28 19 33 41
rect 45 12 50 36
rect 62 19 67 41
rect 79 12 84 36
rect 96 19 101 41
rect 113 12 118 36
rect 130 19 135 41
rect 147 12 152 36
rect 0 0 164 12
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 134 76 142 77
rect 133 70 143 76
rect 134 69 142 70
rect 8 43 18 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
<< labels >>
rlabel metal2 s 8 43 18 51 6 A
port 1 nsew signal input
rlabel metal1 s 8 44 18 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 45 70 50 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 79 70 84 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 113 70 118 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 148 70 153 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 164 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 0 50 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 79 0 84 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 113 0 118 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 147 0 152 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 164 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 134 69 142 77 6 Y
port 2 nsew signal output
rlabel metal2 s 133 70 143 76 6 Y
port 2 nsew signal output
rlabel metal1 s 28 19 33 104 6 Y
port 2 nsew signal output
rlabel metal1 s 62 19 67 104 6 Y
port 2 nsew signal output
rlabel metal1 s 96 19 101 104 6 Y
port 2 nsew signal output
rlabel metal1 s 28 41 135 46 6 Y
port 2 nsew signal output
rlabel metal1 s 28 60 135 65 6 Y
port 2 nsew signal output
rlabel metal1 s 130 19 135 104 6 Y
port 2 nsew signal output
rlabel metal1 s 130 70 143 76 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 164 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 382306
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 369858
<< end >>
