magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -169 461 170 502
rect -169 409 -132 461
rect -80 409 80 461
rect 132 409 170 461
rect -169 244 170 409
rect -169 192 -132 244
rect -80 192 80 244
rect 132 192 170 244
rect -169 26 170 192
rect -169 -26 -132 26
rect -80 -26 80 26
rect 132 -26 170 26
rect -169 -192 170 -26
rect -169 -244 -132 -192
rect -80 -244 80 -192
rect 132 -244 170 -192
rect -169 -409 170 -244
rect -169 -461 -132 -409
rect -80 -461 80 -409
rect 132 -461 170 -409
rect -169 -502 170 -461
<< via1 >>
rect -132 409 -80 461
rect 80 409 132 461
rect -132 192 -80 244
rect 80 192 132 244
rect -132 -26 -80 26
rect 80 -26 132 26
rect -132 -244 -80 -192
rect 80 -244 132 -192
rect -132 -461 -80 -409
rect 80 -461 132 -409
<< metal2 >>
rect -169 461 170 502
rect -169 409 -132 461
rect -80 409 80 461
rect 132 409 170 461
rect -169 244 170 409
rect -169 192 -132 244
rect -80 192 80 244
rect 132 192 170 244
rect -169 26 170 192
rect -169 -26 -132 26
rect -80 -26 80 26
rect 132 -26 170 26
rect -169 -192 170 -26
rect -169 -244 -132 -192
rect -80 -244 80 -192
rect 132 -244 170 -192
rect -169 -409 170 -244
rect -169 -461 -132 -409
rect -80 -461 80 -409
rect 132 -461 170 -409
rect -169 -502 170 -461
<< properties >>
string GDS_END 623054
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 622282
<< end >>
