magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 568 35
<< polysilicon >>
rect -31 227 89 300
rect 193 227 313 300
rect -31 -74 89 -1
rect 193 -74 313 -1
use pmos_5p0431059054873_128x8m81  pmos_5p0431059054873_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 348
<< properties >>
string GDS_END 312190
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 311748
<< end >>
