magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 2268 89 2341
rect -31 -73 89 -1
use nmos_5p0431059130205_512x8m81  nmos_5p0431059130205_512x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 2312
<< properties >>
string GDS_END 256508
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 256258
<< end >>
