magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -221 -1452 221 1452
<< nsubdiff >>
rect -77 1247 78 1304
rect -77 1201 -23 1247
rect 23 1201 78 1247
rect -77 1084 78 1201
rect -77 1038 -23 1084
rect 23 1038 78 1084
rect -77 921 78 1038
rect -77 875 -23 921
rect 23 875 78 921
rect -77 758 78 875
rect -77 712 -23 758
rect 23 712 78 758
rect -77 595 78 712
rect -77 549 -23 595
rect 23 549 78 595
rect -77 431 78 549
rect -77 385 -23 431
rect 23 385 78 431
rect -77 268 78 385
rect -77 222 -23 268
rect 23 222 78 268
rect -77 105 78 222
rect -77 59 -23 105
rect 23 59 78 105
rect -77 -59 78 59
rect -77 -105 -23 -59
rect 23 -105 78 -59
rect -77 -222 78 -105
rect -77 -268 -23 -222
rect 23 -268 78 -222
rect -77 -385 78 -268
rect -77 -431 -23 -385
rect 23 -431 78 -385
rect -77 -549 78 -431
rect -77 -595 -23 -549
rect 23 -595 78 -549
rect -77 -712 78 -595
rect -77 -758 -23 -712
rect 23 -758 78 -712
rect -77 -875 78 -758
rect -77 -921 -23 -875
rect 23 -921 78 -875
rect -77 -1038 78 -921
rect -77 -1084 -23 -1038
rect 23 -1084 78 -1038
rect -77 -1201 78 -1084
rect -77 -1247 -23 -1201
rect 23 -1247 78 -1201
rect -77 -1305 78 -1247
<< nsubdiffcont >>
rect -23 1201 23 1247
rect -23 1038 23 1084
rect -23 875 23 921
rect -23 712 23 758
rect -23 549 23 595
rect -23 385 23 431
rect -23 222 23 268
rect -23 59 23 105
rect -23 -105 23 -59
rect -23 -268 23 -222
rect -23 -431 23 -385
rect -23 -595 23 -549
rect -23 -758 23 -712
rect -23 -921 23 -875
rect -23 -1084 23 -1038
rect -23 -1247 23 -1201
<< metal1 >>
rect -58 1247 58 1284
rect -58 1201 -23 1247
rect 23 1201 58 1247
rect -58 1084 58 1201
rect -58 1038 -23 1084
rect 23 1038 58 1084
rect -58 921 58 1038
rect -58 875 -23 921
rect 23 875 58 921
rect -58 758 58 875
rect -58 712 -23 758
rect 23 712 58 758
rect -58 595 58 712
rect -58 549 -23 595
rect 23 549 58 595
rect -58 431 58 549
rect -58 385 -23 431
rect 23 385 58 431
rect -58 268 58 385
rect -58 222 -23 268
rect 23 222 58 268
rect -58 105 58 222
rect -58 59 -23 105
rect 23 59 58 105
rect -58 -59 58 59
rect -58 -105 -23 -59
rect 23 -105 58 -59
rect -58 -222 58 -105
rect -58 -268 -23 -222
rect 23 -268 58 -222
rect -58 -385 58 -268
rect -58 -431 -23 -385
rect 23 -431 58 -385
rect -58 -549 58 -431
rect -58 -595 -23 -549
rect 23 -595 58 -549
rect -58 -712 58 -595
rect -58 -758 -23 -712
rect 23 -758 58 -712
rect -58 -875 58 -758
rect -58 -921 -23 -875
rect 23 -921 58 -875
rect -58 -1038 58 -921
rect -58 -1084 -23 -1038
rect 23 -1084 58 -1038
rect -58 -1201 58 -1084
rect -58 -1247 -23 -1201
rect 23 -1247 58 -1201
rect -58 -1284 58 -1247
<< properties >>
string GDS_END 539548
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 538264
<< end >>
