magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3894 1094
<< pwell >>
rect -86 -86 3894 453
<< mvnmos >>
rect 124 156 244 316
rect 484 156 604 316
rect 708 156 828 316
rect 932 156 1052 316
rect 1156 156 1276 316
rect 1380 156 1500 316
rect 1851 156 1971 316
rect 2075 156 2195 316
rect 2443 156 2563 316
rect 2667 156 2787 316
rect 2891 156 3011 316
rect 3115 156 3235 316
rect 3339 156 3459 316
rect 3563 156 3683 316
<< mvpmos >>
rect 144 596 244 852
rect 416 596 516 852
rect 658 596 758 852
rect 884 596 984 852
rect 1176 596 1276 852
rect 1380 596 1480 852
rect 1861 596 1961 852
rect 2107 596 2207 852
rect 2471 596 2571 852
rect 2687 596 2787 852
rect 2905 596 3005 852
rect 3109 596 3209 852
rect 3339 596 3439 852
rect 3563 596 3663 852
<< mvndiff >>
rect 36 297 124 316
rect 36 251 49 297
rect 95 251 124 297
rect 36 156 124 251
rect 244 297 484 316
rect 244 251 273 297
rect 319 251 484 297
rect 244 156 484 251
rect 604 297 708 316
rect 604 251 633 297
rect 679 251 708 297
rect 604 156 708 251
rect 828 297 932 316
rect 828 251 857 297
rect 903 251 932 297
rect 828 156 932 251
rect 1052 297 1156 316
rect 1052 251 1081 297
rect 1127 251 1156 297
rect 1052 156 1156 251
rect 1276 297 1380 316
rect 1276 251 1305 297
rect 1351 251 1380 297
rect 1276 156 1380 251
rect 1500 297 1588 316
rect 1500 251 1529 297
rect 1575 251 1588 297
rect 1500 156 1588 251
rect 1715 299 1851 316
rect 1715 253 1728 299
rect 1774 253 1851 299
rect 1715 156 1851 253
rect 1971 297 2075 316
rect 1971 251 2000 297
rect 2046 251 2075 297
rect 1971 156 2075 251
rect 2195 297 2283 316
rect 2195 251 2224 297
rect 2270 251 2283 297
rect 2195 156 2283 251
rect 2355 297 2443 316
rect 2355 251 2368 297
rect 2414 251 2443 297
rect 2355 156 2443 251
rect 2563 297 2667 316
rect 2563 251 2592 297
rect 2638 251 2667 297
rect 2563 156 2667 251
rect 2787 297 2891 316
rect 2787 251 2816 297
rect 2862 251 2891 297
rect 2787 156 2891 251
rect 3011 297 3115 316
rect 3011 251 3040 297
rect 3086 251 3115 297
rect 3011 156 3115 251
rect 3235 297 3339 316
rect 3235 251 3264 297
rect 3310 251 3339 297
rect 3235 156 3339 251
rect 3459 297 3563 316
rect 3459 251 3488 297
rect 3534 251 3563 297
rect 3459 156 3563 251
rect 3683 297 3771 316
rect 3683 251 3712 297
rect 3758 251 3771 297
rect 3683 156 3771 251
<< mvpdiff >>
rect 1044 871 1116 884
rect 1044 852 1057 871
rect 37 767 144 852
rect 37 627 50 767
rect 96 627 144 767
rect 37 596 144 627
rect 244 767 416 852
rect 244 627 273 767
rect 319 627 416 767
rect 244 596 416 627
rect 516 767 658 852
rect 516 627 545 767
rect 591 627 658 767
rect 516 596 658 627
rect 758 665 884 852
rect 758 619 809 665
rect 855 619 884 665
rect 758 596 884 619
rect 984 825 1057 852
rect 1103 852 1116 871
rect 1103 825 1176 852
rect 984 596 1176 825
rect 1276 665 1380 852
rect 1276 619 1305 665
rect 1351 619 1380 665
rect 1276 596 1380 619
rect 1480 767 1568 852
rect 1480 627 1509 767
rect 1555 627 1568 767
rect 1480 596 1568 627
rect 1742 767 1861 852
rect 1742 627 1755 767
rect 1801 627 1861 767
rect 1742 596 1861 627
rect 1961 767 2107 852
rect 1961 627 1990 767
rect 2036 627 2107 767
rect 1961 596 2107 627
rect 2207 767 2295 852
rect 2207 627 2236 767
rect 2282 627 2295 767
rect 2207 596 2295 627
rect 2383 767 2471 852
rect 2383 627 2396 767
rect 2442 627 2471 767
rect 2383 596 2471 627
rect 2571 767 2687 852
rect 2571 627 2600 767
rect 2646 627 2687 767
rect 2571 596 2687 627
rect 2787 767 2905 852
rect 2787 627 2816 767
rect 2862 627 2905 767
rect 2787 596 2905 627
rect 3005 767 3109 852
rect 3005 627 3034 767
rect 3080 627 3109 767
rect 3005 596 3109 627
rect 3209 767 3339 852
rect 3209 627 3238 767
rect 3284 627 3339 767
rect 3209 596 3339 627
rect 3439 767 3563 852
rect 3439 627 3468 767
rect 3514 627 3563 767
rect 3439 596 3563 627
rect 3663 767 3751 852
rect 3663 627 3692 767
rect 3738 627 3751 767
rect 3663 596 3751 627
<< mvndiffc >>
rect 49 251 95 297
rect 273 251 319 297
rect 633 251 679 297
rect 857 251 903 297
rect 1081 251 1127 297
rect 1305 251 1351 297
rect 1529 251 1575 297
rect 1728 253 1774 299
rect 2000 251 2046 297
rect 2224 251 2270 297
rect 2368 251 2414 297
rect 2592 251 2638 297
rect 2816 251 2862 297
rect 3040 251 3086 297
rect 3264 251 3310 297
rect 3488 251 3534 297
rect 3712 251 3758 297
<< mvpdiffc >>
rect 50 627 96 767
rect 273 627 319 767
rect 545 627 591 767
rect 809 619 855 665
rect 1057 825 1103 871
rect 1305 619 1351 665
rect 1509 627 1555 767
rect 1755 627 1801 767
rect 1990 627 2036 767
rect 2236 627 2282 767
rect 2396 627 2442 767
rect 2600 627 2646 767
rect 2816 627 2862 767
rect 3034 627 3080 767
rect 3238 627 3284 767
rect 3468 627 3514 767
rect 3692 627 3738 767
<< polysilicon >>
rect 658 944 3005 984
rect 144 852 244 896
rect 416 852 516 896
rect 658 852 758 944
rect 884 852 984 896
rect 1176 852 1276 896
rect 1380 852 1480 896
rect 1861 852 1961 896
rect 2107 852 2207 896
rect 2471 852 2571 896
rect 2687 852 2787 896
rect 2905 852 3005 944
rect 3109 944 3663 984
rect 3109 852 3209 944
rect 3339 852 3439 896
rect 3563 852 3663 944
rect 144 467 244 596
rect 144 421 157 467
rect 203 421 244 467
rect 144 360 244 421
rect 416 467 516 596
rect 658 536 758 596
rect 416 421 457 467
rect 503 421 516 467
rect 416 408 516 421
rect 564 502 758 536
rect 564 496 680 502
rect 564 360 604 496
rect 884 467 984 596
rect 704 441 828 454
rect 704 395 717 441
rect 763 395 828 441
rect 884 421 925 467
rect 971 421 984 467
rect 884 408 984 421
rect 704 382 828 395
rect 124 316 244 360
rect 484 316 604 360
rect 708 316 828 382
rect 932 360 984 408
rect 1176 448 1276 596
rect 1380 467 1480 596
rect 1380 448 1421 467
rect 1176 421 1421 448
rect 1467 421 1480 467
rect 1861 536 1961 596
rect 2107 555 2207 596
rect 1861 464 2059 536
rect 2107 509 2120 555
rect 2166 536 2207 555
rect 2471 552 2571 596
rect 2471 536 2563 552
rect 2166 509 2563 536
rect 2107 496 2563 509
rect 1176 376 1480 421
rect 2019 448 2059 464
rect 2019 435 2395 448
rect 1176 360 1276 376
rect 932 316 1052 360
rect 1156 316 1276 360
rect 1380 360 1480 376
rect 1851 395 1971 408
rect 1380 316 1500 360
rect 1851 349 1912 395
rect 1958 349 1971 395
rect 2019 389 2336 435
rect 2382 389 2395 435
rect 2019 376 2395 389
rect 1851 316 1971 349
rect 2075 316 2195 376
rect 2443 316 2563 496
rect 2687 467 2787 596
rect 2687 421 2718 467
rect 2764 421 2787 467
rect 2905 480 3005 596
rect 3109 552 3209 596
rect 2905 467 3291 480
rect 2905 440 3232 467
rect 2687 360 2787 421
rect 3115 421 3232 440
rect 3278 421 3291 467
rect 3115 408 3291 421
rect 3339 408 3439 596
rect 2667 316 2787 360
rect 2891 316 3011 360
rect 3115 316 3235 408
rect 3339 395 3459 408
rect 3339 349 3390 395
rect 3436 349 3459 395
rect 3339 316 3459 349
rect 3563 360 3663 596
rect 3563 316 3683 360
rect 124 112 244 156
rect 484 112 604 156
rect 708 64 828 156
rect 932 112 1052 156
rect 1156 112 1276 156
rect 1380 112 1500 156
rect 1851 112 1971 156
rect 2075 112 2195 156
rect 2443 112 2563 156
rect 2667 112 2787 156
rect 2891 64 3011 156
rect 3115 112 3235 156
rect 3339 112 3459 156
rect 3563 64 3683 156
rect 708 24 3683 64
<< polycontact >>
rect 157 421 203 467
rect 457 421 503 467
rect 717 395 763 441
rect 925 421 971 467
rect 1421 421 1467 467
rect 2120 509 2166 555
rect 1912 349 1958 395
rect 2336 389 2382 435
rect 2718 421 2764 467
rect 3232 421 3278 467
rect 3390 349 3436 395
<< metal1 >>
rect 0 918 3808 1098
rect 50 767 96 918
rect 1057 871 1103 918
rect 1057 814 1103 825
rect 273 767 319 778
rect 50 616 96 627
rect 142 467 203 654
rect 142 421 157 467
rect 142 410 203 421
rect 49 297 95 308
rect 49 90 95 251
rect 273 297 319 627
rect 365 768 591 778
rect 365 767 1463 768
rect 365 722 545 767
rect 365 297 411 722
rect 591 722 1463 767
rect 545 616 591 627
rect 809 665 855 676
rect 457 467 503 478
rect 457 400 503 421
rect 702 441 763 452
rect 702 400 717 441
rect 457 395 717 400
rect 457 354 763 395
rect 809 369 855 619
rect 1262 665 1351 676
rect 1262 619 1305 665
rect 925 467 978 542
rect 971 421 978 467
rect 925 410 978 421
rect 809 323 903 369
rect 857 297 903 323
rect 365 251 633 297
rect 679 251 690 297
rect 273 240 319 251
rect 857 240 903 251
rect 1081 297 1127 308
rect 1081 90 1127 251
rect 1262 297 1351 619
rect 1417 570 1463 722
rect 1509 767 1555 918
rect 2224 824 2554 870
rect 1509 616 1555 627
rect 1728 767 1801 778
rect 1728 627 1755 767
rect 1728 616 1801 627
rect 1847 767 2036 778
rect 1847 732 1990 767
rect 1728 570 1774 616
rect 1417 524 1774 570
rect 1421 467 1467 478
rect 1421 400 1467 421
rect 1421 354 1682 400
rect 1262 251 1305 297
rect 1262 240 1351 251
rect 1529 297 1575 308
rect 1529 90 1575 251
rect 1636 196 1682 354
rect 1728 299 1774 524
rect 1847 514 1893 732
rect 1990 616 2036 627
rect 2224 767 2282 824
rect 2224 627 2236 767
rect 1728 242 1774 253
rect 1820 472 1893 514
rect 2120 555 2166 566
rect 1820 196 1866 472
rect 2120 430 2166 509
rect 1912 395 2166 430
rect 1958 354 2166 395
rect 1912 338 1958 349
rect 2000 297 2046 308
rect 2000 196 2046 251
rect 2224 297 2282 627
rect 2270 251 2282 297
rect 2224 240 2282 251
rect 2336 767 2442 778
rect 2336 627 2396 767
rect 2336 435 2442 627
rect 2508 570 2554 824
rect 2600 767 2646 918
rect 2600 616 2646 627
rect 2692 824 3086 870
rect 2692 570 2738 824
rect 2508 524 2738 570
rect 2816 767 2862 778
rect 2382 389 2442 435
rect 2336 297 2442 389
rect 2718 467 2770 478
rect 2764 421 2770 467
rect 2718 354 2770 421
rect 2336 251 2368 297
rect 2414 251 2442 297
rect 2336 240 2442 251
rect 2592 297 2638 308
rect 1636 150 2046 196
rect 2592 90 2638 251
rect 2816 297 2862 627
rect 2816 240 2862 251
rect 3034 767 3086 824
rect 3080 627 3086 767
rect 3034 297 3086 627
rect 3238 767 3284 778
rect 3238 579 3284 627
rect 3468 767 3514 918
rect 3468 616 3514 627
rect 3692 767 3758 778
rect 3738 627 3758 767
rect 3034 251 3040 297
rect 3140 533 3284 579
rect 3140 297 3186 533
rect 3692 498 3758 627
rect 3314 487 3758 498
rect 3232 467 3758 487
rect 3278 452 3758 467
rect 3278 421 3344 452
rect 3232 410 3344 421
rect 3390 395 3442 406
rect 3436 349 3442 395
rect 3140 251 3264 297
rect 3310 251 3321 297
rect 3034 240 3086 251
rect 3390 242 3442 349
rect 3488 297 3534 308
rect 3488 90 3534 251
rect 3712 297 3758 452
rect 3712 240 3758 251
rect 0 -90 3808 90
<< labels >>
flabel metal1 s 3390 242 3442 406 0 FreeSans 200 0 0 0 I0
port 1 nsew default input
flabel metal1 s 2718 354 2770 478 0 FreeSans 200 0 0 0 I1
port 2 nsew default input
flabel metal1 s 142 410 203 654 0 FreeSans 200 0 0 0 I2
port 3 nsew default input
flabel metal1 s 925 410 978 542 0 FreeSans 200 0 0 0 I3
port 4 nsew default input
flabel metal1 s 457 452 503 478 0 FreeSans 200 0 0 0 S0
port 5 nsew default input
flabel metal1 s 2120 430 2166 566 0 FreeSans 200 0 0 0 S1
port 6 nsew default input
flabel metal1 s 0 918 3808 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 3488 90 3534 308 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1262 240 1351 676 0 FreeSans 200 0 0 0 Z
port 7 nsew default output
rlabel metal1 s 702 400 763 452 1 S0
port 5 nsew default input
rlabel metal1 s 457 400 503 452 1 S0
port 5 nsew default input
rlabel metal1 s 457 354 763 400 1 S0
port 5 nsew default input
rlabel metal1 s 1912 354 2166 430 1 S1
port 6 nsew default input
rlabel metal1 s 1912 338 1958 354 1 S1
port 6 nsew default input
rlabel metal1 s 3468 814 3514 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2600 814 2646 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1509 814 1555 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1057 814 1103 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 50 814 96 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3468 616 3514 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2600 616 2646 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1509 616 1555 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 50 616 96 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2592 90 2638 308 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1529 90 1575 308 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1081 90 1127 308 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 308 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3808 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 1008
string GDS_END 23244
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 14320
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
