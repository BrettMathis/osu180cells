magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -2205 102 2204 159
rect -2205 56 -2145 102
rect -2099 56 -1982 102
rect -1936 56 -1819 102
rect -1773 56 -1656 102
rect -1610 56 -1492 102
rect -1446 56 -1329 102
rect -1283 56 -1166 102
rect -1120 56 -1003 102
rect -957 56 -839 102
rect -793 56 -676 102
rect -630 56 -513 102
rect -467 56 -350 102
rect -304 56 -186 102
rect -140 56 -23 102
rect 23 56 140 102
rect 186 56 304 102
rect 350 56 467 102
rect 513 56 630 102
rect 676 56 793 102
rect 839 56 957 102
rect 1003 56 1120 102
rect 1166 56 1283 102
rect 1329 56 1446 102
rect 1492 56 1610 102
rect 1656 56 1773 102
rect 1819 56 1942 102
rect 1988 56 2105 102
rect 2151 56 2204 102
rect -2205 -56 2204 56
rect -2205 -102 -2145 -56
rect -2099 -102 -1982 -56
rect -1936 -102 -1819 -56
rect -1773 -102 -1656 -56
rect -1610 -102 -1492 -56
rect -1446 -102 -1329 -56
rect -1283 -102 -1166 -56
rect -1120 -102 -1003 -56
rect -957 -102 -839 -56
rect -793 -102 -676 -56
rect -630 -102 -513 -56
rect -467 -102 -350 -56
rect -304 -102 -186 -56
rect -140 -102 -23 -56
rect 23 -102 140 -56
rect 186 -102 304 -56
rect 350 -102 467 -56
rect 513 -102 630 -56
rect 676 -102 793 -56
rect 839 -102 957 -56
rect 1003 -102 1120 -56
rect 1166 -102 1283 -56
rect 1329 -102 1446 -56
rect 1492 -102 1610 -56
rect 1656 -102 1773 -56
rect 1819 -102 1942 -56
rect 1988 -102 2105 -56
rect 2151 -102 2204 -56
rect -2205 -159 2204 -102
<< psubdiffcont >>
rect -2145 56 -2099 102
rect -1982 56 -1936 102
rect -1819 56 -1773 102
rect -1656 56 -1610 102
rect -1492 56 -1446 102
rect -1329 56 -1283 102
rect -1166 56 -1120 102
rect -1003 56 -957 102
rect -839 56 -793 102
rect -676 56 -630 102
rect -513 56 -467 102
rect -350 56 -304 102
rect -186 56 -140 102
rect -23 56 23 102
rect 140 56 186 102
rect 304 56 350 102
rect 467 56 513 102
rect 630 56 676 102
rect 793 56 839 102
rect 957 56 1003 102
rect 1120 56 1166 102
rect 1283 56 1329 102
rect 1446 56 1492 102
rect 1610 56 1656 102
rect 1773 56 1819 102
rect 1942 56 1988 102
rect 2105 56 2151 102
rect -2145 -102 -2099 -56
rect -1982 -102 -1936 -56
rect -1819 -102 -1773 -56
rect -1656 -102 -1610 -56
rect -1492 -102 -1446 -56
rect -1329 -102 -1283 -56
rect -1166 -102 -1120 -56
rect -1003 -102 -957 -56
rect -839 -102 -793 -56
rect -676 -102 -630 -56
rect -513 -102 -467 -56
rect -350 -102 -304 -56
rect -186 -102 -140 -56
rect -23 -102 23 -56
rect 140 -102 186 -56
rect 304 -102 350 -56
rect 467 -102 513 -56
rect 630 -102 676 -56
rect 793 -102 839 -56
rect 957 -102 1003 -56
rect 1120 -102 1166 -56
rect 1283 -102 1329 -56
rect 1446 -102 1492 -56
rect 1610 -102 1656 -56
rect 1773 -102 1819 -56
rect 1942 -102 1988 -56
rect 2105 -102 2151 -56
<< metal1 >>
rect -2195 102 2195 150
rect -2195 56 -2145 102
rect -2099 56 -1982 102
rect -1936 56 -1819 102
rect -1773 56 -1656 102
rect -1610 56 -1492 102
rect -1446 56 -1329 102
rect -1283 56 -1166 102
rect -1120 56 -1003 102
rect -957 56 -839 102
rect -793 56 -676 102
rect -630 56 -513 102
rect -467 56 -350 102
rect -304 56 -186 102
rect -140 56 -23 102
rect 23 56 140 102
rect 186 56 304 102
rect 350 56 467 102
rect 513 56 630 102
rect 676 56 793 102
rect 839 56 957 102
rect 1003 56 1120 102
rect 1166 56 1283 102
rect 1329 56 1446 102
rect 1492 56 1610 102
rect 1656 56 1773 102
rect 1819 56 1942 102
rect 1988 56 2105 102
rect 2151 56 2195 102
rect -2195 -56 2195 56
rect -2195 -102 -2145 -56
rect -2099 -102 -1982 -56
rect -1936 -102 -1819 -56
rect -1773 -102 -1656 -56
rect -1610 -102 -1492 -56
rect -1446 -102 -1329 -56
rect -1283 -102 -1166 -56
rect -1120 -102 -1003 -56
rect -957 -102 -839 -56
rect -793 -102 -676 -56
rect -630 -102 -513 -56
rect -467 -102 -350 -56
rect -304 -102 -186 -56
rect -140 -102 -23 -56
rect 23 -102 140 -56
rect 186 -102 304 -56
rect 350 -102 467 -56
rect 513 -102 630 -56
rect 676 -102 793 -56
rect 839 -102 957 -56
rect 1003 -102 1120 -56
rect 1166 -102 1283 -56
rect 1329 -102 1446 -56
rect 1492 -102 1610 -56
rect 1656 -102 1773 -56
rect 1819 -102 1942 -56
rect 1988 -102 2105 -56
rect 2151 -102 2195 -56
rect -2195 -150 2195 -102
<< properties >>
string GDS_END 640776
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 637124
<< end >>
