magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 457 23867 23908 29129
rect 331 17407 22310 19961
rect 22338 17406 22926 19961
rect 22827 14326 23842 15917
rect 22880 8391 23005 9181
<< mvpmos >>
rect 6089 27950 6209 28632
rect 6314 27950 6434 28632
rect 6780 27950 6900 28632
rect 7005 27950 7125 28632
rect 16889 27950 17009 28632
rect 17114 27950 17234 28632
rect 17580 27950 17700 28632
rect 17805 27950 17925 28632
rect 6089 27175 6209 27857
rect 6314 27175 6434 27857
rect 6780 27175 6900 27857
rect 7005 27175 7125 27857
rect 16889 27175 17009 27857
rect 17114 27175 17234 27857
rect 17580 27175 17700 27857
rect 17805 27175 17925 27857
<< mvpdiff >>
rect 5981 27950 6089 28632
rect 6209 27950 6314 28632
rect 6434 27950 6780 28632
rect 6900 27950 7005 28632
rect 7125 27950 7294 28632
rect 16775 27950 16889 28632
rect 17009 27950 17114 28632
rect 17234 27950 17580 28632
rect 17700 27950 17805 28632
rect 17925 27950 18094 28632
rect 5981 27175 6089 27857
rect 6209 27175 6314 27857
rect 6434 27175 6780 27857
rect 6900 27175 7005 27857
rect 7125 27175 7294 27857
rect 16775 27175 16889 27857
rect 17009 27175 17114 27857
rect 17234 27175 17580 27857
rect 17700 27175 17805 27857
rect 17925 27175 18094 27857
<< metal1 >>
rect 54 30375 130 30387
rect 54 30323 66 30375
rect 118 30323 130 30375
rect 54 30311 130 30323
rect 11739 29839 11919 29851
rect 936 29818 1116 29830
rect 936 29766 948 29818
rect 1104 29766 1116 29818
rect 11739 29787 11751 29839
rect 11907 29787 11919 29839
rect 11739 29775 11919 29787
rect 22286 29793 24936 29890
rect 936 29754 1116 29766
rect 22286 29741 22912 29793
rect 23068 29741 24936 29793
rect 22286 29720 24936 29741
rect 22263 27031 22913 27105
rect 23206 18457 23552 19818
rect 23259 4973 23599 5013
rect 23259 4921 23297 4973
rect 23349 4921 23509 4973
rect 23561 4921 23599 4973
rect 23259 4755 23599 4921
rect 23259 4703 23297 4755
rect 23349 4703 23509 4755
rect 23561 4703 23599 4755
rect 23259 4662 23599 4703
<< via1 >>
rect 66 30323 118 30375
rect 948 29766 1104 29818
rect 11751 29787 11907 29839
rect 22912 29741 23068 29793
rect 23297 4921 23349 4973
rect 23509 4921 23561 4973
rect 23297 4703 23349 4755
rect 23509 4703 23561 4755
<< metal2 >>
rect 23857 51990 23982 52518
rect 54 30375 130 30387
rect 54 30323 66 30375
rect 118 30323 130 30375
rect 54 30311 130 30323
rect 976 29979 1077 31182
rect 976 29923 996 29979
rect 1052 29923 1077 29979
rect 976 29847 1077 29923
rect 976 29830 996 29847
rect 936 29818 996 29830
rect 1052 29830 1077 29847
rect 1052 29818 1116 29830
rect 936 29766 948 29818
rect 1104 29766 1116 29818
rect 936 29754 1116 29766
rect 976 29715 1077 29754
rect 976 29659 996 29715
rect 1052 29659 1077 29715
rect 976 29583 1077 29659
rect 976 29527 996 29583
rect 1052 29527 1077 29583
rect 976 29471 1077 29527
rect 1337 27527 1437 31182
rect 11777 29982 11877 31182
rect 11777 29926 11798 29982
rect 11854 29926 11877 29982
rect 11777 29851 11877 29926
rect 11739 29850 11919 29851
rect 11739 29839 11798 29850
rect 11854 29839 11919 29850
rect 11739 29787 11751 29839
rect 11907 29787 11919 29839
rect 11739 29775 11919 29787
rect 11777 29718 11877 29775
rect 11777 29662 11798 29718
rect 11854 29662 11877 29718
rect 11777 29586 11877 29662
rect 11777 29530 11798 29586
rect 11854 29530 11877 29586
rect 11777 29517 11877 29530
rect 12137 27527 12237 31182
rect 22577 27527 22677 31182
rect 22937 29979 23037 31182
rect 22937 29923 22958 29979
rect 23014 29923 23037 29979
rect 22937 29847 23037 29923
rect 22937 29805 22958 29847
rect 22900 29793 22958 29805
rect 23014 29805 23037 29847
rect 23857 29979 23982 30303
rect 23857 29923 23898 29979
rect 23954 29923 23982 29979
rect 23857 29847 23982 29923
rect 23014 29793 23080 29805
rect 22900 29741 22912 29793
rect 23068 29741 23080 29793
rect 22900 29729 23080 29741
rect 23857 29791 23898 29847
rect 23954 29791 23982 29847
rect 22937 29715 23037 29729
rect 22937 29659 22958 29715
rect 23014 29659 23037 29715
rect 22937 29583 23037 29659
rect 22937 29527 22958 29583
rect 23014 29527 23037 29583
rect 22937 27527 23037 29527
rect 23857 29715 23982 29791
rect 23857 29659 23898 29715
rect 23954 29659 23982 29715
rect 23857 29583 23982 29659
rect 23857 29527 23898 29583
rect 23954 29527 23982 29583
rect 23857 29471 23982 29527
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4757 23599 4919
rect 23259 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 23259 4662 23599 4701
<< via2 >>
rect 996 29923 1052 29979
rect 996 29818 1052 29847
rect 996 29791 1052 29818
rect 996 29659 1052 29715
rect 996 29527 1052 29583
rect 11798 29926 11854 29982
rect 11798 29839 11854 29850
rect 11798 29794 11854 29839
rect 11798 29662 11854 29718
rect 11798 29530 11854 29586
rect 22958 29923 23014 29979
rect 22958 29793 23014 29847
rect 23898 29923 23954 29979
rect 22958 29791 23014 29793
rect 23898 29791 23954 29847
rect 22958 29659 23014 29715
rect 22958 29527 23014 29583
rect 23898 29659 23954 29715
rect 23898 29527 23954 29583
rect 23295 4973 23351 4975
rect 23295 4921 23297 4973
rect 23297 4921 23349 4973
rect 23349 4921 23351 4973
rect 23295 4919 23351 4921
rect 23507 4973 23563 4975
rect 23507 4921 23509 4973
rect 23509 4921 23561 4973
rect 23561 4921 23563 4973
rect 23507 4919 23563 4921
rect 23295 4755 23351 4757
rect 23295 4703 23297 4755
rect 23297 4703 23349 4755
rect 23349 4703 23351 4755
rect 23295 4701 23351 4703
rect 23507 4755 23563 4757
rect 23507 4703 23509 4755
rect 23509 4703 23561 4755
rect 23561 4703 23563 4755
rect 23507 4701 23563 4703
<< metal3 >>
rect -493 60707 23681 60907
rect -229 30537 23681 30897
rect 48 30279 136 30368
rect -229 30139 23681 30279
rect 48 29997 136 30139
rect -229 29982 24087 29997
rect -229 29979 11798 29982
rect -229 29923 996 29979
rect 1052 29926 11798 29979
rect 11854 29979 24087 29982
rect 11854 29926 22958 29979
rect 1052 29923 22958 29926
rect 23014 29923 23898 29979
rect 23954 29923 24087 29979
rect -229 29850 24087 29923
rect -229 29847 11798 29850
rect -229 29791 996 29847
rect 1052 29794 11798 29847
rect 11854 29847 24087 29850
rect 11854 29794 22958 29847
rect 1052 29791 22958 29794
rect 23014 29791 23898 29847
rect 23954 29791 24087 29847
rect -229 29718 24087 29791
rect -229 29715 11798 29718
rect -229 29659 996 29715
rect 1052 29662 11798 29715
rect 11854 29715 24087 29718
rect 11854 29662 22958 29715
rect 1052 29659 22958 29662
rect 23014 29659 23898 29715
rect 23954 29659 24087 29715
rect -229 29586 24087 29659
rect -229 29583 11798 29586
rect -229 29527 996 29583
rect 1052 29530 11798 29583
rect 11854 29583 24087 29586
rect 11854 29530 22958 29583
rect 1052 29527 22958 29530
rect 23014 29527 23898 29583
rect 23954 29527 24087 29583
rect -229 29517 24087 29527
rect -229 27296 24087 29105
rect 314 21089 23252 21304
rect 314 20767 23252 20983
rect 314 20446 23252 20661
rect 314 20124 23252 20339
rect 314 19432 23252 19648
rect 314 19110 23252 19326
rect 314 18789 23252 19004
rect 314 18467 23252 18682
rect 314 17918 23252 18361
rect -336 16807 23252 17263
rect 991 12996 23252 15720
rect 1249 9308 23252 12711
rect 969 8442 23710 9158
rect 173 7016 24488 7827
rect 1314 6471 23971 6474
rect 225 5154 23971 6471
rect 76 4923 22676 5011
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4758 23599 4919
rect 76 4757 23599 4758
rect 76 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 76 4662 23599 4701
rect 225 3133 24166 4495
rect 225 1961 24276 2576
rect 225 1286 23252 1855
rect 225 747 24089 1179
rect 225 155 24508 610
rect 188 -959 24602 -504
rect 188 -1599 23252 -1247
rect 1082 -2041 23252 -1953
rect 188 -2517 23252 -2165
rect 188 -3242 23252 -2787
use M2_M1$$43374636_256x8m81  M2_M1$$43374636_256x8m81_0
timestamp 1669390400
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1669390400
transform -1 0 1026 0 -1 29792
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_1
timestamp 1669390400
transform 1 0 11829 0 1 29813
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_2
timestamp 1669390400
transform 1 0 22990 0 1 29767
box 0 0 1 1
use M2_M14310590878116_256x8m81  M2_M14310590878116_256x8m81_0
timestamp 1669390400
transform 1 0 92 0 1 30349
box 0 0 1 1
use M3_M2$$201416748_256x8m81  M3_M2$$201416748_256x8m81_0
timestamp 1669390400
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_0
timestamp 1669390400
transform 1 0 1024 0 1 29753
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_1
timestamp 1669390400
transform 1 0 23926 0 1 29753
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_2
timestamp 1669390400
transform 1 0 11826 0 1 29756
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_3
timestamp 1669390400
transform 1 0 22986 0 1 29753
box 0 0 1 1
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_0
timestamp 1669390400
transform 1 0 12186 0 1 28317
box -38 -764 38 764
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_1
timestamp 1669390400
transform 1 0 22626 0 1 28317
box -38 -764 38 764
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_2
timestamp 1669390400
transform 1 0 1386 0 1 28317
box -38 -764 38 764
use dcap_103_novia_256x8m81  dcap_103_novia_256x8m81_0
array 0 35 619 0 0 0
timestamp 1669390400
transform 1 0 21 0 1 29009
box -203 -284 822 881
use rarray4_256_256x8m81  rarray4_256_256x8m81_0
timestamp 1669390400
transform 1 0 907 0 1 31107
box 430 -68 22268 28868
use rdummy_256x4_256x8m81  rdummy_256x4_256x8m81_0
timestamp 1669390400
transform 1 0 -5093 0 1 30207
box 5143 -25410 29464 30688
use saout_R_m2_256x8m81  saout_R_m2_256x8m81_0
timestamp 1669390400
transform -1 0 12194 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_256x8m81  saout_R_m2_256x8m81_1
timestamp 1669390400
transform -1 0 22994 0 1 6
box -269 -3400 7633 31133
use saout_m2_256x8m81  saout_m2_256x8m81_0
timestamp 1669390400
transform 1 0 11820 0 1 -1
box -269 -3393 7633 31140
use saout_m2_256x8m81  saout_m2_256x8m81_1
timestamp 1669390400
transform 1 0 1020 0 1 -1
box -269 -3393 7633 31140
<< labels >>
rlabel metal1 s 7342 15928 7342 15928 4 pcb[6]
port 1 nsew
rlabel metal1 s 5921 15928 5921 15928 4 pcb[7]
port 2 nsew
rlabel metal1 s 18209 15928 18209 15928 4 pcb[4]
port 3 nsew
rlabel metal1 s 1827 18163 1827 18163 4 vdd
port 4 nsew
flabel metal1 s 23444 27062 23444 27062 0 FreeSans 100 0 0 0 PCB[8]
port 5 nsew
flabel metal1 s 22465 -3332 22465 -3332 0 FreeSans 600 0 0 0 WEN[4]
port 6 nsew
flabel metal1 s 1584 -3332 1584 -3332 0 FreeSans 600 0 0 0 WEN[7]
port 7 nsew
rlabel metal1 s 16588 15928 16588 15928 4 pcb[5]
port 8 nsew
flabel metal1 s 12358 -3332 12358 -3332 0 FreeSans 600 0 0 0 WEN[5]
port 9 nsew
flabel metal1 s 11643 -3332 11643 -3332 0 FreeSans 600 0 0 0 WEN[6]
port 10 nsew
flabel metal3 s 1659 24526 1659 24526 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
rlabel metal3 s 1607 36968 1607 36968 4 WL[6]
port 12 nsew
rlabel metal3 s 1607 36068 1607 36068 4 WL[5]
port 13 nsew
rlabel metal3 s 1777 1467 1777 1467 4 men
port 14 nsew
rlabel metal3 s 1704 18914 1704 18914 4 ypass[1]
port 15 nsew
rlabel metal3 s 1704 19231 1704 19231 4 ypass[2]
port 16 nsew
rlabel metal3 s 1704 19548 1704 19548 4 ypass[3]
port 17 nsew
rlabel metal3 s 1704 20204 1704 20204 4 ypass[4]
port 18 nsew
rlabel metal3 s 1704 20528 1704 20528 4 ypass[5]
port 19 nsew
rlabel metal3 s 1704 20845 1704 20845 4 ypass[6]
port 20 nsew
rlabel metal3 s 1774 1467 1774 1467 4 men
port 14 nsew
rlabel metal3 s 1592 60357 1592 60357 4 DWL
port 21 nsew
rlabel metal3 s 1346 4726 1346 4726 4 tblhl
port 22 nsew
flabel metal3 s 1659 -2004 1659 -2004 0 FreeSans 1000 0 0 0 GWEN
port 23 nsew
flabel metal3 s 1659 -3019 1659 -3019 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
rlabel metal3 s 1777 8832 1777 8832 4 VDD
port 11 nsew
rlabel metal3 s 1777 5806 1777 5806 4 VSS
port 24 nsew
flabel metal3 s 1659 -781 1659 -781 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 1659 -2347 1659 -2347 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
rlabel metal3 s 240 30277 240 30277 4 VSS
port 24 nsew
rlabel metal3 s 1777 60853 1777 60853 4 VSS
port 24 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 14 nsew
rlabel metal3 s 1704 18591 1704 18591 4 ypass[0]
port 25 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 14 nsew
rlabel metal3 s 1608 57668 1608 57668 4 WL[29]
port 26 nsew
rlabel metal3 s 1608 54068 1608 54068 4 WL[25]
port 27 nsew
rlabel metal3 s 1608 53168 1608 53168 4 WL[24]
port 28 nsew
rlabel metal3 s 1608 52268 1608 52268 4 WL[23]
port 29 nsew
rlabel metal3 s 1608 51368 1608 51368 4 WL[22]
port 30 nsew
rlabel metal3 s 1608 49568 1608 49568 4 WL[20]
port 31 nsew
rlabel metal3 s 1608 55868 1608 55868 4 WL[27]
port 32 nsew
rlabel metal3 s 1608 58568 1608 58568 4 WL[30]
port 33 nsew
rlabel metal3 s 1608 47768 1608 47768 4 WL[18]
port 34 nsew
rlabel metal3 s 1346 4983 1346 4983 4 GWE
port 35 nsew
rlabel metal3 s 1608 41468 1608 41468 4 WL[11]
port 36 nsew
rlabel metal3 s 1608 45068 1608 45068 4 WL[15]
port 37 nsew
rlabel metal3 s 1608 31568 1608 31568 4 WL[0]
port 38 nsew
rlabel metal3 s 1608 33368 1608 33368 4 WL[2]
port 39 nsew
rlabel metal3 s 1608 42368 1608 42368 4 WL[12]
port 40 nsew
rlabel metal3 s 1608 34268 1608 34268 4 WL[3]
port 41 nsew
rlabel metal3 s 1608 35168 1608 35168 4 WL[4]
port 42 nsew
rlabel metal3 s 1608 37868 1608 37868 4 WL[7]
port 43 nsew
rlabel metal3 s 1608 38768 1608 38768 4 WL[8]
port 44 nsew
rlabel metal3 s 1608 39668 1608 39668 4 WL[9]
port 45 nsew
rlabel metal3 s 1608 32468 1608 32468 4 WL[1]
port 46 nsew
rlabel metal3 s 1705 21162 1705 21162 4 ypass[7]
port 47 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 14 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 14 nsew
flabel metal3 s 1659 -1446 1659 -1446 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
rlabel metal3 s 1608 59468 1608 59468 4 WL[31]
port 48 nsew
rlabel metal3 s 1608 40568 1608 40568 4 WL[10]
port 49 nsew
rlabel metal3 s 1608 43268 1608 43268 4 WL[13]
port 50 nsew
rlabel metal3 s 1608 44168 1608 44168 4 WL[14]
port 51 nsew
rlabel metal3 s 1608 45968 1608 45968 4 WL[16]
port 52 nsew
rlabel metal3 s 1608 46868 1608 46868 4 WL[17]
port 53 nsew
rlabel metal3 s 1608 54968 1608 54968 4 WL[26]
port 54 nsew
rlabel metal3 s 1608 48668 1608 48668 4 WL[19]
port 55 nsew
rlabel metal3 s 1608 56768 1608 56768 4 WL[28]
port 56 nsew
rlabel metal3 s 1608 50468 1608 50468 4 WL[21]
port 57 nsew
flabel metal3 s 1659 390 1659 390 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 1659 3623 1659 3623 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 1659 7598 1659 7598 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 1659 18106 1659 18106 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 1659 28191 1659 28191 0 FreeSans 2000 0 0 0 VDD
port 11 nsew
flabel metal3 s 151 29699 151 29699 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 1659 23123 1659 23123 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 436 16976 436 16976 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 1659 12236 1659 12236 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 1659 6155 1659 6155 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 1659 2247 1659 2247 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
flabel metal3 s 1659 949 1659 949 0 FreeSans 2000 0 0 0 VSS
port 24 nsew
rlabel metal2 s 1519 104 1519 104 4 din[4]
port 58 nsew
rlabel metal2 s 22489 104 22489 104 4 din[7]
port 59 nsew
rlabel metal2 s 10835 138 10835 138 4 q[5]
port 60 nsew
rlabel metal2 s 13174 104 13174 104 4 q[6]
port 61 nsew
rlabel metal2 s 21643 104 21643 104 4 q[7]
port 62 nsew
rlabel metal2 s 11696 104 11696 104 4 din[5]
port 63 nsew
rlabel metal2 s 12325 104 12325 104 4 din[6]
port 64 nsew
rlabel metal2 s 2378 104 2378 104 4 q[4]
port 65 nsew
<< properties >>
string GDS_END 2346082
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2334856
<< end >>
