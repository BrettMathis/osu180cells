magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -42 44423 342 44442
rect -42 -23 -23 44423
rect 323 -23 342 44423
rect -42 -42 342 -23
<< psubdiffcont >>
rect -23 -23 323 44423
<< metal1 >>
rect -34 44423 334 44434
rect -34 -23 -23 44423
rect 323 -23 334 44423
rect -34 -34 334 -23
<< properties >>
string GDS_END 1212234
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1098118
<< end >>
