magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -1962 137 1962 176
rect -1962 81 -1926 137
rect -1870 81 -1715 137
rect -1659 81 -1504 137
rect -1448 81 -1293 137
rect -1237 81 -1082 137
rect -1026 81 -872 137
rect -816 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 816 137
rect 872 81 1026 137
rect 1082 81 1237 137
rect 1293 81 1448 137
rect 1504 81 1659 137
rect 1715 81 1870 137
rect 1926 81 1962 137
rect -1962 -81 1962 81
rect -1962 -137 -1926 -81
rect -1870 -137 -1715 -81
rect -1659 -137 -1504 -81
rect -1448 -137 -1293 -81
rect -1237 -137 -1082 -81
rect -1026 -137 -872 -81
rect -816 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 816 -81
rect 872 -137 1026 -81
rect 1082 -137 1237 -81
rect 1293 -137 1448 -81
rect 1504 -137 1659 -81
rect 1715 -137 1870 -81
rect 1926 -137 1962 -81
rect -1962 -175 1962 -137
<< via2 >>
rect -1926 81 -1870 137
rect -1715 81 -1659 137
rect -1504 81 -1448 137
rect -1293 81 -1237 137
rect -1082 81 -1026 137
rect -872 81 -816 137
rect -661 81 -605 137
rect -450 81 -394 137
rect -239 81 -183 137
rect -28 81 28 137
rect 183 81 239 137
rect 394 81 450 137
rect 605 81 661 137
rect 816 81 872 137
rect 1026 81 1082 137
rect 1237 81 1293 137
rect 1448 81 1504 137
rect 1659 81 1715 137
rect 1870 81 1926 137
rect -1926 -137 -1870 -81
rect -1715 -137 -1659 -81
rect -1504 -137 -1448 -81
rect -1293 -137 -1237 -81
rect -1082 -137 -1026 -81
rect -872 -137 -816 -81
rect -661 -137 -605 -81
rect -450 -137 -394 -81
rect -239 -137 -183 -81
rect -28 -137 28 -81
rect 183 -137 239 -81
rect 394 -137 450 -81
rect 605 -137 661 -81
rect 816 -137 872 -81
rect 1026 -137 1082 -81
rect 1237 -137 1293 -81
rect 1448 -137 1504 -81
rect 1659 -137 1715 -81
rect 1870 -137 1926 -81
<< metal3 >>
rect -1962 137 1962 176
rect -1962 81 -1926 137
rect -1870 81 -1715 137
rect -1659 81 -1504 137
rect -1448 81 -1293 137
rect -1237 81 -1082 137
rect -1026 81 -872 137
rect -816 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 816 137
rect 872 81 1026 137
rect 1082 81 1237 137
rect 1293 81 1448 137
rect 1504 81 1659 137
rect 1715 81 1870 137
rect 1926 81 1962 137
rect -1962 -81 1962 81
rect -1962 -137 -1926 -81
rect -1870 -137 -1715 -81
rect -1659 -137 -1504 -81
rect -1448 -137 -1293 -81
rect -1237 -137 -1082 -81
rect -1026 -137 -872 -81
rect -816 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 816 -81
rect 872 -137 1026 -81
rect 1082 -137 1237 -81
rect 1293 -137 1448 -81
rect 1504 -137 1659 -81
rect 1715 -137 1870 -81
rect 1926 -137 1962 -81
rect -1962 -176 1962 -137
<< properties >>
string GDS_END 953794
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 951230
<< end >>
