magic
tech gf180mcuB
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -50 231 50 236
rect -50 203 -45 231
rect -17 203 17 231
rect 45 203 50 231
rect -50 169 50 203
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -203 50 -169
rect -50 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 50 -203
rect -50 -236 50 -231
<< via2 >>
rect -45 203 -17 231
rect 17 203 45 231
rect -45 141 -17 169
rect 17 141 45 169
rect -45 79 -17 107
rect 17 79 45 107
rect -45 17 -17 45
rect 17 17 45 45
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect -45 -169 -17 -141
rect 17 -169 45 -141
rect -45 -231 -17 -203
rect 17 -231 45 -203
<< metal3 >>
rect -50 231 50 236
rect -50 203 -45 231
rect -17 203 17 231
rect 45 203 50 231
rect -50 169 50 203
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -203 50 -169
rect -50 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 50 -203
rect -50 -236 50 -231
<< properties >>
string GDS_END 1105610
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1104454
<< end >>
