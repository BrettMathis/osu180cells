magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 459 3334 1094
rect -86 453 86 459
rect 2663 453 3334 459
<< pwell >>
rect 86 453 2663 459
rect -86 -86 3334 453
<< mvnmos >>
rect 386 267 506 339
rect 124 123 244 195
rect 386 123 506 195
rect 818 212 938 284
rect 1186 212 1306 284
rect 818 68 938 140
rect 1186 68 1306 140
rect 1618 258 1738 330
rect 1986 258 2106 330
rect 1618 114 1738 186
rect 1986 114 2106 186
rect 2418 213 2538 285
rect 2418 69 2538 141
rect 2778 69 2898 333
rect 3002 69 3122 333
<< mvpmos >>
rect 124 783 224 855
rect 386 783 486 855
rect 386 639 486 711
rect 818 783 918 855
rect 1186 783 1286 855
rect 818 639 918 711
rect 1186 639 1286 711
rect 1618 783 1718 855
rect 1986 783 2086 855
rect 1618 639 1718 711
rect 1986 639 2086 711
rect 2418 783 2518 855
rect 2418 639 2518 711
rect 2778 574 2878 940
rect 3002 574 3102 940
<< mvndiff >>
rect 298 326 386 339
rect 298 280 311 326
rect 357 280 386 326
rect 298 267 386 280
rect 506 267 626 339
rect 566 195 626 267
rect 36 182 124 195
rect 36 136 49 182
rect 95 136 124 182
rect 36 123 124 136
rect 244 182 386 195
rect 244 136 273 182
rect 319 136 386 182
rect 244 123 386 136
rect 506 123 626 195
rect 698 212 818 284
rect 938 271 1026 284
rect 938 225 967 271
rect 1013 225 1026 271
rect 938 212 1026 225
rect 1098 271 1186 284
rect 1098 225 1111 271
rect 1157 225 1186 271
rect 1098 212 1186 225
rect 1306 212 1426 284
rect 698 140 758 212
rect 1366 140 1426 212
rect 698 68 818 140
rect 938 127 1186 140
rect 938 81 967 127
rect 1013 81 1186 127
rect 938 68 1186 81
rect 1306 68 1426 140
rect 1498 258 1618 330
rect 1738 317 1826 330
rect 1738 271 1767 317
rect 1813 271 1826 317
rect 1738 258 1826 271
rect 1898 317 1986 330
rect 1898 271 1911 317
rect 1957 271 1986 317
rect 1898 258 1986 271
rect 2106 258 2226 330
rect 1498 186 1558 258
rect 2166 186 2226 258
rect 1498 114 1618 186
rect 1738 173 1986 186
rect 1738 127 1767 173
rect 1813 127 1986 173
rect 1738 114 1986 127
rect 2106 114 2226 186
rect 2298 213 2418 285
rect 2538 272 2626 285
rect 2538 226 2567 272
rect 2613 226 2626 272
rect 2538 213 2626 226
rect 2298 141 2358 213
rect 2698 141 2778 333
rect 2298 69 2418 141
rect 2538 128 2778 141
rect 2538 82 2567 128
rect 2613 82 2778 128
rect 2538 69 2778 82
rect 2898 320 3002 333
rect 2898 180 2927 320
rect 2973 180 3002 320
rect 2898 69 3002 180
rect 3122 276 3210 333
rect 3122 136 3151 276
rect 3197 136 3210 276
rect 3122 69 3210 136
<< mvpdiff >>
rect 2698 855 2778 940
rect 36 842 124 855
rect 36 796 49 842
rect 95 796 124 842
rect 36 783 124 796
rect 224 842 386 855
rect 224 796 253 842
rect 299 796 386 842
rect 224 783 386 796
rect 486 783 606 855
rect 546 711 606 783
rect 298 698 386 711
rect 298 652 311 698
rect 357 652 386 698
rect 298 639 386 652
rect 486 639 606 711
rect 698 783 818 855
rect 918 842 1186 855
rect 918 796 947 842
rect 993 796 1186 842
rect 918 783 1186 796
rect 1286 783 1406 855
rect 698 711 758 783
rect 1346 711 1406 783
rect 698 639 818 711
rect 918 698 1006 711
rect 918 652 947 698
rect 993 652 1006 698
rect 918 639 1006 652
rect 1098 698 1186 711
rect 1098 652 1111 698
rect 1157 652 1186 698
rect 1098 639 1186 652
rect 1286 639 1406 711
rect 1498 783 1618 855
rect 1718 842 1986 855
rect 1718 796 1747 842
rect 1793 796 1986 842
rect 1718 783 1986 796
rect 2086 783 2206 855
rect 1498 711 1558 783
rect 2146 711 2206 783
rect 1498 639 1618 711
rect 1718 698 1806 711
rect 1718 652 1747 698
rect 1793 652 1806 698
rect 1718 639 1806 652
rect 1898 698 1986 711
rect 1898 652 1911 698
rect 1957 652 1986 698
rect 1898 639 1986 652
rect 2086 639 2206 711
rect 2298 783 2418 855
rect 2518 842 2778 855
rect 2518 796 2547 842
rect 2593 796 2778 842
rect 2518 783 2778 796
rect 2298 711 2358 783
rect 2298 639 2418 711
rect 2518 698 2606 711
rect 2518 652 2547 698
rect 2593 652 2606 698
rect 2518 639 2606 652
rect 2698 574 2778 783
rect 2878 861 3002 940
rect 2878 721 2907 861
rect 2953 721 3002 861
rect 2878 574 3002 721
rect 3102 868 3190 940
rect 3102 728 3131 868
rect 3177 728 3190 868
rect 3102 574 3190 728
<< mvndiffc >>
rect 311 280 357 326
rect 49 136 95 182
rect 273 136 319 182
rect 967 225 1013 271
rect 1111 225 1157 271
rect 967 81 1013 127
rect 1767 271 1813 317
rect 1911 271 1957 317
rect 1767 127 1813 173
rect 2567 226 2613 272
rect 2567 82 2613 128
rect 2927 180 2973 320
rect 3151 136 3197 276
<< mvpdiffc >>
rect 49 796 95 842
rect 253 796 299 842
rect 311 652 357 698
rect 947 796 993 842
rect 947 652 993 698
rect 1111 652 1157 698
rect 1747 796 1793 842
rect 1747 652 1793 698
rect 1911 652 1957 698
rect 2547 796 2593 842
rect 2547 652 2593 698
rect 2907 721 2953 861
rect 3131 728 3177 868
<< polysilicon >>
rect 2778 940 2878 984
rect 3002 940 3102 984
rect 124 855 224 899
rect 386 855 486 899
rect 818 855 918 899
rect 1186 855 1286 899
rect 1618 855 1718 899
rect 1986 855 2086 899
rect 2418 855 2518 899
rect 124 514 224 783
rect 386 711 486 783
rect 818 711 918 783
rect 1186 711 1286 783
rect 1618 711 1718 783
rect 1986 711 2086 783
rect 2418 711 2518 783
rect 124 374 141 514
rect 187 374 224 514
rect 124 239 224 374
rect 386 595 486 639
rect 386 455 399 595
rect 445 455 486 595
rect 386 383 486 455
rect 818 514 918 639
rect 386 339 506 383
rect 818 374 831 514
rect 877 374 918 514
rect 818 328 918 374
rect 1186 514 1286 639
rect 1186 374 1199 514
rect 1245 374 1286 514
rect 1186 328 1286 374
rect 1618 514 1718 639
rect 1618 374 1631 514
rect 1677 374 1718 514
rect 1986 514 2086 639
rect 1986 374 1999 514
rect 2045 374 2086 514
rect 2418 514 2518 639
rect 2418 374 2431 514
rect 2477 374 2518 514
rect 1618 330 1738 374
rect 1986 330 2106 374
rect 818 284 938 328
rect 1186 284 1306 328
rect 124 195 244 239
rect 386 195 506 267
rect 818 140 938 212
rect 1186 140 1306 212
rect 124 79 244 123
rect 386 79 506 123
rect 2418 329 2518 374
rect 2778 480 2878 574
rect 3002 480 3102 574
rect 2778 467 3102 480
rect 2778 421 2791 467
rect 3025 421 3102 467
rect 2778 408 3102 421
rect 2778 333 2898 408
rect 3002 377 3102 408
rect 3002 333 3122 377
rect 2418 285 2538 329
rect 1618 186 1738 258
rect 1986 186 2106 258
rect 2418 141 2538 213
rect 1618 70 1738 114
rect 1986 70 2106 114
rect 818 24 938 68
rect 1186 24 1306 68
rect 2418 25 2538 69
rect 2778 25 2898 69
rect 3002 25 3122 69
<< polycontact >>
rect 141 374 187 514
rect 399 455 445 595
rect 831 374 877 514
rect 1199 374 1245 514
rect 1631 374 1677 514
rect 1999 374 2045 514
rect 2431 374 2477 514
rect 2791 421 3025 467
<< metal1 >>
rect 0 918 3248 1098
rect 38 842 95 853
rect 38 796 49 842
rect 38 606 95 796
rect 253 842 299 918
rect 253 785 299 796
rect 947 842 993 918
rect 947 785 993 796
rect 1747 842 1793 918
rect 1747 785 1793 796
rect 2547 842 2593 918
rect 2706 861 2953 872
rect 2706 814 2907 861
rect 2547 785 2593 796
rect 947 698 993 709
rect 300 652 311 698
rect 357 652 877 698
rect 38 595 445 606
rect 38 560 399 595
rect 38 182 84 560
rect 130 374 141 514
rect 187 374 198 514
rect 399 444 445 455
rect 831 514 877 652
rect 130 354 198 374
rect 831 326 877 374
rect 300 280 311 326
rect 357 280 877 326
rect 947 525 993 652
rect 1111 698 1157 709
rect 1111 617 1157 652
rect 1747 698 1793 709
rect 1111 571 1677 617
rect 947 514 1245 525
rect 947 374 1199 514
rect 947 363 1245 374
rect 1631 514 1677 571
rect 947 271 1013 363
rect 1631 317 1677 374
rect 947 225 967 271
rect 947 214 1013 225
rect 1111 271 1677 317
rect 1747 525 1793 652
rect 1911 698 1957 709
rect 1911 617 1957 652
rect 2547 698 2593 709
rect 1911 571 2477 617
rect 1747 514 2045 525
rect 1747 374 1999 514
rect 1747 363 2045 374
rect 2431 514 2477 571
rect 1747 317 1813 363
rect 2431 317 2477 374
rect 1747 271 1767 317
rect 1900 271 1911 317
rect 1957 271 2477 317
rect 2547 478 2593 652
rect 2907 673 2953 721
rect 3131 868 3177 918
rect 3131 717 3177 728
rect 2907 627 3117 673
rect 2547 467 3025 478
rect 2547 421 2791 467
rect 2547 410 3025 421
rect 2547 272 2613 410
rect 3071 364 3117 627
rect 1747 260 1813 271
rect 1111 214 1157 225
rect 2547 226 2567 272
rect 2547 215 2613 226
rect 2927 320 3117 364
rect 273 182 319 193
rect 38 136 49 182
rect 95 136 106 182
rect 1767 173 1813 184
rect 273 90 319 136
rect 967 127 1013 138
rect 0 81 967 90
rect 2973 318 3117 320
rect 2927 169 2973 180
rect 3151 276 3197 287
rect 1767 90 1813 127
rect 2567 128 2613 139
rect 1013 82 2567 90
rect 3151 90 3197 136
rect 2613 82 3248 90
rect 1013 81 3248 82
rect 0 -90 3248 81
<< labels >>
flabel metal1 s 130 354 198 514 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 3248 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 3151 193 3197 287 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2706 814 2953 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
rlabel metal1 s 2907 673 2953 814 1 Z
port 2 nsew default output
rlabel metal1 s 2907 627 3117 673 1 Z
port 2 nsew default output
rlabel metal1 s 3071 364 3117 627 1 Z
port 2 nsew default output
rlabel metal1 s 2927 318 3117 364 1 Z
port 2 nsew default output
rlabel metal1 s 2927 169 2973 318 1 Z
port 2 nsew default output
rlabel metal1 s 3131 785 3177 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2547 785 2593 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1747 785 1793 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 947 785 993 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 253 785 299 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3131 717 3177 785 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3151 184 3197 193 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 184 319 193 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3151 139 3197 184 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1767 139 1813 184 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 139 319 184 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3151 138 3197 139 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2567 138 2613 139 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1767 138 1813 139 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 138 319 139 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3151 90 3197 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2567 90 2613 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1767 90 1813 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 967 90 1013 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3248 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3248 1008
string GDS_END 740868
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 733710
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
