magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 7386 4662 7661 7575
<< metal2 >>
rect 978 11057 1108 11191
rect 1334 11057 1464 11191
rect 2768 11057 2898 11191
rect 3130 11057 3260 11191
rect 4079 10021 4433 12483
rect 5188 11456 5313 11457
rect 12566 11456 12691 11457
rect 5186 11418 5315 11456
rect 5186 11362 5223 11418
rect 5279 11362 5315 11418
rect 5186 11200 5315 11362
rect 5186 11144 5223 11200
rect 5279 11144 5315 11200
rect 12565 11418 12694 11456
rect 12565 11362 12601 11418
rect 12657 11362 12694 11418
rect 12565 11200 12694 11362
rect 14996 11279 15349 12544
rect 5186 10293 5315 11144
rect 8357 11057 8486 11191
rect 8713 11057 8842 11191
rect 10147 11057 10276 11191
rect 10509 11057 10638 11191
rect 12565 11144 12601 11200
rect 12657 11144 12694 11200
rect 12565 10293 12694 11144
rect 12868 10915 15349 11279
rect 12868 10021 13221 10915
rect 15755 10724 15977 11417
rect 16107 10724 16328 11417
rect 17389 10724 17611 11417
rect 17741 10724 17962 11417
rect 19023 10724 19245 11417
rect 19374 10724 19596 11417
rect 20657 10724 20878 11417
rect 21008 10724 21230 11417
rect 21944 10021 22297 12483
rect 23052 11456 23177 11457
rect 23051 11418 23180 11456
rect 23051 11362 23087 11418
rect 23143 11362 23180 11418
rect 23051 11200 23180 11362
rect 23051 11144 23087 11200
rect 23143 11144 23180 11200
rect 23051 10293 23180 11144
rect 5485 212 5614 346
rect 7176 212 7305 346
rect 12863 212 12993 346
rect 14554 212 14683 346
rect 23349 212 23478 346
rect 25040 212 25169 346
rect 26731 212 26860 346
<< via2 >>
rect 5223 11362 5279 11418
rect 5223 11144 5279 11200
rect 12601 11362 12657 11418
rect 12601 11144 12657 11200
rect 23087 11362 23143 11418
rect 23087 11144 23143 11200
<< metal3 >>
rect 47 11636 27260 12544
rect 5188 11456 5314 11457
rect 12566 11456 12692 11457
rect 23052 11456 23178 11457
rect 47 11418 23180 11456
rect 47 11362 5223 11418
rect 5279 11362 12601 11418
rect 12657 11362 23087 11418
rect 23143 11362 23180 11418
rect 47 11200 23180 11362
rect 47 11144 5223 11200
rect 5279 11144 12601 11200
rect 12657 11144 23087 11200
rect 23143 11144 23180 11200
rect 47 11105 23180 11144
rect 7509 2234 8254 2916
rect 7509 1078 8254 1986
rect 7509 -1 8254 907
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_0
timestamp 1669390400
transform 1 0 5251 0 1 11281
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_1
timestamp 1669390400
transform 1 0 12629 0 1 11281
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_2
timestamp 1669390400
transform 1 0 23115 0 1 11281
box 0 0 1 1
use M3_M2$$47115308_64x8m81  M3_M2$$47115308_64x8m81_0
timestamp 1669390400
transform 1 0 4256 0 1 12090
box -170 -393 170 393
use M3_M2$$47115308_64x8m81  M3_M2$$47115308_64x8m81_1
timestamp 1669390400
transform 1 0 22120 0 1 12090
box -170 -393 170 393
use M3_M2$$201412652_64x8m81  M3_M2$$201412652_64x8m81_0
timestamp 1669390400
transform 1 0 15172 0 1 12090
box -170 -393 170 393
use xpredec0_64x8m81  xpredec0_64x8m81_0
timestamp 1669390400
transform 1 0 7704 0 1 0
box -289 -1 7456 11434
use xpredec0_64x8m81  xpredec0_64x8m81_1
timestamp 1669390400
transform 1 0 325 0 1 0
box -289 -1 7456 11434
use xpredec1_64x8m81  xpredec1_64x8m81_0
timestamp 1669390400
transform 1 0 15082 0 1 0
box -1 -1 12233 10971
<< labels >>
rlabel metal3 s 22643 11310 22643 11310 4 clk
port 1 nsew
rlabel metal3 s 25504 12090 25504 12090 4 men
port 2 nsew
rlabel metal2 s 23414 279 23414 279 4 A[2]
port 3 nsew
rlabel metal2 s 5549 279 5549 279 4 A[6]
port 4 nsew
rlabel metal2 s 12928 279 12928 279 4 A[4]
port 5 nsew
rlabel metal2 s 8422 11124 8422 11124 4 xb[3]
port 6 nsew
rlabel metal2 s 21123 11351 21123 11351 4 xa[0]
port 7 nsew
rlabel metal2 s 3195 11120 3195 11120 4 xc[0]
port 8 nsew
rlabel metal2 s 2833 11120 2833 11120 4 xc[1]
port 9 nsew
rlabel metal2 s 1399 11124 1399 11124 4 xc[2]
port 10 nsew
rlabel metal2 s 1043 11124 1043 11124 4 xc[3]
port 11 nsew
rlabel metal2 s 10211 11120 10211 11120 4 xb[1]
port 12 nsew
rlabel metal2 s 8777 11124 8777 11124 4 xb[2]
port 13 nsew
rlabel metal2 s 10574 11120 10574 11120 4 xb[0]
port 14 nsew
rlabel metal2 s 20763 11351 20763 11351 4 xa[1]
port 15 nsew
rlabel metal2 s 19476 11351 19476 11351 4 xa[2]
port 16 nsew
rlabel metal2 s 19134 11351 19134 11351 4 xa[3]
port 17 nsew
rlabel metal2 s 17853 11351 17853 11351 4 xa[4]
port 18 nsew
rlabel metal2 s 17498 11351 17498 11351 4 xa[5]
port 19 nsew
rlabel metal2 s 16215 11351 16215 11351 4 xa[6]
port 20 nsew
rlabel metal2 s 15864 11351 15864 11351 4 xa[7]
port 21 nsew
rlabel metal2 s 26796 279 26796 279 4 A[0]
port 22 nsew
rlabel metal2 s 14619 279 14619 279 4 A[3]
port 23 nsew
rlabel metal2 s 7240 279 7240 279 4 A[5]
port 24 nsew
rlabel metal2 s 25105 279 25105 279 4 A[1]
port 25 nsew
<< properties >>
string GDS_END 1624044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1620322
<< end >>
