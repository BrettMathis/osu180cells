magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 3160 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
rect 1550 190 1610 360
rect 1720 190 1780 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2230 190 2290 360
rect 2400 190 2460 360
rect 2570 190 2630 360
rect 2740 190 2800 360
rect 2910 190 2970 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
rect 870 1090 930 1430
rect 1040 1090 1100 1430
rect 1210 1090 1270 1430
rect 1380 1090 1440 1430
rect 1550 1090 1610 1430
rect 1720 1090 1780 1430
rect 1890 1090 1950 1430
rect 2060 1090 2120 1430
rect 2230 1090 2290 1430
rect 2400 1090 2460 1430
rect 2570 1090 2630 1430
rect 2740 1090 2800 1430
rect 2910 1090 2970 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 870 360
rect 760 252 792 298
rect 838 252 870 298
rect 760 190 870 252
rect 930 298 1040 360
rect 930 252 962 298
rect 1008 252 1040 298
rect 930 190 1040 252
rect 1100 298 1210 360
rect 1100 252 1132 298
rect 1178 252 1210 298
rect 1100 190 1210 252
rect 1270 298 1380 360
rect 1270 252 1302 298
rect 1348 252 1380 298
rect 1270 190 1380 252
rect 1440 298 1550 360
rect 1440 252 1472 298
rect 1518 252 1550 298
rect 1440 190 1550 252
rect 1610 298 1720 360
rect 1610 252 1642 298
rect 1688 252 1720 298
rect 1610 190 1720 252
rect 1780 298 1890 360
rect 1780 252 1812 298
rect 1858 252 1890 298
rect 1780 190 1890 252
rect 1950 298 2060 360
rect 1950 252 1982 298
rect 2028 252 2060 298
rect 1950 190 2060 252
rect 2120 298 2230 360
rect 2120 252 2152 298
rect 2198 252 2230 298
rect 2120 190 2230 252
rect 2290 298 2400 360
rect 2290 252 2322 298
rect 2368 252 2400 298
rect 2290 190 2400 252
rect 2460 298 2570 360
rect 2460 252 2492 298
rect 2538 252 2570 298
rect 2460 190 2570 252
rect 2630 298 2740 360
rect 2630 252 2662 298
rect 2708 252 2740 298
rect 2630 190 2740 252
rect 2800 298 2910 360
rect 2800 252 2832 298
rect 2878 252 2910 298
rect 2800 190 2910 252
rect 2970 298 3070 360
rect 2970 252 3002 298
rect 3048 252 3070 298
rect 2970 190 3070 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 870 1430
rect 760 1143 792 1377
rect 838 1143 870 1377
rect 760 1090 870 1143
rect 930 1377 1040 1430
rect 930 1143 962 1377
rect 1008 1143 1040 1377
rect 930 1090 1040 1143
rect 1100 1377 1210 1430
rect 1100 1143 1132 1377
rect 1178 1143 1210 1377
rect 1100 1090 1210 1143
rect 1270 1377 1380 1430
rect 1270 1143 1302 1377
rect 1348 1143 1380 1377
rect 1270 1090 1380 1143
rect 1440 1377 1550 1430
rect 1440 1143 1472 1377
rect 1518 1143 1550 1377
rect 1440 1090 1550 1143
rect 1610 1377 1720 1430
rect 1610 1143 1642 1377
rect 1688 1143 1720 1377
rect 1610 1090 1720 1143
rect 1780 1377 1890 1430
rect 1780 1143 1812 1377
rect 1858 1143 1890 1377
rect 1780 1090 1890 1143
rect 1950 1377 2060 1430
rect 1950 1143 1982 1377
rect 2028 1143 2060 1377
rect 1950 1090 2060 1143
rect 2120 1377 2230 1430
rect 2120 1143 2152 1377
rect 2198 1143 2230 1377
rect 2120 1090 2230 1143
rect 2290 1377 2400 1430
rect 2290 1143 2322 1377
rect 2368 1143 2400 1377
rect 2290 1090 2400 1143
rect 2460 1377 2570 1430
rect 2460 1143 2492 1377
rect 2538 1143 2570 1377
rect 2460 1090 2570 1143
rect 2630 1377 2740 1430
rect 2630 1143 2662 1377
rect 2708 1143 2740 1377
rect 2630 1090 2740 1143
rect 2800 1377 2910 1430
rect 2800 1143 2832 1377
rect 2878 1143 2910 1377
rect 2800 1090 2910 1143
rect 2970 1377 3070 1430
rect 2970 1143 3002 1377
rect 3048 1143 3070 1377
rect 2970 1090 3070 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
rect 962 252 1008 298
rect 1132 252 1178 298
rect 1302 252 1348 298
rect 1472 252 1518 298
rect 1642 252 1688 298
rect 1812 252 1858 298
rect 1982 252 2028 298
rect 2152 252 2198 298
rect 2322 252 2368 298
rect 2492 252 2538 298
rect 2662 252 2708 298
rect 2832 252 2878 298
rect 3002 252 3048 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
rect 962 1143 1008 1377
rect 1132 1143 1178 1377
rect 1302 1143 1348 1377
rect 1472 1143 1518 1377
rect 1642 1143 1688 1377
rect 1812 1143 1858 1377
rect 1982 1143 2028 1377
rect 2152 1143 2198 1377
rect 2322 1143 2368 1377
rect 2492 1143 2538 1377
rect 2662 1143 2708 1377
rect 2832 1143 2878 1377
rect 3002 1143 3048 1377
<< psubdiff >>
rect 90 98 190 120
rect 90 52 112 98
rect 158 52 190 98
rect 90 30 190 52
rect 330 98 430 120
rect 330 52 352 98
rect 398 52 430 98
rect 330 30 430 52
rect 570 98 670 120
rect 570 52 592 98
rect 638 52 670 98
rect 570 30 670 52
rect 810 98 910 120
rect 810 52 832 98
rect 878 52 910 98
rect 810 30 910 52
rect 1050 98 1150 120
rect 1050 52 1072 98
rect 1118 52 1150 98
rect 1050 30 1150 52
rect 1290 98 1390 120
rect 1290 52 1312 98
rect 1358 52 1390 98
rect 1290 30 1390 52
rect 1530 98 1630 120
rect 1530 52 1552 98
rect 1598 52 1630 98
rect 1530 30 1630 52
rect 1770 98 1870 120
rect 1770 52 1792 98
rect 1838 52 1870 98
rect 1770 30 1870 52
rect 2010 98 2110 120
rect 2010 52 2032 98
rect 2078 52 2110 98
rect 2010 30 2110 52
rect 2250 98 2350 120
rect 2250 52 2272 98
rect 2318 52 2350 98
rect 2250 30 2350 52
rect 2490 98 2590 120
rect 2490 52 2512 98
rect 2558 52 2590 98
rect 2490 30 2590 52
rect 2730 98 2830 120
rect 2730 52 2752 98
rect 2798 52 2830 98
rect 2730 30 2830 52
<< nsubdiff >>
rect 90 1568 190 1590
rect 90 1522 112 1568
rect 158 1522 190 1568
rect 90 1500 190 1522
rect 330 1568 430 1590
rect 330 1522 352 1568
rect 398 1522 430 1568
rect 330 1500 430 1522
rect 570 1568 670 1590
rect 570 1522 592 1568
rect 638 1522 670 1568
rect 570 1500 670 1522
rect 810 1568 910 1590
rect 810 1522 832 1568
rect 878 1522 910 1568
rect 810 1500 910 1522
rect 1050 1568 1150 1590
rect 1050 1522 1072 1568
rect 1118 1522 1150 1568
rect 1050 1500 1150 1522
rect 1290 1568 1390 1590
rect 1290 1522 1312 1568
rect 1358 1522 1390 1568
rect 1290 1500 1390 1522
rect 1530 1568 1630 1590
rect 1530 1522 1552 1568
rect 1598 1522 1630 1568
rect 1530 1500 1630 1522
rect 1770 1568 1870 1590
rect 1770 1522 1792 1568
rect 1838 1522 1870 1568
rect 1770 1500 1870 1522
rect 2010 1568 2110 1590
rect 2010 1522 2032 1568
rect 2078 1522 2110 1568
rect 2010 1500 2110 1522
rect 2250 1568 2350 1590
rect 2250 1522 2272 1568
rect 2318 1522 2350 1568
rect 2250 1500 2350 1522
rect 2490 1568 2590 1590
rect 2490 1522 2512 1568
rect 2558 1522 2590 1568
rect 2490 1500 2590 1522
rect 2730 1568 2830 1590
rect 2730 1522 2752 1568
rect 2798 1522 2830 1568
rect 2730 1500 2830 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
rect 2752 52 2798 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
rect 1552 1522 1598 1568
rect 1792 1522 1838 1568
rect 2032 1522 2078 1568
rect 2272 1522 2318 1568
rect 2512 1522 2558 1568
rect 2752 1522 2798 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 870 1430 930 1480
rect 1040 1430 1100 1480
rect 1210 1430 1270 1480
rect 1380 1430 1440 1480
rect 1550 1430 1610 1480
rect 1720 1430 1780 1480
rect 1890 1430 1950 1480
rect 2060 1430 2120 1480
rect 2230 1430 2290 1480
rect 2400 1430 2460 1480
rect 2570 1430 2630 1480
rect 2740 1430 2800 1480
rect 2910 1430 2970 1480
rect 190 910 250 1090
rect 360 1070 420 1090
rect 530 1070 590 1090
rect 700 1070 760 1090
rect 870 1070 930 1090
rect 1040 1070 1100 1090
rect 1210 1070 1270 1090
rect 1380 1070 1440 1090
rect 1550 1070 1610 1090
rect 1720 1070 1780 1090
rect 1890 1070 1950 1090
rect 2060 1070 2120 1090
rect 2230 1070 2290 1090
rect 2400 1070 2460 1090
rect 2570 1070 2630 1090
rect 2740 1070 2800 1090
rect 2910 1070 2970 1090
rect 360 1010 2970 1070
rect 190 883 310 910
rect 190 837 237 883
rect 283 837 310 883
rect 190 810 310 837
rect 190 360 250 810
rect 360 670 420 1010
rect 300 633 420 670
rect 300 587 327 633
rect 373 587 420 633
rect 300 550 420 587
rect 360 440 420 550
rect 700 440 760 1010
rect 1040 440 1100 1010
rect 1380 440 1440 1010
rect 1720 440 1780 1010
rect 2060 440 2120 1010
rect 2400 440 2460 1010
rect 2740 440 2800 1010
rect 360 380 2970 440
rect 360 360 420 380
rect 530 360 590 380
rect 700 360 760 380
rect 870 360 930 380
rect 1040 360 1100 380
rect 1210 360 1270 380
rect 1380 360 1440 380
rect 1550 360 1610 380
rect 1720 360 1780 380
rect 1890 360 1950 380
rect 2060 360 2120 380
rect 2230 360 2290 380
rect 2400 360 2460 380
rect 2570 360 2630 380
rect 2740 360 2800 380
rect 2910 360 2970 380
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
rect 1550 140 1610 190
rect 1720 140 1780 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2230 140 2290 190
rect 2400 140 2460 190
rect 2570 140 2630 190
rect 2740 140 2800 190
rect 2910 140 2970 190
<< polycontact >>
rect 237 837 283 883
rect 327 587 373 633
<< metal1 >>
rect 0 1590 3160 1620
rect -170 1568 3160 1590
rect -170 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1552 1568
rect 1598 1566 1792 1568
rect 1838 1566 2032 1568
rect 2078 1566 2272 1568
rect 2318 1566 2512 1568
rect 2558 1566 2752 1568
rect 2798 1566 3160 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 1366 1522 1552 1566
rect 1606 1522 1792 1566
rect 1846 1522 2032 1566
rect 2086 1522 2272 1566
rect 2326 1522 2512 1566
rect 2566 1522 2752 1566
rect -170 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1794 1522
rect 1846 1514 2034 1522
rect 2086 1514 2274 1522
rect 2326 1514 2514 1522
rect 2566 1514 2754 1522
rect 2806 1514 3160 1566
rect -170 1500 3160 1514
rect -170 1470 2990 1500
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 860 160 1143
rect 280 1377 330 1470
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 1000 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1030 500 1143
rect 620 1377 670 1470
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 1030 670 1143
rect 790 1377 840 1470
rect 790 1143 792 1377
rect 838 1143 840 1377
rect 790 1030 840 1143
rect 960 1377 1010 1470
rect 960 1143 962 1377
rect 1008 1143 1010 1377
rect 960 1030 1010 1143
rect 1130 1377 1180 1470
rect 1130 1143 1132 1377
rect 1178 1143 1180 1377
rect 1130 1030 1180 1143
rect 1300 1377 1350 1470
rect 1300 1143 1302 1377
rect 1348 1143 1350 1377
rect 1300 1030 1350 1143
rect 1470 1377 1520 1470
rect 1470 1143 1472 1377
rect 1518 1143 1520 1377
rect 1470 1030 1520 1143
rect 1640 1377 1690 1470
rect 1640 1143 1642 1377
rect 1688 1143 1690 1377
rect 1640 1030 1690 1143
rect 1810 1377 1860 1470
rect 1810 1143 1812 1377
rect 1858 1143 1860 1377
rect 1810 1030 1860 1143
rect 1980 1377 2030 1470
rect 1980 1143 1982 1377
rect 2028 1143 2030 1377
rect 1980 1030 2030 1143
rect 2150 1377 2200 1470
rect 2150 1143 2152 1377
rect 2198 1143 2200 1377
rect 2150 1030 2200 1143
rect 2320 1377 2370 1470
rect 2320 1143 2322 1377
rect 2368 1143 2370 1377
rect 2320 1030 2370 1143
rect 2490 1377 2540 1470
rect 2490 1143 2492 1377
rect 2538 1143 2540 1377
rect 2490 1030 2540 1143
rect 2660 1377 2710 1470
rect 2660 1143 2662 1377
rect 2708 1143 2710 1377
rect 2660 1030 2710 1143
rect 2830 1377 2880 1470
rect 2830 1143 2832 1377
rect 2878 1143 2880 1377
rect 2830 1030 2880 1143
rect 3000 1377 3050 1500
rect 3000 1143 3002 1377
rect 3048 1143 3050 1377
rect 3000 1090 3050 1143
rect 450 1026 2910 1030
rect 450 1000 2834 1026
rect 280 974 2834 1000
rect 2886 974 2910 1026
rect 280 970 2910 974
rect 280 940 2740 970
rect 280 890 330 940
rect 40 800 160 860
rect 210 886 330 890
rect 210 834 234 886
rect 286 834 330 886
rect 210 830 330 834
rect 110 640 160 800
rect 280 640 330 830
rect 110 633 400 640
rect 110 587 327 633
rect 373 587 400 633
rect 110 580 400 587
rect 110 298 160 580
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 430 330 580
rect 450 460 500 940
rect 620 460 670 940
rect 790 460 840 940
rect 960 460 1010 940
rect 1130 460 1180 940
rect 1300 460 1350 940
rect 1470 460 1520 940
rect 1640 460 1690 940
rect 1810 460 1860 940
rect 1980 460 2030 940
rect 2150 460 2200 940
rect 2320 460 2370 940
rect 2490 460 2540 940
rect 2660 460 2710 940
rect 2830 460 2880 970
rect 450 430 2880 460
rect 280 410 2880 430
rect 280 380 2710 410
rect 280 298 330 380
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 450 298 500 380
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 380
rect 620 252 622 298
rect 668 252 670 298
rect 620 120 670 252
rect 790 298 840 380
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 960 298 1010 380
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 120 1010 252
rect 1130 298 1180 380
rect 1130 252 1132 298
rect 1178 252 1180 298
rect 1130 120 1180 252
rect 1300 298 1350 380
rect 1300 252 1302 298
rect 1348 252 1350 298
rect 1300 120 1350 252
rect 1470 298 1520 380
rect 1470 252 1472 298
rect 1518 252 1520 298
rect 1470 120 1520 252
rect 1640 298 1690 380
rect 1640 252 1642 298
rect 1688 252 1690 298
rect 1640 120 1690 252
rect 1810 298 1860 380
rect 1810 252 1812 298
rect 1858 252 1860 298
rect 1810 120 1860 252
rect 1980 298 2030 380
rect 1980 252 1982 298
rect 2028 252 2030 298
rect 1980 120 2030 252
rect 2150 298 2200 380
rect 2150 252 2152 298
rect 2198 252 2200 298
rect 2150 120 2200 252
rect 2320 298 2370 380
rect 2320 252 2322 298
rect 2368 252 2370 298
rect 2320 120 2370 252
rect 2490 298 2540 380
rect 2490 252 2492 298
rect 2538 252 2540 298
rect 2490 120 2540 252
rect 2660 298 2710 380
rect 2660 252 2662 298
rect 2708 252 2710 298
rect 2660 120 2710 252
rect 2830 298 2880 410
rect 2830 252 2832 298
rect 2878 252 2880 298
rect 2830 120 2880 252
rect 3000 298 3050 360
rect 3000 252 3002 298
rect 3048 252 3050 298
rect 3000 120 3050 252
rect 0 106 3160 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 2566 98 2754 106
rect 0 90 112 98
rect -170 52 112 90
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2752 98
rect 2806 54 3160 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2752 54
rect 2798 52 3160 54
rect -170 0 3160 52
rect -170 -30 2990 0
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 1554 1522 1598 1566
rect 1598 1522 1606 1566
rect 1794 1522 1838 1566
rect 1838 1522 1846 1566
rect 2034 1522 2078 1566
rect 2078 1522 2086 1566
rect 2274 1522 2318 1566
rect 2318 1522 2326 1566
rect 2514 1522 2558 1566
rect 2558 1522 2566 1566
rect 2754 1522 2798 1566
rect 2798 1522 2806 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 1794 1514 1846 1522
rect 2034 1514 2086 1522
rect 2274 1514 2326 1522
rect 2514 1514 2566 1522
rect 2754 1514 2806 1522
rect 2834 974 2886 1026
rect 234 883 286 886
rect 234 837 237 883
rect 237 837 283 883
rect 283 837 286 883
rect 234 834 286 837
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 2754 98 2806 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
rect 2754 54 2798 98
rect 2798 54 2806 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect 1780 1570 1860 1580
rect 2020 1570 2100 1580
rect 2260 1570 2340 1580
rect 2500 1570 2580 1580
rect 2740 1570 2820 1580
rect 90 1566 190 1570
rect -70 1540 10 1550
rect -80 1480 20 1540
rect 90 1514 114 1566
rect 166 1550 190 1566
rect 330 1566 430 1570
rect 166 1540 250 1550
rect 166 1514 260 1540
rect 90 1510 260 1514
rect 330 1514 354 1566
rect 406 1550 430 1566
rect 570 1566 670 1570
rect 406 1540 490 1550
rect 406 1514 500 1540
rect 330 1510 500 1514
rect 570 1514 594 1566
rect 646 1550 670 1566
rect 810 1566 910 1570
rect 646 1540 730 1550
rect 646 1514 740 1540
rect 570 1510 740 1514
rect 810 1514 834 1566
rect 886 1550 910 1566
rect 1050 1566 1150 1570
rect 886 1540 970 1550
rect 886 1514 980 1540
rect 810 1510 980 1514
rect 1050 1514 1074 1566
rect 1126 1550 1150 1566
rect 1290 1566 1390 1570
rect 1126 1540 1210 1550
rect 1126 1514 1220 1540
rect 1050 1510 1220 1514
rect 1290 1514 1314 1566
rect 1366 1550 1390 1566
rect 1530 1566 1630 1570
rect 1366 1540 1450 1550
rect 1366 1514 1460 1540
rect 1290 1510 1460 1514
rect 1530 1514 1554 1566
rect 1606 1550 1630 1566
rect 1770 1566 1870 1570
rect 1606 1540 1690 1550
rect 1606 1514 1700 1540
rect 1530 1510 1700 1514
rect 1770 1514 1794 1566
rect 1846 1550 1870 1566
rect 2010 1566 2110 1570
rect 1846 1540 1930 1550
rect 1846 1514 1940 1540
rect 1770 1510 1940 1514
rect 2010 1514 2034 1566
rect 2086 1550 2110 1566
rect 2250 1566 2350 1570
rect 2086 1540 2170 1550
rect 2086 1514 2180 1540
rect 2010 1510 2180 1514
rect 2250 1514 2274 1566
rect 2326 1550 2350 1566
rect 2490 1566 2590 1570
rect 2326 1540 2410 1550
rect 2326 1514 2420 1540
rect 2250 1510 2420 1514
rect 2490 1514 2514 1566
rect 2566 1550 2590 1566
rect 2730 1566 2830 1570
rect 2566 1540 2650 1550
rect 2566 1514 2660 1540
rect 2490 1510 2660 1514
rect 2730 1514 2754 1566
rect 2806 1514 2830 1566
rect 2730 1510 2830 1514
rect 100 1500 260 1510
rect 340 1500 500 1510
rect 580 1500 740 1510
rect 820 1500 980 1510
rect 1060 1500 1220 1510
rect 1300 1500 1460 1510
rect 1540 1500 1700 1510
rect 1780 1500 1940 1510
rect 2020 1500 2180 1510
rect 2260 1500 2420 1510
rect 2500 1500 2660 1510
rect 2740 1500 2820 1510
rect 160 1480 260 1500
rect 400 1480 500 1500
rect 640 1480 740 1500
rect 880 1480 980 1500
rect 1120 1480 1220 1500
rect 1360 1480 1460 1500
rect 1600 1480 1700 1500
rect 1840 1480 1940 1500
rect 2080 1480 2180 1500
rect 2320 1480 2420 1500
rect 2560 1480 2660 1500
rect -70 1470 10 1480
rect 170 1470 250 1480
rect 410 1470 490 1480
rect 650 1470 730 1480
rect 890 1470 970 1480
rect 1130 1470 1210 1480
rect 1370 1470 1450 1480
rect 1610 1470 1690 1480
rect 1850 1470 1930 1480
rect 2090 1470 2170 1480
rect 2330 1470 2410 1480
rect 2570 1470 2650 1480
rect 2810 1030 2910 1040
rect 2800 1026 2910 1030
rect 2640 1000 2740 1010
rect 2630 940 2740 1000
rect 2800 974 2834 1026
rect 2886 974 2910 1026
rect 2800 970 2910 974
rect 2810 960 2910 970
rect 2640 930 2740 940
rect 220 890 300 900
rect 210 886 310 890
rect 50 860 130 870
rect 40 800 140 860
rect 210 834 234 886
rect 286 834 310 886
rect 210 830 310 834
rect 220 820 300 830
rect 50 790 130 800
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 2740 110 2820 120
rect 90 106 190 110
rect -70 80 10 90
rect -80 20 20 80
rect 90 54 114 106
rect 166 90 190 106
rect 330 106 430 110
rect 166 80 250 90
rect 166 54 260 80
rect 90 50 260 54
rect 330 54 354 106
rect 406 90 430 106
rect 570 106 670 110
rect 406 80 490 90
rect 406 54 500 80
rect 330 50 500 54
rect 570 54 594 106
rect 646 90 670 106
rect 810 106 910 110
rect 646 80 730 90
rect 646 54 740 80
rect 570 50 740 54
rect 810 54 834 106
rect 886 90 910 106
rect 1050 106 1150 110
rect 886 80 970 90
rect 886 54 980 80
rect 810 50 980 54
rect 1050 54 1074 106
rect 1126 90 1150 106
rect 1290 106 1390 110
rect 1126 80 1210 90
rect 1126 54 1220 80
rect 1050 50 1220 54
rect 1290 54 1314 106
rect 1366 90 1390 106
rect 1530 106 1630 110
rect 1366 80 1450 90
rect 1366 54 1460 80
rect 1290 50 1460 54
rect 1530 54 1554 106
rect 1606 90 1630 106
rect 1770 106 1870 110
rect 1606 80 1690 90
rect 1606 54 1700 80
rect 1530 50 1700 54
rect 1770 54 1794 106
rect 1846 90 1870 106
rect 2010 106 2110 110
rect 1846 80 1930 90
rect 1846 54 1940 80
rect 1770 50 1940 54
rect 2010 54 2034 106
rect 2086 90 2110 106
rect 2250 106 2350 110
rect 2086 80 2170 90
rect 2086 54 2180 80
rect 2010 50 2180 54
rect 2250 54 2274 106
rect 2326 90 2350 106
rect 2490 106 2590 110
rect 2326 80 2410 90
rect 2326 54 2420 80
rect 2250 50 2420 54
rect 2490 54 2514 106
rect 2566 90 2590 106
rect 2730 106 2830 110
rect 2566 80 2650 90
rect 2566 54 2660 80
rect 2490 50 2660 54
rect 2730 54 2754 106
rect 2806 54 2830 106
rect 2730 50 2830 54
rect 100 40 260 50
rect 340 40 500 50
rect 580 40 740 50
rect 820 40 980 50
rect 1060 40 1220 50
rect 1300 40 1460 50
rect 1540 40 1700 50
rect 1780 40 1940 50
rect 2020 40 2180 50
rect 2260 40 2420 50
rect 2500 40 2660 50
rect 2740 40 2820 50
rect 160 20 260 40
rect 400 20 500 40
rect 640 20 740 40
rect 880 20 980 40
rect 1120 20 1220 40
rect 1360 20 1460 40
rect 1600 20 1700 40
rect 1840 20 1940 40
rect 2080 20 2180 40
rect 2320 20 2420 40
rect 2560 20 2660 40
rect -70 10 10 20
rect 170 10 250 20
rect 410 10 490 20
rect 650 10 730 20
rect 890 10 970 20
rect 1130 10 1210 20
rect 1370 10 1450 20
rect 1610 10 1690 20
rect 1850 10 1930 20
rect 2090 10 2170 20
rect 2330 10 2410 20
rect 2570 10 2650 20
<< labels >>
rlabel metal2 s -70 10 10 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s -70 1470 10 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 50 790 130 870 4 A
port 1 nsew signal input
rlabel metal2 s 2630 940 2740 1000 4 Y
port 2 nsew signal output
rlabel metal2 s 40 800 140 860 1 A
port 1 nsew signal input
rlabel metal1 s 40 800 140 860 1 A
port 1 nsew signal input
rlabel metal2 s -80 1480 20 1540 3 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 170 1470 250 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 160 1480 260 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 410 1470 490 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 400 1480 500 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 650 1470 730 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 640 1480 740 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 890 1470 970 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 880 1480 980 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1130 1470 1210 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1120 1480 1220 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1370 1470 1450 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1360 1480 1460 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1610 1470 1690 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1600 1480 1700 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1850 1470 1930 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1840 1480 1940 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2090 1470 2170 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2080 1480 2180 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2330 1470 2410 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2320 1480 2420 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2570 1470 2650 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2560 1480 2660 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 1060 840 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1130 1060 1180 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1470 1060 1520 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1810 1060 1860 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 1060 2200 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2490 1060 2540 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2830 1060 2880 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s -170 1470 2990 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s -80 20 20 80 3 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 170 10 250 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 160 20 260 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 410 10 490 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 400 20 500 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 650 10 730 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 640 20 740 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 890 10 970 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 880 20 980 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1130 10 1210 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1120 20 1220 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1370 10 1450 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1360 20 1460 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1610 10 1690 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1600 20 1700 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1850 10 1930 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1840 20 1940 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2090 10 2170 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2080 20 2180 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2330 10 2410 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2320 20 2420 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2570 10 2650 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2560 20 2660 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 -30 840 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1130 -30 1180 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1470 -30 1520 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1810 -30 1860 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2150 -30 2200 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2490 -30 2540 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2830 -30 2880 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s -170 -30 2990 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2640 930 2740 1010 1 Y
port 2 nsew signal output
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 620 160 670 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 960 160 1010 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 160 1350 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1640 160 1690 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1980 160 2030 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 2320 160 2370 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 380 2710 430 1 Y
port 2 nsew signal output
rlabel metal1 s 2660 160 2710 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 940 2740 1000 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX -170 -30 2990 1590
string GDS_END 110506
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 87498
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
