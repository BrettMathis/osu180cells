magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -295 -137 355 1454
<< polysilicon >>
rect -31 1318 89 1389
rect -31 -71 89 -1
use pmos_5p043105908781101_256x8m81  pmos_5p043105908781101_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 1438
<< properties >>
string GDS_END 2072556
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2072240
<< end >>
