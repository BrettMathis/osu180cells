magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 388 4678 870
rect -86 352 645 388
rect 2851 352 4678 388
<< pwell >>
rect 645 352 2851 388
rect -86 -86 4678 352
<< mvnmos >>
rect 124 151 244 232
rect 348 151 468 232
rect 788 171 908 244
rect 1012 171 1132 244
rect 1236 171 1356 244
rect 1404 171 1524 244
rect 1572 171 1692 244
rect 1916 156 2036 257
rect 2084 156 2204 257
rect 2320 156 2440 257
rect 2544 156 2664 257
rect 3112 156 3232 232
rect 3296 156 3416 232
rect 3520 156 3640 232
rect 3692 156 3812 232
rect 4060 69 4180 232
rect 4284 69 4404 232
<< mvpmos >>
rect 124 472 224 645
rect 328 472 428 645
rect 732 517 832 590
rect 936 517 1036 590
rect 1140 517 1240 590
rect 1344 517 1444 590
rect 1636 526 1736 677
rect 1984 526 2084 677
rect 2276 508 2376 580
rect 2480 508 2580 580
rect 2684 508 2784 580
rect 3132 491 3232 645
rect 3336 491 3436 645
rect 3540 491 3640 645
rect 3744 491 3844 645
rect 4092 472 4192 715
rect 4296 472 4396 715
<< mvndiff >>
rect 1771 244 1916 257
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 151 124 173
rect 244 210 348 232
rect 244 164 273 210
rect 319 164 348 210
rect 244 151 348 164
rect 468 210 556 232
rect 468 164 497 210
rect 543 164 556 210
rect 700 230 788 244
rect 700 184 713 230
rect 759 184 788 230
rect 700 171 788 184
rect 908 230 1012 244
rect 908 184 937 230
rect 983 184 1012 230
rect 908 171 1012 184
rect 1132 230 1236 244
rect 1132 184 1161 230
rect 1207 184 1236 230
rect 1132 171 1236 184
rect 1356 171 1404 244
rect 1524 171 1572 244
rect 1692 183 1916 244
rect 1692 171 1781 183
rect 468 151 556 164
rect 1752 137 1781 171
rect 1827 156 1916 183
rect 2036 156 2084 257
rect 2204 244 2320 257
rect 2204 198 2245 244
rect 2291 198 2320 244
rect 2204 156 2320 198
rect 2440 244 2544 257
rect 2440 198 2469 244
rect 2515 198 2544 244
rect 2440 156 2544 198
rect 2664 244 2752 257
rect 2664 198 2693 244
rect 2739 198 2752 244
rect 2664 156 2752 198
rect 3024 215 3112 232
rect 3024 169 3037 215
rect 3083 169 3112 215
rect 3024 156 3112 169
rect 3232 156 3296 232
rect 3416 215 3520 232
rect 3416 169 3445 215
rect 3491 169 3520 215
rect 3416 156 3520 169
rect 3640 156 3692 232
rect 3812 215 3900 232
rect 3812 169 3841 215
rect 3887 169 3900 215
rect 3812 156 3900 169
rect 1827 137 1856 156
rect 1752 124 1856 137
rect 3972 142 4060 232
rect 3972 96 3985 142
rect 4031 96 4060 142
rect 3972 69 4060 96
rect 4180 218 4284 232
rect 4180 172 4209 218
rect 4255 172 4284 218
rect 4180 69 4284 172
rect 4404 128 4512 232
rect 4404 82 4453 128
rect 4499 82 4512 128
rect 4404 69 4512 82
<< mvpdiff >>
rect 588 647 672 660
rect 36 632 124 645
rect 36 492 49 632
rect 95 492 124 632
rect 36 472 124 492
rect 224 632 328 645
rect 224 586 253 632
rect 299 586 328 632
rect 224 472 328 586
rect 428 632 516 645
rect 428 492 457 632
rect 503 492 516 632
rect 588 601 613 647
rect 659 601 672 647
rect 588 590 672 601
rect 1504 735 1576 748
rect 1504 689 1517 735
rect 1563 689 1576 735
rect 2144 735 2216 748
rect 1504 677 1576 689
rect 2144 689 2157 735
rect 2203 689 2216 735
rect 2144 677 2216 689
rect 1504 590 1636 677
rect 588 517 732 590
rect 832 576 936 590
rect 832 530 861 576
rect 907 530 936 576
rect 832 517 936 530
rect 1036 576 1140 590
rect 1036 530 1065 576
rect 1111 530 1140 576
rect 1036 517 1140 530
rect 1240 576 1344 590
rect 1240 530 1269 576
rect 1315 530 1344 576
rect 1240 517 1344 530
rect 1444 526 1636 590
rect 1736 585 1824 677
rect 1736 539 1765 585
rect 1811 539 1824 585
rect 1736 526 1824 539
rect 1896 585 1984 677
rect 1896 539 1909 585
rect 1955 539 1984 585
rect 1896 526 1984 539
rect 2084 580 2216 677
rect 4004 665 4092 715
rect 3023 632 3132 645
rect 3023 586 3036 632
rect 3082 586 3132 632
rect 2084 526 2276 580
rect 1444 517 1576 526
rect 428 472 516 492
rect 2144 508 2276 526
rect 2376 567 2480 580
rect 2376 521 2405 567
rect 2451 521 2480 567
rect 2376 508 2480 521
rect 2580 567 2684 580
rect 2580 521 2609 567
rect 2655 521 2684 567
rect 2580 508 2684 521
rect 2784 567 2872 580
rect 2784 521 2813 567
rect 2859 521 2872 567
rect 2784 508 2872 521
rect 3023 491 3132 586
rect 3232 550 3336 645
rect 3232 504 3261 550
rect 3307 504 3336 550
rect 3232 491 3336 504
rect 3436 632 3540 645
rect 3436 586 3465 632
rect 3511 586 3540 632
rect 3436 491 3540 586
rect 3640 550 3744 645
rect 3640 504 3669 550
rect 3715 504 3744 550
rect 3640 491 3744 504
rect 3844 619 3932 645
rect 3844 573 3873 619
rect 3919 573 3932 619
rect 3844 491 3932 573
rect 4004 525 4017 665
rect 4063 525 4092 665
rect 4004 472 4092 525
rect 4192 665 4296 715
rect 4192 525 4221 665
rect 4267 525 4296 665
rect 4192 472 4296 525
rect 4396 665 4484 715
rect 4396 525 4425 665
rect 4471 525 4484 665
rect 4396 472 4484 525
<< mvndiffc >>
rect 49 173 95 219
rect 273 164 319 210
rect 497 164 543 210
rect 713 184 759 230
rect 937 184 983 230
rect 1161 184 1207 230
rect 1781 137 1827 183
rect 2245 198 2291 244
rect 2469 198 2515 244
rect 2693 198 2739 244
rect 3037 169 3083 215
rect 3445 169 3491 215
rect 3841 169 3887 215
rect 3985 96 4031 142
rect 4209 172 4255 218
rect 4453 82 4499 128
<< mvpdiffc >>
rect 49 492 95 632
rect 253 586 299 632
rect 457 492 503 632
rect 613 601 659 647
rect 1517 689 1563 735
rect 2157 689 2203 735
rect 861 530 907 576
rect 1065 530 1111 576
rect 1269 530 1315 576
rect 1765 539 1811 585
rect 1909 539 1955 585
rect 3036 586 3082 632
rect 2405 521 2451 567
rect 2609 521 2655 567
rect 2813 521 2859 567
rect 3261 504 3307 550
rect 3465 586 3511 632
rect 3669 504 3715 550
rect 3873 573 3919 619
rect 4017 525 4063 665
rect 4221 525 4267 665
rect 4425 525 4471 665
<< polysilicon >>
rect 328 720 1240 760
rect 124 645 224 690
rect 328 645 428 720
rect 1140 669 1240 720
rect 732 590 832 656
rect 936 590 1036 656
rect 1140 623 1181 669
rect 1227 623 1240 669
rect 1636 677 1736 721
rect 1984 677 2084 721
rect 1140 590 1240 623
rect 1344 590 1444 656
rect 2276 720 3232 760
rect 2276 580 2376 720
rect 2480 659 2580 672
rect 2480 613 2493 659
rect 2539 613 2580 659
rect 3132 645 3232 720
rect 4092 715 4192 760
rect 4296 715 4396 760
rect 3336 645 3436 690
rect 3540 645 3640 690
rect 3744 645 3844 690
rect 2480 580 2580 613
rect 2684 580 2784 630
rect 124 415 224 472
rect 328 416 428 472
rect 124 369 145 415
rect 191 369 224 415
rect 124 288 224 369
rect 348 326 428 416
rect 732 416 832 517
rect 936 436 1036 517
rect 732 415 860 416
rect 732 369 745 415
rect 791 369 860 415
rect 732 356 860 369
rect 124 232 244 288
rect 348 280 365 326
rect 411 288 428 326
rect 788 288 860 356
rect 936 390 973 436
rect 1019 390 1036 436
rect 1140 424 1240 517
rect 1344 416 1444 517
rect 936 376 1036 390
rect 1404 380 1444 416
rect 1636 380 1736 526
rect 1984 466 2084 526
rect 936 336 1312 376
rect 1236 326 1312 336
rect 411 280 468 288
rect 348 232 468 280
rect 788 244 908 288
rect 1012 244 1132 288
rect 1236 280 1253 326
rect 1299 288 1312 326
rect 1404 367 1524 380
rect 1404 321 1417 367
rect 1463 321 1524 367
rect 1299 280 1356 288
rect 1236 244 1356 280
rect 1404 244 1524 321
rect 1572 340 1736 380
rect 1964 459 2084 466
rect 1964 413 1997 459
rect 2043 413 2084 459
rect 2276 448 2376 508
rect 1964 400 2084 413
rect 2164 408 2376 448
rect 2480 448 2580 508
rect 2684 475 2784 508
rect 2480 408 2636 448
rect 1964 344 2036 400
rect 2164 344 2204 408
rect 1572 244 1692 340
rect 1916 257 2036 344
rect 2084 257 2204 344
rect 2320 336 2440 349
rect 2320 290 2352 336
rect 2398 290 2440 336
rect 2320 257 2440 290
rect 2544 321 2636 408
rect 2684 429 2701 475
rect 2747 429 2784 475
rect 2684 407 2784 429
rect 3132 409 3232 491
rect 3336 431 3436 491
rect 3132 363 3145 409
rect 3191 363 3232 409
rect 2544 257 2664 321
rect 3132 293 3232 363
rect 124 107 244 151
rect 348 79 468 151
rect 788 127 908 171
rect 1012 79 1132 171
rect 1236 127 1356 171
rect 1404 127 1524 171
rect 348 39 1132 79
rect 1572 64 1692 171
rect 3112 232 3232 293
rect 3296 416 3436 431
rect 3296 311 3416 416
rect 3296 265 3340 311
rect 3386 265 3416 311
rect 3540 415 3640 491
rect 3540 369 3577 415
rect 3623 369 3640 415
rect 3540 293 3640 369
rect 3744 458 3844 491
rect 3744 412 3761 458
rect 3807 412 3844 458
rect 3744 399 3844 412
rect 3744 293 3812 399
rect 4092 364 4192 472
rect 4296 364 4396 472
rect 3296 232 3416 265
rect 3520 232 3640 293
rect 3692 232 3812 293
rect 4060 351 4396 364
rect 4060 305 4073 351
rect 4213 305 4396 351
rect 4060 292 4396 305
rect 4060 232 4180 292
rect 4284 276 4396 292
rect 4284 232 4404 276
rect 1916 112 2036 156
rect 2084 112 2204 156
rect 2320 112 2440 156
rect 2544 112 2664 156
rect 3112 112 3232 156
rect 3296 112 3416 156
rect 3520 64 3640 156
rect 3692 112 3812 156
rect 1572 24 3640 64
rect 4060 24 4180 69
rect 4284 24 4404 69
<< polycontact >>
rect 1181 623 1227 669
rect 2493 613 2539 659
rect 145 369 191 415
rect 745 369 791 415
rect 365 280 411 326
rect 973 390 1019 436
rect 1253 280 1299 326
rect 1417 321 1463 367
rect 1997 413 2043 459
rect 2352 290 2398 336
rect 2701 429 2747 475
rect 3145 363 3191 409
rect 3340 265 3386 311
rect 3577 369 3623 415
rect 3761 412 3807 458
rect 4073 305 4213 351
<< metal1 >>
rect 0 735 4592 844
rect 0 724 1517 735
rect 49 632 95 645
rect 241 632 311 724
rect 602 647 670 724
rect 1506 689 1517 724
rect 1563 724 2157 735
rect 1563 689 1574 724
rect 2146 689 2157 724
rect 2203 724 4592 735
rect 2203 689 2214 724
rect 241 586 253 632
rect 299 586 311 632
rect 457 632 503 645
rect 95 492 411 518
rect 49 472 411 492
rect 62 415 315 426
rect 62 369 145 415
rect 191 369 315 415
rect 62 354 315 369
rect 365 326 411 472
rect 49 280 365 302
rect 49 256 411 280
rect 602 601 613 647
rect 659 601 670 647
rect 730 622 1019 668
rect 1170 623 1181 669
rect 1227 643 1460 669
rect 1636 643 2096 678
rect 2260 643 2493 659
rect 1227 631 2493 643
rect 1227 623 1682 631
rect 1170 622 1682 623
rect 730 545 776 622
rect 503 498 776 545
rect 850 530 861 576
rect 907 530 918 576
rect 49 219 95 256
rect 457 221 503 492
rect 578 415 792 430
rect 578 369 745 415
rect 791 369 792 415
rect 578 354 792 369
rect 850 241 918 530
rect 973 436 1019 622
rect 1414 597 1682 622
rect 2049 613 2493 631
rect 2539 613 2550 659
rect 2609 624 2963 671
rect 2049 597 2306 613
rect 1065 576 1111 588
rect 1065 459 1111 530
rect 1258 530 1269 576
rect 1315 551 1326 576
rect 1754 551 1765 585
rect 1315 539 1765 551
rect 1811 539 1822 585
rect 1315 530 1822 539
rect 1258 505 1822 530
rect 1898 539 1909 585
rect 1955 551 1966 585
rect 2609 567 2655 624
rect 2394 551 2405 567
rect 1955 539 2405 551
rect 1898 521 2405 539
rect 2451 521 2462 567
rect 1898 505 2462 521
rect 1065 413 1997 459
rect 2043 413 2054 459
rect 1065 408 1207 413
rect 973 379 1019 390
rect 850 230 983 241
rect 457 210 543 221
rect 49 162 95 173
rect 262 164 273 210
rect 319 164 330 210
rect 262 60 330 164
rect 457 164 497 210
rect 457 153 543 164
rect 702 184 713 230
rect 759 184 770 230
rect 702 60 770 184
rect 850 184 937 230
rect 850 173 983 184
rect 1161 230 1207 408
rect 2256 367 2302 505
rect 2609 459 2655 521
rect 2813 567 2859 578
rect 1253 326 1299 337
rect 1406 321 1417 367
rect 1463 321 2302 367
rect 2480 412 2655 459
rect 2701 475 2747 486
rect 1253 275 1299 280
rect 1253 229 2176 275
rect 1161 173 1207 184
rect 1770 137 1781 183
rect 1827 137 1838 183
rect 1770 60 1838 137
rect 2130 152 2176 229
rect 2234 244 2302 321
rect 2234 198 2245 244
rect 2291 198 2302 244
rect 2349 336 2400 347
rect 2349 290 2352 336
rect 2398 290 2400 336
rect 2349 152 2400 290
rect 2480 244 2526 412
rect 2701 366 2747 429
rect 2458 198 2469 244
rect 2515 198 2526 244
rect 2579 320 2747 366
rect 2579 152 2625 320
rect 2813 244 2859 521
rect 2917 540 2963 624
rect 3025 632 3093 724
rect 3025 586 3036 632
rect 3082 586 3093 632
rect 3139 618 3407 665
rect 3139 540 3185 618
rect 2917 493 3185 540
rect 3237 550 3307 561
rect 3237 504 3261 550
rect 3237 493 3307 504
rect 3361 540 3407 618
rect 3454 632 3522 724
rect 3454 586 3465 632
rect 3511 586 3522 632
rect 3577 607 3807 654
rect 3577 540 3623 607
rect 3361 493 3623 540
rect 3669 550 3715 561
rect 2930 409 3191 430
rect 2930 363 3145 409
rect 2930 340 3191 363
rect 2682 198 2693 244
rect 2739 215 2859 244
rect 3237 215 3283 493
rect 3343 415 3623 430
rect 3343 369 3577 415
rect 3343 357 3623 369
rect 3669 311 3715 504
rect 3761 458 3807 607
rect 3873 619 3919 724
rect 3873 562 3919 573
rect 4017 665 4063 724
rect 4017 514 4063 525
rect 4220 665 4351 676
rect 4220 525 4221 665
rect 4267 525 4351 665
rect 4220 466 4351 525
rect 4425 665 4471 724
rect 4425 514 4471 525
rect 3761 401 3807 412
rect 4061 311 4073 351
rect 3329 265 3340 311
rect 3386 305 4073 311
rect 4213 305 4224 351
rect 3386 265 4119 305
rect 3841 215 3887 265
rect 4274 218 4351 466
rect 2739 198 3037 215
rect 2813 169 3037 198
rect 3083 169 3283 215
rect 3434 169 3445 215
rect 3491 169 3502 215
rect 2130 106 2625 152
rect 3434 60 3502 169
rect 4198 172 4209 218
rect 4255 172 4351 218
rect 3841 158 3887 169
rect 3985 142 4031 153
rect 3985 60 4031 96
rect 4442 82 4453 128
rect 4499 82 4510 128
rect 4442 60 4510 82
rect 0 -60 4592 60
<< labels >>
flabel metal1 s 3343 357 3623 430 0 FreeSans 600 0 0 0 RN
port 2 nsew default input
flabel metal1 s 578 354 792 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 4220 466 4351 676 0 FreeSans 600 0 0 0 Q
port 5 nsew default output
flabel metal1 s 62 354 315 426 0 FreeSans 600 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 702 215 770 230 0 FreeSans 600 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 0 724 4592 844 0 FreeSans 600 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2930 340 3191 430 0 FreeSans 600 0 0 0 SETN
port 3 nsew default input
rlabel metal1 s 4274 218 4351 466 1 Q
port 5 nsew default output
rlabel metal1 s 4198 172 4351 218 1 Q
port 5 nsew default output
rlabel metal1 s 4425 689 4471 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 689 4063 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3873 689 3919 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3454 689 3522 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3025 689 3093 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2146 689 2214 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1506 689 1574 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 602 689 670 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 241 689 311 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4425 601 4471 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 601 4063 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3873 601 3919 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3454 601 3522 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3025 601 3093 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 602 601 670 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 241 601 311 689 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4425 586 4471 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 586 4063 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3873 586 3919 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3454 586 3522 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3025 586 3093 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 241 586 311 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4425 562 4471 586 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 562 4063 586 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3873 562 3919 586 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4425 514 4471 562 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 514 4063 562 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3434 210 3502 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 702 210 770 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3434 183 3502 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 702 183 770 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 183 330 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3434 153 3502 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1770 153 1838 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 702 153 770 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 153 330 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3985 128 4031 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3434 128 3502 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1770 128 1838 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 702 128 770 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 128 330 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4442 60 4510 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3985 60 4031 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3434 60 3502 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1770 60 1838 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 702 60 770 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4592 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4592 784
string GDS_END 1018566
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1008420
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
