magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect 0 459 56 549
rect 0 -45 56 45
<< labels >>
rlabel metal1 s 0 459 56 549 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -45 56 45 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 56 504
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 751942
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 750908
<< end >>
