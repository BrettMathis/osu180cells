magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 5600 844
rect 49 646 95 724
rect 477 610 523 724
rect 925 610 971 724
rect 1373 610 1419 724
rect 1877 638 1923 724
rect 2101 600 2147 678
rect 2305 646 2351 724
rect 2529 600 2575 678
rect 2753 646 2799 724
rect 2977 600 3023 678
rect 3201 646 3247 724
rect 3425 600 3471 678
rect 3649 646 3695 724
rect 3873 600 3919 678
rect 4097 646 4143 724
rect 4321 600 4367 678
rect 4545 646 4591 724
rect 4769 600 4815 678
rect 4993 646 5039 724
rect 5217 600 5263 678
rect 74 348 1662 430
rect 2101 484 5263 600
rect 5441 552 5487 724
rect 3597 307 3777 484
rect 486 60 554 208
rect 934 60 1002 208
rect 1382 60 1450 208
rect 2101 243 5283 307
rect 1866 60 1934 192
rect 2101 138 2147 243
rect 2314 60 2382 197
rect 2549 138 2595 243
rect 2762 60 2830 197
rect 2997 138 3043 243
rect 3210 60 3278 197
rect 3445 138 3491 243
rect 3658 60 3726 197
rect 3893 138 3939 243
rect 4106 60 4174 197
rect 4341 138 4387 243
rect 4554 60 4622 197
rect 4789 138 4835 243
rect 5002 60 5070 197
rect 5237 138 5283 243
rect 5450 60 5518 197
rect 0 -60 5600 60
<< obsm1 >>
rect 253 552 299 678
rect 701 552 747 678
rect 1149 552 1195 678
rect 1597 552 1643 678
rect 253 506 1770 552
rect 1724 413 1770 506
rect 1724 353 3432 413
rect 1724 300 1770 353
rect 3948 353 5432 413
rect 273 254 1770 300
rect 273 148 319 254
rect 721 148 767 254
rect 1169 148 1215 254
rect 1617 148 1663 254
<< labels >>
rlabel metal1 s 74 348 1662 430 6 I
port 1 nsew default input
rlabel metal1 s 5217 600 5263 678 6 Z
port 2 nsew default output
rlabel metal1 s 4769 600 4815 678 6 Z
port 2 nsew default output
rlabel metal1 s 4321 600 4367 678 6 Z
port 2 nsew default output
rlabel metal1 s 3873 600 3919 678 6 Z
port 2 nsew default output
rlabel metal1 s 3425 600 3471 678 6 Z
port 2 nsew default output
rlabel metal1 s 2977 600 3023 678 6 Z
port 2 nsew default output
rlabel metal1 s 2529 600 2575 678 6 Z
port 2 nsew default output
rlabel metal1 s 2101 600 2147 678 6 Z
port 2 nsew default output
rlabel metal1 s 2101 484 5263 600 6 Z
port 2 nsew default output
rlabel metal1 s 3597 307 3777 484 6 Z
port 2 nsew default output
rlabel metal1 s 2101 243 5283 307 6 Z
port 2 nsew default output
rlabel metal1 s 5237 138 5283 243 6 Z
port 2 nsew default output
rlabel metal1 s 4789 138 4835 243 6 Z
port 2 nsew default output
rlabel metal1 s 4341 138 4387 243 6 Z
port 2 nsew default output
rlabel metal1 s 3893 138 3939 243 6 Z
port 2 nsew default output
rlabel metal1 s 3445 138 3491 243 6 Z
port 2 nsew default output
rlabel metal1 s 2997 138 3043 243 6 Z
port 2 nsew default output
rlabel metal1 s 2549 138 2595 243 6 Z
port 2 nsew default output
rlabel metal1 s 2101 138 2147 243 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 5600 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5441 646 5487 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4993 646 5039 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4545 646 4591 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4097 646 4143 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3649 646 3695 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3201 646 3247 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2753 646 2799 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2305 646 2351 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1877 646 1923 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5441 638 5487 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1877 638 1923 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 638 1419 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 638 971 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 638 523 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5441 610 5487 638 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 610 1419 638 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 610 971 638 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 610 523 638 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5441 552 5487 610 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1382 197 1450 208 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 197 1002 208 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 197 554 208 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5450 192 5518 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5002 192 5070 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4554 192 4622 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4106 192 4174 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3658 192 3726 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3210 192 3278 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2762 192 2830 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2314 192 2382 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 192 1450 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 192 1002 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 192 554 197 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5450 60 5518 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5002 60 5070 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4554 60 4622 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4106 60 4174 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3658 60 3726 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3210 60 3278 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2762 60 2830 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2314 60 2382 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1866 60 1934 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 192 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5600 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5600 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 785380
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 773856
<< end >>
