magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect 303 3049 496 3094
rect 303 3003 377 3049
rect 423 3003 496 3049
rect 303 2957 496 3003
rect 1423 3049 1616 3094
rect 1423 3003 1497 3049
rect 1543 3003 1616 3049
rect 1423 2957 1616 3003
rect 1936 3049 2129 3094
rect 1936 3003 2010 3049
rect 2056 3003 2129 3049
rect 1936 2957 2129 3003
rect 3056 3049 3249 3094
rect 3056 3003 3130 3049
rect 3176 3003 3249 3049
rect 3056 2957 3249 3003
rect 527 2850 720 2895
rect 527 2804 601 2850
rect 647 2804 720 2850
rect 527 2758 720 2804
rect 1199 2850 1392 2895
rect 1199 2804 1273 2850
rect 1319 2804 1392 2850
rect 1199 2758 1392 2804
rect 3794 2850 3987 2895
rect 3794 2804 3868 2850
rect 3914 2804 3987 2850
rect 3794 2758 3987 2804
rect 4466 2850 4659 2895
rect 4466 2804 4540 2850
rect 4586 2804 4659 2850
rect 4466 2758 4659 2804
rect 751 2646 944 2691
rect 751 2600 825 2646
rect 871 2600 944 2646
rect 751 2554 944 2600
rect 2384 2646 2577 2691
rect 2384 2600 2458 2646
rect 2504 2600 2577 2646
rect 2384 2554 2577 2600
rect 4018 2646 4211 2691
rect 4018 2600 4092 2646
rect 4138 2600 4211 2646
rect 4018 2554 4211 2600
rect 5652 2646 5845 2691
rect 5652 2600 5726 2646
rect 5772 2600 5845 2646
rect 5652 2554 5845 2600
rect 3570 2444 3763 2489
rect 3570 2398 3644 2444
rect 3690 2398 3763 2444
rect 3570 2352 3763 2398
rect 4690 2444 4883 2489
rect 4690 2398 4764 2444
rect 4810 2398 4883 2444
rect 4690 2352 4883 2398
rect 5204 2444 5397 2489
rect 5204 2398 5278 2444
rect 5324 2398 5397 2444
rect 5204 2352 5397 2398
rect 6324 2444 6517 2489
rect 6324 2398 6398 2444
rect 6444 2398 6517 2444
rect 6324 2352 6517 2398
rect 2160 2242 2353 2287
rect 2160 2196 2234 2242
rect 2280 2196 2353 2242
rect 2160 2150 2353 2196
rect 2832 2242 3025 2287
rect 2832 2196 2906 2242
rect 2952 2196 3025 2242
rect 2832 2150 3025 2196
rect 5428 2242 5621 2287
rect 5428 2196 5502 2242
rect 5548 2196 5621 2242
rect 5428 2150 5621 2196
rect 6100 2242 6293 2287
rect 6100 2196 6174 2242
rect 6220 2196 6293 2242
rect 6100 2150 6293 2196
rect 975 2041 1168 2086
rect 975 1995 1049 2041
rect 1095 1995 1168 2041
rect 975 1949 1168 1995
rect 2608 2041 2801 2086
rect 2608 1995 2682 2041
rect 2728 1995 2801 2041
rect 2608 1949 2801 1995
rect 4242 2041 4435 2086
rect 4242 1995 4316 2041
rect 4362 1995 4435 2041
rect 4242 1949 4435 1995
rect 5876 2041 6069 2086
rect 5876 1995 5950 2041
rect 5996 1995 6069 2041
rect 5876 1949 6069 1995
<< polycontact >>
rect 377 3003 423 3049
rect 1497 3003 1543 3049
rect 2010 3003 2056 3049
rect 3130 3003 3176 3049
rect 601 2804 647 2850
rect 1273 2804 1319 2850
rect 3868 2804 3914 2850
rect 4540 2804 4586 2850
rect 825 2600 871 2646
rect 2458 2600 2504 2646
rect 4092 2600 4138 2646
rect 5726 2600 5772 2646
rect 3644 2398 3690 2444
rect 4764 2398 4810 2444
rect 5278 2398 5324 2444
rect 6398 2398 6444 2444
rect 2234 2196 2280 2242
rect 2906 2196 2952 2242
rect 5502 2196 5548 2242
rect 6174 2196 6220 2242
rect 1049 1995 1095 2041
rect 2682 1995 2728 2041
rect 4316 1995 4362 2041
rect 5950 1995 5996 2041
<< metal1 >>
rect 342 3049 457 3085
rect 342 3003 377 3049
rect 423 3003 457 3049
rect 342 2966 457 3003
rect 1462 3049 1577 3085
rect 1462 3003 1497 3049
rect 1543 3003 1577 3049
rect 1462 2966 1577 3003
rect 1975 3049 2090 3085
rect 1975 3003 2010 3049
rect 2056 3003 2090 3049
rect 1975 2966 2090 3003
rect 3095 3049 3210 3085
rect 3095 3003 3130 3049
rect 3176 3003 3210 3049
rect 3095 2966 3210 3003
rect 566 2850 681 2886
rect 566 2804 601 2850
rect 647 2804 681 2850
rect 566 2767 681 2804
rect 1238 2850 1353 2886
rect 1238 2804 1273 2850
rect 1319 2804 1353 2850
rect 1238 2767 1353 2804
rect 3833 2850 3948 2886
rect 3833 2804 3868 2850
rect 3914 2804 3948 2850
rect 3833 2767 3948 2804
rect 4505 2850 4620 2886
rect 4505 2804 4540 2850
rect 4586 2804 4620 2850
rect 4505 2767 4620 2804
rect 790 2646 905 2682
rect 790 2600 825 2646
rect 871 2600 905 2646
rect 790 2563 905 2600
rect 2423 2646 2538 2682
rect 2423 2600 2458 2646
rect 2504 2600 2538 2646
rect 2423 2563 2538 2600
rect 4057 2646 4172 2682
rect 4057 2600 4092 2646
rect 4138 2600 4172 2646
rect 4057 2563 4172 2600
rect 5691 2646 5806 2682
rect 5691 2600 5726 2646
rect 5772 2600 5806 2646
rect 5691 2563 5806 2600
rect 3609 2444 3724 2480
rect 3609 2398 3644 2444
rect 3690 2398 3724 2444
rect 3609 2361 3724 2398
rect 4729 2444 4844 2480
rect 4729 2398 4764 2444
rect 4810 2398 4844 2444
rect 4729 2361 4844 2398
rect 5243 2444 5358 2480
rect 5243 2398 5278 2444
rect 5324 2398 5358 2444
rect 5243 2361 5358 2398
rect 6363 2444 6478 2480
rect 6363 2398 6398 2444
rect 6444 2398 6478 2444
rect 6363 2361 6478 2398
rect 2199 2242 2314 2278
rect 2199 2196 2234 2242
rect 2280 2196 2314 2242
rect 2199 2159 2314 2196
rect 2871 2242 2986 2278
rect 2871 2196 2906 2242
rect 2952 2196 2986 2242
rect 2871 2159 2986 2196
rect 5467 2242 5582 2278
rect 5467 2196 5502 2242
rect 5548 2196 5582 2242
rect 5467 2159 5582 2196
rect 6139 2242 6254 2278
rect 6139 2196 6174 2242
rect 6220 2196 6254 2242
rect 6139 2159 6254 2196
rect 1014 2041 1129 2077
rect 1014 1995 1049 2041
rect 1095 1995 1129 2041
rect 1014 1958 1129 1995
rect 2647 2041 2762 2077
rect 2647 1995 2682 2041
rect 2728 1995 2762 2041
rect 2647 1958 2762 1995
rect 4281 2041 4396 2077
rect 4281 1995 4316 2041
rect 4362 1995 4396 2041
rect 4281 1958 4396 1995
rect 5915 2041 6030 2077
rect 5915 1995 5950 2041
rect 5996 1995 6030 2041
rect 5915 1958 6030 1995
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1669390400
transform 1 0 4563 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1669390400
transform 1 0 3891 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1669390400
transform 1 0 400 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1669390400
transform 1 0 1520 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1669390400
transform 1 0 5749 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1669390400
transform 1 0 5973 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1669390400
transform 1 0 1072 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_7
timestamp 1669390400
transform 1 0 848 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_8
timestamp 1669390400
transform 1 0 4787 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_9
timestamp 1669390400
transform 1 0 3667 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_10
timestamp 1669390400
transform 1 0 5525 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_11
timestamp 1669390400
transform 1 0 6197 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_12
timestamp 1669390400
transform 1 0 2929 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_13
timestamp 1669390400
transform 1 0 2257 0 1 2219
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_14
timestamp 1669390400
transform 1 0 2705 0 1 2018
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_15
timestamp 1669390400
transform 1 0 2481 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_16
timestamp 1669390400
transform 1 0 6421 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_17
timestamp 1669390400
transform 1 0 3153 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_18
timestamp 1669390400
transform 1 0 2033 0 1 3026
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_19
timestamp 1669390400
transform 1 0 5301 0 1 2421
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_20
timestamp 1669390400
transform 1 0 1296 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_21
timestamp 1669390400
transform 1 0 624 0 1 2827
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_22
timestamp 1669390400
transform 1 0 4115 0 1 2623
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_23
timestamp 1669390400
transform 1 0 4339 0 1 2018
box 0 0 1 1
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_0
timestamp 1669390400
transform 1 0 2594 0 1 1002
box -38 -506 38 506
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_1
timestamp 1669390400
transform 1 0 4227 0 1 1002
box -38 -506 38 506
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_2
timestamp 1669390400
transform 1 0 5861 0 1 1002
box -38 -506 38 506
use M2_M14310590878151_256x8m81  M2_M14310590878151_256x8m81_3
timestamp 1669390400
transform 1 0 960 0 1 1002
box -38 -506 38 506
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_0
timestamp 1669390400
transform 1 0 960 0 1 1002
box -38 -506 38 506
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_1
timestamp 1669390400
transform 1 0 4227 0 1 1002
box -38 -506 38 506
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_2
timestamp 1669390400
transform 1 0 5861 0 1 1002
box -38 -506 38 506
use M3_M24310590878152_256x8m81  M3_M24310590878152_256x8m81_3
timestamp 1669390400
transform 1 0 2594 0 1 1002
box -38 -506 38 506
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_0
timestamp 1669390400
transform -1 0 4372 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_1
timestamp 1669390400
transform -1 0 6006 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_2
timestamp 1669390400
transform -1 0 2738 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_3
timestamp 1669390400
transform -1 0 1105 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_4
timestamp 1669390400
transform 1 0 4082 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_5
timestamp 1669390400
transform 1 0 5716 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_6
timestamp 1669390400
transform 1 0 2448 0 1 7069
box -144 -7124 1106 327
use ypredec1_xa_256x8m81  ypredec1_xa_256x8m81_7
timestamp 1669390400
transform 1 0 815 0 1 7069
box -144 -7124 1106 327
<< properties >>
string GDS_END 967878
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 965786
<< end >>
