****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__addf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addf_1 A B CI S CO VDD VSS
X0 a_110_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 S a_161_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 S a_161_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD CI a_195_109# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_195_19# B a_178_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_76_109# B a_59_19# VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_76_109# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_59_19# CI a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_178_19# A a_161_19# VSS nmos_3p3 w=0.85u l=0.3u
X9 a_9_109# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 a_110_19# CI VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VDD A a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X12 a_59_19# CI a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS B a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X14 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 CO a_59_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS CI a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X17 CO a_59_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X18 VSS A a_76_19# VSS nmos_3p3 w=0.85u l=0.3u
X19 a_161_19# a_59_19# a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_76_19# B a_59_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_178_109# A a_161_19# VDD pmos_3p3 w=1.7u l=0.3u
X22 a_195_109# B a_178_109# VDD pmos_3p3 w=1.7u l=0.3u
X23 a_9_19# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X24 a_110_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 a_161_19# a_59_19# a_110_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 VDD B a_110_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_110_109# CI VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__addf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__addh_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addh_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addh_1 A B S CO VDD VSS
X0 VDD B a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_19_14# CO VDD pmos_3p3 w=1.7u l=0.3u
X3 a_19_14# B a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 S a_91_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS a_19_14# CO VSS nmos_3p3 w=0.85u l=0.3u
X6 S a_91_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 a_91_19# B a_91_109# VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_19_14# a_91_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_91_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 a_91_19# A a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_19_14# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_75_19# B a_91_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__addh_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__and2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__and2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__and2_1 A B Y VDD VSS
X0 Y a_12_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD B a_12_19# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_12_19# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_12_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 a_28_19# A a_12_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS B a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__and2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__aoi21_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__aoi21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__aoi21_1 A0 A1 B Y VDD VSS
X0 Y B a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_9_109# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A0 a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS B Y VSS nmos_3p3 w=0.85u l=0.3u
X4 a_28_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 Y A1 a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__aoi21_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__aoi22_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__aoi22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__aoi22_1 Y A0 A1 B0 B1
X0 a_9_109# B1 Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y B0 a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_9_109# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD A0 a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_56_19# B0 Y VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS B1 a_56_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_28_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 Y A1 a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__aoi22_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_1 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_16 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X14 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X17 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X18 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X20 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X21 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X22 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X23 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X24 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X26 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X27 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X29 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X30 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X31 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X32 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X33 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_2 A Y VDD VSS
X0 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_4 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__buf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__buf_8 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X8 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X16 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X17 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__buf_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_1 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_16 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X14 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X17 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X18 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X20 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X21 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X22 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X23 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X24 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X26 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X27 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X29 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X30 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X31 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X32 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X33 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_2 A Y VDD VSS
X0 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_4 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkbuf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_8 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X8 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X16 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X17 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkbuf_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_1 A Y VDD VSS
X0 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_16 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X6 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X11 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X17 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X18 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X20 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X22 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X23 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X24 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X26 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X27 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X28 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X29 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X30 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X31 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_2 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_4 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__clkinv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__clkinv_8 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X8 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X15 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__clkinv_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dff_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dff_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dff_1 D Q QN CLK VDD VSS
X0 a_75_109# a_52_14# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# CLK a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_135_68# a_114_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 a_131_19# a_52_14# a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_42_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 a_135_68# a_114_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_75_19# CLK a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X9 VSS a_135_68# a_131_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 a_19_14# a_52_14# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X12 a_52_14# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 VDD a_135_68# a_131_109# VDD pmos_3p3 w=1.7u l=0.3u
X14 a_131_109# CLK a_114_19# VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS a_135_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X16 a_114_19# a_52_14# a_103_109# VDD pmos_3p3 w=1.7u l=0.3u
X17 a_114_19# CLK a_103_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 a_52_14# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 a_103_109# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X20 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD a_9_19# a_75_109# VDD pmos_3p3 w=1.7u l=0.3u
X22 a_103_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 VDD a_135_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X25 VSS a_9_19# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dff_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffn_1 Q QN D CLK VDD VSS
X0 a_75_109# a_52_14# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# a_52_81# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_131_19# a_52_14# a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 a_42_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_75_19# a_52_81# a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X6 VDD a_135_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X7 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 VSS a_135_68# a_131_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 a_19_14# a_52_14# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_135_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X13 a_52_14# a_52_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD a_135_68# a_131_109# VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS CLK a_52_81# VSS nmos_3p3 w=0.85u l=0.3u
X16 a_131_109# a_52_81# a_114_19# VDD pmos_3p3 w=1.7u l=0.3u
X17 a_114_19# a_52_14# a_103_109# VDD pmos_3p3 w=1.7u l=0.3u
X18 a_135_68# a_114_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 a_114_19# a_52_81# a_103_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_52_14# a_52_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X21 a_103_109# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD a_9_19# a_75_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_103_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 a_135_68# a_114_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X26 VDD CLK a_52_81# VDD pmos_3p3 w=1.7u l=0.3u
X27 VSS a_9_19# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffr_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffr_1 D Q QN CLK RN VDD VSS
X0 VDD a_41_109# a_145_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_173_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_122_14# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_122_14# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_205_68# a_201_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_62_98# CLK a_112_109# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_145_109# a_122_14# a_62_98# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_145_19# CLK a_62_98# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 a_62_98# a_122_14# a_112_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_112_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_205_68# a_184_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 VDD a_205_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X15 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 a_201_19# a_122_14# a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X17 VSS a_205_68# a_201_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 a_205_68# a_25_19# a_273_109# VDD pmos_3p3 w=1.7u l=0.3u
X20 a_273_109# a_184_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X21 VSS a_205_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X22 VSS a_62_98# a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD a_62_98# a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_112_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS a_25_19# a_205_68# VSS nmos_3p3 w=0.85u l=0.3u
X26 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_173_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 a_201_109# CLK a_184_19# VDD pmos_3p3 w=1.7u l=0.3u
X29 a_184_19# a_122_14# a_173_109# VDD pmos_3p3 w=1.7u l=0.3u
X30 VSS a_41_109# a_145_19# VSS nmos_3p3 w=0.85u l=0.3u
X31 a_184_19# CLK a_173_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffr_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffrn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffrn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffrn_1 D Q QN RN CLK VDD VSS
X0 VDD a_41_109# a_145_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_173_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_122_14# a_122_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_122_14# a_122_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_205_68# a_201_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_205_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X6 a_62_98# a_122_81# a_112_109# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_145_109# a_122_14# a_62_98# VDD pmos_3p3 w=1.7u l=0.3u
X8 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD a_205_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X10 a_145_19# a_122_81# a_62_98# VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_25_19# a_205_68# VSS nmos_3p3 w=0.85u l=0.3u
X12 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 a_62_98# a_122_14# a_112_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 VDD CLK a_122_81# VDD pmos_3p3 w=1.7u l=0.3u
X16 VSS CLK a_122_81# VSS nmos_3p3 w=0.85u l=0.3u
X17 a_205_68# a_184_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X18 a_112_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X20 a_201_19# a_122_14# a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 VSS a_205_68# a_201_19# VSS nmos_3p3 w=0.85u l=0.3u
X22 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 a_205_68# a_25_19# a_306_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_306_109# a_184_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X25 VSS a_62_98# a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X26 VDD a_62_98# a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_112_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X29 a_173_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X30 a_201_109# a_122_81# a_184_19# VDD pmos_3p3 w=1.7u l=0.3u
X31 a_184_19# a_122_14# a_173_109# VDD pmos_3p3 w=1.7u l=0.3u
X32 VSS a_41_109# a_145_19# VSS nmos_3p3 w=0.85u l=0.3u
X33 a_184_19# a_122_81# a_173_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffrn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffs_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffs_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffs_1 D Q QN SN CLK VDD VSS
X0 a_75_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_227_19# a_147_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 a_208_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS SN a_108_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD a_147_19# a_208_109# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_85_14# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_168_68# SN a_227_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_75_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 a_85_14# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_168_68# a_164_109# VDD pmos_3p3 w=1.7u l=0.3u
X11 VDD SN SN VDD pmos_3p3 w=1.7u l=0.3u
X12 SN a_34_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 a_147_19# a_85_14# a_136_109# VDD pmos_3p3 w=1.7u l=0.3u
X14 a_164_109# CLK a_147_19# VDD pmos_3p3 w=1.7u l=0.3u
X15 a_136_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 a_136_19# SN VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 VDD SN a_108_109# VDD pmos_3p3 w=1.7u l=0.3u
X18 VSS a_168_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X19 a_108_109# a_85_14# a_34_14# VDD pmos_3p3 w=1.7u l=0.3u
X20 a_164_19# a_85_14# a_147_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 VDD a_168_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X23 a_147_19# CLK a_136_19# VSS nmos_3p3 w=0.85u l=0.3u
X24 VSS a_168_68# a_164_19# VSS nmos_3p3 w=0.85u l=0.3u
X25 a_34_14# CLK a_75_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 a_29_19# SN SN VSS nmos_3p3 w=0.85u l=0.3u
X27 a_34_14# a_85_14# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X28 VSS a_34_14# a_29_19# VSS nmos_3p3 w=0.85u l=0.3u
X29 a_108_19# CLK a_34_14# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffs_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsn_1 D Q QN CLK SN VDD VSS
X0 a_75_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD a_147_19# a_242_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_242_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS SN a_108_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS CLK a_85_81# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_85_14# a_85_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_75_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_85_14# a_85_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_168_68# a_164_109# VDD pmos_3p3 w=1.7u l=0.3u
X9 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 VDD SN SN VDD pmos_3p3 w=1.7u l=0.3u
X11 SN a_34_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_147_19# a_85_14# a_136_109# VDD pmos_3p3 w=1.7u l=0.3u
X13 a_164_109# a_85_81# a_147_19# VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD CLK a_85_81# VDD pmos_3p3 w=1.7u l=0.3u
X15 a_261_19# a_147_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS a_168_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X17 a_136_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X18 a_136_19# SN VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 VDD SN a_108_109# VDD pmos_3p3 w=1.7u l=0.3u
X20 a_108_109# a_85_14# a_34_14# VDD pmos_3p3 w=1.7u l=0.3u
X21 a_164_19# a_85_14# a_147_19# VSS nmos_3p3 w=0.85u l=0.3u
X22 a_168_68# SN a_261_19# VSS nmos_3p3 w=0.85u l=0.3u
X23 a_147_19# a_85_81# a_136_19# VSS nmos_3p3 w=0.85u l=0.3u
X24 VSS a_168_68# a_164_19# VSS nmos_3p3 w=0.85u l=0.3u
X25 a_34_14# a_85_81# a_75_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 a_29_19# SN SN VSS nmos_3p3 w=0.85u l=0.3u
X27 a_34_14# a_85_14# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X28 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X29 VDD a_168_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X30 VSS a_34_14# a_29_19# VSS nmos_3p3 w=0.85u l=0.3u
X31 a_108_19# a_85_81# a_34_14# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsr_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsr_1 D Q QN RN SN CLK VDD VSS
X0 a_156_109# a_133_14# a_82_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_41_109# a_156_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 a_82_14# CLK a_123_109# VDD pmos_3p3 w=1.7u l=0.3u
X3 a_212_109# CLK a_195_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS a_25_19# a_216_68# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_195_19# CLK a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_133_14# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_216_68# SN a_275_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 a_123_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_216_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X11 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 a_82_14# a_133_14# a_123_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 a_256_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 a_275_19# a_195_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 VDD a_195_19# a_256_109# VDD pmos_3p3 w=1.7u l=0.3u
X18 a_212_19# a_133_14# a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X19 a_216_68# a_25_19# a_256_109# VDD pmos_3p3 w=1.7u l=0.3u
X20 VSS a_216_68# a_212_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_77_19# SN a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X22 a_57_109# a_82_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X23 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 VDD SN a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X25 a_195_19# a_133_14# a_184_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X27 a_184_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X28 VSS a_82_14# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X29 a_156_19# CLK a_82_14# VSS nmos_3p3 w=0.85u l=0.3u
X30 VDD a_41_109# a_156_109# VDD pmos_3p3 w=1.7u l=0.3u
X31 a_133_14# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X32 a_123_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X33 VDD a_216_68# a_212_109# VDD pmos_3p3 w=1.7u l=0.3u
X34 a_184_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X35 VSS a_216_68# QN VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsr_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsrn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsrn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsrn_1 D Q QN CLK RN SN VDD VSS
X0 a_156_109# a_133_14# a_82_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_41_109# a_156_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 a_82_14# a_133_81# a_123_109# VDD pmos_3p3 w=1.7u l=0.3u
X3 a_212_109# a_133_81# a_195_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD CLK a_133_81# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_195_19# a_133_81# a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_133_14# a_133_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 a_123_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS a_216_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X11 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_310_19# a_195_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 VDD a_216_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X14 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 a_82_14# a_133_14# a_123_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS CLK a_133_81# VSS nmos_3p3 w=0.85u l=0.3u
X17 a_216_68# SN a_310_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 a_212_19# a_133_14# a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X19 VSS a_216_68# a_212_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_77_19# SN a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_57_109# a_82_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 a_216_68# a_25_19# a_291_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X25 VDD SN a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 a_195_19# a_133_14# a_184_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_291_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X28 VDD a_195_19# a_291_109# VDD pmos_3p3 w=1.7u l=0.3u
X29 a_184_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X30 VSS a_82_14# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X31 a_156_19# a_133_81# a_82_14# VSS nmos_3p3 w=0.85u l=0.3u
X32 VDD a_41_109# a_156_109# VDD pmos_3p3 w=1.7u l=0.3u
X33 a_133_14# a_133_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X34 a_123_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X35 VDD a_216_68# a_212_109# VDD pmos_3p3 w=1.7u l=0.3u
X36 a_184_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X37 VSS a_25_19# a_216_68# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dffsrn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dlat_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dlat_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dlat_1 D Q CLK VDD VSS
X0 a_52_92# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_46_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_20_14# CLK a_46_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS a_10_19# a_127_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_10_19# a_77_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_77_109# CLK a_20_14# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_20_14# a_52_92# a_43_109# VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD a_20_14# a_10_19# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_43_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 Q a_127_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_10_19# a_127_19# VDD pmos_3p3 w=1.7u l=0.3u
X11 a_77_19# a_52_92# a_20_14# VSS nmos_3p3 w=0.85u l=0.3u
X12 Q a_127_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS a_10_19# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X14 a_52_92# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS a_20_14# a_10_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dlat_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__dlatn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dlatn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dlatn_1 D Q CLK VDD VSS
X0 VDD CLK a_54_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 Q a_161_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_52_92# a_54_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS CLK a_54_14# VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS a_10_19# a_161_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_46_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_20_14# a_54_14# a_46_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_10_19# a_77_109# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_77_109# a_54_14# a_20_14# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_20_14# a_52_92# a_43_109# VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_20_14# a_10_19# VDD pmos_3p3 w=1.7u l=0.3u
X11 a_43_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 VDD a_10_19# a_161_19# VDD pmos_3p3 w=1.7u l=0.3u
X13 Q a_161_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 a_77_19# a_52_92# a_20_14# VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS a_10_19# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 a_52_92# a_54_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 VSS a_20_14# a_10_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__dlatn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_1 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_16 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_2 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_4 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__fill_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__fill_8 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__fill_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_1 A Y VDD VSS
X0 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_16 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X6 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X11 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X17 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X18 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X20 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X22 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X23 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X24 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X26 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X27 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X28 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X29 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X30 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X31 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_2 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_4 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_8 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X8 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X13 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X15 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__inv_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__lshifdown.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__lshifdown.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__lshifdown A Y VDDH VDD VSS
X0 a_26_19# A VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X1 Y a_26_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y a_26_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_26_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__lshifdown.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__lshifup.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__lshifup.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__lshifup A Y VDDH VDD VSS
X0 a_26_19# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS A a_67_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 Y a_67_19# VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X3 Y a_67_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 VDDH a_78_82# a_67_19# VDDH pmos_3p3 w=1.7u l=0.3u
X5 a_78_82# a_67_19# VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X6 a_26_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_78_82# a_26_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__lshifup.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__mux2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__mux2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__mux2_1 A B Y Sel VDD VSS
X0 B a_25_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y Sel A VDD pmos_3p3 w=1.7u l=0.3u
X2 a_25_19# Sel VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_25_19# A VSS nmos_3p3 w=0.85u l=0.3u
X4 a_25_19# Sel VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 B Sel Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__mux2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__nand2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nand2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__nand2_1 A B Y VDD VSS
X0 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_28_19# A Y VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS B a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__nand2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__nor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__nor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__nor2_1 A B Y VDD VSS
X0 Y B a_25_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_25_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS B Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__nor2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__oai21_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai21_1 A0 A1 B Y VDD VSS
X0 Y B a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 VSS A0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 a_27_109# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A1 a_27_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_8_19# A1 VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__oai21_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__oai22_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai22_1 A0 A1 B0 B1 Y VDD VSS
X0 a_8_19# B1 Y VSS nmos_3p3 w=0.85u l=0.3u
X1 Y B0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 VSS A0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD B1 a_56_109# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_27_109# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 a_56_109# B0 Y VDD pmos_3p3 w=1.7u l=0.3u
X6 Y A1 a_27_109# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_8_19# A1 VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__oai22_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__oai31_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__oai31_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__oai31_1 A0 A1 A2 B Y VDD VSS
X0 a_35_109# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_25_19# A2 VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_25_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 Y B a_25_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 Y A2 a_46_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X6 VSS A1 a_25_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 a_46_109# A1 a_35_109# VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__oai31_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__or2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__or2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__or2_1 A B Y VDD VSS
X0 VDD B a_25_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_25_109# A a_9_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 a_9_109# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y a_9_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS B a_9_109# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__or2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__tbuf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tbuf_1 A Y EN VDD VSS
X0 Y EN a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 Y a_47_94# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_42_109# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_47_94# EN VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_47_94# EN VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 a_42_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__tbuf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__tieh.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tieh.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tieh Y VDD VSS
X0 Y a_19_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# a_19_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__tieh.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__tiel.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tiel.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tiel Y VDD VSS
X0 a_19_14# a_19_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_19_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__tiel.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__tinv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__tinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__tinv_1 A Y EN VDD VSS
X0 Y EN a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 Y a_9_19# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_42_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD EN a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS EN a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__tinv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__xnor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__xnor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__xnor2_1 A B Y VDD VSS
X0 Y a_47_14# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 VDD B a_76_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_47_14# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_47_14# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_76_109# A Y VDD pmos_3p3 w=1.7u l=0.3u
X5 a_42_109# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_76_19# a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X9 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 a_47_14# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS B a_76_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__xnor2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp12t3v3__xor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__xor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__xor2_1 A B Y VDD VSS
X0 Y B a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 VDD B a_76_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_47_94# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_47_94# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_76_109# a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X5 a_42_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_76_19# a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X9 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 a_47_94# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_47_94# a_76_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp12t3v3__xor2_1.spice
