magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 448 300
<< mvpmos >>
rect 0 0 240 180
<< mvpdiff >>
rect -88 167 0 180
rect -88 121 -75 167
rect -29 121 0 167
rect -88 59 0 121
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 240 167 328 180
rect 240 121 269 167
rect 315 121 328 167
rect 240 59 328 121
rect 240 13 269 59
rect 315 13 328 59
rect 240 0 328 13
<< mvpdiffc >>
rect -75 121 -29 167
rect -75 13 -29 59
rect 269 121 315 167
rect 269 13 315 59
<< polysilicon >>
rect 0 180 240 224
rect 0 -44 240 0
<< metal1 >>
rect -75 167 -29 180
rect -75 59 -29 121
rect -75 0 -29 13
rect 269 167 315 180
rect 269 59 315 121
rect 269 0 315 13
<< labels >>
flabel metal1 s -52 90 -52 90 0 FreeSans 400 0 0 0 S
flabel metal1 s 292 90 292 90 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 1066092
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1064876
<< end >>
