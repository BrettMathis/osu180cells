magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
use 3LM_METAL_RAIL  3LM_METAL_RAIL_0
timestamp 1669390400
transform 1 0 0 0 1 0
box -32 13097 15032 69968
use Bondpad_3LM  Bondpad_3LM_0
timestamp 1669390400
transform 1 0 1100 0 1 0
box -400 0 13200 13065
<< properties >>
string GDS_END 148204
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 148126
<< end >>
