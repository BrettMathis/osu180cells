magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 2206
<< mvpmos >>
rect 0 0 120 2086
<< mvpdiff >>
rect -88 2073 0 2086
rect -88 13 -75 2073
rect -29 13 0 2073
rect -88 0 0 13
rect 120 2073 208 2086
rect 120 13 149 2073
rect 195 13 208 2073
rect 120 0 208 13
<< mvpdiffc >>
rect -75 13 -29 2073
rect 149 13 195 2073
<< polysilicon >>
rect 0 2086 120 2130
rect 0 -44 120 0
<< metal1 >>
rect -75 2073 -29 2086
rect -75 0 -29 13
rect 149 2073 195 2086
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1043 -52 1043 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1043 172 1043 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 169732
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 166084
<< end >>
