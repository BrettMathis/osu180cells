magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 3792 28769 6188 28903
rect 3761 23673 5873 23868
<< metal2 >>
rect 4045 2101 5045 52645
<< metal3 >>
rect 3339 36945 6351 37145
rect 3339 36835 4353 36945
rect 3339 36355 6350 36835
rect 3339 34134 6350 35944
rect 3339 31533 5045 34134
rect 3339 31249 6632 31533
rect 3339 28254 6350 30235
rect 3339 25199 5045 25757
rect 3339 24757 6350 25199
rect 3339 23646 6350 24101
rect 3339 23101 4353 23646
rect 3339 19835 6350 22558
rect 3339 16147 6350 19549
rect 3339 15280 6350 15997
rect 3339 14665 5045 15280
rect 3339 13855 6350 14665
rect 3339 11995 6350 13312
rect 3339 9971 6350 11333
rect 3339 8801 6350 9415
rect 3339 8018 4353 8801
rect 3339 7585 6350 8018
rect 3339 6992 6350 7448
rect 3339 6334 5051 6992
rect 3339 5879 6350 6334
rect 3339 5239 6350 5591
rect 3339 4673 4339 5239
rect 3339 4321 6350 4673
rect 3339 3051 6350 4051
use M2_M14310590878181_256x8m81  M2_M14310590878181_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 36745
box -162 -348 162 348
use M2_M14310590878183_256x8m81  M2_M14310590878183_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 4942
box -162 -596 162 596
use M2_M14310590878183_256x8m81  M2_M14310590878183_256x8m81_1
timestamp 1669390400
transform 1 0 3783 0 1 12642
box -162 -596 162 596
use M2_M14310590878184_256x8m81  M2_M14310590878184_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 23602
box -162 -472 162 472
use M2_M14310590878193_256x8m81  M2_M14310590878193_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 17867
box -162 -1650 162 1650
use M2_M14310590878194_256x8m81  M2_M14310590878194_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 8496
box -162 -906 162 906
use M2_M14310590878194_256x8m81  M2_M14310590878194_256x8m81_1
timestamp 1669390400
transform 1 0 3783 0 1 29263
box -162 -906 162 906
use M3_M24310590878180_256x8m81  M3_M24310590878180_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 3548
box -472 -472 472 472
use M3_M24310590878180_256x8m81  M3_M24310590878180_256x8m81_1
timestamp 1669390400
transform 1 0 4557 0 1 25229
box -472 -472 472 472
use M3_M24310590878182_256x8m81  M3_M24310590878182_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 36745
box -162 -348 162 348
use M3_M24310590878185_256x8m81  M3_M24310590878185_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 6663
box -472 -782 472 782
use M3_M24310590878186_256x8m81  M3_M24310590878186_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 33607
box -472 -2332 472 2332
use M3_M24310590878187_256x8m81  M3_M24310590878187_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 17867
box -162 -1650 162 1650
use M3_M24310590878188_256x8m81  M3_M24310590878188_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 23602
box -162 -472 162 472
use M3_M24310590878189_256x8m81  M3_M24310590878189_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 8496
box -162 -906 162 906
use M3_M24310590878189_256x8m81  M3_M24310590878189_256x8m81_1
timestamp 1669390400
transform 1 0 3783 0 1 29263
box -162 -906 162 906
use M3_M24310590878190_256x8m81  M3_M24310590878190_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 14922
box -472 -1030 472 1030
use M3_M24310590878191_256x8m81  M3_M24310590878191_256x8m81_0
timestamp 1669390400
transform 1 0 3783 0 1 4942
box -162 -596 162 596
use M3_M24310590878191_256x8m81  M3_M24310590878191_256x8m81_1
timestamp 1669390400
transform 1 0 3783 0 1 12642
box -162 -596 162 596
use M3_M24310590878192_256x8m81  M3_M24310590878192_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 10644
box -472 -658 472 658
use M3_M24310590878195_256x8m81  M3_M24310590878195_256x8m81_0
timestamp 1669390400
transform 1 0 4557 0 1 21182
box -472 -1340 472 1340
<< properties >>
string GDS_END 1798900
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1796252
<< end >>
