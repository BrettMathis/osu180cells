magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -80 2553 80 2612
rect -80 2507 -23 2553
rect 23 2507 80 2553
rect -80 2390 80 2507
rect -80 2344 -23 2390
rect 23 2344 80 2390
rect -80 2227 80 2344
rect -80 2181 -23 2227
rect 23 2181 80 2227
rect -80 2064 80 2181
rect -80 2018 -23 2064
rect 23 2018 80 2064
rect -80 1900 80 2018
rect -80 1854 -23 1900
rect 23 1854 80 1900
rect -80 1737 80 1854
rect -80 1691 -23 1737
rect 23 1691 80 1737
rect -80 1574 80 1691
rect -80 1528 -23 1574
rect 23 1528 80 1574
rect -80 1411 80 1528
rect -80 1365 -23 1411
rect 23 1365 80 1411
rect -80 1247 80 1365
rect -80 1201 -23 1247
rect 23 1201 80 1247
rect -80 1084 80 1201
rect -80 1038 -23 1084
rect 23 1038 80 1084
rect -80 921 80 1038
rect -80 875 -23 921
rect 23 875 80 921
rect -80 758 80 875
rect -80 712 -23 758
rect 23 712 80 758
rect -80 595 80 712
rect -80 549 -23 595
rect 23 549 80 595
rect -80 431 80 549
rect -80 385 -23 431
rect 23 385 80 431
rect -80 268 80 385
rect -80 222 -23 268
rect 23 222 80 268
rect -80 105 80 222
rect -80 59 -23 105
rect 23 59 80 105
rect -80 -59 80 59
rect -80 -105 -23 -59
rect 23 -105 80 -59
rect -80 -222 80 -105
rect -80 -268 -23 -222
rect 23 -268 80 -222
rect -80 -385 80 -268
rect -80 -431 -23 -385
rect 23 -431 80 -385
rect -80 -549 80 -431
rect -80 -595 -23 -549
rect 23 -595 80 -549
rect -80 -712 80 -595
rect -80 -758 -23 -712
rect 23 -758 80 -712
rect -80 -875 80 -758
rect -80 -921 -23 -875
rect 23 -921 80 -875
rect -80 -1038 80 -921
rect -80 -1084 -23 -1038
rect 23 -1084 80 -1038
rect -80 -1201 80 -1084
rect -80 -1247 -23 -1201
rect 23 -1247 80 -1201
rect -80 -1365 80 -1247
rect -80 -1411 -23 -1365
rect 23 -1411 80 -1365
rect -80 -1528 80 -1411
rect -80 -1574 -23 -1528
rect 23 -1574 80 -1528
rect -80 -1691 80 -1574
rect -80 -1737 -23 -1691
rect 23 -1737 80 -1691
rect -80 -1854 80 -1737
rect -80 -1900 -23 -1854
rect 23 -1900 80 -1854
rect -80 -2018 80 -1900
rect -80 -2064 -23 -2018
rect 23 -2064 80 -2018
rect -80 -2181 80 -2064
rect -80 -2227 -23 -2181
rect 23 -2227 80 -2181
rect -80 -2344 80 -2227
rect -80 -2390 -23 -2344
rect 23 -2390 80 -2344
rect -80 -2507 80 -2390
rect -80 -2553 -23 -2507
rect 23 -2553 80 -2507
rect -80 -2613 80 -2553
<< psubdiffcont >>
rect -23 2507 23 2553
rect -23 2344 23 2390
rect -23 2181 23 2227
rect -23 2018 23 2064
rect -23 1854 23 1900
rect -23 1691 23 1737
rect -23 1528 23 1574
rect -23 1365 23 1411
rect -23 1201 23 1247
rect -23 1038 23 1084
rect -23 875 23 921
rect -23 712 23 758
rect -23 549 23 595
rect -23 385 23 431
rect -23 222 23 268
rect -23 59 23 105
rect -23 -105 23 -59
rect -23 -268 23 -222
rect -23 -431 23 -385
rect -23 -595 23 -549
rect -23 -758 23 -712
rect -23 -921 23 -875
rect -23 -1084 23 -1038
rect -23 -1247 23 -1201
rect -23 -1411 23 -1365
rect -23 -1574 23 -1528
rect -23 -1737 23 -1691
rect -23 -1900 23 -1854
rect -23 -2064 23 -2018
rect -23 -2227 23 -2181
rect -23 -2390 23 -2344
rect -23 -2553 23 -2507
<< metal1 >>
rect -71 2553 71 2603
rect -71 2507 -23 2553
rect 23 2507 71 2553
rect -71 2390 71 2507
rect -71 2344 -23 2390
rect 23 2344 71 2390
rect -71 2227 71 2344
rect -71 2181 -23 2227
rect 23 2181 71 2227
rect -71 2064 71 2181
rect -71 2018 -23 2064
rect 23 2018 71 2064
rect -71 1900 71 2018
rect -71 1854 -23 1900
rect 23 1854 71 1900
rect -71 1737 71 1854
rect -71 1691 -23 1737
rect 23 1691 71 1737
rect -71 1574 71 1691
rect -71 1528 -23 1574
rect 23 1528 71 1574
rect -71 1411 71 1528
rect -71 1365 -23 1411
rect 23 1365 71 1411
rect -71 1247 71 1365
rect -71 1201 -23 1247
rect 23 1201 71 1247
rect -71 1084 71 1201
rect -71 1038 -23 1084
rect 23 1038 71 1084
rect -71 921 71 1038
rect -71 875 -23 921
rect 23 875 71 921
rect -71 758 71 875
rect -71 712 -23 758
rect 23 712 71 758
rect -71 595 71 712
rect -71 549 -23 595
rect 23 549 71 595
rect -71 431 71 549
rect -71 385 -23 431
rect 23 385 71 431
rect -71 268 71 385
rect -71 222 -23 268
rect 23 222 71 268
rect -71 105 71 222
rect -71 59 -23 105
rect 23 59 71 105
rect -71 -59 71 59
rect -71 -105 -23 -59
rect 23 -105 71 -59
rect -71 -222 71 -105
rect -71 -268 -23 -222
rect 23 -268 71 -222
rect -71 -385 71 -268
rect -71 -431 -23 -385
rect 23 -431 71 -385
rect -71 -549 71 -431
rect -71 -595 -23 -549
rect 23 -595 71 -549
rect -71 -712 71 -595
rect -71 -758 -23 -712
rect 23 -758 71 -712
rect -71 -875 71 -758
rect -71 -921 -23 -875
rect 23 -921 71 -875
rect -71 -1038 71 -921
rect -71 -1084 -23 -1038
rect 23 -1084 71 -1038
rect -71 -1201 71 -1084
rect -71 -1247 -23 -1201
rect 23 -1247 71 -1201
rect -71 -1365 71 -1247
rect -71 -1411 -23 -1365
rect 23 -1411 71 -1365
rect -71 -1528 71 -1411
rect -71 -1574 -23 -1528
rect 23 -1574 71 -1528
rect -71 -1691 71 -1574
rect -71 -1737 -23 -1691
rect 23 -1737 71 -1691
rect -71 -1854 71 -1737
rect -71 -1900 -23 -1854
rect 23 -1900 71 -1854
rect -71 -2018 71 -1900
rect -71 -2064 -23 -2018
rect 23 -2064 71 -2018
rect -71 -2181 71 -2064
rect -71 -2227 -23 -2181
rect 23 -2227 71 -2181
rect -71 -2344 71 -2227
rect -71 -2390 -23 -2344
rect 23 -2390 71 -2344
rect -71 -2507 71 -2390
rect -71 -2553 -23 -2507
rect 23 -2553 71 -2507
rect -71 -2604 71 -2553
<< properties >>
string GDS_END 365990
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 363746
<< end >>
