magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 620 1620
<< nmos >>
rect 220 190 280 360
rect 330 190 390 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
<< ndiff >>
rect 120 298 220 360
rect 120 252 142 298
rect 188 252 220 298
rect 120 190 220 252
rect 280 190 330 360
rect 390 298 490 360
rect 390 252 422 298
rect 468 252 490 298
rect 390 190 490 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 520 1430
rect 420 1143 452 1377
rect 498 1143 520 1377
rect 420 1090 520 1143
<< ndiffc >>
rect 142 252 188 298
rect 422 252 468 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 190 780 250 1090
rect 110 753 250 780
rect 110 707 147 753
rect 193 707 250 753
rect 110 680 250 707
rect 190 450 250 680
rect 360 650 420 1090
rect 360 623 480 650
rect 360 577 407 623
rect 453 577 480 623
rect 360 550 480 577
rect 360 450 420 550
rect 190 410 280 450
rect 220 360 280 410
rect 330 410 420 450
rect 330 360 390 410
rect 220 140 280 190
rect 330 140 390 190
<< polycontact >>
rect 147 707 193 753
rect 407 577 453 623
<< metal1 >>
rect 0 1568 620 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 620 1568
rect 166 1522 352 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 620 1566
rect 0 1470 620 1514
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1060 160 1143
rect 280 1377 330 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 890 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1060 500 1143
rect 260 886 360 890
rect 260 834 284 886
rect 336 834 360 886
rect 260 800 360 834
rect 120 756 220 760
rect 120 704 144 756
rect 196 704 220 756
rect 120 670 220 704
rect 280 430 330 800
rect 380 626 480 630
rect 380 574 404 626
rect 456 574 480 626
rect 380 540 480 574
rect 140 350 330 430
rect 140 298 190 350
rect 140 252 142 298
rect 188 252 190 298
rect 140 160 190 252
rect 420 298 470 360
rect 420 252 422 298
rect 468 252 470 298
rect 420 120 470 252
rect 0 106 620 120
rect 0 98 114 106
rect 166 98 354 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 620 106
rect 158 52 352 54
rect 398 52 620 54
rect 0 -30 620 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 284 834 336 886
rect 144 753 196 756
rect 144 707 147 753
rect 147 707 193 753
rect 193 707 196 753
rect 144 704 196 707
rect 404 623 456 626
rect 404 577 407 623
rect 407 577 453 623
rect 453 577 456 623
rect 404 574 456 577
rect 114 98 166 106
rect 354 98 406 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 260 886 360 900
rect 260 834 284 886
rect 336 834 360 886
rect 260 790 360 834
rect 120 756 220 770
rect 120 704 144 756
rect 196 704 220 756
rect 120 660 220 704
rect 380 626 480 640
rect 380 574 404 626
rect 456 574 480 626
rect 380 530 480 574
rect 100 110 180 120
rect 340 110 420 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 100 10 180 20
rect 340 10 420 20
<< labels >>
rlabel metal2 s 100 1470 180 1550 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 100 10 180 90 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 120 660 220 740 4 A
port 1 nsew signal input
rlabel metal2 s 380 530 480 610 4 B
port 2 nsew signal input
rlabel metal2 s 260 790 360 870 4 Y
port 3 nsew signal output
rlabel metal1 s 120 670 220 730 1 A
port 1 nsew signal input
rlabel metal1 s 380 540 480 600 1 B
port 2 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1470 620 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 420 -30 470 330 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 -30 620 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 140 160 190 400 1 Y
port 3 nsew signal output
rlabel metal1 s 140 350 330 400 1 Y
port 3 nsew signal output
rlabel metal1 s 280 350 330 1400 1 Y
port 3 nsew signal output
rlabel metal1 s 260 800 360 860 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 620 1590
string GDS_END 406470
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 401152
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
