magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -296 -137 853 1235
<< polysilicon >>
rect -31 1099 89 1169
rect 193 1099 313 1169
rect -31 -71 89 -1
rect 193 -71 313 -1
use pmos_5p043105899832105_64x8m81  pmos_5p043105899832105_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 1220
<< properties >>
string GDS_END 524386
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 523944
<< end >>
