magic
tech gf180mcuB
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -236 230 236 236
rect -236 204 -230 230
rect -204 204 -168 230
rect -142 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 142 230
rect 168 204 204 230
rect 230 204 236 230
rect -236 168 236 204
rect -236 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 236 168
rect -236 106 236 142
rect -236 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 236 106
rect -236 44 236 80
rect -236 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 236 44
rect -236 -18 236 18
rect -236 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 236 -18
rect -236 -80 236 -44
rect -236 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 236 -80
rect -236 -142 236 -106
rect -236 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 236 -142
rect -236 -204 236 -168
rect -236 -230 -230 -204
rect -204 -230 -168 -204
rect -142 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 142 -204
rect 168 -230 204 -204
rect 230 -230 236 -204
rect -236 -236 236 -230
<< via1 >>
rect -230 204 -204 230
rect -168 204 -142 230
rect -106 204 -80 230
rect -44 204 -18 230
rect 18 204 44 230
rect 80 204 106 230
rect 142 204 168 230
rect 204 204 230 230
rect -230 142 -204 168
rect -168 142 -142 168
rect -106 142 -80 168
rect -44 142 -18 168
rect 18 142 44 168
rect 80 142 106 168
rect 142 142 168 168
rect 204 142 230 168
rect -230 80 -204 106
rect -168 80 -142 106
rect -106 80 -80 106
rect -44 80 -18 106
rect 18 80 44 106
rect 80 80 106 106
rect 142 80 168 106
rect 204 80 230 106
rect -230 18 -204 44
rect -168 18 -142 44
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect 142 18 168 44
rect 204 18 230 44
rect -230 -44 -204 -18
rect -168 -44 -142 -18
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect 142 -44 168 -18
rect 204 -44 230 -18
rect -230 -106 -204 -80
rect -168 -106 -142 -80
rect -106 -106 -80 -80
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect 80 -106 106 -80
rect 142 -106 168 -80
rect 204 -106 230 -80
rect -230 -168 -204 -142
rect -168 -168 -142 -142
rect -106 -168 -80 -142
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect 80 -168 106 -142
rect 142 -168 168 -142
rect 204 -168 230 -142
rect -230 -230 -204 -204
rect -168 -230 -142 -204
rect -106 -230 -80 -204
rect -44 -230 -18 -204
rect 18 -230 44 -204
rect 80 -230 106 -204
rect 142 -230 168 -204
rect 204 -230 230 -204
<< metal2 >>
rect -236 230 236 236
rect -236 204 -230 230
rect -204 204 -168 230
rect -142 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 142 230
rect 168 204 204 230
rect 230 204 236 230
rect -236 168 236 204
rect -236 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 236 168
rect -236 106 236 142
rect -236 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 236 106
rect -236 44 236 80
rect -236 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 236 44
rect -236 -18 236 18
rect -236 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 236 -18
rect -236 -80 236 -44
rect -236 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 236 -80
rect -236 -142 236 -106
rect -236 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 236 -142
rect -236 -204 236 -168
rect -236 -230 -230 -204
rect -204 -230 -168 -204
rect -142 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 142 -204
rect 168 -230 204 -204
rect 230 -230 236 -204
rect -236 -236 236 -230
<< properties >>
string GDS_END 2111526
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2107298
<< end >>
