magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect 0 111 410 123
rect 11 70 16 111
rect 16 55 22 65
rect 77 85 82 111
rect 114 95 119 111
rect 186 82 191 111
rect 258 95 263 111
rect 310 85 315 111
rect 68 60 78 66
rect 136 63 274 66
rect 121 57 131 63
rect 136 60 276 63
rect 164 49 170 60
rect 207 49 213 60
rect 266 57 276 60
rect 11 12 16 36
rect 162 43 172 49
rect 205 44 215 49
rect 318 57 328 63
rect 359 76 364 104
rect 376 81 381 111
rect 393 91 398 104
rect 392 81 398 91
rect 359 70 388 76
rect 380 69 386 70
rect 46 12 51 28
rect 91 12 96 29
rect 114 12 119 30
rect 186 12 191 28
rect 258 12 263 34
rect 381 42 386 69
rect 296 12 301 36
rect 359 37 386 42
rect 341 12 346 28
rect 359 19 364 37
rect 376 12 381 32
rect 393 19 398 81
rect 0 0 410 12
<< obsm1 >>
rect 28 51 33 104
rect 28 50 34 51
rect 28 44 36 50
rect 28 38 34 44
rect 43 38 48 104
rect 60 80 65 104
rect 94 80 99 104
rect 152 90 163 104
rect 60 75 99 80
rect 108 84 163 90
rect 108 66 114 84
rect 214 74 225 104
rect 247 84 257 90
rect 249 82 255 84
rect 275 77 280 104
rect 293 80 298 104
rect 327 80 332 104
rect 214 71 220 74
rect 275 72 286 77
rect 293 75 332 80
rect 344 82 349 104
rect 344 77 350 82
rect 88 60 114 66
rect 108 50 114 60
rect 53 44 63 50
rect 108 44 131 50
rect 77 38 103 44
rect 28 19 33 38
rect 43 33 82 38
rect 63 32 82 33
rect 125 33 131 44
rect 140 43 150 49
rect 180 46 186 47
rect 178 40 188 46
rect 228 44 234 54
rect 247 49 257 55
rect 281 50 286 72
rect 291 57 313 63
rect 345 57 350 77
rect 275 44 286 50
rect 228 39 280 44
rect 292 41 302 47
rect 214 33 220 39
rect 63 19 68 32
rect 125 28 163 33
rect 152 19 163 28
rect 214 19 225 33
rect 275 19 280 39
rect 307 38 313 57
rect 345 51 372 57
rect 330 43 340 49
rect 345 38 350 51
rect 307 33 350 38
rect 324 19 329 33
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 274 118 282 119
rect 298 118 306 119
rect 322 118 330 119
rect 346 118 354 119
rect 370 118 378 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 177 112 187 118
rect 201 112 211 118
rect 225 112 235 118
rect 249 112 259 118
rect 273 112 283 118
rect 297 112 307 118
rect 321 112 331 118
rect 345 112 355 118
rect 369 112 379 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 274 111 282 112
rect 298 111 306 112
rect 322 111 330 112
rect 346 111 354 112
rect 370 111 378 112
rect 70 99 326 105
rect 70 67 76 99
rect 15 63 23 64
rect 14 57 24 63
rect 68 59 78 67
rect 121 63 131 64
rect 120 57 132 63
rect 15 56 23 57
rect 121 56 131 57
rect 320 64 326 99
rect 391 89 399 90
rect 390 83 400 89
rect 391 82 399 83
rect 379 76 387 77
rect 378 70 388 76
rect 379 69 387 70
rect 267 63 275 64
rect 266 57 276 63
rect 267 56 275 57
rect 318 56 328 64
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 274 11 282 12
rect 298 11 306 12
rect 322 11 330 12
rect 346 11 354 12
rect 370 11 378 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 273 5 283 11
rect 297 5 307 11
rect 321 5 331 11
rect 345 5 355 11
rect 369 5 379 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
rect 274 4 282 5
rect 298 4 306 5
rect 322 4 330 5
rect 346 4 354 5
rect 370 4 378 5
<< obsm2 >>
rect 142 87 234 93
rect 248 90 256 91
rect 88 59 98 67
rect 27 50 35 51
rect 53 50 63 51
rect 142 50 148 87
rect 214 80 220 81
rect 213 72 221 80
rect 26 44 63 50
rect 141 49 150 50
rect 27 43 35 44
rect 53 43 63 44
rect 93 44 103 45
rect 55 24 61 43
rect 93 38 132 44
rect 140 43 150 49
rect 180 47 186 48
rect 141 42 150 43
rect 179 46 187 47
rect 93 37 103 38
rect 126 36 132 38
rect 179 40 188 46
rect 179 39 187 40
rect 179 36 186 39
rect 214 38 220 72
rect 228 52 234 87
rect 247 84 290 90
rect 248 83 256 84
rect 249 56 255 83
rect 284 64 290 84
rect 284 57 301 64
rect 291 56 301 57
rect 363 57 371 58
rect 248 55 256 56
rect 227 44 235 52
rect 247 49 257 55
rect 360 51 372 57
rect 332 50 338 51
rect 363 50 371 51
rect 248 48 256 49
rect 228 43 234 44
rect 292 40 302 48
rect 331 41 339 50
rect 213 37 221 38
rect 292 37 300 40
rect 126 30 186 36
rect 212 31 300 37
rect 213 30 221 31
rect 331 24 337 41
rect 55 18 337 24
<< labels >>
rlabel metal2 s 267 56 275 64 6 CLK
port 4 nsew clock input
rlabel metal2 s 266 57 276 63 6 CLK
port 4 nsew clock input
rlabel metal1 s 164 43 170 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 162 43 172 49 6 CLK
port 4 nsew clock input
rlabel metal1 s 207 44 213 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 205 44 215 49 6 CLK
port 4 nsew clock input
rlabel metal1 s 136 60 274 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 266 57 276 63 6 CLK
port 4 nsew clock input
rlabel metal2 s 121 56 131 64 6 D
port 1 nsew signal input
rlabel metal2 s 120 57 132 63 6 D
port 1 nsew signal input
rlabel metal1 s 121 57 131 63 6 D
port 1 nsew signal input
rlabel metal2 s 391 82 399 90 6 Q
port 2 nsew signal output
rlabel metal2 s 390 83 400 89 6 Q
port 2 nsew signal output
rlabel metal1 s 392 81 398 91 6 Q
port 2 nsew signal output
rlabel metal1 s 393 19 398 104 6 Q
port 2 nsew signal output
rlabel metal2 s 379 69 387 77 6 QN
port 3 nsew signal output
rlabel metal2 s 378 70 388 76 6 QN
port 3 nsew signal output
rlabel metal1 s 359 19 364 42 6 QN
port 3 nsew signal output
rlabel metal1 s 359 70 364 104 6 QN
port 3 nsew signal output
rlabel metal1 s 359 37 386 42 6 QN
port 3 nsew signal output
rlabel metal1 s 381 37 386 76 6 QN
port 3 nsew signal output
rlabel metal1 s 380 69 386 76 6 QN
port 3 nsew signal output
rlabel metal1 s 359 70 388 76 6 QN
port 3 nsew signal output
rlabel metal2 s 15 56 23 64 6 RN
port 5 nsew signal input
rlabel metal2 s 14 57 24 63 6 RN
port 5 nsew signal input
rlabel metal1 s 16 55 22 65 6 RN
port 5 nsew signal input
rlabel metal2 s 70 59 76 105 6 SN
port 6 nsew signal output
rlabel metal2 s 68 59 78 67 6 SN
port 6 nsew signal output
rlabel metal2 s 320 56 326 105 6 SN
port 6 nsew signal output
rlabel metal2 s 70 99 326 105 6 SN
port 6 nsew signal output
rlabel metal2 s 318 56 328 64 6 SN
port 6 nsew signal output
rlabel metal1 s 68 60 78 66 6 SN
port 6 nsew signal output
rlabel metal1 s 318 57 328 63 6 SN
port 6 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 178 111 186 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 177 112 187 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 202 111 210 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 201 112 211 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 226 111 234 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 225 112 235 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 250 111 258 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 249 112 259 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 274 111 282 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 273 112 283 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 298 111 306 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 297 112 307 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 322 111 330 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 321 112 331 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 346 111 354 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 345 112 355 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 370 111 378 119 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 369 112 379 118 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 77 85 82 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 114 95 119 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 186 82 191 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 258 95 263 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 310 85 315 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 376 81 381 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 0 111 410 123 6 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 274 4 282 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 273 5 283 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 298 4 306 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 297 5 307 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 322 4 330 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 321 5 331 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 346 4 354 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 345 5 355 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 370 4 378 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 369 5 379 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 46 0 51 28 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 91 0 96 29 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 114 0 119 30 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 186 0 191 28 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 258 0 263 34 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 296 0 301 36 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 341 0 346 28 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 376 0 381 32 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 410 12 6 VSS
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 410 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 316728
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 277374
<< end >>
