magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 5798 870
rect -86 352 1890 377
rect 5479 352 5798 377
<< pwell >>
rect -86 -86 5798 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 2060 93 2180 257
rect 2284 93 2404 257
rect 2508 93 2628 257
rect 2732 93 2852 257
rect 2956 93 3076 257
rect 3180 93 3300 257
rect 3404 93 3524 257
rect 3628 93 3748 257
rect 3852 93 3972 257
rect 4076 93 4196 257
rect 4300 93 4420 257
rect 4524 93 4644 257
rect 4748 93 4868 257
rect 4972 93 5092 257
rect 5196 93 5316 257
rect 5464 68 5584 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 572 497 672 716
rect 816 497 916 716
rect 1020 497 1120 716
rect 1264 497 1364 716
rect 1468 497 1568 716
rect 1712 497 1812 716
rect 2080 497 2180 716
rect 2304 497 2404 716
rect 2508 497 2608 716
rect 2752 497 2852 716
rect 2956 497 3056 716
rect 3200 497 3300 716
rect 3404 497 3504 716
rect 3628 497 3728 716
rect 3872 497 3972 716
rect 4096 497 4196 716
rect 4300 497 4400 716
rect 4544 497 4644 716
rect 4748 497 4848 716
rect 4992 497 5092 716
rect 5196 497 5296 716
rect 5464 497 5564 716
<< mvndiff >>
rect 36 127 124 232
rect 36 81 49 127
rect 95 81 124 127
rect 36 68 124 81
rect 244 219 348 232
rect 244 173 273 219
rect 319 173 348 219
rect 244 68 348 173
rect 468 127 572 232
rect 468 81 497 127
rect 543 81 572 127
rect 468 68 572 81
rect 692 219 796 232
rect 692 173 721 219
rect 767 173 796 219
rect 692 68 796 173
rect 916 127 1020 232
rect 916 81 945 127
rect 991 81 1020 127
rect 916 68 1020 81
rect 1140 219 1244 232
rect 1140 173 1169 219
rect 1215 173 1244 219
rect 1140 68 1244 173
rect 1364 127 1468 232
rect 1364 81 1393 127
rect 1439 81 1468 127
rect 1364 68 1468 81
rect 1588 219 1692 232
rect 1588 173 1617 219
rect 1663 173 1692 219
rect 1588 68 1692 173
rect 1812 127 1900 232
rect 1812 81 1841 127
rect 1887 81 1900 127
rect 1972 152 2060 257
rect 1972 106 1985 152
rect 2031 106 2060 152
rect 1972 93 2060 106
rect 2180 244 2284 257
rect 2180 198 2209 244
rect 2255 198 2284 244
rect 2180 93 2284 198
rect 2404 152 2508 257
rect 2404 106 2433 152
rect 2479 106 2508 152
rect 2404 93 2508 106
rect 2628 244 2732 257
rect 2628 198 2657 244
rect 2703 198 2732 244
rect 2628 93 2732 198
rect 2852 152 2956 257
rect 2852 106 2881 152
rect 2927 106 2956 152
rect 2852 93 2956 106
rect 3076 244 3180 257
rect 3076 198 3105 244
rect 3151 198 3180 244
rect 3076 93 3180 198
rect 3300 152 3404 257
rect 3300 106 3329 152
rect 3375 106 3404 152
rect 3300 93 3404 106
rect 3524 244 3628 257
rect 3524 198 3553 244
rect 3599 198 3628 244
rect 3524 93 3628 198
rect 3748 152 3852 257
rect 3748 106 3777 152
rect 3823 106 3852 152
rect 3748 93 3852 106
rect 3972 244 4076 257
rect 3972 198 4001 244
rect 4047 198 4076 244
rect 3972 93 4076 198
rect 4196 152 4300 257
rect 4196 106 4225 152
rect 4271 106 4300 152
rect 4196 93 4300 106
rect 4420 244 4524 257
rect 4420 198 4449 244
rect 4495 198 4524 244
rect 4420 93 4524 198
rect 4644 152 4748 257
rect 4644 106 4673 152
rect 4719 106 4748 152
rect 4644 93 4748 106
rect 4868 244 4972 257
rect 4868 198 4897 244
rect 4943 198 4972 244
rect 4868 93 4972 198
rect 5092 152 5196 257
rect 5092 106 5121 152
rect 5167 106 5196 152
rect 5092 93 5196 106
rect 5316 244 5404 257
rect 5316 198 5345 244
rect 5391 232 5404 244
rect 5391 198 5464 232
rect 5316 93 5464 198
rect 1812 68 1900 81
rect 5384 68 5464 93
rect 5584 152 5672 232
rect 5584 106 5613 152
rect 5659 106 5672 152
rect 5584 68 5672 106
<< mvpdiff >>
rect 46 665 144 716
rect 46 525 59 665
rect 105 525 144 665
rect 46 497 144 525
rect 244 497 368 716
rect 468 702 572 716
rect 468 656 497 702
rect 543 656 572 702
rect 468 497 572 656
rect 672 497 816 716
rect 916 665 1020 716
rect 916 525 945 665
rect 991 525 1020 665
rect 916 497 1020 525
rect 1120 497 1264 716
rect 1364 703 1468 716
rect 1364 657 1393 703
rect 1439 657 1468 703
rect 1364 497 1468 657
rect 1568 497 1712 716
rect 1812 610 2080 716
rect 1812 564 1841 610
rect 1887 564 2005 610
rect 2051 564 2080 610
rect 1812 497 2080 564
rect 2180 497 2304 716
rect 2404 703 2508 716
rect 2404 657 2433 703
rect 2479 657 2508 703
rect 2404 497 2508 657
rect 2608 497 2752 716
rect 2852 639 2956 716
rect 2852 593 2881 639
rect 2927 593 2956 639
rect 2852 497 2956 593
rect 3056 497 3200 716
rect 3300 703 3404 716
rect 3300 657 3329 703
rect 3375 657 3404 703
rect 3300 497 3404 657
rect 3504 497 3628 716
rect 3728 665 3872 716
rect 3728 525 3777 665
rect 3823 525 3872 665
rect 3728 497 3872 525
rect 3972 497 4096 716
rect 4196 703 4300 716
rect 4196 657 4225 703
rect 4271 657 4300 703
rect 4196 497 4300 657
rect 4400 497 4544 716
rect 4644 639 4748 716
rect 4644 593 4673 639
rect 4719 593 4748 639
rect 4644 497 4748 593
rect 4848 497 4992 716
rect 5092 703 5196 716
rect 5092 657 5121 703
rect 5167 657 5196 703
rect 5092 497 5196 657
rect 5296 497 5464 716
rect 5564 665 5652 716
rect 5564 525 5593 665
rect 5639 525 5652 665
rect 5564 497 5652 525
<< mvndiffc >>
rect 49 81 95 127
rect 273 173 319 219
rect 497 81 543 127
rect 721 173 767 219
rect 945 81 991 127
rect 1169 173 1215 219
rect 1393 81 1439 127
rect 1617 173 1663 219
rect 1841 81 1887 127
rect 1985 106 2031 152
rect 2209 198 2255 244
rect 2433 106 2479 152
rect 2657 198 2703 244
rect 2881 106 2927 152
rect 3105 198 3151 244
rect 3329 106 3375 152
rect 3553 198 3599 244
rect 3777 106 3823 152
rect 4001 198 4047 244
rect 4225 106 4271 152
rect 4449 198 4495 244
rect 4673 106 4719 152
rect 4897 198 4943 244
rect 5121 106 5167 152
rect 5345 198 5391 244
rect 5613 106 5659 152
<< mvpdiffc >>
rect 59 525 105 665
rect 497 656 543 702
rect 945 525 991 665
rect 1393 657 1439 703
rect 1841 564 1887 610
rect 2005 564 2051 610
rect 2433 657 2479 703
rect 2881 593 2927 639
rect 3329 657 3375 703
rect 3777 525 3823 665
rect 4225 657 4271 703
rect 4673 593 4719 639
rect 5121 657 5167 703
rect 5593 525 5639 665
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 1020 716 1120 760
rect 1264 716 1364 760
rect 1468 716 1568 760
rect 1712 716 1812 760
rect 2080 716 2180 760
rect 2304 716 2404 760
rect 2508 716 2608 760
rect 2752 716 2852 760
rect 2956 716 3056 760
rect 3200 716 3300 760
rect 3404 716 3504 760
rect 3628 716 3728 760
rect 3872 716 3972 760
rect 4096 716 4196 760
rect 4300 716 4400 760
rect 4544 716 4644 760
rect 4748 716 4848 760
rect 4992 716 5092 760
rect 5196 716 5296 760
rect 5464 716 5564 760
rect 144 415 244 497
rect 144 402 171 415
rect 124 369 171 402
rect 217 369 244 415
rect 368 415 468 497
rect 368 402 395 415
rect 124 232 244 369
rect 348 369 395 402
rect 441 394 468 415
rect 572 415 672 497
rect 572 394 599 415
rect 441 369 599 394
rect 645 402 672 415
rect 816 402 916 497
rect 645 369 692 402
rect 348 348 692 369
rect 348 232 468 348
rect 572 232 692 348
rect 796 394 916 402
rect 1020 402 1120 497
rect 1264 415 1364 497
rect 1264 402 1291 415
rect 1020 394 1140 402
rect 796 348 1140 394
rect 796 312 916 348
rect 796 266 833 312
rect 879 266 916 312
rect 796 232 916 266
rect 1020 312 1140 348
rect 1020 266 1057 312
rect 1103 266 1140 312
rect 1020 232 1140 266
rect 1244 369 1291 402
rect 1337 394 1364 415
rect 1468 415 1568 497
rect 1468 394 1495 415
rect 1337 369 1495 394
rect 1541 402 1568 415
rect 1712 415 1812 497
rect 1712 402 1739 415
rect 1541 369 1588 402
rect 1244 348 1588 369
rect 1244 232 1364 348
rect 1468 232 1588 348
rect 1692 369 1739 402
rect 1785 369 1812 415
rect 2080 415 2180 497
rect 2080 402 2107 415
rect 1692 232 1812 369
rect 2060 369 2107 402
rect 2153 369 2180 415
rect 2304 415 2404 497
rect 2304 402 2331 415
rect 2060 257 2180 369
rect 2284 369 2331 402
rect 2377 394 2404 415
rect 2508 415 2608 497
rect 2508 394 2535 415
rect 2377 369 2535 394
rect 2581 402 2608 415
rect 2752 436 2852 497
rect 2752 402 2779 436
rect 2581 369 2628 402
rect 2284 348 2628 369
rect 2284 257 2404 348
rect 2508 257 2628 348
rect 2732 390 2779 402
rect 2825 394 2852 436
rect 2956 436 3056 497
rect 2956 394 2983 436
rect 2825 390 2983 394
rect 3029 402 3056 436
rect 3200 415 3300 497
rect 3200 402 3227 415
rect 3029 390 3076 402
rect 2732 348 3076 390
rect 2732 257 2852 348
rect 2956 257 3076 348
rect 3180 369 3227 402
rect 3273 394 3300 415
rect 3404 415 3504 497
rect 3404 394 3431 415
rect 3273 369 3431 394
rect 3477 402 3504 415
rect 3628 436 3728 497
rect 3477 369 3524 402
rect 3180 348 3524 369
rect 3180 257 3300 348
rect 3404 257 3524 348
rect 3628 390 3655 436
rect 3701 402 3728 436
rect 3872 415 3972 497
rect 3872 402 3899 415
rect 3701 390 3748 402
rect 3628 257 3748 390
rect 3852 369 3899 402
rect 3945 369 3972 415
rect 4096 415 4196 497
rect 4096 402 4123 415
rect 3852 257 3972 369
rect 4076 369 4123 402
rect 4169 394 4196 415
rect 4300 415 4400 497
rect 4300 394 4327 415
rect 4169 369 4327 394
rect 4373 402 4400 415
rect 4544 436 4644 497
rect 4544 402 4571 436
rect 4373 369 4420 402
rect 4076 348 4420 369
rect 4076 257 4196 348
rect 4300 257 4420 348
rect 4524 390 4571 402
rect 4617 394 4644 436
rect 4748 436 4848 497
rect 4748 394 4775 436
rect 4617 390 4775 394
rect 4821 402 4848 436
rect 4992 415 5092 497
rect 4992 402 5019 415
rect 4821 390 4868 402
rect 4524 348 4868 390
rect 4524 257 4644 348
rect 4748 257 4868 348
rect 4972 369 5019 402
rect 5065 394 5092 415
rect 5196 415 5296 497
rect 5196 394 5223 415
rect 5065 369 5223 394
rect 5269 402 5296 415
rect 5464 415 5564 497
rect 5269 369 5316 402
rect 4972 348 5316 369
rect 4972 257 5092 348
rect 5196 257 5316 348
rect 5464 369 5491 415
rect 5537 402 5564 415
rect 5537 369 5584 402
rect 5464 232 5584 369
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 2060 24 2180 93
rect 2284 24 2404 93
rect 2508 24 2628 93
rect 2732 24 2852 93
rect 2956 24 3076 93
rect 3180 24 3300 93
rect 3404 24 3524 93
rect 3628 24 3748 93
rect 3852 24 3972 93
rect 4076 24 4196 93
rect 4300 24 4420 93
rect 4524 24 4644 93
rect 4748 24 4868 93
rect 4972 24 5092 93
rect 5196 24 5316 93
rect 5464 24 5584 68
<< polycontact >>
rect 171 369 217 415
rect 395 369 441 415
rect 599 369 645 415
rect 833 266 879 312
rect 1057 266 1103 312
rect 1291 369 1337 415
rect 1495 369 1541 415
rect 1739 369 1785 415
rect 2107 369 2153 415
rect 2331 369 2377 415
rect 2535 369 2581 415
rect 2779 390 2825 436
rect 2983 390 3029 436
rect 3227 369 3273 415
rect 3431 369 3477 415
rect 3655 390 3701 436
rect 3899 369 3945 415
rect 4123 369 4169 415
rect 4327 369 4373 415
rect 4571 390 4617 436
rect 4775 390 4821 436
rect 5019 369 5065 415
rect 5223 369 5269 415
rect 5491 369 5537 415
<< metal1 >>
rect 0 724 5712 844
rect 486 702 554 724
rect 59 665 105 676
rect 486 656 497 702
rect 543 656 554 702
rect 1382 703 1450 724
rect 945 665 991 676
rect 604 610 945 648
rect 105 564 945 610
rect 59 506 105 525
rect 1382 657 1393 703
rect 1439 657 1450 703
rect 2422 703 2490 724
rect 2422 657 2433 703
rect 2479 657 2490 703
rect 3318 703 3386 724
rect 3318 657 3329 703
rect 3375 657 3386 703
rect 4214 703 4282 724
rect 3762 665 3824 676
rect 991 610 1332 648
rect 2540 639 3268 648
rect 2540 610 2881 639
rect 991 564 1841 610
rect 1887 564 2005 610
rect 2051 593 2881 610
rect 2927 610 3268 639
rect 3762 610 3777 665
rect 2927 593 3777 610
rect 2051 584 3777 593
rect 2051 564 2590 584
rect 3218 564 3777 584
rect 945 506 991 525
rect 2640 516 3168 536
rect 3762 525 3777 564
rect 3823 610 3824 665
rect 4214 657 4225 703
rect 4271 657 4282 703
rect 5110 703 5178 724
rect 5110 657 5121 703
rect 5167 657 5178 703
rect 5593 665 5639 676
rect 4332 639 5060 648
rect 4332 610 4673 639
rect 3823 593 4673 610
rect 4719 610 5060 639
rect 4719 593 5593 610
rect 3823 584 5593 593
rect 3823 564 4382 584
rect 5010 564 5593 584
rect 3823 525 3824 564
rect 2172 470 3712 516
rect 2172 430 2218 470
rect 56 415 314 430
rect 56 369 171 415
rect 217 369 314 415
rect 56 354 314 369
rect 384 415 1568 424
rect 384 369 395 415
rect 441 369 599 415
rect 645 369 1291 415
rect 1337 369 1495 415
rect 1541 369 1568 415
rect 384 360 1568 369
rect 1640 415 1880 430
rect 1640 369 1739 415
rect 1785 369 1880 415
rect 251 312 314 354
rect 1640 354 1880 369
rect 1926 415 2218 430
rect 2768 436 2836 470
rect 1926 369 2107 415
rect 2153 369 2218 415
rect 1926 354 2218 369
rect 2264 415 2678 424
rect 2264 369 2331 415
rect 2377 369 2535 415
rect 2581 369 2678 415
rect 2768 390 2779 436
rect 2825 390 2836 436
rect 2972 436 3040 470
rect 2972 390 2983 436
rect 3029 390 3040 436
rect 3644 436 3712 470
rect 3124 415 3574 424
rect 2264 360 2678 369
rect 1640 312 1703 354
rect 251 266 833 312
rect 879 266 1057 312
rect 1103 266 1703 312
rect 2586 340 2678 360
rect 3124 369 3227 415
rect 3273 369 3431 415
rect 3477 369 3574 415
rect 3644 390 3655 436
rect 3701 390 3712 436
rect 3124 360 3574 369
rect 3124 340 3170 360
rect 2586 294 3170 340
rect 3762 244 3824 525
rect 4432 516 4960 536
rect 3898 470 5543 516
rect 5593 506 5639 525
rect 3898 415 3946 470
rect 4560 436 4628 470
rect 3898 369 3899 415
rect 3945 369 3946 415
rect 3898 358 3946 369
rect 4042 415 4470 424
rect 4042 369 4123 415
rect 4169 369 4327 415
rect 4373 369 4470 415
rect 4560 390 4571 436
rect 4617 390 4628 436
rect 4764 436 4832 470
rect 4764 390 4775 436
rect 4821 390 4832 436
rect 4938 415 5366 424
rect 4042 360 4470 369
rect 4414 340 4470 360
rect 4938 369 5019 415
rect 5065 369 5223 415
rect 5269 369 5366 415
rect 4938 360 5366 369
rect 5484 415 5543 470
rect 5484 369 5491 415
rect 5537 369 5543 415
rect 4938 340 4994 360
rect 5484 344 5543 369
rect 4414 294 4994 340
rect 1853 219 2209 244
rect 262 173 273 219
rect 319 173 721 219
rect 767 173 1169 219
rect 1215 173 1617 219
rect 1663 198 2209 219
rect 2255 198 2657 244
rect 2703 198 3105 244
rect 3151 198 3553 244
rect 3599 198 3610 244
rect 3762 198 4001 244
rect 4047 198 4449 244
rect 4495 198 4897 244
rect 4943 198 5345 244
rect 5391 198 5402 244
rect 1663 173 1899 198
rect 38 81 49 127
rect 95 81 106 127
rect 38 60 106 81
rect 486 81 497 127
rect 543 81 554 127
rect 486 60 554 81
rect 934 81 945 127
rect 991 81 1002 127
rect 934 60 1002 81
rect 1382 81 1393 127
rect 1439 81 1450 127
rect 1382 60 1450 81
rect 1830 81 1841 127
rect 1887 81 1898 127
rect 1972 106 1985 152
rect 2031 106 2433 152
rect 2479 106 2881 152
rect 2927 106 3329 152
rect 3375 106 3777 152
rect 3823 106 4225 152
rect 4271 106 4673 152
rect 4719 106 5121 152
rect 5167 106 5613 152
rect 5659 106 5672 152
rect 1830 60 1898 81
rect 0 -60 5712 60
<< labels >>
flabel metal1 s 2640 516 3168 536 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 3124 360 3574 424 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel metal1 s 1640 354 1880 430 0 FreeSans 400 0 0 0 C1
port 5 nsew default input
flabel metal1 s 384 360 1568 424 0 FreeSans 400 0 0 0 C2
port 6 nsew default input
flabel metal1 s 0 724 5712 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 1830 60 1898 127 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 5593 648 5639 676 0 FreeSans 400 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 4432 516 4960 536 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 4938 360 5366 424 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
rlabel metal1 s 3898 470 5543 516 1 A1
port 1 nsew default input
rlabel metal1 s 5484 390 5543 470 1 A1
port 1 nsew default input
rlabel metal1 s 4764 390 4832 470 1 A1
port 1 nsew default input
rlabel metal1 s 4560 390 4628 470 1 A1
port 1 nsew default input
rlabel metal1 s 3898 390 3946 470 1 A1
port 1 nsew default input
rlabel metal1 s 5484 358 5543 390 1 A1
port 1 nsew default input
rlabel metal1 s 3898 358 3946 390 1 A1
port 1 nsew default input
rlabel metal1 s 5484 344 5543 358 1 A1
port 1 nsew default input
rlabel metal1 s 4042 360 4470 424 1 A2
port 2 nsew default input
rlabel metal1 s 4938 340 4994 360 1 A2
port 2 nsew default input
rlabel metal1 s 4414 340 4470 360 1 A2
port 2 nsew default input
rlabel metal1 s 4414 294 4994 340 1 A2
port 2 nsew default input
rlabel metal1 s 2172 470 3712 516 1 B1
port 3 nsew default input
rlabel metal1 s 3644 430 3712 470 1 B1
port 3 nsew default input
rlabel metal1 s 2972 430 3040 470 1 B1
port 3 nsew default input
rlabel metal1 s 2768 430 2836 470 1 B1
port 3 nsew default input
rlabel metal1 s 2172 430 2218 470 1 B1
port 3 nsew default input
rlabel metal1 s 3644 390 3712 430 1 B1
port 3 nsew default input
rlabel metal1 s 2972 390 3040 430 1 B1
port 3 nsew default input
rlabel metal1 s 2768 390 2836 430 1 B1
port 3 nsew default input
rlabel metal1 s 1926 390 2218 430 1 B1
port 3 nsew default input
rlabel metal1 s 1926 354 2218 390 1 B1
port 3 nsew default input
rlabel metal1 s 2264 360 2678 424 1 B2
port 4 nsew default input
rlabel metal1 s 3124 340 3170 360 1 B2
port 4 nsew default input
rlabel metal1 s 2586 340 2678 360 1 B2
port 4 nsew default input
rlabel metal1 s 2586 294 3170 340 1 B2
port 4 nsew default input
rlabel metal1 s 56 354 314 430 1 C1
port 5 nsew default input
rlabel metal1 s 1640 312 1703 354 1 C1
port 5 nsew default input
rlabel metal1 s 251 312 314 354 1 C1
port 5 nsew default input
rlabel metal1 s 251 266 1703 312 1 C1
port 5 nsew default input
rlabel metal1 s 3762 648 3824 676 1 ZN
port 7 nsew default output
rlabel metal1 s 945 648 991 676 1 ZN
port 7 nsew default output
rlabel metal1 s 59 648 105 676 1 ZN
port 7 nsew default output
rlabel metal1 s 5593 610 5639 648 1 ZN
port 7 nsew default output
rlabel metal1 s 4332 610 5060 648 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 610 3824 648 1 ZN
port 7 nsew default output
rlabel metal1 s 2540 610 3268 648 1 ZN
port 7 nsew default output
rlabel metal1 s 604 610 1332 648 1 ZN
port 7 nsew default output
rlabel metal1 s 59 610 105 648 1 ZN
port 7 nsew default output
rlabel metal1 s 59 584 5639 610 1 ZN
port 7 nsew default output
rlabel metal1 s 5010 564 5639 584 1 ZN
port 7 nsew default output
rlabel metal1 s 3218 564 4382 584 1 ZN
port 7 nsew default output
rlabel metal1 s 59 564 2590 584 1 ZN
port 7 nsew default output
rlabel metal1 s 5593 506 5639 564 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 506 3824 564 1 ZN
port 7 nsew default output
rlabel metal1 s 945 506 991 564 1 ZN
port 7 nsew default output
rlabel metal1 s 59 506 105 564 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 244 3824 506 1 ZN
port 7 nsew default output
rlabel metal1 s 3762 198 5402 244 1 ZN
port 7 nsew default output
rlabel metal1 s 5110 657 5178 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4214 657 4282 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3318 657 3386 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2422 657 2490 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1382 657 1450 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 486 657 554 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 486 656 554 657 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1382 60 1450 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5712 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5712 784
string GDS_END 140516
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 130730
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
