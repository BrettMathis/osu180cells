magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 792 979
<< polysilicon >>
rect -31 908 89 980
rect 193 908 313 980
rect 417 908 537 980
rect -31 -73 89 -1
rect 193 -73 313 -1
rect 417 -73 537 -1
use pmos_5p04310590548725_128x8m81  pmos_5p04310590548725_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 776 1028
<< properties >>
string GDS_END 258512
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 257942
<< end >>
