magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -19 377 19 382
rect -19 349 -14 377
rect 14 349 19 377
rect -19 311 19 349
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -349 19 -311
rect -19 -377 -14 -349
rect 14 -377 19 -349
rect -19 -382 19 -377
<< via2 >>
rect -14 349 14 377
rect -14 283 14 311
rect -14 217 14 245
rect -14 151 14 179
rect -14 85 14 113
rect -14 19 14 47
rect -14 -47 14 -19
rect -14 -113 14 -85
rect -14 -179 14 -151
rect -14 -245 14 -217
rect -14 -311 14 -283
rect -14 -377 14 -349
<< metal3 >>
rect -19 377 19 382
rect -19 349 -14 377
rect 14 349 19 377
rect -19 311 19 349
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -349 19 -311
rect -19 -377 -14 -349
rect 14 -377 19 -349
rect -19 -382 19 -377
<< properties >>
string GDS_END 660708
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 659808
<< end >>
