magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -1273 112 1273 118
rect -1273 86 -1267 112
rect -1241 86 -1201 112
rect -1175 86 -1135 112
rect -1109 86 -1069 112
rect -1043 86 -1003 112
rect -977 86 -937 112
rect -911 86 -871 112
rect -845 86 -805 112
rect -779 86 -739 112
rect -713 86 -673 112
rect -647 86 -607 112
rect -581 86 -541 112
rect -515 86 -475 112
rect -449 86 -409 112
rect -383 86 -343 112
rect -317 86 -277 112
rect -251 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 251 112
rect 277 86 317 112
rect 343 86 383 112
rect 409 86 449 112
rect 475 86 515 112
rect 541 86 581 112
rect 607 86 647 112
rect 673 86 713 112
rect 739 86 779 112
rect 805 86 845 112
rect 871 86 911 112
rect 937 86 977 112
rect 1003 86 1043 112
rect 1069 86 1109 112
rect 1135 86 1175 112
rect 1201 86 1241 112
rect 1267 86 1273 112
rect -1273 46 1273 86
rect -1273 20 -1267 46
rect -1241 20 -1201 46
rect -1175 20 -1135 46
rect -1109 20 -1069 46
rect -1043 20 -1003 46
rect -977 20 -937 46
rect -911 20 -871 46
rect -845 20 -805 46
rect -779 20 -739 46
rect -713 20 -673 46
rect -647 20 -607 46
rect -581 20 -541 46
rect -515 20 -475 46
rect -449 20 -409 46
rect -383 20 -343 46
rect -317 20 -277 46
rect -251 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 251 46
rect 277 20 317 46
rect 343 20 383 46
rect 409 20 449 46
rect 475 20 515 46
rect 541 20 581 46
rect 607 20 647 46
rect 673 20 713 46
rect 739 20 779 46
rect 805 20 845 46
rect 871 20 911 46
rect 937 20 977 46
rect 1003 20 1043 46
rect 1069 20 1109 46
rect 1135 20 1175 46
rect 1201 20 1241 46
rect 1267 20 1273 46
rect -1273 -20 1273 20
rect -1273 -46 -1267 -20
rect -1241 -46 -1201 -20
rect -1175 -46 -1135 -20
rect -1109 -46 -1069 -20
rect -1043 -46 -1003 -20
rect -977 -46 -937 -20
rect -911 -46 -871 -20
rect -845 -46 -805 -20
rect -779 -46 -739 -20
rect -713 -46 -673 -20
rect -647 -46 -607 -20
rect -581 -46 -541 -20
rect -515 -46 -475 -20
rect -449 -46 -409 -20
rect -383 -46 -343 -20
rect -317 -46 -277 -20
rect -251 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 251 -20
rect 277 -46 317 -20
rect 343 -46 383 -20
rect 409 -46 449 -20
rect 475 -46 515 -20
rect 541 -46 581 -20
rect 607 -46 647 -20
rect 673 -46 713 -20
rect 739 -46 779 -20
rect 805 -46 845 -20
rect 871 -46 911 -20
rect 937 -46 977 -20
rect 1003 -46 1043 -20
rect 1069 -46 1109 -20
rect 1135 -46 1175 -20
rect 1201 -46 1241 -20
rect 1267 -46 1273 -20
rect -1273 -86 1273 -46
rect -1273 -112 -1267 -86
rect -1241 -112 -1201 -86
rect -1175 -112 -1135 -86
rect -1109 -112 -1069 -86
rect -1043 -112 -1003 -86
rect -977 -112 -937 -86
rect -911 -112 -871 -86
rect -845 -112 -805 -86
rect -779 -112 -739 -86
rect -713 -112 -673 -86
rect -647 -112 -607 -86
rect -581 -112 -541 -86
rect -515 -112 -475 -86
rect -449 -112 -409 -86
rect -383 -112 -343 -86
rect -317 -112 -277 -86
rect -251 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 251 -86
rect 277 -112 317 -86
rect 343 -112 383 -86
rect 409 -112 449 -86
rect 475 -112 515 -86
rect 541 -112 581 -86
rect 607 -112 647 -86
rect 673 -112 713 -86
rect 739 -112 779 -86
rect 805 -112 845 -86
rect 871 -112 911 -86
rect 937 -112 977 -86
rect 1003 -112 1043 -86
rect 1069 -112 1109 -86
rect 1135 -112 1175 -86
rect 1201 -112 1241 -86
rect 1267 -112 1273 -86
rect -1273 -118 1273 -112
<< via1 >>
rect -1267 86 -1241 112
rect -1201 86 -1175 112
rect -1135 86 -1109 112
rect -1069 86 -1043 112
rect -1003 86 -977 112
rect -937 86 -911 112
rect -871 86 -845 112
rect -805 86 -779 112
rect -739 86 -713 112
rect -673 86 -647 112
rect -607 86 -581 112
rect -541 86 -515 112
rect -475 86 -449 112
rect -409 86 -383 112
rect -343 86 -317 112
rect -277 86 -251 112
rect -211 86 -185 112
rect -145 86 -119 112
rect -79 86 -53 112
rect -13 86 13 112
rect 53 86 79 112
rect 119 86 145 112
rect 185 86 211 112
rect 251 86 277 112
rect 317 86 343 112
rect 383 86 409 112
rect 449 86 475 112
rect 515 86 541 112
rect 581 86 607 112
rect 647 86 673 112
rect 713 86 739 112
rect 779 86 805 112
rect 845 86 871 112
rect 911 86 937 112
rect 977 86 1003 112
rect 1043 86 1069 112
rect 1109 86 1135 112
rect 1175 86 1201 112
rect 1241 86 1267 112
rect -1267 20 -1241 46
rect -1201 20 -1175 46
rect -1135 20 -1109 46
rect -1069 20 -1043 46
rect -1003 20 -977 46
rect -937 20 -911 46
rect -871 20 -845 46
rect -805 20 -779 46
rect -739 20 -713 46
rect -673 20 -647 46
rect -607 20 -581 46
rect -541 20 -515 46
rect -475 20 -449 46
rect -409 20 -383 46
rect -343 20 -317 46
rect -277 20 -251 46
rect -211 20 -185 46
rect -145 20 -119 46
rect -79 20 -53 46
rect -13 20 13 46
rect 53 20 79 46
rect 119 20 145 46
rect 185 20 211 46
rect 251 20 277 46
rect 317 20 343 46
rect 383 20 409 46
rect 449 20 475 46
rect 515 20 541 46
rect 581 20 607 46
rect 647 20 673 46
rect 713 20 739 46
rect 779 20 805 46
rect 845 20 871 46
rect 911 20 937 46
rect 977 20 1003 46
rect 1043 20 1069 46
rect 1109 20 1135 46
rect 1175 20 1201 46
rect 1241 20 1267 46
rect -1267 -46 -1241 -20
rect -1201 -46 -1175 -20
rect -1135 -46 -1109 -20
rect -1069 -46 -1043 -20
rect -1003 -46 -977 -20
rect -937 -46 -911 -20
rect -871 -46 -845 -20
rect -805 -46 -779 -20
rect -739 -46 -713 -20
rect -673 -46 -647 -20
rect -607 -46 -581 -20
rect -541 -46 -515 -20
rect -475 -46 -449 -20
rect -409 -46 -383 -20
rect -343 -46 -317 -20
rect -277 -46 -251 -20
rect -211 -46 -185 -20
rect -145 -46 -119 -20
rect -79 -46 -53 -20
rect -13 -46 13 -20
rect 53 -46 79 -20
rect 119 -46 145 -20
rect 185 -46 211 -20
rect 251 -46 277 -20
rect 317 -46 343 -20
rect 383 -46 409 -20
rect 449 -46 475 -20
rect 515 -46 541 -20
rect 581 -46 607 -20
rect 647 -46 673 -20
rect 713 -46 739 -20
rect 779 -46 805 -20
rect 845 -46 871 -20
rect 911 -46 937 -20
rect 977 -46 1003 -20
rect 1043 -46 1069 -20
rect 1109 -46 1135 -20
rect 1175 -46 1201 -20
rect 1241 -46 1267 -20
rect -1267 -112 -1241 -86
rect -1201 -112 -1175 -86
rect -1135 -112 -1109 -86
rect -1069 -112 -1043 -86
rect -1003 -112 -977 -86
rect -937 -112 -911 -86
rect -871 -112 -845 -86
rect -805 -112 -779 -86
rect -739 -112 -713 -86
rect -673 -112 -647 -86
rect -607 -112 -581 -86
rect -541 -112 -515 -86
rect -475 -112 -449 -86
rect -409 -112 -383 -86
rect -343 -112 -317 -86
rect -277 -112 -251 -86
rect -211 -112 -185 -86
rect -145 -112 -119 -86
rect -79 -112 -53 -86
rect -13 -112 13 -86
rect 53 -112 79 -86
rect 119 -112 145 -86
rect 185 -112 211 -86
rect 251 -112 277 -86
rect 317 -112 343 -86
rect 383 -112 409 -86
rect 449 -112 475 -86
rect 515 -112 541 -86
rect 581 -112 607 -86
rect 647 -112 673 -86
rect 713 -112 739 -86
rect 779 -112 805 -86
rect 845 -112 871 -86
rect 911 -112 937 -86
rect 977 -112 1003 -86
rect 1043 -112 1069 -86
rect 1109 -112 1135 -86
rect 1175 -112 1201 -86
rect 1241 -112 1267 -86
<< metal2 >>
rect -1273 112 1273 118
rect -1273 86 -1267 112
rect -1241 86 -1201 112
rect -1175 86 -1135 112
rect -1109 86 -1069 112
rect -1043 86 -1003 112
rect -977 86 -937 112
rect -911 86 -871 112
rect -845 86 -805 112
rect -779 86 -739 112
rect -713 86 -673 112
rect -647 86 -607 112
rect -581 86 -541 112
rect -515 86 -475 112
rect -449 86 -409 112
rect -383 86 -343 112
rect -317 86 -277 112
rect -251 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 251 112
rect 277 86 317 112
rect 343 86 383 112
rect 409 86 449 112
rect 475 86 515 112
rect 541 86 581 112
rect 607 86 647 112
rect 673 86 713 112
rect 739 86 779 112
rect 805 86 845 112
rect 871 86 911 112
rect 937 86 977 112
rect 1003 86 1043 112
rect 1069 86 1109 112
rect 1135 86 1175 112
rect 1201 86 1241 112
rect 1267 86 1273 112
rect -1273 46 1273 86
rect -1273 20 -1267 46
rect -1241 20 -1201 46
rect -1175 20 -1135 46
rect -1109 20 -1069 46
rect -1043 20 -1003 46
rect -977 20 -937 46
rect -911 20 -871 46
rect -845 20 -805 46
rect -779 20 -739 46
rect -713 20 -673 46
rect -647 20 -607 46
rect -581 20 -541 46
rect -515 20 -475 46
rect -449 20 -409 46
rect -383 20 -343 46
rect -317 20 -277 46
rect -251 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 251 46
rect 277 20 317 46
rect 343 20 383 46
rect 409 20 449 46
rect 475 20 515 46
rect 541 20 581 46
rect 607 20 647 46
rect 673 20 713 46
rect 739 20 779 46
rect 805 20 845 46
rect 871 20 911 46
rect 937 20 977 46
rect 1003 20 1043 46
rect 1069 20 1109 46
rect 1135 20 1175 46
rect 1201 20 1241 46
rect 1267 20 1273 46
rect -1273 -20 1273 20
rect -1273 -46 -1267 -20
rect -1241 -46 -1201 -20
rect -1175 -46 -1135 -20
rect -1109 -46 -1069 -20
rect -1043 -46 -1003 -20
rect -977 -46 -937 -20
rect -911 -46 -871 -20
rect -845 -46 -805 -20
rect -779 -46 -739 -20
rect -713 -46 -673 -20
rect -647 -46 -607 -20
rect -581 -46 -541 -20
rect -515 -46 -475 -20
rect -449 -46 -409 -20
rect -383 -46 -343 -20
rect -317 -46 -277 -20
rect -251 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 251 -20
rect 277 -46 317 -20
rect 343 -46 383 -20
rect 409 -46 449 -20
rect 475 -46 515 -20
rect 541 -46 581 -20
rect 607 -46 647 -20
rect 673 -46 713 -20
rect 739 -46 779 -20
rect 805 -46 845 -20
rect 871 -46 911 -20
rect 937 -46 977 -20
rect 1003 -46 1043 -20
rect 1069 -46 1109 -20
rect 1135 -46 1175 -20
rect 1201 -46 1241 -20
rect 1267 -46 1273 -20
rect -1273 -86 1273 -46
rect -1273 -112 -1267 -86
rect -1241 -112 -1201 -86
rect -1175 -112 -1135 -86
rect -1109 -112 -1069 -86
rect -1043 -112 -1003 -86
rect -977 -112 -937 -86
rect -911 -112 -871 -86
rect -845 -112 -805 -86
rect -779 -112 -739 -86
rect -713 -112 -673 -86
rect -647 -112 -607 -86
rect -581 -112 -541 -86
rect -515 -112 -475 -86
rect -449 -112 -409 -86
rect -383 -112 -343 -86
rect -317 -112 -277 -86
rect -251 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 251 -86
rect 277 -112 317 -86
rect 343 -112 383 -86
rect 409 -112 449 -86
rect 475 -112 515 -86
rect 541 -112 581 -86
rect 607 -112 647 -86
rect 673 -112 713 -86
rect 739 -112 779 -86
rect 805 -112 845 -86
rect 871 -112 911 -86
rect 937 -112 977 -86
rect 1003 -112 1043 -86
rect 1069 -112 1109 -86
rect 1135 -112 1175 -86
rect 1201 -112 1241 -86
rect 1267 -112 1273 -86
rect -1273 -118 1273 -112
<< properties >>
string GDS_END 978236
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 968120
<< end >>
