magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect 0 111 96 123
rect 11 70 16 111
rect 28 65 33 104
rect 45 70 50 111
rect 62 76 67 104
rect 62 70 75 76
rect 80 70 85 111
rect 62 65 67 70
rect 28 60 67 65
rect 8 44 18 50
rect 28 46 33 60
rect 62 46 67 60
rect 28 41 67 46
rect 11 12 16 36
rect 28 19 33 41
rect 45 12 50 36
rect 62 19 67 41
rect 79 12 84 36
rect 0 0 96 12
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 66 76 74 77
rect 65 70 75 76
rect 66 69 74 70
rect 8 43 18 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 s 8 43 18 51 6 A
port 1 nsew signal input
rlabel metal1 s 8 44 18 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 45 70 50 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 80 70 85 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 96 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 0 50 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 79 0 84 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 96 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 66 69 74 77 6 Y
port 2 nsew signal output
rlabel metal2 s 65 70 75 76 6 Y
port 2 nsew signal output
rlabel metal1 s 28 19 33 104 6 Y
port 2 nsew signal output
rlabel metal1 s 28 41 67 46 6 Y
port 2 nsew signal output
rlabel metal1 s 28 60 67 65 6 Y
port 2 nsew signal output
rlabel metal1 s 62 19 67 104 6 Y
port 2 nsew signal output
rlabel metal1 s 62 70 75 76 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 96 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 186686
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 179294
<< end >>
