magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -747 23 747 42
rect -747 -23 -728 23
rect 728 -23 747 23
rect -747 -42 747 -23
<< psubdiffcont >>
rect -728 -23 728 23
<< metal1 >>
rect -739 23 739 34
rect -739 -23 -728 23
rect 728 -23 739 23
rect -739 -34 739 -23
<< properties >>
string GDS_END 432576
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 431356
<< end >>
