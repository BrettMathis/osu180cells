magic
tech gf180mcuB
timestamp 1669390400
<< properties >>
string GDS_END 7678182
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7677154
<< end >>
