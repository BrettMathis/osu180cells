magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -50 200 50 205
rect -50 172 -45 200
rect -17 172 17 200
rect 45 172 50 200
rect -50 138 50 172
rect -50 110 -45 138
rect -17 110 17 138
rect 45 110 50 138
rect -50 76 50 110
rect -50 48 -45 76
rect -17 48 17 76
rect 45 48 50 76
rect -50 14 50 48
rect -50 -14 -45 14
rect -17 -14 17 14
rect 45 -14 50 14
rect -50 -48 50 -14
rect -50 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 50 -48
rect -50 -110 50 -76
rect -50 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 50 -110
rect -50 -172 50 -138
rect -50 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 50 -172
rect -50 -205 50 -200
<< via2 >>
rect -45 172 -17 200
rect 17 172 45 200
rect -45 110 -17 138
rect 17 110 45 138
rect -45 48 -17 76
rect 17 48 45 76
rect -45 -14 -17 14
rect 17 -14 45 14
rect -45 -76 -17 -48
rect 17 -76 45 -48
rect -45 -138 -17 -110
rect 17 -138 45 -110
rect -45 -200 -17 -172
rect 17 -200 45 -172
<< metal3 >>
rect -50 200 50 205
rect -50 172 -45 200
rect -17 172 17 200
rect 45 172 50 200
rect -50 138 50 172
rect -50 110 -45 138
rect -17 110 17 138
rect 45 110 50 138
rect -50 76 50 110
rect -50 48 -45 76
rect -17 48 17 76
rect 45 48 50 76
rect -50 14 50 48
rect -50 -14 -45 14
rect -17 -14 17 14
rect 45 -14 50 14
rect -50 -48 50 -14
rect -50 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 50 -48
rect -50 -110 50 -76
rect -50 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 50 -110
rect -50 -172 50 -138
rect -50 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 50 -172
rect -50 -205 50 -200
<< properties >>
string GDS_END 992328
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 991300
<< end >>
