magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -64 1878 65 1917
rect -64 1822 -28 1878
rect 28 1822 65 1878
rect -64 1660 65 1822
rect -64 1604 -28 1660
rect 28 1604 65 1660
rect -64 1443 65 1604
rect -64 1387 -28 1443
rect 28 1387 65 1443
rect -64 1225 65 1387
rect -64 1169 -28 1225
rect 28 1169 65 1225
rect -64 1007 65 1169
rect -64 951 -28 1007
rect 28 951 65 1007
rect -64 790 65 951
rect -64 734 -28 790
rect 28 734 65 790
rect -64 572 65 734
rect -64 516 -28 572
rect 28 516 65 572
rect -64 355 65 516
rect -64 299 -28 355
rect 28 299 65 355
rect -64 137 65 299
rect -64 81 -28 137
rect 28 81 65 137
rect -64 -81 65 81
rect -64 -137 -28 -81
rect 28 -137 65 -81
rect -64 -299 65 -137
rect -64 -355 -28 -299
rect 28 -355 65 -299
rect -64 -516 65 -355
rect -64 -572 -28 -516
rect 28 -572 65 -516
rect -64 -734 65 -572
rect -64 -790 -28 -734
rect 28 -790 65 -734
rect -64 -951 65 -790
rect -64 -1007 -28 -951
rect 28 -1007 65 -951
rect -64 -1169 65 -1007
rect -64 -1225 -28 -1169
rect 28 -1225 65 -1169
rect -64 -1387 65 -1225
rect -64 -1443 -28 -1387
rect 28 -1443 65 -1387
rect -64 -1604 65 -1443
rect -64 -1660 -28 -1604
rect 28 -1660 65 -1604
rect -64 -1822 65 -1660
rect -64 -1878 -28 -1822
rect 28 -1878 65 -1822
rect -64 -1916 65 -1878
<< via2 >>
rect -28 1822 28 1878
rect -28 1604 28 1660
rect -28 1387 28 1443
rect -28 1169 28 1225
rect -28 951 28 1007
rect -28 734 28 790
rect -28 516 28 572
rect -28 299 28 355
rect -28 81 28 137
rect -28 -137 28 -81
rect -28 -355 28 -299
rect -28 -572 28 -516
rect -28 -790 28 -734
rect -28 -1007 28 -951
rect -28 -1225 28 -1169
rect -28 -1443 28 -1387
rect -28 -1660 28 -1604
rect -28 -1878 28 -1822
<< metal3 >>
rect -65 1878 65 1917
rect -65 1822 -28 1878
rect 28 1822 65 1878
rect -65 1660 65 1822
rect -65 1604 -28 1660
rect 28 1604 65 1660
rect -65 1443 65 1604
rect -65 1387 -28 1443
rect 28 1387 65 1443
rect -65 1225 65 1387
rect -65 1169 -28 1225
rect 28 1169 65 1225
rect -65 1007 65 1169
rect -65 951 -28 1007
rect 28 951 65 1007
rect -65 790 65 951
rect -65 734 -28 790
rect 28 734 65 790
rect -65 572 65 734
rect -65 516 -28 572
rect 28 516 65 572
rect -65 355 65 516
rect -65 299 -28 355
rect 28 299 65 355
rect -65 137 65 299
rect -65 81 -28 137
rect 28 81 65 137
rect -65 -81 65 81
rect -65 -137 -28 -81
rect 28 -137 65 -81
rect -65 -299 65 -137
rect -65 -355 -28 -299
rect 28 -355 65 -299
rect -65 -516 65 -355
rect -65 -572 -28 -516
rect 28 -572 65 -516
rect -65 -734 65 -572
rect -65 -790 -28 -734
rect 28 -790 65 -734
rect -65 -951 65 -790
rect -65 -1007 -28 -951
rect 28 -1007 65 -951
rect -65 -1169 65 -1007
rect -65 -1225 -28 -1169
rect 28 -1225 65 -1169
rect -65 -1387 65 -1225
rect -65 -1443 -28 -1387
rect 28 -1443 65 -1387
rect -65 -1604 65 -1443
rect -65 -1660 -28 -1604
rect 28 -1660 65 -1604
rect -65 -1822 65 -1660
rect -65 -1878 -28 -1822
rect 28 -1878 65 -1822
rect -65 -1917 65 -1878
<< properties >>
string GDS_END 861096
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 859812
<< end >>
