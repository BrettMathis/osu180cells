magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 644
<< mvpmos >>
rect 0 0 120 524
<< mvpdiff >>
rect -88 511 0 524
rect -88 465 -75 511
rect -29 465 0 511
rect -88 398 0 465
rect -88 352 -75 398
rect -29 352 0 398
rect -88 285 0 352
rect -88 239 -75 285
rect -29 239 0 285
rect -88 172 0 239
rect -88 126 -75 172
rect -29 126 0 172
rect -88 59 0 126
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 511 208 524
rect 120 465 149 511
rect 195 465 208 511
rect 120 398 208 465
rect 120 352 149 398
rect 195 352 208 398
rect 120 285 208 352
rect 120 239 149 285
rect 195 239 208 285
rect 120 172 208 239
rect 120 126 149 172
rect 195 126 208 172
rect 120 59 208 126
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 465 -29 511
rect -75 352 -29 398
rect -75 239 -29 285
rect -75 126 -29 172
rect -75 13 -29 59
rect 149 465 195 511
rect 149 352 195 398
rect 149 239 195 285
rect 149 126 195 172
rect 149 13 195 59
<< polysilicon >>
rect 0 524 120 568
rect 0 -44 120 0
<< metal1 >>
rect -75 511 -29 524
rect -75 398 -29 465
rect -75 285 -29 352
rect -75 172 -29 239
rect -75 59 -29 126
rect -75 0 -29 13
rect 149 511 195 524
rect 149 398 195 465
rect 149 285 195 352
rect 149 172 195 239
rect 149 59 195 126
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 262 -52 262 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 262 172 262 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 322214
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 320614
<< end >>
