magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect 0 0 1000 1000
<< metal3 >>
rect 0 -282 1000 650
use M2_M143105899832110_64x8m81  M2_M143105899832110_64x8m81_0
timestamp 1669390400
transform 1 0 500 0 1 485
box -472 -472 472 472
use M3_M243105899832111_64x8m81  M3_M243105899832111_64x8m81_0
timestamp 1669390400
transform 1 0 500 0 1 299
box -472 -286 472 286
<< properties >>
string GDS_END 2258784
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2258548
<< end >>
