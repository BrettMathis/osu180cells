magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -381 246 381 284
rect -381 190 -345 246
rect -289 190 -134 246
rect -78 190 78 246
rect 134 190 289 246
rect 345 190 381 246
rect -381 28 381 190
rect -381 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 381 28
rect -381 -190 381 -28
rect -381 -246 -345 -190
rect -289 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 289 -190
rect 345 -246 381 -190
rect -381 -284 381 -246
<< via2 >>
rect -345 190 -289 246
rect -134 190 -78 246
rect 78 190 134 246
rect 289 190 345 246
rect -345 -28 -289 28
rect -134 -28 -78 28
rect 78 -28 134 28
rect 289 -28 345 28
rect -345 -246 -289 -190
rect -134 -246 -78 -190
rect 78 -246 134 -190
rect 289 -246 345 -190
<< metal3 >>
rect -381 246 381 284
rect -381 190 -345 246
rect -289 190 -134 246
rect -78 190 78 246
rect 134 190 289 246
rect 345 190 381 246
rect -381 28 381 190
rect -381 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 381 28
rect -381 -190 381 -28
rect -381 -246 -345 -190
rect -289 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 289 -190
rect 345 -246 381 -190
rect -381 -284 381 -246
<< properties >>
string GDS_END 2225066
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2224166
<< end >>
