magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 344 595
<< polysilicon >>
rect -31 454 89 527
rect -31 -73 89 -1
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 574
<< properties >>
string GDS_END 208224
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 207910
<< end >>
