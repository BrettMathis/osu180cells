magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 92 93 128
rect 0 40 20 92
rect 72 40 93 92
rect 0 0 93 40
<< via1 >>
rect 20 40 72 92
<< metal2 >>
rect 0 94 93 127
rect 0 66 18 94
rect -1 54 18 66
rect 0 38 18 54
rect 74 38 93 94
rect 0 -1 93 38
<< via2 >>
rect 18 92 74 94
rect 18 40 20 92
rect 20 40 72 92
rect 72 40 74 92
rect 18 38 74 40
<< metal3 >>
rect 0 94 93 128
rect 0 38 18 94
rect 74 38 93 94
rect 0 -1 93 38
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 0
box 0 0 1 1
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 35662
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 35574
<< end >>
