magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect 0 111 128 123
rect 28 92 33 111
rect 61 95 66 104
rect 60 81 66 95
rect 94 92 99 111
rect 70 60 80 66
rect 25 44 35 50
rect 91 44 101 50
rect 28 12 33 36
rect 60 28 66 39
rect 61 19 66 28
rect 94 12 99 36
rect 0 0 128 12
<< obsm1 >>
rect 11 66 16 104
rect 111 76 116 104
rect 55 71 116 76
rect 11 60 48 66
rect 11 19 16 60
rect 42 50 48 60
rect 55 58 61 71
rect 42 44 70 50
rect 111 19 116 71
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 60 90 66 95
rect 59 82 67 90
rect 59 81 66 82
rect 27 51 33 52
rect 26 43 34 51
rect 27 24 33 43
rect 59 38 65 81
rect 72 67 79 68
rect 71 59 80 67
rect 72 58 80 59
rect 58 30 68 38
rect 74 24 80 58
rect 93 51 99 52
rect 92 50 100 51
rect 91 44 101 50
rect 92 43 100 44
rect 93 42 99 43
rect 27 18 80 24
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
<< labels >>
rlabel metal2 s 27 18 33 52 6 A
port 1 nsew signal input
rlabel metal2 s 26 43 34 51 6 A
port 1 nsew signal input
rlabel metal2 s 27 18 80 24 6 A
port 1 nsew signal input
rlabel metal2 s 72 58 79 68 6 A
port 1 nsew signal input
rlabel metal2 s 74 18 80 67 6 A
port 1 nsew signal input
rlabel metal2 s 71 59 80 67 6 A
port 1 nsew signal input
rlabel metal1 s 25 44 35 50 6 A
port 1 nsew signal input
rlabel metal1 s 70 60 80 66 6 A
port 1 nsew signal input
rlabel metal2 s 93 42 99 52 6 B
port 3 nsew signal input
rlabel metal2 s 92 43 100 51 6 B
port 3 nsew signal input
rlabel metal2 s 91 44 101 50 6 B
port 3 nsew signal input
rlabel metal1 s 91 44 101 50 6 B
port 3 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 28 92 33 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 94 92 99 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 111 128 123 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 94 0 99 36 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 0 0 128 12 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 59 30 65 90 6 Y
port 2 nsew signal output
rlabel metal2 s 60 81 66 95 6 Y
port 2 nsew signal output
rlabel metal2 s 59 82 67 90 6 Y
port 2 nsew signal output
rlabel metal2 s 58 30 68 38 6 Y
port 2 nsew signal output
rlabel metal1 s 60 81 66 95 6 Y
port 2 nsew signal output
rlabel metal1 s 61 81 66 104 6 Y
port 2 nsew signal output
rlabel metal1 s 61 19 66 39 6 Y
port 2 nsew signal output
rlabel metal1 s 60 28 66 39 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 128 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 456236
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 445158
<< end >>
