magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 11116 28588 11245 28628
rect 11116 28536 11154 28588
rect 11206 28536 11245 28588
rect 11116 28509 11245 28536
rect 11116 28496 11244 28509
rect 11871 28357 12000 28397
rect 11871 28305 11909 28357
rect 11961 28305 12000 28357
rect 11871 28278 12000 28305
rect 11871 28265 11999 28278
rect 15156 28248 15285 28288
rect 15156 28196 15194 28248
rect 15246 28196 15285 28248
rect 15156 28169 15285 28196
rect 15156 28156 15284 28169
rect 15534 27604 15663 27644
rect 15534 27552 15572 27604
rect 15624 27552 15663 27604
rect 11871 27495 12000 27535
rect 15534 27525 15663 27552
rect 15534 27512 15662 27525
rect 11871 27443 11909 27495
rect 11961 27443 12000 27495
rect 11871 27416 12000 27443
rect 11871 27403 11999 27416
rect 11116 27264 11245 27304
rect 11116 27212 11154 27264
rect 11206 27212 11245 27264
rect 11116 27185 11245 27212
rect 11116 27172 11244 27185
rect 11116 26788 11245 26828
rect 11116 26736 11154 26788
rect 11206 26736 11245 26788
rect 11116 26709 11245 26736
rect 11116 26696 11244 26709
rect 11871 26557 12000 26597
rect 11871 26505 11909 26557
rect 11961 26505 12000 26557
rect 11871 26478 12000 26505
rect 11871 26465 11999 26478
rect 15912 26448 16041 26488
rect 15912 26396 15950 26448
rect 16002 26396 16041 26448
rect 15912 26369 16041 26396
rect 15912 26356 16040 26369
rect 16290 25804 16419 25844
rect 16290 25752 16328 25804
rect 16380 25752 16419 25804
rect 11871 25695 12000 25735
rect 16290 25725 16419 25752
rect 16290 25712 16418 25725
rect 11871 25643 11909 25695
rect 11961 25643 12000 25695
rect 11871 25616 12000 25643
rect 11871 25603 11999 25616
rect 11116 25464 11245 25504
rect 11116 25412 11154 25464
rect 11206 25412 11245 25464
rect 11116 25385 11245 25412
rect 11116 25372 11244 25385
rect 11116 24988 11245 25028
rect 11116 24936 11154 24988
rect 11206 24936 11245 24988
rect 11116 24909 11245 24936
rect 11116 24896 11244 24909
rect 11871 24757 12000 24797
rect 11871 24705 11909 24757
rect 11961 24705 12000 24757
rect 11871 24678 12000 24705
rect 11871 24665 11999 24678
rect 16667 24648 16796 24688
rect 16667 24596 16705 24648
rect 16757 24596 16796 24648
rect 16667 24569 16796 24596
rect 16667 24556 16795 24569
rect 17045 24004 17174 24044
rect 17045 23952 17083 24004
rect 17135 23952 17174 24004
rect 11871 23895 12000 23935
rect 17045 23925 17174 23952
rect 17045 23912 17173 23925
rect 11871 23843 11909 23895
rect 11961 23843 12000 23895
rect 11871 23816 12000 23843
rect 11871 23803 11999 23816
rect 11116 23664 11245 23704
rect 11116 23612 11154 23664
rect 11206 23612 11245 23664
rect 11116 23585 11245 23612
rect 11116 23572 11244 23585
rect 11116 23188 11245 23228
rect 11116 23136 11154 23188
rect 11206 23136 11245 23188
rect 11116 23109 11245 23136
rect 11116 23096 11244 23109
rect 11871 22957 12000 22997
rect 11871 22905 11909 22957
rect 11961 22905 12000 22957
rect 11871 22878 12000 22905
rect 11871 22865 11999 22878
rect 17423 22848 17552 22888
rect 17423 22796 17461 22848
rect 17513 22796 17552 22848
rect 17423 22769 17552 22796
rect 17423 22756 17551 22769
rect 17800 22204 17929 22244
rect 17800 22152 17838 22204
rect 17890 22152 17929 22204
rect 11871 22095 12000 22135
rect 17800 22125 17929 22152
rect 17800 22112 17928 22125
rect 11871 22043 11909 22095
rect 11961 22043 12000 22095
rect 11871 22016 12000 22043
rect 11871 22003 11999 22016
rect 11116 21864 11245 21904
rect 11116 21812 11154 21864
rect 11206 21812 11245 21864
rect 11116 21785 11245 21812
rect 11116 21772 11244 21785
rect 11116 21388 11245 21428
rect 11116 21336 11154 21388
rect 11206 21336 11245 21388
rect 11116 21309 11245 21336
rect 11116 21296 11244 21309
rect 12249 21157 12378 21197
rect 12249 21105 12287 21157
rect 12339 21105 12378 21157
rect 12249 21078 12378 21105
rect 12249 21065 12377 21078
rect 15156 21048 15285 21088
rect 15156 20996 15194 21048
rect 15246 20996 15285 21048
rect 15156 20969 15285 20996
rect 15156 20956 15284 20969
rect 15534 20404 15663 20444
rect 15534 20352 15572 20404
rect 15624 20352 15663 20404
rect 12249 20295 12378 20335
rect 15534 20325 15663 20352
rect 15534 20312 15662 20325
rect 12249 20243 12287 20295
rect 12339 20243 12378 20295
rect 12249 20216 12378 20243
rect 12249 20203 12377 20216
rect 11116 20064 11245 20104
rect 11116 20012 11154 20064
rect 11206 20012 11245 20064
rect 11116 19985 11245 20012
rect 11116 19972 11244 19985
rect 11116 19588 11245 19628
rect 11116 19536 11154 19588
rect 11206 19536 11245 19588
rect 11116 19509 11245 19536
rect 11116 19496 11244 19509
rect 12249 19357 12378 19397
rect 12249 19305 12287 19357
rect 12339 19305 12378 19357
rect 12249 19278 12378 19305
rect 12249 19265 12377 19278
rect 15912 19248 16041 19288
rect 15912 19196 15950 19248
rect 16002 19196 16041 19248
rect 15912 19169 16041 19196
rect 15912 19156 16040 19169
rect 16290 18604 16419 18644
rect 16290 18552 16328 18604
rect 16380 18552 16419 18604
rect 12249 18495 12378 18535
rect 16290 18525 16419 18552
rect 16290 18512 16418 18525
rect 12249 18443 12287 18495
rect 12339 18443 12378 18495
rect 12249 18416 12378 18443
rect 12249 18403 12377 18416
rect 11116 18264 11245 18304
rect 11116 18212 11154 18264
rect 11206 18212 11245 18264
rect 11116 18185 11245 18212
rect 11116 18172 11244 18185
rect 11116 17788 11245 17828
rect 11116 17736 11154 17788
rect 11206 17736 11245 17788
rect 11116 17709 11245 17736
rect 11116 17696 11244 17709
rect 12249 17557 12378 17597
rect 12249 17505 12287 17557
rect 12339 17505 12378 17557
rect 12249 17478 12378 17505
rect 12249 17465 12377 17478
rect 16667 17448 16796 17488
rect 16667 17396 16705 17448
rect 16757 17396 16796 17448
rect 16667 17369 16796 17396
rect 16667 17356 16795 17369
rect 17045 16804 17174 16844
rect 17045 16752 17083 16804
rect 17135 16752 17174 16804
rect 12249 16695 12378 16735
rect 17045 16725 17174 16752
rect 17045 16712 17173 16725
rect 12249 16643 12287 16695
rect 12339 16643 12378 16695
rect 12249 16616 12378 16643
rect 12249 16603 12377 16616
rect 11116 16464 11245 16504
rect 11116 16412 11154 16464
rect 11206 16412 11245 16464
rect 11116 16385 11245 16412
rect 11116 16372 11244 16385
rect 11116 15988 11245 16028
rect 11116 15936 11154 15988
rect 11206 15936 11245 15988
rect 11116 15909 11245 15936
rect 11116 15896 11244 15909
rect 12249 15757 12378 15797
rect 12249 15705 12287 15757
rect 12339 15705 12378 15757
rect 12249 15678 12378 15705
rect 12249 15665 12377 15678
rect 17423 15648 17552 15688
rect 17423 15596 17461 15648
rect 17513 15596 17552 15648
rect 17423 15569 17552 15596
rect 17423 15556 17551 15569
rect 17800 15004 17929 15044
rect 17800 14952 17838 15004
rect 17890 14952 17929 15004
rect 12249 14895 12378 14935
rect 17800 14925 17929 14952
rect 17800 14912 17928 14925
rect 12249 14843 12287 14895
rect 12339 14843 12378 14895
rect 12249 14816 12378 14843
rect 12249 14803 12377 14816
rect 11116 14664 11245 14704
rect 11116 14612 11154 14664
rect 11206 14612 11245 14664
rect 11116 14585 11245 14612
rect 11116 14572 11244 14585
rect 11116 14188 11245 14228
rect 11116 14136 11154 14188
rect 11206 14136 11245 14188
rect 11116 14109 11245 14136
rect 11116 14096 11244 14109
rect 12627 13957 12756 13997
rect 12627 13905 12665 13957
rect 12717 13905 12756 13957
rect 12627 13878 12756 13905
rect 12627 13865 12755 13878
rect 15156 13848 15285 13888
rect 15156 13796 15194 13848
rect 15246 13796 15285 13848
rect 15156 13769 15285 13796
rect 15156 13756 15284 13769
rect 15534 13204 15663 13244
rect 15534 13152 15572 13204
rect 15624 13152 15663 13204
rect 12627 13095 12756 13135
rect 15534 13125 15663 13152
rect 15534 13112 15662 13125
rect 12627 13043 12665 13095
rect 12717 13043 12756 13095
rect 12627 13016 12756 13043
rect 12627 13003 12755 13016
rect 11116 12864 11245 12904
rect 11116 12812 11154 12864
rect 11206 12812 11245 12864
rect 11116 12785 11245 12812
rect 11116 12772 11244 12785
rect 11116 12388 11245 12428
rect 11116 12336 11154 12388
rect 11206 12336 11245 12388
rect 11116 12309 11245 12336
rect 11116 12296 11244 12309
rect 12627 12157 12756 12197
rect 12627 12105 12665 12157
rect 12717 12105 12756 12157
rect 12627 12078 12756 12105
rect 12627 12065 12755 12078
rect 15912 12048 16041 12088
rect 15912 11996 15950 12048
rect 16002 11996 16041 12048
rect 15912 11969 16041 11996
rect 15912 11956 16040 11969
rect 16290 11404 16419 11444
rect 16290 11352 16328 11404
rect 16380 11352 16419 11404
rect 12627 11295 12756 11335
rect 16290 11325 16419 11352
rect 16290 11312 16418 11325
rect 12627 11243 12665 11295
rect 12717 11243 12756 11295
rect 12627 11216 12756 11243
rect 12627 11203 12755 11216
rect 11116 11064 11245 11104
rect 11116 11012 11154 11064
rect 11206 11012 11245 11064
rect 11116 10985 11245 11012
rect 11116 10972 11244 10985
rect 11116 10588 11245 10628
rect 11116 10536 11154 10588
rect 11206 10536 11245 10588
rect 11116 10509 11245 10536
rect 11116 10496 11244 10509
rect 12627 10357 12756 10397
rect 12627 10305 12665 10357
rect 12717 10305 12756 10357
rect 12627 10278 12756 10305
rect 12627 10265 12755 10278
rect 16667 10248 16796 10288
rect 16667 10196 16705 10248
rect 16757 10196 16796 10248
rect 16667 10169 16796 10196
rect 16667 10156 16795 10169
rect 17045 9604 17174 9644
rect 17045 9552 17083 9604
rect 17135 9552 17174 9604
rect 12627 9495 12756 9535
rect 17045 9525 17174 9552
rect 17045 9512 17173 9525
rect 12627 9443 12665 9495
rect 12717 9443 12756 9495
rect 12627 9416 12756 9443
rect 12627 9403 12755 9416
rect 11116 9264 11245 9304
rect 11116 9212 11154 9264
rect 11206 9212 11245 9264
rect 11116 9185 11245 9212
rect 11116 9172 11244 9185
rect 11116 8788 11245 8828
rect 11116 8736 11154 8788
rect 11206 8736 11245 8788
rect 11116 8709 11245 8736
rect 11116 8696 11244 8709
rect 12627 8557 12756 8597
rect 12627 8505 12665 8557
rect 12717 8505 12756 8557
rect 12627 8478 12756 8505
rect 12627 8465 12755 8478
rect 17423 8448 17552 8488
rect 17423 8396 17461 8448
rect 17513 8396 17552 8448
rect 17423 8369 17552 8396
rect 17423 8356 17551 8369
rect 17800 7804 17929 7844
rect 17800 7752 17838 7804
rect 17890 7752 17929 7804
rect 12627 7695 12756 7735
rect 17800 7725 17929 7752
rect 17800 7712 17928 7725
rect 12627 7643 12665 7695
rect 12717 7643 12756 7695
rect 12627 7616 12756 7643
rect 12627 7603 12755 7616
rect 11116 7464 11245 7504
rect 11116 7412 11154 7464
rect 11206 7412 11245 7464
rect 11116 7385 11245 7412
rect 11116 7372 11244 7385
rect 11116 6988 11245 7028
rect 11116 6936 11154 6988
rect 11206 6936 11245 6988
rect 11116 6909 11245 6936
rect 11116 6896 11244 6909
rect 13004 6757 13133 6797
rect 13004 6705 13042 6757
rect 13094 6705 13133 6757
rect 13004 6678 13133 6705
rect 13004 6665 13132 6678
rect 15156 6648 15285 6688
rect 15156 6596 15194 6648
rect 15246 6596 15285 6648
rect 15156 6569 15285 6596
rect 15156 6556 15284 6569
rect 15534 6004 15663 6044
rect 15534 5952 15572 6004
rect 15624 5952 15663 6004
rect 13004 5895 13133 5935
rect 15534 5925 15663 5952
rect 15534 5912 15662 5925
rect 13004 5843 13042 5895
rect 13094 5843 13133 5895
rect 13004 5816 13133 5843
rect 13004 5803 13132 5816
rect 11116 5664 11245 5704
rect 11116 5612 11154 5664
rect 11206 5612 11245 5664
rect 11116 5585 11245 5612
rect 11116 5572 11244 5585
rect 11116 5188 11245 5228
rect 11116 5136 11154 5188
rect 11206 5136 11245 5188
rect 11116 5109 11245 5136
rect 11116 5096 11244 5109
rect 13004 4957 13133 4997
rect 13004 4905 13042 4957
rect 13094 4905 13133 4957
rect 13004 4878 13133 4905
rect 13004 4865 13132 4878
rect 15912 4848 16041 4888
rect 15912 4796 15950 4848
rect 16002 4796 16041 4848
rect 15912 4769 16041 4796
rect 15912 4756 16040 4769
rect 16290 4204 16419 4244
rect 16290 4152 16328 4204
rect 16380 4152 16419 4204
rect 13004 4095 13133 4135
rect 16290 4125 16419 4152
rect 16290 4112 16418 4125
rect 13004 4043 13042 4095
rect 13094 4043 13133 4095
rect 13004 4016 13133 4043
rect 13004 4003 13132 4016
rect 11116 3864 11245 3904
rect 11116 3812 11154 3864
rect 11206 3812 11245 3864
rect 11116 3785 11245 3812
rect 11116 3772 11244 3785
rect 11116 3388 11245 3428
rect 11116 3336 11154 3388
rect 11206 3336 11245 3388
rect 11116 3309 11245 3336
rect 11116 3296 11244 3309
rect 13004 3157 13133 3197
rect 13004 3105 13042 3157
rect 13094 3105 13133 3157
rect 13004 3078 13133 3105
rect 13004 3065 13132 3078
rect 16667 3048 16796 3088
rect 16667 2996 16705 3048
rect 16757 2996 16796 3048
rect 16667 2969 16796 2996
rect 16667 2956 16795 2969
rect 17045 2404 17174 2444
rect 17045 2352 17083 2404
rect 17135 2352 17174 2404
rect 13004 2295 13133 2335
rect 17045 2325 17174 2352
rect 17045 2312 17173 2325
rect 13004 2243 13042 2295
rect 13094 2243 13133 2295
rect 13004 2216 13133 2243
rect 13004 2203 13132 2216
rect 11116 2064 11245 2104
rect 11116 2012 11154 2064
rect 11206 2012 11245 2064
rect 11116 1985 11245 2012
rect 11116 1972 11244 1985
rect 11116 1588 11245 1628
rect 11116 1536 11154 1588
rect 11206 1536 11245 1588
rect 11116 1509 11245 1536
rect 11116 1496 11244 1509
rect 13004 1357 13133 1397
rect 13004 1305 13042 1357
rect 13094 1305 13133 1357
rect 13004 1278 13133 1305
rect 13004 1265 13132 1278
rect 17423 1248 17552 1288
rect 17423 1196 17461 1248
rect 17513 1196 17552 1248
rect 17423 1169 17552 1196
rect 17423 1156 17551 1169
rect 17800 604 17929 644
rect 17800 552 17838 604
rect 17890 552 17929 604
rect 13004 495 13133 535
rect 17800 525 17929 552
rect 17800 512 17928 525
rect 13004 443 13042 495
rect 13094 443 13133 495
rect 13004 416 13133 443
rect 13004 403 13132 416
rect 11116 264 11245 304
rect 11116 212 11154 264
rect 11206 212 11245 264
rect 11116 185 11245 212
rect 11116 172 11244 185
<< via1 >>
rect 11154 28536 11206 28588
rect 11909 28305 11961 28357
rect 15194 28196 15246 28248
rect 15572 27552 15624 27604
rect 11909 27443 11961 27495
rect 11154 27212 11206 27264
rect 11154 26736 11206 26788
rect 11909 26505 11961 26557
rect 15950 26396 16002 26448
rect 16328 25752 16380 25804
rect 11909 25643 11961 25695
rect 11154 25412 11206 25464
rect 11154 24936 11206 24988
rect 11909 24705 11961 24757
rect 16705 24596 16757 24648
rect 17083 23952 17135 24004
rect 11909 23843 11961 23895
rect 11154 23612 11206 23664
rect 11154 23136 11206 23188
rect 11909 22905 11961 22957
rect 17461 22796 17513 22848
rect 17838 22152 17890 22204
rect 11909 22043 11961 22095
rect 11154 21812 11206 21864
rect 11154 21336 11206 21388
rect 12287 21105 12339 21157
rect 15194 20996 15246 21048
rect 15572 20352 15624 20404
rect 12287 20243 12339 20295
rect 11154 20012 11206 20064
rect 11154 19536 11206 19588
rect 12287 19305 12339 19357
rect 15950 19196 16002 19248
rect 16328 18552 16380 18604
rect 12287 18443 12339 18495
rect 11154 18212 11206 18264
rect 11154 17736 11206 17788
rect 12287 17505 12339 17557
rect 16705 17396 16757 17448
rect 17083 16752 17135 16804
rect 12287 16643 12339 16695
rect 11154 16412 11206 16464
rect 11154 15936 11206 15988
rect 12287 15705 12339 15757
rect 17461 15596 17513 15648
rect 17838 14952 17890 15004
rect 12287 14843 12339 14895
rect 11154 14612 11206 14664
rect 11154 14136 11206 14188
rect 12665 13905 12717 13957
rect 15194 13796 15246 13848
rect 15572 13152 15624 13204
rect 12665 13043 12717 13095
rect 11154 12812 11206 12864
rect 11154 12336 11206 12388
rect 12665 12105 12717 12157
rect 15950 11996 16002 12048
rect 16328 11352 16380 11404
rect 12665 11243 12717 11295
rect 11154 11012 11206 11064
rect 11154 10536 11206 10588
rect 12665 10305 12717 10357
rect 16705 10196 16757 10248
rect 17083 9552 17135 9604
rect 12665 9443 12717 9495
rect 11154 9212 11206 9264
rect 11154 8736 11206 8788
rect 12665 8505 12717 8557
rect 17461 8396 17513 8448
rect 17838 7752 17890 7804
rect 12665 7643 12717 7695
rect 11154 7412 11206 7464
rect 11154 6936 11206 6988
rect 13042 6705 13094 6757
rect 15194 6596 15246 6648
rect 15572 5952 15624 6004
rect 13042 5843 13094 5895
rect 11154 5612 11206 5664
rect 11154 5136 11206 5188
rect 13042 4905 13094 4957
rect 15950 4796 16002 4848
rect 16328 4152 16380 4204
rect 13042 4043 13094 4095
rect 11154 3812 11206 3864
rect 11154 3336 11206 3388
rect 13042 3105 13094 3157
rect 16705 2996 16757 3048
rect 17083 2352 17135 2404
rect 13042 2243 13094 2295
rect 11154 2012 11206 2064
rect 11154 1536 11206 1588
rect 13042 1305 13094 1357
rect 17461 1196 17513 1248
rect 17838 552 17890 604
rect 13042 443 13094 495
rect 11154 212 11206 264
<< metal2 >>
rect 11116 28588 11244 28629
rect 11116 28536 11154 28588
rect 11206 28536 11244 28588
rect 11116 28495 11244 28536
rect 11871 28357 11999 28398
rect 11871 28305 11909 28357
rect 11961 28305 11999 28357
rect 11871 28264 11999 28305
rect 15156 28248 15284 28289
rect 15156 28196 15194 28248
rect 15246 28196 15284 28248
rect 15156 28155 15284 28196
rect 15534 27604 15662 27645
rect 15534 27552 15572 27604
rect 15624 27552 15662 27604
rect 11871 27495 11999 27536
rect 15534 27511 15662 27552
rect 11871 27443 11909 27495
rect 11961 27443 11999 27495
rect 11871 27402 11999 27443
rect 11116 27264 11244 27305
rect 11116 27212 11154 27264
rect 11206 27212 11244 27264
rect 11116 27171 11244 27212
rect 11116 26788 11244 26829
rect 11116 26736 11154 26788
rect 11206 26736 11244 26788
rect 11116 26695 11244 26736
rect 11871 26557 11999 26598
rect 11871 26505 11909 26557
rect 11961 26505 11999 26557
rect 11871 26464 11999 26505
rect 15912 26448 16040 26489
rect 15912 26396 15950 26448
rect 16002 26396 16040 26448
rect 15912 26355 16040 26396
rect 16290 25804 16418 25845
rect 16290 25752 16328 25804
rect 16380 25752 16418 25804
rect 11871 25695 11999 25736
rect 16290 25711 16418 25752
rect 11871 25643 11909 25695
rect 11961 25643 11999 25695
rect 11871 25602 11999 25643
rect 11116 25464 11244 25505
rect 11116 25412 11154 25464
rect 11206 25412 11244 25464
rect 11116 25371 11244 25412
rect 11116 24988 11244 25029
rect 11116 24936 11154 24988
rect 11206 24936 11244 24988
rect 11116 24895 11244 24936
rect 11871 24757 11999 24798
rect 11871 24705 11909 24757
rect 11961 24705 11999 24757
rect 11871 24664 11999 24705
rect 16667 24648 16795 24689
rect 16667 24596 16705 24648
rect 16757 24596 16795 24648
rect 16667 24555 16795 24596
rect 17045 24004 17173 24045
rect 17045 23952 17083 24004
rect 17135 23952 17173 24004
rect 11871 23895 11999 23936
rect 17045 23911 17173 23952
rect 11871 23843 11909 23895
rect 11961 23843 11999 23895
rect 11871 23802 11999 23843
rect 11116 23664 11244 23705
rect 11116 23612 11154 23664
rect 11206 23612 11244 23664
rect 11116 23571 11244 23612
rect 11116 23188 11244 23229
rect 11116 23136 11154 23188
rect 11206 23136 11244 23188
rect 11116 23095 11244 23136
rect 11871 22957 11999 22998
rect 11871 22905 11909 22957
rect 11961 22905 11999 22957
rect 11871 22864 11999 22905
rect 17423 22848 17551 22889
rect 17423 22796 17461 22848
rect 17513 22796 17551 22848
rect 17423 22755 17551 22796
rect 17800 22204 17928 22245
rect 17800 22152 17838 22204
rect 17890 22152 17928 22204
rect 11871 22095 11999 22136
rect 17800 22111 17928 22152
rect 11871 22043 11909 22095
rect 11961 22043 11999 22095
rect 11871 22002 11999 22043
rect 11116 21864 11244 21905
rect 11116 21812 11154 21864
rect 11206 21812 11244 21864
rect 11116 21771 11244 21812
rect 11116 21388 11244 21429
rect 11116 21336 11154 21388
rect 11206 21336 11244 21388
rect 11116 21295 11244 21336
rect 12249 21157 12377 21198
rect 12249 21105 12287 21157
rect 12339 21105 12377 21157
rect 12249 21064 12377 21105
rect 15156 21048 15284 21089
rect 15156 20996 15194 21048
rect 15246 20996 15284 21048
rect 15156 20955 15284 20996
rect 15534 20404 15662 20445
rect 15534 20352 15572 20404
rect 15624 20352 15662 20404
rect 12249 20295 12377 20336
rect 15534 20311 15662 20352
rect 12249 20243 12287 20295
rect 12339 20243 12377 20295
rect 12249 20202 12377 20243
rect 11116 20064 11244 20105
rect 11116 20012 11154 20064
rect 11206 20012 11244 20064
rect 11116 19971 11244 20012
rect 11116 19588 11244 19629
rect 11116 19536 11154 19588
rect 11206 19536 11244 19588
rect 11116 19495 11244 19536
rect 12249 19357 12377 19398
rect 12249 19305 12287 19357
rect 12339 19305 12377 19357
rect 12249 19264 12377 19305
rect 15912 19248 16040 19289
rect 15912 19196 15950 19248
rect 16002 19196 16040 19248
rect 15912 19155 16040 19196
rect 16290 18604 16418 18645
rect 16290 18552 16328 18604
rect 16380 18552 16418 18604
rect 12249 18495 12377 18536
rect 16290 18511 16418 18552
rect 12249 18443 12287 18495
rect 12339 18443 12377 18495
rect 12249 18402 12377 18443
rect 11116 18264 11244 18305
rect 11116 18212 11154 18264
rect 11206 18212 11244 18264
rect 11116 18171 11244 18212
rect 11116 17788 11244 17829
rect 11116 17736 11154 17788
rect 11206 17736 11244 17788
rect 11116 17695 11244 17736
rect 12249 17557 12377 17598
rect 12249 17505 12287 17557
rect 12339 17505 12377 17557
rect 12249 17464 12377 17505
rect 16667 17448 16795 17489
rect 16667 17396 16705 17448
rect 16757 17396 16795 17448
rect 16667 17355 16795 17396
rect 17045 16804 17173 16845
rect 17045 16752 17083 16804
rect 17135 16752 17173 16804
rect 12249 16695 12377 16736
rect 17045 16711 17173 16752
rect 12249 16643 12287 16695
rect 12339 16643 12377 16695
rect 12249 16602 12377 16643
rect 11116 16464 11244 16505
rect 11116 16412 11154 16464
rect 11206 16412 11244 16464
rect 11116 16371 11244 16412
rect 11116 15988 11244 16029
rect 11116 15936 11154 15988
rect 11206 15936 11244 15988
rect 11116 15895 11244 15936
rect 12249 15757 12377 15798
rect 12249 15705 12287 15757
rect 12339 15705 12377 15757
rect 12249 15664 12377 15705
rect 17423 15648 17551 15689
rect 17423 15596 17461 15648
rect 17513 15596 17551 15648
rect 17423 15555 17551 15596
rect 17800 15004 17928 15045
rect 17800 14952 17838 15004
rect 17890 14952 17928 15004
rect 12249 14895 12377 14936
rect 17800 14911 17928 14952
rect 12249 14843 12287 14895
rect 12339 14843 12377 14895
rect 12249 14802 12377 14843
rect 11116 14664 11244 14705
rect 11116 14612 11154 14664
rect 11206 14612 11244 14664
rect 11116 14571 11244 14612
rect 11116 14188 11244 14229
rect 11116 14136 11154 14188
rect 11206 14136 11244 14188
rect 11116 14095 11244 14136
rect 12627 13957 12755 13998
rect 12627 13905 12665 13957
rect 12717 13905 12755 13957
rect 12627 13864 12755 13905
rect 15156 13848 15284 13889
rect 15156 13796 15194 13848
rect 15246 13796 15284 13848
rect 15156 13755 15284 13796
rect 15534 13204 15662 13245
rect 15534 13152 15572 13204
rect 15624 13152 15662 13204
rect 12627 13095 12755 13136
rect 15534 13111 15662 13152
rect 12627 13043 12665 13095
rect 12717 13043 12755 13095
rect 12627 13002 12755 13043
rect 11116 12864 11244 12905
rect 11116 12812 11154 12864
rect 11206 12812 11244 12864
rect 11116 12771 11244 12812
rect 11116 12388 11244 12429
rect 11116 12336 11154 12388
rect 11206 12336 11244 12388
rect 11116 12295 11244 12336
rect 12627 12157 12755 12198
rect 12627 12105 12665 12157
rect 12717 12105 12755 12157
rect 12627 12064 12755 12105
rect 15912 12048 16040 12089
rect 15912 11996 15950 12048
rect 16002 11996 16040 12048
rect 15912 11955 16040 11996
rect 16290 11404 16418 11445
rect 16290 11352 16328 11404
rect 16380 11352 16418 11404
rect 12627 11295 12755 11336
rect 16290 11311 16418 11352
rect 12627 11243 12665 11295
rect 12717 11243 12755 11295
rect 12627 11202 12755 11243
rect 11116 11064 11244 11105
rect 11116 11012 11154 11064
rect 11206 11012 11244 11064
rect 11116 10971 11244 11012
rect 11116 10588 11244 10629
rect 11116 10536 11154 10588
rect 11206 10536 11244 10588
rect 11116 10495 11244 10536
rect 12627 10357 12755 10398
rect 12627 10305 12665 10357
rect 12717 10305 12755 10357
rect 12627 10264 12755 10305
rect 16667 10248 16795 10289
rect 16667 10196 16705 10248
rect 16757 10196 16795 10248
rect 16667 10155 16795 10196
rect 17045 9604 17173 9645
rect 17045 9552 17083 9604
rect 17135 9552 17173 9604
rect 12627 9495 12755 9536
rect 17045 9511 17173 9552
rect 12627 9443 12665 9495
rect 12717 9443 12755 9495
rect 12627 9402 12755 9443
rect 11116 9264 11244 9305
rect 11116 9212 11154 9264
rect 11206 9212 11244 9264
rect 11116 9171 11244 9212
rect 11116 8788 11244 8829
rect 11116 8736 11154 8788
rect 11206 8736 11244 8788
rect 11116 8695 11244 8736
rect 12627 8557 12755 8598
rect 12627 8505 12665 8557
rect 12717 8505 12755 8557
rect 12627 8464 12755 8505
rect 17423 8448 17551 8489
rect 17423 8396 17461 8448
rect 17513 8396 17551 8448
rect 17423 8355 17551 8396
rect 17800 7804 17928 7845
rect 17800 7752 17838 7804
rect 17890 7752 17928 7804
rect 12627 7695 12755 7736
rect 17800 7711 17928 7752
rect 12627 7643 12665 7695
rect 12717 7643 12755 7695
rect 12627 7602 12755 7643
rect 11116 7464 11244 7505
rect 11116 7412 11154 7464
rect 11206 7412 11244 7464
rect 11116 7371 11244 7412
rect 11116 6988 11244 7029
rect 11116 6936 11154 6988
rect 11206 6936 11244 6988
rect 11116 6895 11244 6936
rect 13004 6757 13132 6798
rect 13004 6705 13042 6757
rect 13094 6705 13132 6757
rect 13004 6664 13132 6705
rect 15156 6648 15284 6689
rect 15156 6596 15194 6648
rect 15246 6596 15284 6648
rect 15156 6555 15284 6596
rect 15534 6004 15662 6045
rect 15534 5952 15572 6004
rect 15624 5952 15662 6004
rect 13004 5895 13132 5936
rect 15534 5911 15662 5952
rect 13004 5843 13042 5895
rect 13094 5843 13132 5895
rect 13004 5802 13132 5843
rect 11116 5664 11244 5705
rect 11116 5612 11154 5664
rect 11206 5612 11244 5664
rect 11116 5571 11244 5612
rect 11116 5188 11244 5229
rect 11116 5136 11154 5188
rect 11206 5136 11244 5188
rect 11116 5095 11244 5136
rect 13004 4957 13132 4998
rect 13004 4905 13042 4957
rect 13094 4905 13132 4957
rect 13004 4864 13132 4905
rect 15912 4848 16040 4889
rect 15912 4796 15950 4848
rect 16002 4796 16040 4848
rect 15912 4755 16040 4796
rect 16290 4204 16418 4245
rect 16290 4152 16328 4204
rect 16380 4152 16418 4204
rect 13004 4095 13132 4136
rect 16290 4111 16418 4152
rect 13004 4043 13042 4095
rect 13094 4043 13132 4095
rect 13004 4002 13132 4043
rect 11116 3864 11244 3905
rect 11116 3812 11154 3864
rect 11206 3812 11244 3864
rect 11116 3771 11244 3812
rect 11116 3388 11244 3429
rect 11116 3336 11154 3388
rect 11206 3336 11244 3388
rect 11116 3295 11244 3336
rect 13004 3157 13132 3198
rect 13004 3105 13042 3157
rect 13094 3105 13132 3157
rect 13004 3064 13132 3105
rect 16667 3048 16795 3089
rect 16667 2996 16705 3048
rect 16757 2996 16795 3048
rect 16667 2955 16795 2996
rect 17045 2404 17173 2445
rect 17045 2352 17083 2404
rect 17135 2352 17173 2404
rect 13004 2295 13132 2336
rect 17045 2311 17173 2352
rect 13004 2243 13042 2295
rect 13094 2243 13132 2295
rect 13004 2202 13132 2243
rect 11116 2064 11244 2105
rect 11116 2012 11154 2064
rect 11206 2012 11244 2064
rect 11116 1971 11244 2012
rect 11116 1588 11244 1629
rect 11116 1536 11154 1588
rect 11206 1536 11244 1588
rect 11116 1495 11244 1536
rect 13004 1357 13132 1398
rect 13004 1305 13042 1357
rect 13094 1305 13132 1357
rect 13004 1264 13132 1305
rect 17423 1248 17551 1289
rect 17423 1196 17461 1248
rect 17513 1196 17551 1248
rect 17423 1155 17551 1196
rect 17800 604 17928 645
rect 17800 552 17838 604
rect 17890 552 17928 604
rect 13004 495 13132 536
rect 17800 511 17928 552
rect 13004 443 13042 495
rect 13094 443 13132 495
rect 13004 402 13132 443
rect 11115 264 11245 305
rect 11115 212 11154 264
rect 11206 212 11245 264
rect 11115 171 11245 212
rect 6835 -21 6965 112
rect 11871 -164 12000 -31
rect 12248 -164 12378 -31
rect 12626 -164 12755 -31
rect 13004 -164 13133 -31
rect 15156 -164 15285 -31
rect 15534 -164 15663 -31
rect 15911 -164 16041 -31
rect 16289 -164 16418 -31
rect 16667 -164 16796 -31
rect 17044 -164 17174 -31
rect 17422 -164 17551 -31
rect 17800 -164 17929 -31
<< metal3 >>
rect 131 28733 260 28867
rect 765 28293 895 28427
rect 23358 28293 23487 28427
rect 131 27833 260 27967
rect 765 27373 895 27507
rect 23358 27373 23487 27507
rect 765 26493 895 26627
rect 23358 26493 23487 26627
rect 765 25573 895 25707
rect 23358 25573 23487 25707
rect 765 24693 895 24827
rect 23358 24693 23487 24827
rect 765 23773 895 23907
rect 23358 23773 23487 23907
rect 765 22893 895 23027
rect 23358 22893 23487 23027
rect 765 21973 895 22107
rect 23358 21973 23487 22107
rect 765 21093 895 21227
rect 23358 21093 23487 21227
rect 765 20173 895 20307
rect 23358 20173 23487 20307
rect 765 19293 895 19427
rect 23358 19293 23487 19427
rect 765 18373 895 18507
rect 23358 18373 23487 18507
rect 765 17493 895 17627
rect 23358 17493 23487 17627
rect 765 16573 895 16707
rect 23358 16573 23487 16707
rect 765 15693 895 15827
rect 23358 15693 23487 15827
rect 765 14773 895 14907
rect 23358 14773 23487 14907
rect 765 13893 895 14027
rect 23358 13893 23487 14027
rect 765 12973 895 13107
rect 23358 12973 23487 13107
rect 765 12093 895 12227
rect 23358 12093 23487 12227
rect 765 11173 895 11307
rect 23358 11173 23487 11307
rect 765 10293 895 10427
rect 23358 10293 23487 10427
rect 765 9373 895 9507
rect 23358 9373 23487 9507
rect 765 8493 895 8627
rect 23358 8493 23487 8627
rect 765 7573 895 7707
rect 23358 7573 23487 7707
rect 765 6693 895 6827
rect 23358 6693 23487 6827
rect 765 5773 895 5907
rect 23358 5773 23487 5907
rect 765 4893 895 5027
rect 23358 4893 23487 5027
rect 765 3973 895 4107
rect 23358 3973 23487 4107
rect 765 3093 895 3227
rect 23358 3093 23487 3227
rect 765 2173 895 2307
rect 23358 2173 23487 2307
rect 765 1293 895 1427
rect 23358 1293 23487 1427
rect 765 373 895 507
rect 23358 373 23487 507
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_0
timestamp 1669390400
transform 1 0 11180 0 1 238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_1
timestamp 1669390400
transform 1 0 11180 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_2
timestamp 1669390400
transform 1 0 11180 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_3
timestamp 1669390400
transform 1 0 11935 0 1 22931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_4
timestamp 1669390400
transform 1 0 11935 0 1 23869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_5
timestamp 1669390400
transform 1 0 11935 0 1 24731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_6
timestamp 1669390400
transform 1 0 11935 0 1 25669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_7
timestamp 1669390400
transform 1 0 11935 0 1 26531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_8
timestamp 1669390400
transform 1 0 12313 0 1 21131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_9
timestamp 1669390400
transform 1 0 11935 0 1 28331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_10
timestamp 1669390400
transform 1 0 11935 0 1 27469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_11
timestamp 1669390400
transform 1 0 12691 0 1 7669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_12
timestamp 1669390400
transform 1 0 12691 0 1 8531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_13
timestamp 1669390400
transform 1 0 12691 0 1 9469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_14
timestamp 1669390400
transform 1 0 12691 0 1 10331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_15
timestamp 1669390400
transform 1 0 12691 0 1 11269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_16
timestamp 1669390400
transform 1 0 12691 0 1 12131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_17
timestamp 1669390400
transform 1 0 11180 0 1 28562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_18
timestamp 1669390400
transform 1 0 11180 0 1 26762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_19
timestamp 1669390400
transform 1 0 11180 0 1 24962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_20
timestamp 1669390400
transform 1 0 11180 0 1 23162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_21
timestamp 1669390400
transform 1 0 11180 0 1 21362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_22
timestamp 1669390400
transform 1 0 11180 0 1 19562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_23
timestamp 1669390400
transform 1 0 11180 0 1 17762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_24
timestamp 1669390400
transform 1 0 11180 0 1 15962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_25
timestamp 1669390400
transform 1 0 11180 0 1 14162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_26
timestamp 1669390400
transform 1 0 11180 0 1 12362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_27
timestamp 1669390400
transform 1 0 11180 0 1 10562
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_28
timestamp 1669390400
transform 1 0 11180 0 1 8762
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_29
timestamp 1669390400
transform 1 0 11180 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_30
timestamp 1669390400
transform 1 0 11180 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_31
timestamp 1669390400
transform 1 0 11180 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_32
timestamp 1669390400
transform 1 0 12313 0 1 14869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_33
timestamp 1669390400
transform 1 0 12313 0 1 15731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_34
timestamp 1669390400
transform 1 0 13068 0 1 6731
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_35
timestamp 1669390400
transform 1 0 12313 0 1 16669
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_36
timestamp 1669390400
transform 1 0 12691 0 1 13931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_37
timestamp 1669390400
transform 1 0 12691 0 1 13069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_38
timestamp 1669390400
transform 1 0 12313 0 1 17531
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_39
timestamp 1669390400
transform 1 0 12313 0 1 18469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_40
timestamp 1669390400
transform 1 0 12313 0 1 19331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_41
timestamp 1669390400
transform 1 0 13068 0 1 469
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_42
timestamp 1669390400
transform 1 0 13068 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_43
timestamp 1669390400
transform 1 0 13068 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_44
timestamp 1669390400
transform 1 0 13068 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_45
timestamp 1669390400
transform 1 0 13068 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_46
timestamp 1669390400
transform 1 0 13068 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_47
timestamp 1669390400
transform 1 0 13068 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_48
timestamp 1669390400
transform 1 0 11180 0 1 27238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_49
timestamp 1669390400
transform 1 0 11180 0 1 25438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_50
timestamp 1669390400
transform 1 0 11180 0 1 23638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_51
timestamp 1669390400
transform 1 0 11180 0 1 21838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_52
timestamp 1669390400
transform 1 0 11180 0 1 20038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_53
timestamp 1669390400
transform 1 0 11180 0 1 18238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_54
timestamp 1669390400
transform 1 0 11180 0 1 16438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_55
timestamp 1669390400
transform 1 0 11180 0 1 14638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_56
timestamp 1669390400
transform 1 0 11180 0 1 12838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_57
timestamp 1669390400
transform 1 0 11180 0 1 11038
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_58
timestamp 1669390400
transform 1 0 11180 0 1 9238
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_59
timestamp 1669390400
transform 1 0 11180 0 1 7438
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_60
timestamp 1669390400
transform 1 0 11180 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_61
timestamp 1669390400
transform 1 0 11180 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_62
timestamp 1669390400
transform 1 0 12313 0 1 20269
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_63
timestamp 1669390400
transform 1 0 11935 0 1 22069
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_64
timestamp 1669390400
transform 1 0 17864 0 1 578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_65
timestamp 1669390400
transform 1 0 17487 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_66
timestamp 1669390400
transform 1 0 17109 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_67
timestamp 1669390400
transform 1 0 16731 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_68
timestamp 1669390400
transform 1 0 16354 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_69
timestamp 1669390400
transform 1 0 15976 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_70
timestamp 1669390400
transform 1 0 15598 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_71
timestamp 1669390400
transform 1 0 15220 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_72
timestamp 1669390400
transform 1 0 15220 0 1 13822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_73
timestamp 1669390400
transform 1 0 15220 0 1 21022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_74
timestamp 1669390400
transform 1 0 15220 0 1 28222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_75
timestamp 1669390400
transform 1 0 15598 0 1 13178
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_76
timestamp 1669390400
transform 1 0 15598 0 1 20378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_77
timestamp 1669390400
transform 1 0 15598 0 1 27578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_78
timestamp 1669390400
transform 1 0 15976 0 1 12022
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_79
timestamp 1669390400
transform 1 0 15976 0 1 19222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_80
timestamp 1669390400
transform 1 0 15976 0 1 26422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_81
timestamp 1669390400
transform 1 0 16354 0 1 11378
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_82
timestamp 1669390400
transform 1 0 16354 0 1 18578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_83
timestamp 1669390400
transform 1 0 16354 0 1 25778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_84
timestamp 1669390400
transform 1 0 16731 0 1 10222
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_85
timestamp 1669390400
transform 1 0 16731 0 1 17422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_86
timestamp 1669390400
transform 1 0 16731 0 1 24622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_87
timestamp 1669390400
transform 1 0 17109 0 1 9578
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_88
timestamp 1669390400
transform 1 0 17109 0 1 16778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_89
timestamp 1669390400
transform 1 0 17109 0 1 23978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_90
timestamp 1669390400
transform 1 0 17487 0 1 8422
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_91
timestamp 1669390400
transform 1 0 17487 0 1 15622
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_92
timestamp 1669390400
transform 1 0 17487 0 1 22822
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_93
timestamp 1669390400
transform 1 0 17864 0 1 7778
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_94
timestamp 1669390400
transform 1 0 17864 0 1 14978
box 0 0 1 1
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_95
timestamp 1669390400
transform 1 0 17864 0 1 22178
box 0 0 1 1
use xdec8_512x8m81  xdec8_512x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 21600
box 0 -228 24219 7428
use xdec8_512x8m81  xdec8_512x8m81_1
timestamp 1669390400
transform 1 0 0 0 1 0
box 0 -228 24219 7428
use xdec8_512x8m81  xdec8_512x8m81_2
timestamp 1669390400
transform 1 0 0 0 1 7200
box 0 -228 24219 7428
use xdec8_512x8m81  xdec8_512x8m81_3
timestamp 1669390400
transform 1 0 0 0 1 14400
box 0 -228 24219 7428
<< labels >>
rlabel metal3 s 830 5840 830 5840 4 LWL[6]
port 1 nsew
rlabel metal3 s 830 6760 830 6760 4 LWL[7]
port 2 nsew
rlabel metal3 s 23423 16640 23423 16640 4 RWL[18]
port 3 nsew
rlabel metal3 s 23423 15760 23423 15760 4 RWL[17]
port 4 nsew
rlabel metal3 s 23423 14840 23423 14840 4 RWL[16]
port 5 nsew
rlabel metal3 s 23423 13960 23423 13960 4 RWL[15]
port 6 nsew
rlabel metal3 s 23423 13040 23423 13040 4 RWL[14]
port 7 nsew
rlabel metal3 s 23423 12160 23423 12160 4 RWL[13]
port 8 nsew
rlabel metal3 s 23423 11240 23423 11240 4 RWL[12]
port 9 nsew
rlabel metal3 s 830 8560 830 8560 4 LWL[9]
port 10 nsew
rlabel metal3 s 830 7640 830 7640 4 LWL[8]
port 11 nsew
rlabel metal3 s 830 440 830 440 4 LWL[0]
port 12 nsew
rlabel metal3 s 830 1360 830 1360 4 LWL[1]
port 13 nsew
rlabel metal3 s 830 2240 830 2240 4 LWL[2]
port 14 nsew
rlabel metal3 s 830 3160 830 3160 4 LWL[3]
port 15 nsew
rlabel metal3 s 830 4040 830 4040 4 LWL[4]
port 16 nsew
rlabel metal3 s 830 4960 830 4960 4 LWL[5]
port 17 nsew
rlabel metal3 s 23423 10360 23423 10360 4 RWL[11]
port 18 nsew
rlabel metal3 s 23423 9440 23423 9440 4 RWL[10]
port 19 nsew
rlabel metal3 s 23423 8560 23423 8560 4 RWL[9]
port 20 nsew
rlabel metal3 s 23423 7640 23423 7640 4 RWL[8]
port 21 nsew
rlabel metal3 s 23423 6760 23423 6760 4 RWL[7]
port 22 nsew
rlabel metal3 s 23423 4960 23423 4960 4 RWL[5]
port 23 nsew
rlabel metal3 s 23423 3160 23423 3160 4 RWL[3]
port 24 nsew
rlabel metal3 s 23423 1360 23423 1360 4 RWL[1]
port 25 nsew
rlabel metal3 s 23423 440 23423 440 4 RWL[0]
port 26 nsew
rlabel metal3 s 23423 2240 23423 2240 4 RWL[2]
port 27 nsew
rlabel metal3 s 830 16640 830 16640 4 LWL[18]
port 28 nsew
rlabel metal3 s 830 15760 830 15760 4 LWL[17]
port 29 nsew
rlabel metal3 s 830 14840 830 14840 4 LWL[16]
port 30 nsew
rlabel metal3 s 830 13960 830 13960 4 LWL[15]
port 31 nsew
rlabel metal3 s 830 13040 830 13040 4 LWL[14]
port 32 nsew
rlabel metal3 s 830 12160 830 12160 4 LWL[13]
port 33 nsew
rlabel metal3 s 830 11240 830 11240 4 LWL[12]
port 34 nsew
rlabel metal3 s 830 10360 830 10360 4 LWL[11]
port 35 nsew
rlabel metal3 s 830 9440 830 9440 4 LWL[10]
port 36 nsew
rlabel metal3 s 23423 4040 23423 4040 4 RWL[4]
port 37 nsew
rlabel metal3 s 23423 5840 23423 5840 4 RWL[6]
port 38 nsew
rlabel metal3 s 830 25640 830 25640 4 LWL[28]
port 39 nsew
rlabel metal3 s 830 24760 830 24760 4 LWL[27]
port 40 nsew
rlabel metal3 s 830 23840 830 23840 4 LWL[26]
port 41 nsew
rlabel metal3 s 830 22960 830 22960 4 LWL[25]
port 42 nsew
rlabel metal3 s 830 22040 830 22040 4 LWL[24]
port 43 nsew
rlabel metal3 s 830 21160 830 21160 4 LWL[23]
port 44 nsew
rlabel metal3 s 830 20240 830 20240 4 LWL[22]
port 45 nsew
rlabel metal3 s 830 19360 830 19360 4 LWL[21]
port 46 nsew
rlabel metal3 s 830 18440 830 18440 4 LWL[20]
port 47 nsew
rlabel metal3 s 830 17560 830 17560 4 LWL[19]
port 48 nsew
rlabel metal3 s 23423 18440 23423 18440 4 RWL[20]
port 49 nsew
rlabel metal3 s 23423 19360 23423 19360 4 RWL[21]
port 50 nsew
rlabel metal3 s 23423 20240 23423 20240 4 RWL[22]
port 51 nsew
rlabel metal3 s 23423 21160 23423 21160 4 RWL[23]
port 52 nsew
rlabel metal3 s 23423 22040 23423 22040 4 RWL[24]
port 53 nsew
rlabel metal3 s 23423 22960 23423 22960 4 RWL[25]
port 54 nsew
rlabel metal3 s 23423 23840 23423 23840 4 RWL[26]
port 55 nsew
rlabel metal3 s 23423 24760 23423 24760 4 RWL[27]
port 56 nsew
rlabel metal3 s 23423 25640 23423 25640 4 RWL[28]
port 57 nsew
rlabel metal3 s 23423 26560 23423 26560 4 RWL[29]
port 58 nsew
rlabel metal3 s 23423 27440 23423 27440 4 RWL[30]
port 59 nsew
rlabel metal3 s 23423 28360 23423 28360 4 RWL[31]
port 60 nsew
rlabel metal3 s 830 28360 830 28360 4 LWL[31]
port 61 nsew
rlabel metal3 s 830 27440 830 27440 4 LWL[30]
port 62 nsew
rlabel metal3 s 830 26560 830 26560 4 LWL[29]
port 63 nsew
rlabel metal3 s 195 28800 195 28800 4 vdd
port 64 nsew
rlabel metal3 s 195 27900 195 27900 4 vss
port 65 nsew
rlabel metal3 s 23423 17560 23423 17560 4 RWL[19]
port 66 nsew
rlabel metal2 s 17109 -97 17109 -97 4 xa[2]
port 67 nsew
rlabel metal2 s 6900 45 6900 45 4 men
port 68 nsew
rlabel metal2 s 17864 -97 17864 -97 4 xa[0]
port 69 nsew
rlabel metal2 s 16731 -97 16731 -97 4 xa[3]
port 70 nsew
rlabel metal2 s 16354 -97 16354 -97 4 xa[4]
port 71 nsew
rlabel metal2 s 15976 -97 15976 -97 4 xa[5]
port 72 nsew
rlabel metal2 s 15598 -97 15598 -97 4 xa[6]
port 73 nsew
rlabel metal2 s 15220 -97 15220 -97 4 xa[7]
port 74 nsew
rlabel metal2 s 11935 -97 11935 -97 4 xb[3]
port 75 nsew
rlabel metal2 s 12313 -97 12313 -97 4 xb[2]
port 76 nsew
rlabel metal2 s 12691 -97 12691 -97 4 xb[1]
port 77 nsew
rlabel metal2 s 13068 -97 13068 -97 4 xb[0]
port 78 nsew
rlabel metal2 s 11180 238 11180 238 4 xc
port 79 nsew
rlabel metal2 s 17487 -97 17487 -97 4 xa[1]
port 80 nsew
<< properties >>
string GDS_END 2020672
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2007158
<< end >>
