magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 22162 -6340 22775 -1078
rect 22448 -12800 22838 -10246
rect 22671 -14848 23429 -14394
rect 22650 -15879 23535 -14848
rect 22681 -15880 23535 -15879
rect 22685 -22093 23539 -19542
rect 22554 -23170 23539 -22714
<< pwell >>
rect -68 16256 23468 16288
rect -68 -88 23468 -56
<< psubdiff >>
rect 22869 -16594 23345 -16534
rect 22869 -16640 22926 -16594
rect 22972 -16640 23084 -16594
rect 23130 -16640 23242 -16594
rect 23288 -16640 23345 -16594
rect 22869 -16700 23345 -16640
<< nsubdiff >>
rect 22814 -14599 23286 -14542
rect 22814 -14645 22869 -14599
rect 22915 -14645 23027 -14599
rect 23073 -14645 23185 -14599
rect 23231 -14645 23286 -14599
rect 22814 -14702 23286 -14645
rect 22697 -22919 22852 -22862
rect 22697 -22965 22751 -22919
rect 22797 -22965 22852 -22919
rect 22697 -23022 22852 -22965
rect 23241 -22919 23396 -22862
rect 23241 -22965 23295 -22919
rect 23341 -22965 23396 -22919
rect 23241 -23022 23396 -22965
<< psubdiffcont >>
rect 22926 -16640 22972 -16594
rect 23084 -16640 23130 -16594
rect 23242 -16640 23288 -16594
<< nsubdiffcont >>
rect 22869 -14645 22915 -14599
rect 23027 -14645 23073 -14599
rect 23185 -14645 23231 -14599
rect 22751 -22965 22797 -22919
rect 23295 -22965 23341 -22919
<< polysilicon >>
rect -257 16129 57 16148
rect -257 15989 -238 16129
rect -192 15994 57 16129
rect 23341 16065 23711 16148
rect 23341 16019 23592 16065
rect 23638 16019 23711 16065
rect 23341 15994 23711 16019
rect -192 15989 -173 15994
rect -257 15970 -173 15989
rect 23519 15901 23711 15994
rect 23519 15855 23592 15901
rect 23638 15855 23711 15901
rect 23519 15809 23711 15855
rect -257 14470 57 14606
rect -257 14330 -238 14470
rect -192 14452 57 14470
rect 23341 14505 23711 14606
rect 23341 14459 23592 14505
rect 23638 14459 23711 14505
rect 23341 14452 23711 14459
rect -192 14348 -173 14452
rect 23519 14348 23711 14452
rect -192 14330 57 14348
rect -257 14194 57 14330
rect 23341 14341 23711 14348
rect 23341 14295 23592 14341
rect 23638 14295 23711 14341
rect 23341 14194 23711 14295
rect -257 12670 57 12806
rect -257 12530 -238 12670
rect -192 12652 57 12670
rect 23341 12705 23711 12806
rect 23341 12659 23592 12705
rect 23638 12659 23711 12705
rect 23341 12652 23711 12659
rect -192 12548 -173 12652
rect 23519 12548 23711 12652
rect -192 12530 57 12548
rect -257 12394 57 12530
rect 23341 12541 23711 12548
rect 23341 12495 23592 12541
rect 23638 12495 23711 12541
rect 23341 12394 23711 12495
rect -257 10870 57 11006
rect -257 10730 -238 10870
rect -192 10852 57 10870
rect 23341 10905 23711 11006
rect 23341 10859 23592 10905
rect 23638 10859 23711 10905
rect 23341 10852 23711 10859
rect -192 10748 -173 10852
rect 23519 10748 23711 10852
rect -192 10730 57 10748
rect -257 10594 57 10730
rect 23341 10741 23711 10748
rect 23341 10695 23592 10741
rect 23638 10695 23711 10741
rect 23341 10594 23711 10695
rect -257 9070 57 9206
rect -257 8930 -238 9070
rect -192 9052 57 9070
rect 23341 9105 23711 9206
rect 23341 9059 23592 9105
rect 23638 9059 23711 9105
rect 23341 9052 23711 9059
rect -192 8948 -173 9052
rect 23519 8948 23711 9052
rect -192 8930 57 8948
rect -257 8794 57 8930
rect 23341 8941 23711 8948
rect 23341 8895 23592 8941
rect 23638 8895 23711 8941
rect 23341 8794 23711 8895
rect -257 7270 57 7406
rect -257 7130 -238 7270
rect -192 7252 57 7270
rect 23341 7305 23711 7406
rect 23341 7259 23592 7305
rect 23638 7259 23711 7305
rect 23341 7252 23711 7259
rect -192 7148 -173 7252
rect 23519 7148 23711 7252
rect -192 7130 57 7148
rect -257 6994 57 7130
rect 23341 7141 23711 7148
rect 23341 7095 23592 7141
rect 23638 7095 23711 7141
rect 23341 6994 23711 7095
rect -257 5470 57 5606
rect -257 5330 -238 5470
rect -192 5452 57 5470
rect 23341 5505 23711 5606
rect 23341 5459 23592 5505
rect 23638 5459 23711 5505
rect 23341 5452 23711 5459
rect -192 5348 -173 5452
rect 23519 5348 23711 5452
rect -192 5330 57 5348
rect -257 5194 57 5330
rect 23341 5341 23711 5348
rect 23341 5295 23592 5341
rect 23638 5295 23711 5341
rect 23341 5194 23711 5295
rect -257 3670 57 3806
rect -257 3530 -238 3670
rect -192 3652 57 3670
rect 23341 3705 23711 3806
rect 23341 3659 23592 3705
rect 23638 3659 23711 3705
rect 23341 3652 23711 3659
rect -192 3548 -173 3652
rect 23519 3548 23711 3652
rect -192 3530 57 3548
rect -257 3394 57 3530
rect 23341 3541 23711 3548
rect 23341 3495 23592 3541
rect 23638 3495 23711 3541
rect 23341 3394 23711 3495
rect -257 1870 57 2006
rect -257 1730 -238 1870
rect -192 1852 57 1870
rect 23341 1905 23711 2006
rect 23341 1859 23592 1905
rect 23638 1859 23711 1905
rect 23341 1852 23711 1859
rect -192 1748 -173 1852
rect 23519 1748 23711 1852
rect -192 1730 57 1748
rect -257 1594 57 1730
rect 23341 1741 23711 1748
rect 23341 1695 23592 1741
rect 23638 1695 23711 1741
rect 23341 1594 23711 1695
rect 23519 345 23711 391
rect 23519 299 23592 345
rect 23638 299 23711 345
rect -257 211 -173 230
rect -257 71 -238 211
rect -192 206 -173 211
rect 23519 206 23711 299
rect -192 71 57 206
rect -257 52 57 71
rect 23395 181 23711 206
rect 23395 135 23592 181
rect 23638 135 23711 181
rect 23395 52 23711 135
rect 22957 -15781 23034 -15739
rect 23181 -15781 23258 -15739
rect 22936 -15798 23056 -15781
rect 23160 -15798 23280 -15781
rect 22936 -15814 23280 -15798
rect 22936 -15860 23569 -15814
rect 22936 -15906 23291 -15860
rect 23337 -15906 23449 -15860
rect 23495 -15906 23569 -15860
rect 22936 -15952 23569 -15906
rect 22936 -15961 23280 -15952
rect 22936 -16022 23056 -15961
rect 23160 -16022 23280 -15961
rect 22936 -16401 23056 -16319
rect 23160 -16401 23280 -16319
rect 22940 -19466 23060 -19404
rect 23164 -19466 23284 -19404
rect 22940 -19475 23284 -19466
rect 22633 -19521 23284 -19475
rect 22633 -19567 22707 -19521
rect 22753 -19567 22865 -19521
rect 22911 -19567 23284 -19521
rect 22633 -19613 23284 -19567
rect 22940 -19624 23284 -19613
rect 22940 -19640 23060 -19624
rect 23164 -19640 23284 -19624
rect 22961 -19683 23038 -19640
rect 23185 -19683 23262 -19640
<< polycontact >>
rect -238 15989 -192 16129
rect 23592 16019 23638 16065
rect 23592 15855 23638 15901
rect -238 14330 -192 14470
rect 23592 14459 23638 14505
rect 23592 14295 23638 14341
rect -238 12530 -192 12670
rect 23592 12659 23638 12705
rect 23592 12495 23638 12541
rect -238 10730 -192 10870
rect 23592 10859 23638 10905
rect 23592 10695 23638 10741
rect -238 8930 -192 9070
rect 23592 9059 23638 9105
rect 23592 8895 23638 8941
rect -238 7130 -192 7270
rect 23592 7259 23638 7305
rect 23592 7095 23638 7141
rect -238 5330 -192 5470
rect 23592 5459 23638 5505
rect 23592 5295 23638 5341
rect -238 3530 -192 3670
rect 23592 3659 23638 3705
rect 23592 3495 23638 3541
rect -238 1730 -192 1870
rect 23592 1859 23638 1905
rect 23592 1695 23638 1741
rect 23592 299 23638 345
rect -238 71 -192 211
rect 23592 135 23638 181
rect 23291 -15906 23337 -15860
rect 23449 -15906 23495 -15860
rect 22707 -19567 22753 -19521
rect 22865 -19567 22911 -19521
<< metal1 >>
rect -253 16129 -177 16140
rect -253 16128 -238 16129
rect -192 16128 -177 16129
rect -253 15868 -241 16128
rect -189 15868 -177 16128
rect -253 15856 -177 15868
rect 23551 16070 23675 16110
rect 23551 16018 23587 16070
rect 23639 16018 23675 16070
rect 23551 15901 23675 16018
rect 23551 15855 23592 15901
rect 23638 15855 23675 15901
rect 23551 15852 23675 15855
rect 23551 15800 23587 15852
rect 23639 15800 23675 15852
rect 23551 15760 23675 15800
rect -253 14530 -177 14542
rect -253 14270 -241 14530
rect -189 14270 -177 14530
rect -253 14258 -177 14270
rect 23551 14537 23675 14577
rect 23551 14485 23587 14537
rect 23639 14485 23675 14537
rect 23551 14459 23592 14485
rect 23638 14459 23675 14485
rect 23551 14341 23675 14459
rect 23551 14319 23592 14341
rect 23638 14319 23675 14341
rect 23551 14267 23587 14319
rect 23639 14267 23675 14319
rect 23551 14227 23675 14267
rect -253 12730 -177 12742
rect -253 12470 -241 12730
rect -189 12470 -177 12730
rect -253 12458 -177 12470
rect 23551 12733 23675 12773
rect 23551 12681 23587 12733
rect 23639 12681 23675 12733
rect 23551 12659 23592 12681
rect 23638 12659 23675 12681
rect 23551 12541 23675 12659
rect 23551 12515 23592 12541
rect 23638 12515 23675 12541
rect 23551 12463 23587 12515
rect 23639 12463 23675 12515
rect 23551 12423 23675 12463
rect -253 10930 -177 10942
rect -253 10670 -241 10930
rect -189 10670 -177 10930
rect -253 10658 -177 10670
rect 23551 10937 23675 10977
rect 23551 10885 23587 10937
rect 23639 10885 23675 10937
rect 23551 10859 23592 10885
rect 23638 10859 23675 10885
rect 23551 10741 23675 10859
rect 23551 10719 23592 10741
rect 23638 10719 23675 10741
rect 23551 10667 23587 10719
rect 23639 10667 23675 10719
rect 23551 10627 23675 10667
rect -253 9130 -177 9142
rect -253 8870 -241 9130
rect -189 8870 -177 9130
rect -253 8858 -177 8870
rect 23551 9133 23675 9173
rect 23551 9081 23587 9133
rect 23639 9081 23675 9133
rect 23551 9059 23592 9081
rect 23638 9059 23675 9081
rect 23551 8941 23675 9059
rect 23551 8915 23592 8941
rect 23638 8915 23675 8941
rect 23551 8863 23587 8915
rect 23639 8863 23675 8915
rect 23551 8823 23675 8863
rect -253 7330 -177 7342
rect -253 7070 -241 7330
rect -189 7070 -177 7330
rect -253 7058 -177 7070
rect 23551 7337 23675 7377
rect 23551 7285 23587 7337
rect 23639 7285 23675 7337
rect 23551 7259 23592 7285
rect 23638 7259 23675 7285
rect 23551 7141 23675 7259
rect 23551 7119 23592 7141
rect 23638 7119 23675 7141
rect 23551 7067 23587 7119
rect 23639 7067 23675 7119
rect 23551 7027 23675 7067
rect -253 5530 -177 5542
rect -253 5270 -241 5530
rect -189 5270 -177 5530
rect -253 5258 -177 5270
rect 23551 5533 23675 5573
rect 23551 5481 23587 5533
rect 23639 5481 23675 5533
rect 23551 5459 23592 5481
rect 23638 5459 23675 5481
rect 23551 5341 23675 5459
rect 23551 5315 23592 5341
rect 23638 5315 23675 5341
rect 23551 5263 23587 5315
rect 23639 5263 23675 5315
rect 23551 5223 23675 5263
rect -253 3730 -177 3742
rect -253 3470 -241 3730
rect -189 3470 -177 3730
rect -253 3458 -177 3470
rect 23551 3737 23675 3777
rect 23551 3685 23587 3737
rect 23639 3685 23675 3737
rect 23551 3659 23592 3685
rect 23638 3659 23675 3685
rect 23551 3541 23675 3659
rect 23551 3519 23592 3541
rect 23638 3519 23675 3541
rect 23551 3467 23587 3519
rect 23639 3467 23675 3519
rect 23551 3427 23675 3467
rect -253 1930 -177 1942
rect -253 1670 -241 1930
rect -189 1670 -177 1930
rect -253 1658 -177 1670
rect 23551 1933 23675 1973
rect 23551 1881 23587 1933
rect 23639 1881 23675 1933
rect 23551 1859 23592 1881
rect 23638 1859 23675 1881
rect 23551 1741 23675 1859
rect 23551 1715 23592 1741
rect 23638 1715 23675 1741
rect 23551 1663 23587 1715
rect 23639 1663 23675 1715
rect 23551 1623 23675 1663
rect 23551 400 23675 440
rect 23551 348 23587 400
rect 23639 348 23675 400
rect 23551 345 23675 348
rect 23551 299 23592 345
rect 23638 299 23675 345
rect -249 211 -181 222
rect -249 71 -238 211
rect -192 71 -181 211
rect 23551 182 23675 299
rect 23551 130 23587 182
rect 23639 130 23675 182
rect 23551 90 23675 130
rect -249 60 -181 71
rect 22970 -6200 23184 -4838
rect 22472 -11894 23031 -11774
rect 22472 -13621 22588 -11894
rect 23211 -12293 23453 -11996
rect 22472 -13741 23603 -13621
rect 22834 -14599 23266 -14562
rect 22834 -14645 22869 -14599
rect 22915 -14645 23027 -14599
rect 23073 -14645 23185 -14599
rect 23231 -14645 23266 -14599
rect 22834 -14682 23266 -14645
rect 23049 -15809 23166 -15424
rect 22648 -15884 23166 -15809
rect 23486 -15823 23603 -13741
rect 22648 -19484 22720 -15884
rect 23049 -16147 23166 -15884
rect 23256 -15860 23603 -15823
rect 23256 -15906 23291 -15860
rect 23337 -15906 23449 -15860
rect 23495 -15906 23603 -15860
rect 23256 -15943 23603 -15906
rect 22825 -16543 22942 -16269
rect 23273 -16543 23390 -16269
rect 22825 -16594 23390 -16543
rect 22825 -16640 22926 -16594
rect 22972 -16640 23084 -16594
rect 23130 -16640 23242 -16594
rect 23288 -16640 23390 -16594
rect 22825 -16691 23390 -16640
rect 22825 -18488 22942 -16691
rect 22648 -19521 22946 -19484
rect 22648 -19567 22707 -19521
rect 22753 -19567 22865 -19521
rect 22911 -19567 22946 -19521
rect 22648 -19604 22946 -19567
rect 23054 -19830 23170 -18443
rect 23273 -18488 23390 -16691
rect 22830 -22882 22946 -21688
rect 23278 -22882 23394 -21688
rect 22717 -22919 22946 -22882
rect 22717 -22965 22751 -22919
rect 22797 -22965 22946 -22919
rect 22717 -23002 22946 -22965
rect 23049 -23165 23179 -22898
rect 23261 -22919 23394 -22882
rect 23261 -22965 23295 -22919
rect 23341 -22965 23394 -22919
rect 23261 -23002 23394 -22965
rect 23001 -25410 23223 -23165
<< via1 >>
rect -241 15989 -238 16128
rect -238 15989 -192 16128
rect -192 15989 -189 16128
rect -241 15868 -189 15989
rect 23587 16065 23639 16070
rect 23587 16019 23592 16065
rect 23592 16019 23638 16065
rect 23638 16019 23639 16065
rect 23587 16018 23639 16019
rect 23587 15800 23639 15852
rect -241 14470 -189 14530
rect -241 14330 -238 14470
rect -238 14330 -192 14470
rect -192 14330 -189 14470
rect -241 14270 -189 14330
rect 23587 14505 23639 14537
rect 23587 14485 23592 14505
rect 23592 14485 23638 14505
rect 23638 14485 23639 14505
rect 23587 14295 23592 14319
rect 23592 14295 23638 14319
rect 23638 14295 23639 14319
rect 23587 14267 23639 14295
rect -241 12670 -189 12730
rect -241 12530 -238 12670
rect -238 12530 -192 12670
rect -192 12530 -189 12670
rect -241 12470 -189 12530
rect 23587 12705 23639 12733
rect 23587 12681 23592 12705
rect 23592 12681 23638 12705
rect 23638 12681 23639 12705
rect 23587 12495 23592 12515
rect 23592 12495 23638 12515
rect 23638 12495 23639 12515
rect 23587 12463 23639 12495
rect -241 10870 -189 10930
rect -241 10730 -238 10870
rect -238 10730 -192 10870
rect -192 10730 -189 10870
rect -241 10670 -189 10730
rect 23587 10905 23639 10937
rect 23587 10885 23592 10905
rect 23592 10885 23638 10905
rect 23638 10885 23639 10905
rect 23587 10695 23592 10719
rect 23592 10695 23638 10719
rect 23638 10695 23639 10719
rect 23587 10667 23639 10695
rect -241 9070 -189 9130
rect -241 8930 -238 9070
rect -238 8930 -192 9070
rect -192 8930 -189 9070
rect -241 8870 -189 8930
rect 23587 9105 23639 9133
rect 23587 9081 23592 9105
rect 23592 9081 23638 9105
rect 23638 9081 23639 9105
rect 23587 8895 23592 8915
rect 23592 8895 23638 8915
rect 23638 8895 23639 8915
rect 23587 8863 23639 8895
rect -241 7270 -189 7330
rect -241 7130 -238 7270
rect -238 7130 -192 7270
rect -192 7130 -189 7270
rect -241 7070 -189 7130
rect 23587 7305 23639 7337
rect 23587 7285 23592 7305
rect 23592 7285 23638 7305
rect 23638 7285 23639 7305
rect 23587 7095 23592 7119
rect 23592 7095 23638 7119
rect 23638 7095 23639 7119
rect 23587 7067 23639 7095
rect -241 5470 -189 5530
rect -241 5330 -238 5470
rect -238 5330 -192 5470
rect -192 5330 -189 5470
rect -241 5270 -189 5330
rect 23587 5505 23639 5533
rect 23587 5481 23592 5505
rect 23592 5481 23638 5505
rect 23638 5481 23639 5505
rect 23587 5295 23592 5315
rect 23592 5295 23638 5315
rect 23638 5295 23639 5315
rect 23587 5263 23639 5295
rect -241 3670 -189 3730
rect -241 3530 -238 3670
rect -238 3530 -192 3670
rect -192 3530 -189 3670
rect -241 3470 -189 3530
rect 23587 3705 23639 3737
rect 23587 3685 23592 3705
rect 23592 3685 23638 3705
rect 23638 3685 23639 3705
rect 23587 3495 23592 3519
rect 23592 3495 23638 3519
rect 23638 3495 23639 3519
rect 23587 3467 23639 3495
rect -241 1870 -189 1930
rect -241 1730 -238 1870
rect -238 1730 -192 1870
rect -192 1730 -189 1870
rect -241 1670 -189 1730
rect 23587 1905 23639 1933
rect 23587 1881 23592 1905
rect 23592 1881 23638 1905
rect 23638 1881 23639 1905
rect 23587 1695 23592 1715
rect 23592 1695 23638 1715
rect 23638 1695 23639 1715
rect 23587 1663 23639 1695
rect 23587 348 23639 400
rect 23587 181 23639 182
rect 23587 135 23592 181
rect 23592 135 23638 181
rect 23638 135 23639 181
rect 23587 130 23639 135
<< metal2 >>
rect -253 16128 -177 16140
rect -253 15868 -241 16128
rect -189 15868 -177 16128
rect -253 14530 -177 15868
rect -253 14270 -241 14530
rect -189 14270 -177 14530
rect -253 12730 -177 14270
rect 23550 16070 23675 16268
rect 23550 16018 23587 16070
rect 23639 16018 23675 16070
rect 23550 15852 23675 16018
rect 23550 15800 23587 15852
rect 23639 15800 23675 15852
rect 23550 14537 23675 15800
rect 23550 14485 23587 14537
rect 23639 14485 23675 14537
rect 23550 14319 23675 14485
rect 23550 14267 23587 14319
rect 23639 14267 23675 14319
rect 23550 14062 23675 14267
rect -253 12470 -241 12730
rect -189 12470 -177 12730
rect -253 10930 -177 12470
rect -253 10670 -241 10930
rect -189 10670 -177 10930
rect -253 9130 -177 10670
rect -253 8870 -241 9130
rect -189 8870 -177 9130
rect -253 7330 -177 8870
rect -253 7070 -241 7330
rect -189 7070 -177 7330
rect -253 5530 -177 7070
rect -253 5270 -241 5530
rect -189 5270 -177 5530
rect -253 3730 -177 5270
rect -253 3470 -241 3730
rect -189 3470 -177 3730
rect -253 1930 -177 3470
rect -253 1670 -241 1930
rect -189 1670 -177 1930
rect -253 42 -177 1670
rect 23550 12733 23675 13839
rect 23550 12681 23587 12733
rect 23639 12681 23675 12733
rect 23550 12515 23675 12681
rect 23550 12463 23587 12515
rect 23639 12463 23675 12515
rect 23550 10937 23675 12463
rect 23550 10885 23587 10937
rect 23639 10885 23675 10937
rect 23550 10719 23675 10885
rect 23550 10667 23587 10719
rect 23639 10667 23675 10719
rect 23550 9133 23675 10667
rect 23550 9081 23587 9133
rect 23639 9081 23675 9133
rect 23550 8915 23675 9081
rect 23550 8863 23587 8915
rect 23639 8863 23675 8915
rect 23550 7337 23675 8863
rect 23550 7285 23587 7337
rect 23639 7285 23675 7337
rect 23550 7119 23675 7285
rect 23550 7067 23587 7119
rect 23639 7067 23675 7119
rect 23550 5533 23675 7067
rect 23550 5481 23587 5533
rect 23639 5481 23675 5533
rect 23550 5315 23675 5481
rect 23550 5263 23587 5315
rect 23639 5263 23675 5315
rect 23550 3737 23675 5263
rect 23550 3685 23587 3737
rect 23639 3685 23675 3737
rect 23550 3519 23675 3685
rect 23550 3467 23587 3519
rect 23639 3467 23675 3519
rect 23550 1933 23675 3467
rect 23550 1881 23587 1933
rect 23639 1881 23675 1933
rect 23550 1715 23675 1881
rect 23550 1663 23587 1715
rect 23639 1663 23675 1715
rect 23550 400 23675 1663
rect 23550 348 23587 400
rect 23639 348 23675 400
rect -357 32 -73 42
rect -357 -24 -347 32
rect -83 -24 -73 32
rect -357 -34 -73 -24
rect 22890 -857 23010 326
rect 22847 -955 23010 -857
rect 23190 -857 23310 326
rect 23550 182 23675 348
rect 23550 130 23587 182
rect 23639 130 23675 182
rect 23550 90 23675 130
rect 23190 -955 23318 -857
rect 22847 -1250 22903 -955
rect 23262 -1250 23318 -955
rect 23049 -25410 23179 -17598
<< via2 >>
rect -347 -24 -83 32
<< metal3 >>
rect -357 32 -73 72
rect -357 -24 -347 32
rect -83 -24 -73 32
rect -357 -68 -73 -24
rect 22329 -2911 23899 -1101
rect 22384 -8791 23899 -6810
rect 22279 -9117 23899 -8902
rect 22279 -9439 23899 -9223
rect 22279 -9760 23899 -9545
rect 22279 -10082 23899 -9867
rect 22279 -10774 23634 -10559
rect 22279 -11096 23634 -10881
rect 22279 -11418 23634 -11203
rect 22279 -11740 23634 -11524
rect 22384 -12288 23899 -11846
rect 22384 -13399 23899 -12944
rect 22426 -17210 23403 -14487
rect 22426 -20898 23403 -17496
rect 22351 -21764 23403 -21047
rect 22351 -23190 23403 -22379
rect 22426 -25051 23051 -23735
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_0
timestamp 1669390400
transform -1 0 600 0 1 6300
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_1
timestamp 1669390400
transform -1 0 600 0 1 900
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_2
timestamp 1669390400
transform -1 0 600 0 1 11700
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_3
timestamp 1669390400
transform -1 0 600 0 1 4500
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_4
timestamp 1669390400
transform -1 0 600 0 1 8100
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_5
timestamp 1669390400
transform -1 0 600 0 1 9900
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_6
timestamp 1669390400
transform -1 0 600 0 1 13500
box -68 -68 668 1868
use 018SRAM_cell1_2x_128x8m81  018SRAM_cell1_2x_128x8m81_7
timestamp 1669390400
transform -1 0 600 0 1 2700
box -68 -68 668 1868
use 018SRAM_cell1_128x8m81  018SRAM_cell1_128x8m81_0
timestamp 1669390400
transform -1 0 600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_128x8m81  018SRAM_cell1_128x8m81_1
timestamp 1669390400
transform -1 0 600 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_0
timestamp 1669390400
transform -1 0 7800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_1
timestamp 1669390400
transform -1 0 9000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_2
timestamp 1669390400
transform -1 0 8400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_3
timestamp 1669390400
transform -1 0 9600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_4
timestamp 1669390400
transform -1 0 10200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_5
timestamp 1669390400
transform -1 0 10800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_6
timestamp 1669390400
transform -1 0 11400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_7
timestamp 1669390400
transform -1 0 6000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_8
timestamp 1669390400
transform -1 0 5400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_9
timestamp 1669390400
transform -1 0 4800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_10
timestamp 1669390400
transform -1 0 4200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_11
timestamp 1669390400
transform -1 0 3000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_12
timestamp 1669390400
transform -1 0 3600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_13
timestamp 1669390400
transform -1 0 2400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_14
timestamp 1669390400
transform -1 0 1800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_15
timestamp 1669390400
transform -1 0 7200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_16
timestamp 1669390400
transform -1 0 7800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_17
timestamp 1669390400
transform -1 0 9000 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_18
timestamp 1669390400
transform -1 0 8400 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_19
timestamp 1669390400
transform -1 0 9600 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_20
timestamp 1669390400
transform -1 0 10200 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_21
timestamp 1669390400
transform -1 0 10800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_22
timestamp 1669390400
transform -1 0 11400 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_23
timestamp 1669390400
transform -1 0 6000 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_24
timestamp 1669390400
transform -1 0 5400 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_25
timestamp 1669390400
transform -1 0 4800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_26
timestamp 1669390400
transform -1 0 4200 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_27
timestamp 1669390400
transform -1 0 3000 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_28
timestamp 1669390400
transform -1 0 3600 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_29
timestamp 1669390400
transform -1 0 2400 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_30
timestamp 1669390400
transform -1 0 1800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_31
timestamp 1669390400
transform -1 0 7200 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_32
timestamp 1669390400
transform -1 0 18000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_33
timestamp 1669390400
transform -1 0 18600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_34
timestamp 1669390400
transform -1 0 19800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_35
timestamp 1669390400
transform -1 0 19200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_36
timestamp 1669390400
transform -1 0 20400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_37
timestamp 1669390400
transform -1 0 21000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_38
timestamp 1669390400
transform -1 0 21600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_39
timestamp 1669390400
transform -1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_40
timestamp 1669390400
transform -1 0 16800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_41
timestamp 1669390400
transform -1 0 16200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_42
timestamp 1669390400
transform -1 0 15600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_43
timestamp 1669390400
transform -1 0 15000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_44
timestamp 1669390400
transform -1 0 13800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_45
timestamp 1669390400
transform -1 0 14400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_46
timestamp 1669390400
transform -1 0 13200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_47
timestamp 1669390400
transform -1 0 12600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_0
timestamp 1669390400
transform 1 0 22800 0 -1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_1
timestamp 1669390400
transform 1 0 22800 0 -1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_2
timestamp 1669390400
transform 1 0 22800 0 -1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_3
timestamp 1669390400
transform 1 0 22800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_4
timestamp 1669390400
transform 1 0 22800 0 -1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_5
timestamp 1669390400
transform 1 0 22800 0 -1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_6
timestamp 1669390400
transform 1 0 22800 0 -1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_7
timestamp 1669390400
transform 1 0 22800 0 -1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_8
timestamp 1669390400
transform 1 0 22800 0 -1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_9
timestamp 1669390400
transform 1 0 22800 0 1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_10
timestamp 1669390400
transform 1 0 22800 0 1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_11
timestamp 1669390400
transform 1 0 22800 0 1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_12
timestamp 1669390400
transform 1 0 22800 0 1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_13
timestamp 1669390400
transform 1 0 22800 0 1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_14
timestamp 1669390400
transform 1 0 22800 0 1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_15
timestamp 1669390400
transform 1 0 22800 0 1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_16
timestamp 1669390400
transform 1 0 22800 0 1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_128x8m81  018SRAM_cell1_dummy_R_128x8m81_17
timestamp 1669390400
transform 1 0 22800 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_0
timestamp 1669390400
transform -1 0 6600 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_1
timestamp 1669390400
transform -1 0 1200 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_2
timestamp 1669390400
transform -1 0 6600 0 -1 16200
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_3
timestamp 1669390400
transform -1 0 17400 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_4
timestamp 1669390400
transform -1 0 12000 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_5
timestamp 1669390400
transform -1 0 12000 0 -1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_128x8m81  018SRAM_strap1_bndry_128x8m81_0
timestamp 1669390400
transform -1 0 1200 0 -1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_128x8m81  018SRAM_strap1_bndry_128x8m81_1
timestamp 1669390400
transform 1 0 22200 0 1 0
box -68 -68 668 968
use M1_NWELL$$44998700_128x8m81_0  M1_NWELL$$44998700_128x8m81_0_0
timestamp 1669390400
transform 1 0 23318 0 1 -22942
box 0 0 1 1
use M1_NWELL$$44998700_128x8m81_0  M1_NWELL$$44998700_128x8m81_0_1
timestamp 1669390400
transform 1 0 22774 0 1 -22942
box 0 0 1 1
use M1_NWELL$$46277676_128x8m81_0  M1_NWELL$$46277676_128x8m81_0_0
timestamp 1669390400
transform 1 0 23050 0 1 -14622
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_0
timestamp 1669390400
transform 1 0 23615 0 -1 1800
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_1
timestamp 1669390400
transform 1 0 23615 0 -1 15960
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_2
timestamp 1669390400
transform 1 0 23615 0 -1 240
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_3
timestamp 1669390400
transform 1 0 23615 0 -1 3600
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_4
timestamp 1669390400
transform 1 0 23615 0 -1 12600
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_5
timestamp 1669390400
transform 1 0 23615 0 -1 9000
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_6
timestamp 1669390400
transform 1 0 23615 0 -1 14400
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_7
timestamp 1669390400
transform 1 0 23615 0 -1 10800
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_8
timestamp 1669390400
transform 1 0 23615 0 -1 7200
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_9
timestamp 1669390400
transform 1 0 23615 0 -1 5400
box 0 0 1 1
use M1_POLY2$$46559276_128x8m81  M1_POLY2$$46559276_128x8m81_0
timestamp 1669390400
transform -1 0 22809 0 1 -19544
box 0 0 1 1
use M1_POLY2$$46559276_128x8m81  M1_POLY2$$46559276_128x8m81_1
timestamp 1669390400
transform 1 0 23393 0 1 -15883
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1669390400
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1669390400
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1669390400
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_3
timestamp 1669390400
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_4
timestamp 1669390400
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_5
timestamp 1669390400
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_6
timestamp 1669390400
transform 1 0 -215 0 1 16059
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_7
timestamp 1669390400
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_8
timestamp 1669390400
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_9
timestamp 1669390400
transform 1 0 -215 0 1 141
box 0 0 1 1
use M1_PSUB$$46274604_128x8m81  M1_PSUB$$46274604_128x8m81_0
timestamp 1669390400
transform 1 0 23107 0 1 -16617
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1669390400
transform 1 0 23613 0 -1 8998
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1669390400
transform 1 0 23613 0 -1 5398
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1669390400
transform 1 0 23613 0 -1 1798
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_3
timestamp 1669390400
transform 1 0 23613 0 -1 10802
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_4
timestamp 1669390400
transform 1 0 23613 0 -1 3602
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_5
timestamp 1669390400
transform 1 0 23613 0 -1 265
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_6
timestamp 1669390400
transform 1 0 23613 0 -1 14402
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_7
timestamp 1669390400
transform 1 0 23613 0 -1 7202
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_8
timestamp 1669390400
transform 1 0 23613 0 -1 15935
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_9
timestamp 1669390400
transform 1 0 23613 0 -1 12598
box 0 0 1 1
use M2_M1$$47117356_128x8m81  M2_M1$$47117356_128x8m81_0
timestamp 1669390400
transform 1 0 23114 0 1 -20269
box -65 -2678 65 2678
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_0
timestamp 1669390400
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_1
timestamp 1669390400
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_2
timestamp 1669390400
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_3
timestamp 1669390400
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_4
timestamp 1669390400
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_5
timestamp 1669390400
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_6
timestamp 1669390400
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_7
timestamp 1669390400
transform 1 0 -215 0 1 15998
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_8
timestamp 1669390400
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M3_M24310590548730_128x8m81  M3_M24310590548730_128x8m81_0
timestamp 1669390400
transform 0 -1 -215 1 0 4
box 0 0 1 1
use new_dummyrow_unit_128x8m81  new_dummyrow_unit_128x8m81_0
timestamp 1669390400
transform 1 0 11938 0 -1 16377
box -6 109 10930 1145
use nmos_5p04310590548754_128x8m81  nmos_5p04310590548754_128x8m81_0
timestamp 1669390400
transform 1 0 22940 0 1 -19403
box -88 -44 432 1744
use nmos_5p04310590548755_128x8m81  nmos_5p04310590548755_128x8m81_0
timestamp 1669390400
transform 1 0 22936 0 1 -16318
box -88 -44 432 320
use pmos_5p04310590548753_128x8m81  pmos_5p04310590548753_128x8m81_0
timestamp 1669390400
transform 1 0 22936 0 1 -15738
box -208 -120 552 822
use pmos_5p04310590548756_128x8m81  pmos_5p04310590548756_128x8m81_0
timestamp 1669390400
transform 1 0 22940 0 -1 -19684
box -208 -120 552 2248
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_0
timestamp 1669390400
transform -1 0 1200 0 1 2680
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_1
timestamp 1669390400
transform -1 0 1200 0 1 4480
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_2
timestamp 1669390400
transform -1 0 1200 0 1 8080
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_3
timestamp 1669390400
transform -1 0 1200 0 1 6280
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_4
timestamp 1669390400
transform -1 0 1200 0 1 9880
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_5
timestamp 1669390400
transform -1 0 1200 0 1 11680
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_6
timestamp 1669390400
transform -1 0 1200 0 1 13480
box -68 -48 668 1888
use strapx2b_bndry_128x8m81  strapx2b_bndry_128x8m81_7
timestamp 1669390400
transform -1 0 1200 0 1 880
box -68 -48 668 1888
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_0
timestamp 1669390400
transform 1 0 22842 0 1 -19052
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_1
timestamp 1669390400
transform 1 0 22837 0 1 -15470
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_2
timestamp 1669390400
transform 1 0 23288 0 1 -22711
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_3
timestamp 1669390400
transform 1 0 22842 0 1 -18447
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_4
timestamp 1669390400
transform 1 0 22846 0 1 -22897
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_5
timestamp 1669390400
transform 1 0 23283 0 1 -17909
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_6
timestamp 1669390400
transform 1 0 23283 0 1 -19052
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_7
timestamp 1669390400
transform 1 0 23283 0 1 -18447
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_8
timestamp 1669390400
transform 1 0 23285 0 1 -15470
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_9
timestamp 1669390400
transform 1 0 23288 0 1 -22897
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_10
timestamp 1669390400
transform 1 0 22846 0 1 -22711
box 0 -1 93 308
use via1_2_x2_128x8m81_0  via1_2_x2_128x8m81_0_11
timestamp 1669390400
transform 1 0 22842 0 1 -17909
box 0 -1 93 308
use via1_2_x2_R90_128x8m81_0  via1_2_x2_R90_128x8m81_0_0
timestamp 1669390400
transform 0 -1 23187 1 0 -14670
box 0 -1 93 308
use via1_2_x2_R270_128x8m81_0  via1_2_x2_R270_128x8m81_0_0
timestamp 1669390400
transform 0 1 22794 -1 0 -12002
box -1 -1 96 308
use ypass_gate_128x8m81_0  ypass_gate_128x8m81_0_0
timestamp 1669390400
transform -1 0 23395 0 1 -13448
box -221 -1 930 12370
<< labels >>
rlabel metal2 s 902 880 902 880 4 VDD
rlabel metal3 s 22866 1818 22866 1818 4 VSS
rlabel metal3 s 534 1818 534 1818 4 VSS
rlabel metal3 s 22866 893 22866 893 4 VDD
rlabel metal3 s 534 893 534 893 4 VDD
rlabel metal3 s 162 15742 162 15742 4 DWL
rlabel metal3 s 22541 -21185 22541 -21185 4 vdd
port 1 nsew
rlabel metal3 s 22541 -14704 22541 -14704 4 vdd
port 1 nsew
rlabel metal3 s 22644 -13162 22644 -13162 4 vss
port 2 nsew
rlabel metal3 s 22541 -12038 22541 -12038 4 vdd
port 1 nsew
rlabel metal3 s 22541 -6717 22541 -6717 4 vss
port 2 nsew
rlabel metal3 s 22541 -1276 22541 -1276 4 vdd
port 1 nsew
rlabel metal1 s 23127 -25252 23127 -25252 4 tblhl
port 3 nsew
rlabel metal1 s 23039 -16606 23039 -16606 4 vss
port 2 nsew
rlabel metal1 s 23037 -3126 23037 -3126 4 pcb
port 4 nsew
rlabel metal1 s 23037 -3126 23037 -3126 4 pcb
port 4 nsew
<< properties >>
string GDS_END 1723352
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1706070
<< end >>
