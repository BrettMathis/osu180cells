magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 2457 52160 12521 52716
rect 2457 48116 3013 52160
rect 11965 48116 12521 52160
rect 2457 47560 12521 48116
<< pwell >>
rect 747 53655 3923 56655
rect 4183 53655 7359 56655
rect 7619 53655 10795 56655
rect 11055 53655 14231 56655
<< mvnmos >>
rect 835 53655 3835 56655
rect 4271 53655 7271 56655
rect 7707 53655 10707 56655
rect 11143 53655 14143 56655
<< mvndiff >>
rect 747 56618 835 56655
rect 747 53692 760 56618
rect 806 53692 835 56618
rect 747 53655 835 53692
rect 3835 56618 3923 56655
rect 3835 53692 3864 56618
rect 3910 53692 3923 56618
rect 3835 53655 3923 53692
rect 4183 56618 4271 56655
rect 4183 53692 4196 56618
rect 4242 53692 4271 56618
rect 4183 53655 4271 53692
rect 7271 56618 7359 56655
rect 7271 53692 7300 56618
rect 7346 53692 7359 56618
rect 7271 53655 7359 53692
rect 7619 56618 7707 56655
rect 7619 53692 7632 56618
rect 7678 53692 7707 56618
rect 7619 53655 7707 53692
rect 10707 56618 10795 56655
rect 10707 53692 10736 56618
rect 10782 53692 10795 56618
rect 10707 53655 10795 53692
rect 11055 56618 11143 56655
rect 11055 53692 11068 56618
rect 11114 53692 11143 56618
rect 11055 53655 11143 53692
rect 14143 56618 14231 56655
rect 14143 53692 14172 56618
rect 14218 53692 14231 56618
rect 14143 53655 14231 53692
<< mvndiffc >>
rect 760 53692 806 56618
rect 3864 53692 3910 56618
rect 4196 53692 4242 56618
rect 7300 53692 7346 56618
rect 7632 53692 7678 56618
rect 10736 53692 10782 56618
rect 11068 53692 11114 56618
rect 14172 53692 14218 56618
<< psubdiff >>
rect 334 57105 14644 57127
rect 334 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57037 14576 57059
rect 402 53273 424 57037
rect 14554 53273 14576 57037
rect 402 53251 14576 53273
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14644 57105
rect 334 53183 14644 53205
rect 246 52611 2236 52633
rect 246 47665 268 52611
rect 2214 47665 2236 52611
rect 246 47643 2236 47665
rect 3094 52029 11884 52051
rect 3094 51983 3142 52029
rect 11836 51983 11884 52029
rect 3094 51900 11884 51983
rect 3094 48376 3116 51900
rect 3162 51875 11816 51900
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51807 11662 51829
rect 3316 51271 3338 51807
rect 11640 51271 11662 51807
rect 3316 51249 11662 51271
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51095 11816 51203
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 50941 11816 51049
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50873 11662 50895
rect 3316 50337 3338 50873
rect 11640 50337 11662 50873
rect 3316 50315 11662 50337
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50161 11816 50269
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50007 11816 50115
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49939 11662 49961
rect 3316 49403 3338 49939
rect 11640 49403 11662 49939
rect 3316 49381 11662 49403
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49227 11816 49335
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49073 11816 49181
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49005 11662 49027
rect 3316 48469 3338 49005
rect 11640 48469 11662 49005
rect 3316 48447 11662 48469
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48376 11816 48401
rect 11862 48376 11884 51900
rect 3094 48293 11884 48376
rect 3094 48247 3142 48293
rect 11836 48247 11884 48293
rect 3094 48225 11884 48247
rect 12742 52611 14732 52633
rect 12742 47665 12764 52611
rect 14710 47665 14732 52611
rect 12742 47643 14732 47665
rect 246 42647 736 42669
rect 246 1201 268 42647
rect 714 1201 736 42647
rect 13001 42647 13991 42669
rect 13001 27201 13023 42647
rect 13969 27201 13991 42647
rect 13001 27179 13991 27201
rect 14242 42647 14732 42669
rect 246 1179 736 1201
rect 14242 1201 14264 42647
rect 14710 1201 14732 42647
rect 14242 1179 14732 1201
<< nsubdiff >>
rect 2540 52611 12438 52633
rect 2540 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52243 12070 52265
rect 2908 48033 2930 52243
rect 12048 48033 12070 52243
rect 2908 48011 12070 48033
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12438 52611
rect 2540 47643 12438 47665
<< psubdiffcont >>
rect 356 53205 402 57105
rect 510 57059 14468 57105
rect 510 53205 14468 53251
rect 14576 53205 14622 57105
rect 268 47665 2214 52611
rect 3142 51983 11836 52029
rect 3116 48376 3162 51900
rect 3270 51234 3316 51844
rect 3424 51829 11554 51875
rect 3424 51203 11554 51249
rect 11662 51234 11708 51844
rect 3330 51049 11648 51095
rect 3270 50300 3316 50910
rect 3424 50895 11554 50941
rect 3424 50269 11554 50315
rect 11662 50300 11708 50910
rect 3330 50115 11648 50161
rect 3270 49366 3316 49976
rect 3424 49961 11554 50007
rect 3424 49335 11554 49381
rect 11662 49366 11708 49976
rect 3330 49181 11648 49227
rect 3270 48432 3316 49042
rect 3424 49027 11554 49073
rect 3424 48401 11554 48447
rect 11662 48432 11708 49042
rect 11816 48376 11862 51900
rect 3142 48247 11836 48293
rect 12764 47665 14710 52611
rect 268 1201 714 42647
rect 13023 27201 13969 42647
rect 14264 1201 14710 42647
<< nsubdiffcont >>
rect 2562 47665 2908 52611
rect 3016 52265 11962 52611
rect 3016 47665 11962 48011
rect 12070 47665 12416 52611
<< polysilicon >>
rect 835 56734 3835 56747
rect 835 56688 888 56734
rect 3782 56688 3835 56734
rect 835 56655 3835 56688
rect 4271 56734 7271 56747
rect 4271 56688 4324 56734
rect 7218 56688 7271 56734
rect 4271 56655 7271 56688
rect 7707 56734 10707 56747
rect 7707 56688 7760 56734
rect 10654 56688 10707 56734
rect 7707 56655 10707 56688
rect 11143 56734 14143 56747
rect 11143 56688 11196 56734
rect 14090 56688 14143 56734
rect 11143 56655 14143 56688
rect 835 53622 3835 53655
rect 835 53576 888 53622
rect 3782 53576 3835 53622
rect 835 53563 3835 53576
rect 4271 53622 7271 53655
rect 4271 53576 4324 53622
rect 7218 53576 7271 53622
rect 4271 53563 7271 53576
rect 7707 53622 10707 53655
rect 7707 53576 7760 53622
rect 10654 53576 10707 53622
rect 7707 53563 10707 53576
rect 11143 53622 14143 53655
rect 11143 53576 11196 53622
rect 14090 53576 14143 53622
rect 11143 53563 14143 53576
<< polycontact >>
rect 888 56688 3782 56734
rect 4324 56688 7218 56734
rect 7760 56688 10654 56734
rect 11196 56688 14090 56734
rect 888 53576 3782 53622
rect 4324 53576 7218 53622
rect 7760 53576 10654 53622
rect 11196 53576 14090 53622
<< mvndiode >>
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51498 11489 51580
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50564 11489 50646
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49630 11489 49712
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48696 11489 48778
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
<< mvndiodec >>
rect 3502 51580 11476 51626
rect 3502 51452 11476 51498
rect 3502 50646 11476 50692
rect 3502 50518 11476 50564
rect 3502 49712 11476 49758
rect 3502 49584 11476 49630
rect 3502 48778 11476 48824
rect 3502 48650 11476 48696
<< metal1 >>
rect 309 57499 2113 57511
rect 309 57447 321 57499
rect 373 57447 429 57499
rect 481 57447 537 57499
rect 589 57447 645 57499
rect 697 57447 753 57499
rect 805 57447 861 57499
rect 913 57447 969 57499
rect 1021 57447 1077 57499
rect 1129 57447 1185 57499
rect 1237 57447 1293 57499
rect 1345 57447 1401 57499
rect 1453 57447 1509 57499
rect 1561 57447 1617 57499
rect 1669 57447 1725 57499
rect 1777 57447 1833 57499
rect 1885 57447 1941 57499
rect 1993 57447 2049 57499
rect 2101 57447 2113 57499
rect 309 57435 2113 57447
rect 2864 57499 4668 57511
rect 2864 57447 2876 57499
rect 2928 57447 2984 57499
rect 3036 57447 3092 57499
rect 3144 57447 3200 57499
rect 3252 57447 3308 57499
rect 3360 57447 3416 57499
rect 3468 57447 3524 57499
rect 3576 57447 3632 57499
rect 3684 57447 3740 57499
rect 3792 57447 3848 57499
rect 3900 57447 3956 57499
rect 4008 57447 4064 57499
rect 4116 57447 4172 57499
rect 4224 57447 4280 57499
rect 4332 57447 4388 57499
rect 4440 57447 4496 57499
rect 4548 57447 4604 57499
rect 4656 57447 4668 57499
rect 2864 57435 4668 57447
rect 5234 57499 7038 57511
rect 5234 57447 5246 57499
rect 5298 57447 5354 57499
rect 5406 57447 5462 57499
rect 5514 57447 5570 57499
rect 5622 57447 5678 57499
rect 5730 57447 5786 57499
rect 5838 57447 5894 57499
rect 5946 57447 6002 57499
rect 6054 57447 6110 57499
rect 6162 57447 6218 57499
rect 6270 57447 6326 57499
rect 6378 57447 6434 57499
rect 6486 57447 6542 57499
rect 6594 57447 6650 57499
rect 6702 57447 6758 57499
rect 6810 57447 6866 57499
rect 6918 57447 6974 57499
rect 7026 57447 7038 57499
rect 5234 57435 7038 57447
rect 7940 57499 9744 57511
rect 7940 57447 7952 57499
rect 8004 57447 8060 57499
rect 8112 57447 8168 57499
rect 8220 57447 8276 57499
rect 8328 57447 8384 57499
rect 8436 57447 8492 57499
rect 8544 57447 8600 57499
rect 8652 57447 8708 57499
rect 8760 57447 8816 57499
rect 8868 57447 8924 57499
rect 8976 57447 9032 57499
rect 9084 57447 9140 57499
rect 9192 57447 9248 57499
rect 9300 57447 9356 57499
rect 9408 57447 9464 57499
rect 9516 57447 9572 57499
rect 9624 57447 9680 57499
rect 9732 57447 9744 57499
rect 7940 57435 9744 57447
rect 10310 57499 12114 57511
rect 10310 57447 10322 57499
rect 10374 57447 10430 57499
rect 10482 57447 10538 57499
rect 10590 57447 10646 57499
rect 10698 57447 10754 57499
rect 10806 57447 10862 57499
rect 10914 57447 10970 57499
rect 11022 57447 11078 57499
rect 11130 57447 11186 57499
rect 11238 57447 11294 57499
rect 11346 57447 11402 57499
rect 11454 57447 11510 57499
rect 11562 57447 11618 57499
rect 11670 57447 11726 57499
rect 11778 57447 11834 57499
rect 11886 57447 11942 57499
rect 11994 57447 12050 57499
rect 12102 57447 12114 57499
rect 10310 57435 12114 57447
rect 12865 57499 14669 57511
rect 12865 57447 12877 57499
rect 12929 57447 12985 57499
rect 13037 57447 13093 57499
rect 13145 57447 13201 57499
rect 13253 57447 13309 57499
rect 13361 57447 13417 57499
rect 13469 57447 13525 57499
rect 13577 57447 13633 57499
rect 13685 57447 13741 57499
rect 13793 57447 13849 57499
rect 13901 57447 13957 57499
rect 14009 57447 14065 57499
rect 14117 57447 14173 57499
rect 14225 57447 14281 57499
rect 14333 57447 14389 57499
rect 14441 57447 14497 57499
rect 14549 57447 14605 57499
rect 14657 57447 14669 57499
rect 12865 57435 14669 57447
rect 10 57259 86 57271
rect 10 57207 22 57259
rect 74 57207 86 57259
rect 10 57151 86 57207
rect 10 57099 22 57151
rect 74 57099 86 57151
rect 14892 57259 14968 57271
rect 14892 57207 14904 57259
rect 14956 57207 14968 57259
rect 14892 57151 14968 57207
rect 10 57043 86 57099
rect 10 56991 22 57043
rect 74 56991 86 57043
rect 10 56935 86 56991
rect 10 56883 22 56935
rect 74 56883 86 56935
rect 10 56827 86 56883
rect 10 56775 22 56827
rect 74 56775 86 56827
rect 10 56719 86 56775
rect 10 56667 22 56719
rect 74 56667 86 56719
rect 10 56611 86 56667
rect 10 56559 22 56611
rect 74 56559 86 56611
rect 10 56503 86 56559
rect 10 56451 22 56503
rect 74 56451 86 56503
rect 10 56395 86 56451
rect 10 56343 22 56395
rect 74 56343 86 56395
rect 10 56287 86 56343
rect 10 56235 22 56287
rect 74 56235 86 56287
rect 10 56179 86 56235
rect 10 56127 22 56179
rect 74 56127 86 56179
rect 10 56071 86 56127
rect 10 56019 22 56071
rect 74 56019 86 56071
rect 10 56007 86 56019
rect 345 57105 14633 57116
rect 10 54174 86 54186
rect 10 54122 22 54174
rect 74 54122 86 54174
rect 10 54066 86 54122
rect 10 54014 22 54066
rect 74 54014 86 54066
rect 10 53958 86 54014
rect 10 53906 22 53958
rect 74 53906 86 53958
rect 10 53850 86 53906
rect 10 53798 22 53850
rect 74 53798 86 53850
rect 10 53742 86 53798
rect 10 53690 22 53742
rect 74 53690 86 53742
rect 10 53634 86 53690
rect 10 53582 22 53634
rect 74 53582 86 53634
rect 10 53526 86 53582
rect 10 53474 22 53526
rect 74 53474 86 53526
rect 10 53418 86 53474
rect 10 53366 22 53418
rect 74 53366 86 53418
rect 10 53310 86 53366
rect 10 53258 22 53310
rect 74 53258 86 53310
rect 10 53202 86 53258
rect 10 53150 22 53202
rect 74 53150 86 53202
rect 345 53205 356 57105
rect 402 57104 510 57105
rect 14468 57104 14576 57105
rect 427 57052 483 57104
rect 535 57052 591 57059
rect 643 57052 699 57059
rect 751 57052 807 57059
rect 859 57052 915 57059
rect 967 57052 1023 57059
rect 1075 57052 1131 57059
rect 1183 57052 1239 57059
rect 1291 57052 1347 57059
rect 1399 57052 1455 57059
rect 1507 57052 1563 57059
rect 1615 57052 1671 57059
rect 1723 57052 1779 57059
rect 1831 57052 1887 57059
rect 1939 57052 1995 57059
rect 2047 57052 2768 57059
rect 2820 57052 2876 57059
rect 2928 57052 2984 57059
rect 3036 57052 3092 57059
rect 3144 57052 3200 57059
rect 3252 57052 3308 57059
rect 3360 57052 3416 57059
rect 3468 57052 3524 57059
rect 3576 57052 3632 57059
rect 3684 57052 3740 57059
rect 3792 57052 3848 57059
rect 3900 57052 3956 57059
rect 4008 57052 4064 57059
rect 4116 57052 4172 57059
rect 4224 57052 4280 57059
rect 4332 57052 4388 57059
rect 4440 57052 4496 57059
rect 4548 57052 4604 57059
rect 4656 57052 4712 57059
rect 4764 57052 5138 57059
rect 5190 57052 5246 57059
rect 5298 57052 5354 57059
rect 5406 57052 5462 57059
rect 5514 57052 5570 57059
rect 5622 57052 5678 57059
rect 5730 57052 5786 57059
rect 5838 57052 5894 57059
rect 5946 57052 6002 57059
rect 6054 57052 6110 57059
rect 6162 57052 6218 57059
rect 6270 57052 6326 57059
rect 6378 57052 6434 57059
rect 6486 57052 6542 57059
rect 6594 57052 6650 57059
rect 6702 57052 6758 57059
rect 6810 57052 6866 57059
rect 6918 57052 6974 57059
rect 7026 57052 7082 57059
rect 7134 57052 7844 57059
rect 7896 57052 7952 57059
rect 8004 57052 8060 57059
rect 8112 57052 8168 57059
rect 8220 57052 8276 57059
rect 8328 57052 8384 57059
rect 8436 57052 8492 57059
rect 8544 57052 8600 57059
rect 8652 57052 8708 57059
rect 8760 57052 8816 57059
rect 8868 57052 8924 57059
rect 8976 57052 9032 57059
rect 9084 57052 9140 57059
rect 9192 57052 9248 57059
rect 9300 57052 9356 57059
rect 9408 57052 9464 57059
rect 9516 57052 9572 57059
rect 9624 57052 9680 57059
rect 9732 57052 9788 57059
rect 9840 57052 10214 57059
rect 10266 57052 10322 57059
rect 10374 57052 10430 57059
rect 10482 57052 10538 57059
rect 10590 57052 10646 57059
rect 10698 57052 10754 57059
rect 10806 57052 10862 57059
rect 10914 57052 10970 57059
rect 11022 57052 11078 57059
rect 11130 57052 11186 57059
rect 11238 57052 11294 57059
rect 11346 57052 11402 57059
rect 11454 57052 11510 57059
rect 11562 57052 11618 57059
rect 11670 57052 11726 57059
rect 11778 57052 11834 57059
rect 11886 57052 11942 57059
rect 11994 57052 12050 57059
rect 12102 57052 12158 57059
rect 12210 57052 12931 57059
rect 12983 57052 13039 57059
rect 13091 57052 13147 57059
rect 13199 57052 13255 57059
rect 13307 57052 13363 57059
rect 13415 57052 13471 57059
rect 13523 57052 13579 57059
rect 13631 57052 13687 57059
rect 13739 57052 13795 57059
rect 13847 57052 13903 57059
rect 13955 57052 14011 57059
rect 14063 57052 14119 57059
rect 14171 57052 14227 57059
rect 14279 57052 14335 57059
rect 14387 57052 14443 57059
rect 14495 57052 14551 57104
rect 402 57048 14576 57052
rect 402 57040 2059 57048
rect 2756 57040 4776 57048
rect 5126 57040 7146 57048
rect 7832 57040 9852 57048
rect 10202 57040 12222 57048
rect 12919 57040 14576 57048
rect 402 56655 413 57040
rect 2489 56745 2673 56753
rect 12305 56745 12489 56753
rect 877 56741 3793 56745
rect 877 56734 2501 56741
rect 2553 56734 2609 56741
rect 2661 56734 3793 56741
rect 877 56688 888 56734
rect 3782 56688 3793 56734
rect 877 56677 3793 56688
rect 402 56643 817 56655
rect 421 56591 493 56643
rect 545 56591 617 56643
rect 669 56591 741 56643
rect 793 56618 817 56643
rect 402 56519 760 56591
rect 421 56467 493 56519
rect 545 56467 617 56519
rect 669 56467 741 56519
rect 402 56395 760 56467
rect 421 56343 493 56395
rect 545 56343 617 56395
rect 669 56343 741 56395
rect 402 56271 760 56343
rect 421 56219 493 56271
rect 545 56219 617 56271
rect 669 56219 741 56271
rect 402 56147 760 56219
rect 421 56095 493 56147
rect 545 56095 617 56147
rect 669 56095 741 56147
rect 402 56023 760 56095
rect 421 55971 493 56023
rect 545 55971 617 56023
rect 669 55971 741 56023
rect 402 55899 760 55971
rect 421 55847 493 55899
rect 545 55847 617 55899
rect 669 55847 741 55899
rect 402 55775 760 55847
rect 421 55723 493 55775
rect 545 55723 617 55775
rect 669 55723 741 55775
rect 402 55651 760 55723
rect 421 55599 493 55651
rect 545 55599 617 55651
rect 669 55599 741 55651
rect 402 55527 760 55599
rect 421 55475 493 55527
rect 545 55475 617 55527
rect 669 55475 741 55527
rect 402 55403 760 55475
rect 421 55351 493 55403
rect 545 55351 617 55403
rect 669 55351 741 55403
rect 402 55279 760 55351
rect 421 55227 493 55279
rect 545 55227 617 55279
rect 669 55227 741 55279
rect 402 55155 760 55227
rect 421 55103 493 55155
rect 545 55103 617 55155
rect 669 55103 741 55155
rect 402 55031 760 55103
rect 421 54979 493 55031
rect 545 54979 617 55031
rect 669 54979 741 55031
rect 402 54907 760 54979
rect 421 54855 493 54907
rect 545 54855 617 54907
rect 669 54855 741 54907
rect 402 54783 760 54855
rect 421 54731 493 54783
rect 545 54731 617 54783
rect 669 54731 741 54783
rect 402 54659 760 54731
rect 421 54607 493 54659
rect 545 54607 617 54659
rect 669 54607 741 54659
rect 402 54535 760 54607
rect 421 54483 493 54535
rect 545 54483 617 54535
rect 669 54483 741 54535
rect 402 54411 760 54483
rect 421 54359 493 54411
rect 545 54359 617 54411
rect 669 54359 741 54411
rect 402 54287 760 54359
rect 421 54235 493 54287
rect 545 54235 617 54287
rect 669 54235 741 54287
rect 402 54163 760 54235
rect 421 54111 493 54163
rect 545 54111 617 54163
rect 669 54111 741 54163
rect 402 54039 760 54111
rect 421 53987 493 54039
rect 545 53987 617 54039
rect 669 53987 741 54039
rect 402 53915 760 53987
rect 421 53863 493 53915
rect 545 53863 617 53915
rect 669 53863 741 53915
rect 402 53791 760 53863
rect 421 53739 493 53791
rect 545 53739 617 53791
rect 669 53739 741 53791
rect 402 53692 760 53739
rect 806 53692 817 56618
rect 402 53667 817 53692
rect 421 53615 493 53667
rect 545 53615 617 53667
rect 669 53615 741 53667
rect 793 53615 817 53667
rect 402 53543 817 53615
rect 877 53633 1877 56677
rect 2793 53633 3793 56677
rect 4313 56734 7229 56745
rect 4313 56688 4324 56734
rect 7218 56688 7229 56734
rect 877 53622 3793 53633
rect 877 53576 888 53622
rect 3782 53576 3793 53622
rect 877 53569 2501 53576
rect 2553 53569 2609 53576
rect 2661 53569 3793 53576
rect 877 53565 3793 53569
rect 3853 56643 4253 56655
rect 3853 56618 3903 56643
rect 3853 53692 3864 56618
rect 3955 56591 4027 56643
rect 4079 56591 4151 56643
rect 4203 56618 4253 56643
rect 3910 56519 4196 56591
rect 3955 56467 4027 56519
rect 4079 56467 4151 56519
rect 3910 56395 4196 56467
rect 3955 56343 4027 56395
rect 4079 56343 4151 56395
rect 3910 56271 4196 56343
rect 3955 56219 4027 56271
rect 4079 56219 4151 56271
rect 3910 56147 4196 56219
rect 3955 56095 4027 56147
rect 4079 56095 4151 56147
rect 3910 56023 4196 56095
rect 3955 55971 4027 56023
rect 4079 55971 4151 56023
rect 3910 55899 4196 55971
rect 3955 55847 4027 55899
rect 4079 55847 4151 55899
rect 3910 55775 4196 55847
rect 3955 55723 4027 55775
rect 4079 55723 4151 55775
rect 3910 55651 4196 55723
rect 3955 55599 4027 55651
rect 4079 55599 4151 55651
rect 3910 55527 4196 55599
rect 3955 55475 4027 55527
rect 4079 55475 4151 55527
rect 3910 55403 4196 55475
rect 3955 55351 4027 55403
rect 4079 55351 4151 55403
rect 3910 55279 4196 55351
rect 3955 55227 4027 55279
rect 4079 55227 4151 55279
rect 3910 55155 4196 55227
rect 3955 55103 4027 55155
rect 4079 55103 4151 55155
rect 3910 55031 4196 55103
rect 3955 54979 4027 55031
rect 4079 54979 4151 55031
rect 3910 54907 4196 54979
rect 3955 54855 4027 54907
rect 4079 54855 4151 54907
rect 3910 54783 4196 54855
rect 3955 54731 4027 54783
rect 4079 54731 4151 54783
rect 3910 54659 4196 54731
rect 3955 54607 4027 54659
rect 4079 54607 4151 54659
rect 3910 54535 4196 54607
rect 3955 54483 4027 54535
rect 4079 54483 4151 54535
rect 3910 54411 4196 54483
rect 3955 54359 4027 54411
rect 4079 54359 4151 54411
rect 3910 54287 4196 54359
rect 3955 54235 4027 54287
rect 4079 54235 4151 54287
rect 3910 54163 4196 54235
rect 3955 54111 4027 54163
rect 4079 54111 4151 54163
rect 3910 54039 4196 54111
rect 3955 53987 4027 54039
rect 4079 53987 4151 54039
rect 3910 53915 4196 53987
rect 3955 53863 4027 53915
rect 4079 53863 4151 53915
rect 3910 53791 4196 53863
rect 3955 53739 4027 53791
rect 4079 53739 4151 53791
rect 3910 53692 4196 53739
rect 4242 53692 4253 56618
rect 3853 53667 4253 53692
rect 3853 53615 3903 53667
rect 3955 53615 4027 53667
rect 4079 53615 4151 53667
rect 4203 53615 4253 53667
rect 2489 53557 2673 53565
rect 421 53491 493 53543
rect 545 53491 617 53543
rect 669 53491 741 53543
rect 793 53505 817 53543
rect 3853 53543 4253 53615
rect 4313 56641 4871 56688
rect 4923 56641 4979 56688
rect 5031 56677 7229 56688
rect 5031 56641 5313 56677
rect 4313 56585 5313 56641
rect 4313 56533 4871 56585
rect 4923 56533 4979 56585
rect 5031 56533 5313 56585
rect 4313 56477 5313 56533
rect 4313 56425 4871 56477
rect 4923 56425 4979 56477
rect 5031 56425 5313 56477
rect 4313 56369 5313 56425
rect 4313 56317 4871 56369
rect 4923 56317 4979 56369
rect 5031 56317 5313 56369
rect 4313 56261 5313 56317
rect 4313 56209 4871 56261
rect 4923 56209 4979 56261
rect 5031 56209 5313 56261
rect 4313 56153 5313 56209
rect 4313 56101 4871 56153
rect 4923 56101 4979 56153
rect 5031 56101 5313 56153
rect 4313 56045 5313 56101
rect 4313 55993 4871 56045
rect 4923 55993 4979 56045
rect 5031 55993 5313 56045
rect 4313 55937 5313 55993
rect 4313 55885 4871 55937
rect 4923 55885 4979 55937
rect 5031 55885 5313 55937
rect 4313 55829 5313 55885
rect 4313 55777 4871 55829
rect 4923 55777 4979 55829
rect 5031 55777 5313 55829
rect 4313 55721 5313 55777
rect 4313 55669 4871 55721
rect 4923 55669 4979 55721
rect 5031 55669 5313 55721
rect 4313 55613 5313 55669
rect 4313 55561 4871 55613
rect 4923 55561 4979 55613
rect 5031 55561 5313 55613
rect 4313 55505 5313 55561
rect 4313 55453 4871 55505
rect 4923 55453 4979 55505
rect 5031 55453 5313 55505
rect 4313 55397 5313 55453
rect 4313 55345 4871 55397
rect 4923 55345 4979 55397
rect 5031 55345 5313 55397
rect 4313 55289 5313 55345
rect 4313 55237 4871 55289
rect 4923 55237 4979 55289
rect 5031 55237 5313 55289
rect 4313 55181 5313 55237
rect 4313 55129 4871 55181
rect 4923 55129 4979 55181
rect 5031 55129 5313 55181
rect 4313 55073 5313 55129
rect 4313 55021 4871 55073
rect 4923 55021 4979 55073
rect 5031 55021 5313 55073
rect 4313 54965 5313 55021
rect 4313 54913 4871 54965
rect 4923 54913 4979 54965
rect 5031 54913 5313 54965
rect 4313 54857 5313 54913
rect 4313 54805 4871 54857
rect 4923 54805 4979 54857
rect 5031 54805 5313 54857
rect 4313 54749 5313 54805
rect 4313 54697 4871 54749
rect 4923 54697 4979 54749
rect 5031 54697 5313 54749
rect 4313 54641 5313 54697
rect 4313 54589 4871 54641
rect 4923 54589 4979 54641
rect 5031 54589 5313 54641
rect 4313 54533 5313 54589
rect 4313 54481 4871 54533
rect 4923 54481 4979 54533
rect 5031 54481 5313 54533
rect 4313 54425 5313 54481
rect 4313 54373 4871 54425
rect 4923 54373 4979 54425
rect 5031 54373 5313 54425
rect 4313 54317 5313 54373
rect 4313 54265 4871 54317
rect 4923 54265 4979 54317
rect 5031 54265 5313 54317
rect 4313 54209 5313 54265
rect 4313 54157 4871 54209
rect 4923 54157 4979 54209
rect 5031 54157 5313 54209
rect 4313 54101 5313 54157
rect 4313 54049 4871 54101
rect 4923 54049 4979 54101
rect 5031 54049 5313 54101
rect 4313 53993 5313 54049
rect 4313 53941 4871 53993
rect 4923 53941 4979 53993
rect 5031 53941 5313 53993
rect 4313 53885 5313 53941
rect 4313 53833 4871 53885
rect 4923 53833 4979 53885
rect 5031 53833 5313 53885
rect 4313 53777 5313 53833
rect 4313 53725 4871 53777
rect 4923 53725 4979 53777
rect 5031 53725 5313 53777
rect 4313 53669 5313 53725
rect 4313 53622 4871 53669
rect 4923 53622 4979 53669
rect 5031 53633 5313 53669
rect 6229 53633 7229 56677
rect 7749 56734 10665 56745
rect 7749 56688 7760 56734
rect 10654 56688 10665 56734
rect 7749 56677 9947 56688
rect 5031 53622 7229 53633
rect 4313 53576 4324 53622
rect 7218 53576 7229 53622
rect 4313 53565 7229 53576
rect 7289 56618 7689 56655
rect 7289 53692 7300 56618
rect 7346 53692 7632 56618
rect 7678 53692 7689 56618
rect 3853 53505 3903 53543
rect 793 53491 3903 53505
rect 3955 53491 4027 53543
rect 4079 53491 4151 53543
rect 4203 53505 4253 53543
rect 7289 53505 7689 53692
rect 7749 53633 8749 56677
rect 9665 56641 9947 56677
rect 9999 56641 10055 56688
rect 10107 56641 10665 56688
rect 11185 56741 14101 56745
rect 11185 56734 12317 56741
rect 12369 56734 12425 56741
rect 12477 56734 14101 56741
rect 11185 56688 11196 56734
rect 14090 56688 14101 56734
rect 11185 56677 14101 56688
rect 9665 56585 10665 56641
rect 9665 56533 9947 56585
rect 9999 56533 10055 56585
rect 10107 56533 10665 56585
rect 9665 56477 10665 56533
rect 9665 56425 9947 56477
rect 9999 56425 10055 56477
rect 10107 56425 10665 56477
rect 9665 56369 10665 56425
rect 9665 56317 9947 56369
rect 9999 56317 10055 56369
rect 10107 56317 10665 56369
rect 9665 56261 10665 56317
rect 9665 56209 9947 56261
rect 9999 56209 10055 56261
rect 10107 56209 10665 56261
rect 9665 56153 10665 56209
rect 9665 56101 9947 56153
rect 9999 56101 10055 56153
rect 10107 56101 10665 56153
rect 9665 56045 10665 56101
rect 9665 55993 9947 56045
rect 9999 55993 10055 56045
rect 10107 55993 10665 56045
rect 9665 55937 10665 55993
rect 9665 55885 9947 55937
rect 9999 55885 10055 55937
rect 10107 55885 10665 55937
rect 9665 55829 10665 55885
rect 9665 55777 9947 55829
rect 9999 55777 10055 55829
rect 10107 55777 10665 55829
rect 9665 55721 10665 55777
rect 9665 55669 9947 55721
rect 9999 55669 10055 55721
rect 10107 55669 10665 55721
rect 9665 55613 10665 55669
rect 9665 55561 9947 55613
rect 9999 55561 10055 55613
rect 10107 55561 10665 55613
rect 9665 55505 10665 55561
rect 9665 55453 9947 55505
rect 9999 55453 10055 55505
rect 10107 55453 10665 55505
rect 9665 55397 10665 55453
rect 9665 55345 9947 55397
rect 9999 55345 10055 55397
rect 10107 55345 10665 55397
rect 9665 55289 10665 55345
rect 9665 55237 9947 55289
rect 9999 55237 10055 55289
rect 10107 55237 10665 55289
rect 9665 55181 10665 55237
rect 9665 55129 9947 55181
rect 9999 55129 10055 55181
rect 10107 55129 10665 55181
rect 9665 55073 10665 55129
rect 9665 55021 9947 55073
rect 9999 55021 10055 55073
rect 10107 55021 10665 55073
rect 9665 54965 10665 55021
rect 9665 54913 9947 54965
rect 9999 54913 10055 54965
rect 10107 54913 10665 54965
rect 9665 54857 10665 54913
rect 9665 54805 9947 54857
rect 9999 54805 10055 54857
rect 10107 54805 10665 54857
rect 9665 54749 10665 54805
rect 9665 54697 9947 54749
rect 9999 54697 10055 54749
rect 10107 54697 10665 54749
rect 9665 54641 10665 54697
rect 9665 54589 9947 54641
rect 9999 54589 10055 54641
rect 10107 54589 10665 54641
rect 9665 54533 10665 54589
rect 9665 54481 9947 54533
rect 9999 54481 10055 54533
rect 10107 54481 10665 54533
rect 9665 54425 10665 54481
rect 9665 54373 9947 54425
rect 9999 54373 10055 54425
rect 10107 54373 10665 54425
rect 9665 54317 10665 54373
rect 9665 54265 9947 54317
rect 9999 54265 10055 54317
rect 10107 54265 10665 54317
rect 9665 54209 10665 54265
rect 9665 54157 9947 54209
rect 9999 54157 10055 54209
rect 10107 54157 10665 54209
rect 9665 54101 10665 54157
rect 9665 54049 9947 54101
rect 9999 54049 10055 54101
rect 10107 54049 10665 54101
rect 9665 53993 10665 54049
rect 9665 53941 9947 53993
rect 9999 53941 10055 53993
rect 10107 53941 10665 53993
rect 9665 53885 10665 53941
rect 9665 53833 9947 53885
rect 9999 53833 10055 53885
rect 10107 53833 10665 53885
rect 9665 53777 10665 53833
rect 9665 53725 9947 53777
rect 9999 53725 10055 53777
rect 10107 53725 10665 53777
rect 9665 53669 10665 53725
rect 9665 53633 9947 53669
rect 7749 53622 9947 53633
rect 9999 53622 10055 53669
rect 10107 53622 10665 53669
rect 7749 53576 7760 53622
rect 10654 53576 10665 53622
rect 7749 53565 10665 53576
rect 10725 56643 11125 56655
rect 10725 56618 10775 56643
rect 10725 53692 10736 56618
rect 10827 56591 10899 56643
rect 10951 56591 11023 56643
rect 11075 56618 11125 56643
rect 10782 56519 11068 56591
rect 10827 56467 10899 56519
rect 10951 56467 11023 56519
rect 10782 56395 11068 56467
rect 10827 56343 10899 56395
rect 10951 56343 11023 56395
rect 10782 56271 11068 56343
rect 10827 56219 10899 56271
rect 10951 56219 11023 56271
rect 10782 56147 11068 56219
rect 10827 56095 10899 56147
rect 10951 56095 11023 56147
rect 10782 56023 11068 56095
rect 10827 55971 10899 56023
rect 10951 55971 11023 56023
rect 10782 55899 11068 55971
rect 10827 55847 10899 55899
rect 10951 55847 11023 55899
rect 10782 55775 11068 55847
rect 10827 55723 10899 55775
rect 10951 55723 11023 55775
rect 10782 55651 11068 55723
rect 10827 55599 10899 55651
rect 10951 55599 11023 55651
rect 10782 55527 11068 55599
rect 10827 55475 10899 55527
rect 10951 55475 11023 55527
rect 10782 55403 11068 55475
rect 10827 55351 10899 55403
rect 10951 55351 11023 55403
rect 10782 55279 11068 55351
rect 10827 55227 10899 55279
rect 10951 55227 11023 55279
rect 10782 55155 11068 55227
rect 10827 55103 10899 55155
rect 10951 55103 11023 55155
rect 10782 55031 11068 55103
rect 10827 54979 10899 55031
rect 10951 54979 11023 55031
rect 10782 54907 11068 54979
rect 10827 54855 10899 54907
rect 10951 54855 11023 54907
rect 10782 54783 11068 54855
rect 10827 54731 10899 54783
rect 10951 54731 11023 54783
rect 10782 54659 11068 54731
rect 10827 54607 10899 54659
rect 10951 54607 11023 54659
rect 10782 54535 11068 54607
rect 10827 54483 10899 54535
rect 10951 54483 11023 54535
rect 10782 54411 11068 54483
rect 10827 54359 10899 54411
rect 10951 54359 11023 54411
rect 10782 54287 11068 54359
rect 10827 54235 10899 54287
rect 10951 54235 11023 54287
rect 10782 54163 11068 54235
rect 10827 54111 10899 54163
rect 10951 54111 11023 54163
rect 10782 54039 11068 54111
rect 10827 53987 10899 54039
rect 10951 53987 11023 54039
rect 10782 53915 11068 53987
rect 10827 53863 10899 53915
rect 10951 53863 11023 53915
rect 10782 53791 11068 53863
rect 10827 53739 10899 53791
rect 10951 53739 11023 53791
rect 10782 53692 11068 53739
rect 11114 53692 11125 56618
rect 10725 53667 11125 53692
rect 10725 53615 10775 53667
rect 10827 53615 10899 53667
rect 10951 53615 11023 53667
rect 11075 53615 11125 53667
rect 10725 53543 11125 53615
rect 11185 53633 12185 56677
rect 13101 53633 14101 56677
rect 14565 56655 14576 57040
rect 11185 53622 14101 53633
rect 11185 53576 11196 53622
rect 14090 53576 14101 53622
rect 11185 53569 12317 53576
rect 12369 53569 12425 53576
rect 12477 53569 14101 53576
rect 11185 53565 14101 53569
rect 14161 56643 14576 56655
rect 14161 56618 14185 56643
rect 14161 53692 14172 56618
rect 14237 56591 14309 56643
rect 14361 56591 14433 56643
rect 14485 56591 14557 56643
rect 14218 56519 14576 56591
rect 14237 56467 14309 56519
rect 14361 56467 14433 56519
rect 14485 56467 14557 56519
rect 14218 56395 14576 56467
rect 14237 56343 14309 56395
rect 14361 56343 14433 56395
rect 14485 56343 14557 56395
rect 14218 56271 14576 56343
rect 14237 56219 14309 56271
rect 14361 56219 14433 56271
rect 14485 56219 14557 56271
rect 14218 56147 14576 56219
rect 14237 56095 14309 56147
rect 14361 56095 14433 56147
rect 14485 56095 14557 56147
rect 14218 56023 14576 56095
rect 14237 55971 14309 56023
rect 14361 55971 14433 56023
rect 14485 55971 14557 56023
rect 14218 55899 14576 55971
rect 14237 55847 14309 55899
rect 14361 55847 14433 55899
rect 14485 55847 14557 55899
rect 14218 55775 14576 55847
rect 14237 55723 14309 55775
rect 14361 55723 14433 55775
rect 14485 55723 14557 55775
rect 14218 55651 14576 55723
rect 14237 55599 14309 55651
rect 14361 55599 14433 55651
rect 14485 55599 14557 55651
rect 14218 55527 14576 55599
rect 14237 55475 14309 55527
rect 14361 55475 14433 55527
rect 14485 55475 14557 55527
rect 14218 55403 14576 55475
rect 14237 55351 14309 55403
rect 14361 55351 14433 55403
rect 14485 55351 14557 55403
rect 14218 55279 14576 55351
rect 14237 55227 14309 55279
rect 14361 55227 14433 55279
rect 14485 55227 14557 55279
rect 14218 55155 14576 55227
rect 14237 55103 14309 55155
rect 14361 55103 14433 55155
rect 14485 55103 14557 55155
rect 14218 55031 14576 55103
rect 14237 54979 14309 55031
rect 14361 54979 14433 55031
rect 14485 54979 14557 55031
rect 14218 54907 14576 54979
rect 14237 54855 14309 54907
rect 14361 54855 14433 54907
rect 14485 54855 14557 54907
rect 14218 54783 14576 54855
rect 14237 54731 14309 54783
rect 14361 54731 14433 54783
rect 14485 54731 14557 54783
rect 14218 54659 14576 54731
rect 14237 54607 14309 54659
rect 14361 54607 14433 54659
rect 14485 54607 14557 54659
rect 14218 54535 14576 54607
rect 14237 54483 14309 54535
rect 14361 54483 14433 54535
rect 14485 54483 14557 54535
rect 14218 54411 14576 54483
rect 14237 54359 14309 54411
rect 14361 54359 14433 54411
rect 14485 54359 14557 54411
rect 14218 54287 14576 54359
rect 14237 54235 14309 54287
rect 14361 54235 14433 54287
rect 14485 54235 14557 54287
rect 14218 54163 14576 54235
rect 14237 54111 14309 54163
rect 14361 54111 14433 54163
rect 14485 54111 14557 54163
rect 14218 54039 14576 54111
rect 14237 53987 14309 54039
rect 14361 53987 14433 54039
rect 14485 53987 14557 54039
rect 14218 53915 14576 53987
rect 14237 53863 14309 53915
rect 14361 53863 14433 53915
rect 14485 53863 14557 53915
rect 14218 53791 14576 53863
rect 14237 53739 14309 53791
rect 14361 53739 14433 53791
rect 14485 53739 14557 53791
rect 14218 53692 14576 53739
rect 14161 53667 14576 53692
rect 14161 53615 14185 53667
rect 14237 53615 14309 53667
rect 14361 53615 14433 53667
rect 14485 53615 14557 53667
rect 12305 53557 12489 53565
rect 10725 53505 10775 53543
rect 4203 53491 10775 53505
rect 10827 53491 10899 53543
rect 10951 53491 11023 53543
rect 11075 53505 11125 53543
rect 14161 53543 14576 53615
rect 14161 53505 14185 53543
rect 11075 53491 14185 53505
rect 14237 53491 14309 53543
rect 14361 53491 14433 53543
rect 14485 53491 14557 53543
rect 402 53483 14576 53491
rect 402 53431 869 53483
rect 921 53431 977 53483
rect 1029 53431 1085 53483
rect 1137 53431 1193 53483
rect 1245 53431 1301 53483
rect 1353 53431 1409 53483
rect 1461 53431 1517 53483
rect 1569 53431 1625 53483
rect 1677 53431 1733 53483
rect 1785 53431 1841 53483
rect 1893 53431 1949 53483
rect 2001 53431 2057 53483
rect 2109 53431 2763 53483
rect 2815 53431 2871 53483
rect 2923 53431 2979 53483
rect 3031 53431 3087 53483
rect 3139 53431 3195 53483
rect 3247 53431 3303 53483
rect 3355 53431 3411 53483
rect 3463 53431 3519 53483
rect 3571 53431 3627 53483
rect 3679 53431 3735 53483
rect 3787 53431 5138 53483
rect 5190 53431 5246 53483
rect 5298 53431 5354 53483
rect 5406 53431 5462 53483
rect 5514 53431 5570 53483
rect 5622 53431 5678 53483
rect 5730 53431 5786 53483
rect 5838 53431 5894 53483
rect 5946 53431 6002 53483
rect 6054 53431 6110 53483
rect 6162 53431 6218 53483
rect 6270 53431 6326 53483
rect 6378 53431 6434 53483
rect 6486 53431 6542 53483
rect 6594 53431 6650 53483
rect 6702 53431 6758 53483
rect 6810 53431 6866 53483
rect 6918 53431 6974 53483
rect 7026 53431 7082 53483
rect 7134 53431 7844 53483
rect 7896 53431 7952 53483
rect 8004 53431 8060 53483
rect 8112 53431 8168 53483
rect 8220 53431 8276 53483
rect 8328 53431 8384 53483
rect 8436 53431 8492 53483
rect 8544 53431 8600 53483
rect 8652 53431 8708 53483
rect 8760 53431 8816 53483
rect 8868 53431 8924 53483
rect 8976 53431 9032 53483
rect 9084 53431 9140 53483
rect 9192 53431 9248 53483
rect 9300 53431 9356 53483
rect 9408 53431 9464 53483
rect 9516 53431 9572 53483
rect 9624 53431 9680 53483
rect 9732 53431 9788 53483
rect 9840 53431 11191 53483
rect 11243 53431 11299 53483
rect 11351 53431 11407 53483
rect 11459 53431 11515 53483
rect 11567 53431 11623 53483
rect 11675 53431 11731 53483
rect 11783 53431 11839 53483
rect 11891 53431 11947 53483
rect 11999 53431 12055 53483
rect 12107 53431 12163 53483
rect 12215 53431 12869 53483
rect 12921 53431 12977 53483
rect 13029 53431 13085 53483
rect 13137 53431 13193 53483
rect 13245 53431 13301 53483
rect 13353 53431 13409 53483
rect 13461 53431 13517 53483
rect 13569 53431 13625 53483
rect 13677 53431 13733 53483
rect 13785 53431 13841 53483
rect 13893 53431 13949 53483
rect 14001 53431 14057 53483
rect 14109 53431 14576 53483
rect 402 53419 14576 53431
rect 421 53367 493 53419
rect 545 53367 617 53419
rect 669 53367 741 53419
rect 793 53375 3903 53419
rect 793 53367 869 53375
rect 402 53323 869 53367
rect 921 53323 977 53375
rect 1029 53323 1085 53375
rect 1137 53323 1193 53375
rect 1245 53323 1301 53375
rect 1353 53323 1409 53375
rect 1461 53323 1517 53375
rect 1569 53323 1625 53375
rect 1677 53323 1733 53375
rect 1785 53323 1841 53375
rect 1893 53323 1949 53375
rect 2001 53323 2057 53375
rect 2109 53323 2763 53375
rect 2815 53323 2871 53375
rect 2923 53323 2979 53375
rect 3031 53323 3087 53375
rect 3139 53323 3195 53375
rect 3247 53323 3303 53375
rect 3355 53323 3411 53375
rect 3463 53323 3519 53375
rect 3571 53323 3627 53375
rect 3679 53323 3735 53375
rect 3787 53367 3903 53375
rect 3955 53367 4027 53419
rect 4079 53367 4151 53419
rect 4203 53375 10775 53419
rect 4203 53367 5138 53375
rect 3787 53323 5138 53367
rect 5190 53323 5246 53375
rect 5298 53323 5354 53375
rect 5406 53323 5462 53375
rect 5514 53323 5570 53375
rect 5622 53323 5678 53375
rect 5730 53323 5786 53375
rect 5838 53323 5894 53375
rect 5946 53323 6002 53375
rect 6054 53323 6110 53375
rect 6162 53323 6218 53375
rect 6270 53323 6326 53375
rect 6378 53323 6434 53375
rect 6486 53323 6542 53375
rect 6594 53323 6650 53375
rect 6702 53323 6758 53375
rect 6810 53323 6866 53375
rect 6918 53323 6974 53375
rect 7026 53323 7082 53375
rect 7134 53323 7844 53375
rect 7896 53323 7952 53375
rect 8004 53323 8060 53375
rect 8112 53323 8168 53375
rect 8220 53323 8276 53375
rect 8328 53323 8384 53375
rect 8436 53323 8492 53375
rect 8544 53323 8600 53375
rect 8652 53323 8708 53375
rect 8760 53323 8816 53375
rect 8868 53323 8924 53375
rect 8976 53323 9032 53375
rect 9084 53323 9140 53375
rect 9192 53323 9248 53375
rect 9300 53323 9356 53375
rect 9408 53323 9464 53375
rect 9516 53323 9572 53375
rect 9624 53323 9680 53375
rect 9732 53323 9788 53375
rect 9840 53367 10775 53375
rect 10827 53367 10899 53419
rect 10951 53367 11023 53419
rect 11075 53375 14185 53419
rect 11075 53367 11191 53375
rect 9840 53323 11191 53367
rect 11243 53323 11299 53375
rect 11351 53323 11407 53375
rect 11459 53323 11515 53375
rect 11567 53323 11623 53375
rect 11675 53323 11731 53375
rect 11783 53323 11839 53375
rect 11891 53323 11947 53375
rect 11999 53323 12055 53375
rect 12107 53323 12163 53375
rect 12215 53323 12869 53375
rect 12921 53323 12977 53375
rect 13029 53323 13085 53375
rect 13137 53323 13193 53375
rect 13245 53323 13301 53375
rect 13353 53323 13409 53375
rect 13461 53323 13517 53375
rect 13569 53323 13625 53375
rect 13677 53323 13733 53375
rect 13785 53323 13841 53375
rect 13893 53323 13949 53375
rect 14001 53323 14057 53375
rect 14109 53367 14185 53375
rect 14237 53367 14309 53419
rect 14361 53367 14433 53419
rect 14485 53367 14557 53419
rect 14109 53323 14576 53367
rect 402 53295 14576 53323
rect 421 53243 493 53295
rect 545 53251 617 53295
rect 669 53251 741 53295
rect 793 53267 3903 53295
rect 793 53251 869 53267
rect 921 53251 977 53267
rect 1029 53251 1085 53267
rect 1137 53251 1193 53267
rect 1245 53251 1301 53267
rect 1353 53251 1409 53267
rect 1461 53251 1517 53267
rect 1569 53251 1625 53267
rect 1677 53251 1733 53267
rect 1785 53251 1841 53267
rect 1893 53251 1949 53267
rect 2001 53251 2057 53267
rect 2109 53251 2763 53267
rect 2815 53251 2871 53267
rect 2923 53251 2979 53267
rect 3031 53251 3087 53267
rect 3139 53251 3195 53267
rect 3247 53251 3303 53267
rect 3355 53251 3411 53267
rect 3463 53251 3519 53267
rect 3571 53251 3627 53267
rect 3679 53251 3735 53267
rect 3787 53251 3903 53267
rect 3955 53251 4027 53295
rect 4079 53251 4151 53295
rect 4203 53267 10775 53295
rect 4203 53251 5138 53267
rect 5190 53251 5246 53267
rect 5298 53251 5354 53267
rect 5406 53251 5462 53267
rect 5514 53251 5570 53267
rect 5622 53251 5678 53267
rect 5730 53251 5786 53267
rect 5838 53251 5894 53267
rect 5946 53251 6002 53267
rect 6054 53251 6110 53267
rect 6162 53251 6218 53267
rect 6270 53251 6326 53267
rect 6378 53251 6434 53267
rect 6486 53251 6542 53267
rect 6594 53251 6650 53267
rect 6702 53251 6758 53267
rect 6810 53251 6866 53267
rect 6918 53251 6974 53267
rect 7026 53251 7082 53267
rect 7134 53251 7844 53267
rect 7896 53251 7952 53267
rect 8004 53251 8060 53267
rect 8112 53251 8168 53267
rect 8220 53251 8276 53267
rect 8328 53251 8384 53267
rect 8436 53251 8492 53267
rect 8544 53251 8600 53267
rect 8652 53251 8708 53267
rect 8760 53251 8816 53267
rect 8868 53251 8924 53267
rect 8976 53251 9032 53267
rect 9084 53251 9140 53267
rect 9192 53251 9248 53267
rect 9300 53251 9356 53267
rect 9408 53251 9464 53267
rect 9516 53251 9572 53267
rect 9624 53251 9680 53267
rect 9732 53251 9788 53267
rect 9840 53251 10775 53267
rect 10827 53251 10899 53295
rect 10951 53251 11023 53295
rect 11075 53267 14185 53295
rect 11075 53251 11191 53267
rect 11243 53251 11299 53267
rect 11351 53251 11407 53267
rect 11459 53251 11515 53267
rect 11567 53251 11623 53267
rect 11675 53251 11731 53267
rect 11783 53251 11839 53267
rect 11891 53251 11947 53267
rect 11999 53251 12055 53267
rect 12107 53251 12163 53267
rect 12215 53251 12869 53267
rect 12921 53251 12977 53267
rect 13029 53251 13085 53267
rect 13137 53251 13193 53267
rect 13245 53251 13301 53267
rect 13353 53251 13409 53267
rect 13461 53251 13517 53267
rect 13569 53251 13625 53267
rect 13677 53251 13733 53267
rect 13785 53251 13841 53267
rect 13893 53251 13949 53267
rect 14001 53251 14057 53267
rect 14109 53251 14185 53267
rect 14237 53251 14309 53295
rect 14361 53251 14433 53295
rect 402 53205 510 53243
rect 14485 53243 14557 53295
rect 14468 53205 14576 53243
rect 14622 53205 14633 57105
rect 14892 57099 14904 57151
rect 14956 57099 14968 57151
rect 14892 57043 14968 57099
rect 14892 56991 14904 57043
rect 14956 56991 14968 57043
rect 14892 56935 14968 56991
rect 14892 56883 14904 56935
rect 14956 56883 14968 56935
rect 14892 56827 14968 56883
rect 14892 56775 14904 56827
rect 14956 56775 14968 56827
rect 14892 56719 14968 56775
rect 14892 56667 14904 56719
rect 14956 56667 14968 56719
rect 14892 56611 14968 56667
rect 14892 56559 14904 56611
rect 14956 56559 14968 56611
rect 14892 56503 14968 56559
rect 14892 56451 14904 56503
rect 14956 56451 14968 56503
rect 14892 56395 14968 56451
rect 14892 56343 14904 56395
rect 14956 56343 14968 56395
rect 14892 56287 14968 56343
rect 14892 56235 14904 56287
rect 14956 56235 14968 56287
rect 14892 56179 14968 56235
rect 14892 56127 14904 56179
rect 14956 56127 14968 56179
rect 14892 56071 14968 56127
rect 14892 56019 14904 56071
rect 14956 56019 14968 56071
rect 14892 56007 14968 56019
rect 345 53194 14633 53205
rect 14892 54174 14968 54186
rect 14892 54122 14904 54174
rect 14956 54122 14968 54174
rect 14892 54066 14968 54122
rect 14892 54014 14904 54066
rect 14956 54014 14968 54066
rect 14892 53958 14968 54014
rect 14892 53906 14904 53958
rect 14956 53906 14968 53958
rect 14892 53850 14968 53906
rect 14892 53798 14904 53850
rect 14956 53798 14968 53850
rect 14892 53742 14968 53798
rect 14892 53690 14904 53742
rect 14956 53690 14968 53742
rect 14892 53634 14968 53690
rect 14892 53582 14904 53634
rect 14956 53582 14968 53634
rect 14892 53526 14968 53582
rect 14892 53474 14904 53526
rect 14956 53474 14968 53526
rect 14892 53418 14968 53474
rect 14892 53366 14904 53418
rect 14956 53366 14968 53418
rect 14892 53310 14968 53366
rect 14892 53258 14904 53310
rect 14956 53258 14968 53310
rect 14892 53202 14968 53258
rect 10 53094 86 53150
rect 10 53042 22 53094
rect 74 53042 86 53094
rect 10 52986 86 53042
rect 10 52934 22 52986
rect 74 52934 86 52986
rect 10 52878 86 52934
rect 10 52826 22 52878
rect 74 52826 86 52878
rect 10 52814 86 52826
rect 14892 53150 14904 53202
rect 14956 53150 14968 53202
rect 14892 53094 14968 53150
rect 14892 53042 14904 53094
rect 14956 53042 14968 53094
rect 14892 52986 14968 53042
rect 14892 52934 14904 52986
rect 14956 52934 14968 52986
rect 14892 52878 14968 52934
rect 14892 52826 14904 52878
rect 14956 52826 14968 52878
rect 14892 52814 14968 52826
rect 71 52611 2225 52622
rect 71 52586 268 52611
rect 10 52574 268 52586
rect 10 52522 22 52574
rect 74 52522 268 52574
rect 10 52466 268 52522
rect 10 52414 22 52466
rect 74 52414 268 52466
rect 10 52358 268 52414
rect 10 52306 22 52358
rect 74 52306 268 52358
rect 10 52250 268 52306
rect 10 52198 22 52250
rect 74 52198 268 52250
rect 10 52142 268 52198
rect 10 52090 22 52142
rect 74 52090 268 52142
rect 10 52034 268 52090
rect 10 51982 22 52034
rect 74 51982 268 52034
rect 10 51926 268 51982
rect 10 51874 22 51926
rect 74 51874 268 51926
rect 10 51818 268 51874
rect 10 51766 22 51818
rect 74 51766 268 51818
rect 10 51710 268 51766
rect 10 51658 22 51710
rect 74 51658 268 51710
rect 10 51622 268 51658
rect 10 51602 86 51622
rect 10 51550 22 51602
rect 74 51550 86 51602
rect 10 51494 86 51550
rect 10 51442 22 51494
rect 74 51442 86 51494
rect 10 51422 86 51442
rect 257 51422 268 51622
rect 10 51386 268 51422
rect 10 51334 22 51386
rect 74 51334 268 51386
rect 10 51278 268 51334
rect 10 51226 22 51278
rect 74 51226 268 51278
rect 10 51214 268 51226
rect 71 50422 268 51214
rect 257 49854 268 50422
rect 71 49386 268 49854
rect 10 49374 268 49386
rect 10 49322 22 49374
rect 74 49322 268 49374
rect 10 49266 268 49322
rect 10 49214 22 49266
rect 74 49214 268 49266
rect 10 49158 268 49214
rect 10 49106 22 49158
rect 74 49106 268 49158
rect 10 49050 268 49106
rect 10 48998 22 49050
rect 74 48998 268 49050
rect 10 48942 268 48998
rect 10 48890 22 48942
rect 74 48890 268 48942
rect 10 48854 268 48890
rect 10 48834 86 48854
rect 10 48782 22 48834
rect 74 48782 86 48834
rect 10 48726 86 48782
rect 10 48674 22 48726
rect 74 48674 86 48726
rect 10 48654 86 48674
rect 257 48654 268 48854
rect 10 48618 268 48654
rect 10 48566 22 48618
rect 74 48566 268 48618
rect 10 48510 268 48566
rect 10 48458 22 48510
rect 74 48458 268 48510
rect 10 48402 268 48458
rect 10 48350 22 48402
rect 74 48350 268 48402
rect 10 48294 268 48350
rect 10 48242 22 48294
rect 74 48242 268 48294
rect 10 48186 268 48242
rect 10 48134 22 48186
rect 74 48134 268 48186
rect 10 48078 268 48134
rect 10 48026 22 48078
rect 74 48026 268 48078
rect 10 48014 268 48026
rect 71 47665 268 48014
rect 2214 47665 2225 52611
rect 71 47654 2225 47665
rect 2551 52611 12427 52622
rect 2551 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52254 12070 52265
rect 2908 48022 2919 52254
rect 3105 52029 11873 52040
rect 3105 51983 3142 52029
rect 11836 51983 11873 52029
rect 3105 51957 3161 51983
rect 3213 51957 3269 51983
rect 3321 51957 3377 51983
rect 3429 51957 3485 51983
rect 3537 51957 3593 51983
rect 3645 51957 3701 51983
rect 3753 51957 3809 51983
rect 3861 51957 3917 51983
rect 3969 51957 4025 51983
rect 4077 51957 4133 51983
rect 4185 51957 4241 51983
rect 4293 51957 4349 51983
rect 4401 51957 4457 51983
rect 4509 51957 4565 51983
rect 4617 51957 4673 51983
rect 4725 51957 5138 51983
rect 5190 51957 5246 51983
rect 5298 51957 5354 51983
rect 5406 51957 5462 51983
rect 5514 51957 5570 51983
rect 5622 51957 5678 51983
rect 5730 51957 5786 51983
rect 5838 51957 5894 51983
rect 5946 51957 6002 51983
rect 6054 51957 6110 51983
rect 6162 51957 6218 51983
rect 6270 51957 6326 51983
rect 6378 51957 6434 51983
rect 6486 51957 6542 51983
rect 6594 51957 6650 51983
rect 6702 51957 6758 51983
rect 6810 51957 6866 51983
rect 6918 51957 6974 51983
rect 7026 51957 7082 51983
rect 7134 51957 7844 51983
rect 7896 51957 7952 51983
rect 8004 51957 8060 51983
rect 8112 51957 8168 51983
rect 8220 51957 8276 51983
rect 8328 51957 8384 51983
rect 8436 51957 8492 51983
rect 8544 51957 8600 51983
rect 8652 51957 8708 51983
rect 8760 51957 8816 51983
rect 8868 51957 8924 51983
rect 8976 51957 9032 51983
rect 9084 51957 9140 51983
rect 9192 51957 9248 51983
rect 9300 51957 9356 51983
rect 9408 51957 9464 51983
rect 9516 51957 9572 51983
rect 9624 51957 9680 51983
rect 9732 51957 9788 51983
rect 9840 51957 10253 51983
rect 10305 51957 10361 51983
rect 10413 51957 10469 51983
rect 10521 51957 10577 51983
rect 10629 51957 10685 51983
rect 10737 51957 10793 51983
rect 10845 51957 10901 51983
rect 10953 51957 11009 51983
rect 11061 51957 11117 51983
rect 11169 51957 11225 51983
rect 11277 51957 11333 51983
rect 11385 51957 11441 51983
rect 11493 51957 11549 51983
rect 11601 51957 11657 51983
rect 11709 51957 11765 51983
rect 11817 51957 11873 51983
rect 3105 51901 11873 51957
rect 3105 51900 3161 51901
rect 3105 48376 3116 51900
rect 3213 51849 3269 51901
rect 3321 51849 3377 51901
rect 3429 51875 3485 51901
rect 3537 51875 3593 51901
rect 3645 51875 3701 51901
rect 3753 51875 3809 51901
rect 3861 51875 3917 51901
rect 3969 51875 4025 51901
rect 4077 51875 4133 51901
rect 4185 51875 4241 51901
rect 4293 51875 4349 51901
rect 4401 51875 4457 51901
rect 4509 51875 4565 51901
rect 4617 51875 4673 51901
rect 4725 51875 5138 51901
rect 5190 51875 5246 51901
rect 5298 51875 5354 51901
rect 5406 51875 5462 51901
rect 5514 51875 5570 51901
rect 5622 51875 5678 51901
rect 5730 51875 5786 51901
rect 5838 51875 5894 51901
rect 5946 51875 6002 51901
rect 6054 51875 6110 51901
rect 6162 51875 6218 51901
rect 6270 51875 6326 51901
rect 6378 51875 6434 51901
rect 6486 51875 6542 51901
rect 6594 51875 6650 51901
rect 6702 51875 6758 51901
rect 6810 51875 6866 51901
rect 6918 51875 6974 51901
rect 7026 51875 7082 51901
rect 7134 51875 7844 51901
rect 7896 51875 7952 51901
rect 8004 51875 8060 51901
rect 8112 51875 8168 51901
rect 8220 51875 8276 51901
rect 8328 51875 8384 51901
rect 8436 51875 8492 51901
rect 8544 51875 8600 51901
rect 8652 51875 8708 51901
rect 8760 51875 8816 51901
rect 8868 51875 8924 51901
rect 8976 51875 9032 51901
rect 9084 51875 9140 51901
rect 9192 51875 9248 51901
rect 9300 51875 9356 51901
rect 9408 51875 9464 51901
rect 9516 51875 9572 51901
rect 9624 51875 9680 51901
rect 9732 51875 9788 51901
rect 9840 51875 10253 51901
rect 10305 51875 10361 51901
rect 10413 51875 10469 51901
rect 10521 51875 10577 51901
rect 10629 51875 10685 51901
rect 10737 51875 10793 51901
rect 10845 51875 10901 51901
rect 10953 51875 11009 51901
rect 11061 51875 11117 51901
rect 11169 51875 11225 51901
rect 11277 51875 11333 51901
rect 11385 51875 11441 51901
rect 11493 51875 11549 51901
rect 11601 51849 11657 51901
rect 11709 51849 11765 51901
rect 11817 51900 11873 51901
rect 3162 51844 3424 51849
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51849
rect 11554 51829 11662 51844
rect 3316 51818 11662 51829
rect 3316 51260 3327 51818
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51567 4871 51580
rect 4923 51567 4979 51580
rect 5031 51567 7247 51580
rect 7299 51567 7355 51580
rect 7407 51567 7463 51580
rect 7515 51567 7571 51580
rect 7623 51567 7679 51580
rect 7731 51567 9947 51580
rect 9999 51567 10055 51580
rect 10107 51567 11489 51580
rect 3489 51511 11489 51567
rect 3489 51498 4871 51511
rect 4923 51498 4979 51511
rect 5031 51498 7247 51511
rect 7299 51498 7355 51511
rect 7407 51498 7463 51511
rect 7515 51498 7571 51511
rect 7623 51498 7679 51511
rect 7731 51498 9947 51511
rect 9999 51498 10055 51511
rect 10107 51498 11489 51511
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 11651 51260 11662 51818
rect 3316 51249 11662 51260
rect 3316 51234 3424 51249
rect 3162 51206 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51206 11816 51234
rect 3213 51154 3269 51206
rect 3321 51154 3377 51206
rect 3429 51154 3485 51203
rect 3537 51154 3593 51203
rect 3645 51154 3701 51203
rect 3753 51154 3809 51203
rect 3861 51154 3917 51203
rect 3969 51154 4025 51203
rect 4077 51154 4133 51203
rect 4185 51154 4241 51203
rect 4293 51154 4349 51203
rect 4401 51154 4457 51203
rect 4509 51154 4565 51203
rect 4617 51154 4673 51203
rect 4725 51154 5138 51203
rect 5190 51154 5246 51203
rect 5298 51154 5354 51203
rect 5406 51154 5462 51203
rect 5514 51154 5570 51203
rect 5622 51154 5678 51203
rect 5730 51154 5786 51203
rect 5838 51154 5894 51203
rect 5946 51154 6002 51203
rect 6054 51154 6110 51203
rect 6162 51154 6218 51203
rect 6270 51154 6326 51203
rect 6378 51154 6434 51203
rect 6486 51154 6542 51203
rect 6594 51154 6650 51203
rect 6702 51154 6758 51203
rect 6810 51154 6866 51203
rect 6918 51154 6974 51203
rect 7026 51154 7082 51203
rect 7134 51154 7844 51203
rect 7896 51154 7952 51203
rect 8004 51154 8060 51203
rect 8112 51154 8168 51203
rect 8220 51154 8276 51203
rect 8328 51154 8384 51203
rect 8436 51154 8492 51203
rect 8544 51154 8600 51203
rect 8652 51154 8708 51203
rect 8760 51154 8816 51203
rect 8868 51154 8924 51203
rect 8976 51154 9032 51203
rect 9084 51154 9140 51203
rect 9192 51154 9248 51203
rect 9300 51154 9356 51203
rect 9408 51154 9464 51203
rect 9516 51154 9572 51203
rect 9624 51154 9680 51203
rect 9732 51154 9788 51203
rect 9840 51154 10253 51203
rect 10305 51154 10361 51203
rect 10413 51154 10469 51203
rect 10521 51154 10577 51203
rect 10629 51154 10685 51203
rect 10737 51154 10793 51203
rect 10845 51154 10901 51203
rect 10953 51154 11009 51203
rect 11061 51154 11117 51203
rect 11169 51154 11225 51203
rect 11277 51154 11333 51203
rect 11385 51154 11441 51203
rect 11493 51154 11549 51203
rect 11601 51154 11657 51206
rect 11709 51154 11765 51206
rect 3162 51098 11816 51154
rect 3213 51046 3269 51098
rect 3321 51095 3377 51098
rect 3429 51095 3485 51098
rect 3537 51095 3593 51098
rect 3645 51095 3701 51098
rect 3753 51095 3809 51098
rect 3861 51095 3917 51098
rect 3969 51095 4025 51098
rect 4077 51095 4133 51098
rect 4185 51095 4241 51098
rect 4293 51095 4349 51098
rect 4401 51095 4457 51098
rect 4509 51095 4565 51098
rect 4617 51095 4673 51098
rect 4725 51095 5138 51098
rect 5190 51095 5246 51098
rect 5298 51095 5354 51098
rect 5406 51095 5462 51098
rect 5514 51095 5570 51098
rect 5622 51095 5678 51098
rect 5730 51095 5786 51098
rect 5838 51095 5894 51098
rect 5946 51095 6002 51098
rect 6054 51095 6110 51098
rect 6162 51095 6218 51098
rect 6270 51095 6326 51098
rect 6378 51095 6434 51098
rect 6486 51095 6542 51098
rect 6594 51095 6650 51098
rect 6702 51095 6758 51098
rect 6810 51095 6866 51098
rect 6918 51095 6974 51098
rect 7026 51095 7082 51098
rect 7134 51095 7844 51098
rect 7896 51095 7952 51098
rect 8004 51095 8060 51098
rect 8112 51095 8168 51098
rect 8220 51095 8276 51098
rect 8328 51095 8384 51098
rect 8436 51095 8492 51098
rect 8544 51095 8600 51098
rect 8652 51095 8708 51098
rect 8760 51095 8816 51098
rect 8868 51095 8924 51098
rect 8976 51095 9032 51098
rect 9084 51095 9140 51098
rect 9192 51095 9248 51098
rect 9300 51095 9356 51098
rect 9408 51095 9464 51098
rect 9516 51095 9572 51098
rect 9624 51095 9680 51098
rect 9732 51095 9788 51098
rect 9840 51095 10253 51098
rect 10305 51095 10361 51098
rect 10413 51095 10469 51098
rect 10521 51095 10577 51098
rect 10629 51095 10685 51098
rect 10737 51095 10793 51098
rect 10845 51095 10901 51098
rect 10953 51095 11009 51098
rect 11061 51095 11117 51098
rect 11169 51095 11225 51098
rect 11277 51095 11333 51098
rect 11385 51095 11441 51098
rect 11493 51095 11549 51098
rect 11601 51095 11657 51098
rect 3321 51049 3330 51095
rect 11648 51049 11657 51095
rect 3321 51046 3377 51049
rect 3429 51046 3485 51049
rect 3537 51046 3593 51049
rect 3645 51046 3701 51049
rect 3753 51046 3809 51049
rect 3861 51046 3917 51049
rect 3969 51046 4025 51049
rect 4077 51046 4133 51049
rect 4185 51046 4241 51049
rect 4293 51046 4349 51049
rect 4401 51046 4457 51049
rect 4509 51046 4565 51049
rect 4617 51046 4673 51049
rect 4725 51046 5138 51049
rect 5190 51046 5246 51049
rect 5298 51046 5354 51049
rect 5406 51046 5462 51049
rect 5514 51046 5570 51049
rect 5622 51046 5678 51049
rect 5730 51046 5786 51049
rect 5838 51046 5894 51049
rect 5946 51046 6002 51049
rect 6054 51046 6110 51049
rect 6162 51046 6218 51049
rect 6270 51046 6326 51049
rect 6378 51046 6434 51049
rect 6486 51046 6542 51049
rect 6594 51046 6650 51049
rect 6702 51046 6758 51049
rect 6810 51046 6866 51049
rect 6918 51046 6974 51049
rect 7026 51046 7082 51049
rect 7134 51046 7844 51049
rect 7896 51046 7952 51049
rect 8004 51046 8060 51049
rect 8112 51046 8168 51049
rect 8220 51046 8276 51049
rect 8328 51046 8384 51049
rect 8436 51046 8492 51049
rect 8544 51046 8600 51049
rect 8652 51046 8708 51049
rect 8760 51046 8816 51049
rect 8868 51046 8924 51049
rect 8976 51046 9032 51049
rect 9084 51046 9140 51049
rect 9192 51046 9248 51049
rect 9300 51046 9356 51049
rect 9408 51046 9464 51049
rect 9516 51046 9572 51049
rect 9624 51046 9680 51049
rect 9732 51046 9788 51049
rect 9840 51046 10253 51049
rect 10305 51046 10361 51049
rect 10413 51046 10469 51049
rect 10521 51046 10577 51049
rect 10629 51046 10685 51049
rect 10737 51046 10793 51049
rect 10845 51046 10901 51049
rect 10953 51046 11009 51049
rect 11061 51046 11117 51049
rect 11169 51046 11225 51049
rect 11277 51046 11333 51049
rect 11385 51046 11441 51049
rect 11493 51046 11549 51049
rect 11601 51046 11657 51049
rect 11709 51046 11765 51098
rect 3162 50990 11816 51046
rect 3213 50938 3269 50990
rect 3321 50938 3377 50990
rect 3429 50941 3485 50990
rect 3537 50941 3593 50990
rect 3645 50941 3701 50990
rect 3753 50941 3809 50990
rect 3861 50941 3917 50990
rect 3969 50941 4025 50990
rect 4077 50941 4133 50990
rect 4185 50941 4241 50990
rect 4293 50941 4349 50990
rect 4401 50941 4457 50990
rect 4509 50941 4565 50990
rect 4617 50941 4673 50990
rect 4725 50941 5138 50990
rect 5190 50941 5246 50990
rect 5298 50941 5354 50990
rect 5406 50941 5462 50990
rect 5514 50941 5570 50990
rect 5622 50941 5678 50990
rect 5730 50941 5786 50990
rect 5838 50941 5894 50990
rect 5946 50941 6002 50990
rect 6054 50941 6110 50990
rect 6162 50941 6218 50990
rect 6270 50941 6326 50990
rect 6378 50941 6434 50990
rect 6486 50941 6542 50990
rect 6594 50941 6650 50990
rect 6702 50941 6758 50990
rect 6810 50941 6866 50990
rect 6918 50941 6974 50990
rect 7026 50941 7082 50990
rect 7134 50941 7844 50990
rect 7896 50941 7952 50990
rect 8004 50941 8060 50990
rect 8112 50941 8168 50990
rect 8220 50941 8276 50990
rect 8328 50941 8384 50990
rect 8436 50941 8492 50990
rect 8544 50941 8600 50990
rect 8652 50941 8708 50990
rect 8760 50941 8816 50990
rect 8868 50941 8924 50990
rect 8976 50941 9032 50990
rect 9084 50941 9140 50990
rect 9192 50941 9248 50990
rect 9300 50941 9356 50990
rect 9408 50941 9464 50990
rect 9516 50941 9572 50990
rect 9624 50941 9680 50990
rect 9732 50941 9788 50990
rect 9840 50941 10253 50990
rect 10305 50941 10361 50990
rect 10413 50941 10469 50990
rect 10521 50941 10577 50990
rect 10629 50941 10685 50990
rect 10737 50941 10793 50990
rect 10845 50941 10901 50990
rect 10953 50941 11009 50990
rect 11061 50941 11117 50990
rect 11169 50941 11225 50990
rect 11277 50941 11333 50990
rect 11385 50941 11441 50990
rect 11493 50941 11549 50990
rect 11601 50938 11657 50990
rect 11709 50938 11765 50990
rect 3162 50910 3424 50938
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50938
rect 11554 50895 11662 50910
rect 3316 50884 11662 50895
rect 3316 50326 3327 50884
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50633 4871 50646
rect 4923 50633 4979 50646
rect 5031 50633 7247 50646
rect 7299 50633 7355 50646
rect 7407 50633 7463 50646
rect 7515 50633 7571 50646
rect 7623 50633 7679 50646
rect 7731 50633 9947 50646
rect 9999 50633 10055 50646
rect 10107 50633 11489 50646
rect 3489 50577 11489 50633
rect 3489 50564 4871 50577
rect 4923 50564 4979 50577
rect 5031 50564 7247 50577
rect 7299 50564 7355 50577
rect 7407 50564 7463 50577
rect 7515 50564 7571 50577
rect 7623 50564 7679 50577
rect 7731 50564 9947 50577
rect 9999 50564 10055 50577
rect 10107 50564 11489 50577
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 11651 50326 11662 50884
rect 3316 50315 11662 50326
rect 3316 50300 3424 50315
rect 3162 50272 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50272 11816 50300
rect 3213 50220 3269 50272
rect 3321 50220 3377 50272
rect 3429 50220 3485 50269
rect 3537 50220 3593 50269
rect 3645 50220 3701 50269
rect 3753 50220 3809 50269
rect 3861 50220 3917 50269
rect 3969 50220 4025 50269
rect 4077 50220 4133 50269
rect 4185 50220 4241 50269
rect 4293 50220 4349 50269
rect 4401 50220 4457 50269
rect 4509 50220 4565 50269
rect 4617 50220 4673 50269
rect 4725 50220 5138 50269
rect 5190 50220 5246 50269
rect 5298 50220 5354 50269
rect 5406 50220 5462 50269
rect 5514 50220 5570 50269
rect 5622 50220 5678 50269
rect 5730 50220 5786 50269
rect 5838 50220 5894 50269
rect 5946 50220 6002 50269
rect 6054 50220 6110 50269
rect 6162 50220 6218 50269
rect 6270 50220 6326 50269
rect 6378 50220 6434 50269
rect 6486 50220 6542 50269
rect 6594 50220 6650 50269
rect 6702 50220 6758 50269
rect 6810 50220 6866 50269
rect 6918 50220 6974 50269
rect 7026 50220 7082 50269
rect 7134 50220 7844 50269
rect 7896 50220 7952 50269
rect 8004 50220 8060 50269
rect 8112 50220 8168 50269
rect 8220 50220 8276 50269
rect 8328 50220 8384 50269
rect 8436 50220 8492 50269
rect 8544 50220 8600 50269
rect 8652 50220 8708 50269
rect 8760 50220 8816 50269
rect 8868 50220 8924 50269
rect 8976 50220 9032 50269
rect 9084 50220 9140 50269
rect 9192 50220 9248 50269
rect 9300 50220 9356 50269
rect 9408 50220 9464 50269
rect 9516 50220 9572 50269
rect 9624 50220 9680 50269
rect 9732 50220 9788 50269
rect 9840 50220 10253 50269
rect 10305 50220 10361 50269
rect 10413 50220 10469 50269
rect 10521 50220 10577 50269
rect 10629 50220 10685 50269
rect 10737 50220 10793 50269
rect 10845 50220 10901 50269
rect 10953 50220 11009 50269
rect 11061 50220 11117 50269
rect 11169 50220 11225 50269
rect 11277 50220 11333 50269
rect 11385 50220 11441 50269
rect 11493 50220 11549 50269
rect 11601 50220 11657 50272
rect 11709 50220 11765 50272
rect 3162 50164 11816 50220
rect 3213 50112 3269 50164
rect 3321 50161 3377 50164
rect 3429 50161 3485 50164
rect 3537 50161 3593 50164
rect 3645 50161 3701 50164
rect 3753 50161 3809 50164
rect 3861 50161 3917 50164
rect 3969 50161 4025 50164
rect 4077 50161 4133 50164
rect 4185 50161 4241 50164
rect 4293 50161 4349 50164
rect 4401 50161 4457 50164
rect 4509 50161 4565 50164
rect 4617 50161 4673 50164
rect 4725 50161 5138 50164
rect 5190 50161 5246 50164
rect 5298 50161 5354 50164
rect 5406 50161 5462 50164
rect 5514 50161 5570 50164
rect 5622 50161 5678 50164
rect 5730 50161 5786 50164
rect 5838 50161 5894 50164
rect 5946 50161 6002 50164
rect 6054 50161 6110 50164
rect 6162 50161 6218 50164
rect 6270 50161 6326 50164
rect 6378 50161 6434 50164
rect 6486 50161 6542 50164
rect 6594 50161 6650 50164
rect 6702 50161 6758 50164
rect 6810 50161 6866 50164
rect 6918 50161 6974 50164
rect 7026 50161 7082 50164
rect 7134 50161 7844 50164
rect 7896 50161 7952 50164
rect 8004 50161 8060 50164
rect 8112 50161 8168 50164
rect 8220 50161 8276 50164
rect 8328 50161 8384 50164
rect 8436 50161 8492 50164
rect 8544 50161 8600 50164
rect 8652 50161 8708 50164
rect 8760 50161 8816 50164
rect 8868 50161 8924 50164
rect 8976 50161 9032 50164
rect 9084 50161 9140 50164
rect 9192 50161 9248 50164
rect 9300 50161 9356 50164
rect 9408 50161 9464 50164
rect 9516 50161 9572 50164
rect 9624 50161 9680 50164
rect 9732 50161 9788 50164
rect 9840 50161 10253 50164
rect 10305 50161 10361 50164
rect 10413 50161 10469 50164
rect 10521 50161 10577 50164
rect 10629 50161 10685 50164
rect 10737 50161 10793 50164
rect 10845 50161 10901 50164
rect 10953 50161 11009 50164
rect 11061 50161 11117 50164
rect 11169 50161 11225 50164
rect 11277 50161 11333 50164
rect 11385 50161 11441 50164
rect 11493 50161 11549 50164
rect 11601 50161 11657 50164
rect 3321 50115 3330 50161
rect 11648 50115 11657 50161
rect 3321 50112 3377 50115
rect 3429 50112 3485 50115
rect 3537 50112 3593 50115
rect 3645 50112 3701 50115
rect 3753 50112 3809 50115
rect 3861 50112 3917 50115
rect 3969 50112 4025 50115
rect 4077 50112 4133 50115
rect 4185 50112 4241 50115
rect 4293 50112 4349 50115
rect 4401 50112 4457 50115
rect 4509 50112 4565 50115
rect 4617 50112 4673 50115
rect 4725 50112 5138 50115
rect 5190 50112 5246 50115
rect 5298 50112 5354 50115
rect 5406 50112 5462 50115
rect 5514 50112 5570 50115
rect 5622 50112 5678 50115
rect 5730 50112 5786 50115
rect 5838 50112 5894 50115
rect 5946 50112 6002 50115
rect 6054 50112 6110 50115
rect 6162 50112 6218 50115
rect 6270 50112 6326 50115
rect 6378 50112 6434 50115
rect 6486 50112 6542 50115
rect 6594 50112 6650 50115
rect 6702 50112 6758 50115
rect 6810 50112 6866 50115
rect 6918 50112 6974 50115
rect 7026 50112 7082 50115
rect 7134 50112 7844 50115
rect 7896 50112 7952 50115
rect 8004 50112 8060 50115
rect 8112 50112 8168 50115
rect 8220 50112 8276 50115
rect 8328 50112 8384 50115
rect 8436 50112 8492 50115
rect 8544 50112 8600 50115
rect 8652 50112 8708 50115
rect 8760 50112 8816 50115
rect 8868 50112 8924 50115
rect 8976 50112 9032 50115
rect 9084 50112 9140 50115
rect 9192 50112 9248 50115
rect 9300 50112 9356 50115
rect 9408 50112 9464 50115
rect 9516 50112 9572 50115
rect 9624 50112 9680 50115
rect 9732 50112 9788 50115
rect 9840 50112 10253 50115
rect 10305 50112 10361 50115
rect 10413 50112 10469 50115
rect 10521 50112 10577 50115
rect 10629 50112 10685 50115
rect 10737 50112 10793 50115
rect 10845 50112 10901 50115
rect 10953 50112 11009 50115
rect 11061 50112 11117 50115
rect 11169 50112 11225 50115
rect 11277 50112 11333 50115
rect 11385 50112 11441 50115
rect 11493 50112 11549 50115
rect 11601 50112 11657 50115
rect 11709 50112 11765 50164
rect 3162 50056 11816 50112
rect 3213 50004 3269 50056
rect 3321 50004 3377 50056
rect 3429 50007 3485 50056
rect 3537 50007 3593 50056
rect 3645 50007 3701 50056
rect 3753 50007 3809 50056
rect 3861 50007 3917 50056
rect 3969 50007 4025 50056
rect 4077 50007 4133 50056
rect 4185 50007 4241 50056
rect 4293 50007 4349 50056
rect 4401 50007 4457 50056
rect 4509 50007 4565 50056
rect 4617 50007 4673 50056
rect 4725 50007 5138 50056
rect 5190 50007 5246 50056
rect 5298 50007 5354 50056
rect 5406 50007 5462 50056
rect 5514 50007 5570 50056
rect 5622 50007 5678 50056
rect 5730 50007 5786 50056
rect 5838 50007 5894 50056
rect 5946 50007 6002 50056
rect 6054 50007 6110 50056
rect 6162 50007 6218 50056
rect 6270 50007 6326 50056
rect 6378 50007 6434 50056
rect 6486 50007 6542 50056
rect 6594 50007 6650 50056
rect 6702 50007 6758 50056
rect 6810 50007 6866 50056
rect 6918 50007 6974 50056
rect 7026 50007 7082 50056
rect 7134 50007 7844 50056
rect 7896 50007 7952 50056
rect 8004 50007 8060 50056
rect 8112 50007 8168 50056
rect 8220 50007 8276 50056
rect 8328 50007 8384 50056
rect 8436 50007 8492 50056
rect 8544 50007 8600 50056
rect 8652 50007 8708 50056
rect 8760 50007 8816 50056
rect 8868 50007 8924 50056
rect 8976 50007 9032 50056
rect 9084 50007 9140 50056
rect 9192 50007 9248 50056
rect 9300 50007 9356 50056
rect 9408 50007 9464 50056
rect 9516 50007 9572 50056
rect 9624 50007 9680 50056
rect 9732 50007 9788 50056
rect 9840 50007 10253 50056
rect 10305 50007 10361 50056
rect 10413 50007 10469 50056
rect 10521 50007 10577 50056
rect 10629 50007 10685 50056
rect 10737 50007 10793 50056
rect 10845 50007 10901 50056
rect 10953 50007 11009 50056
rect 11061 50007 11117 50056
rect 11169 50007 11225 50056
rect 11277 50007 11333 50056
rect 11385 50007 11441 50056
rect 11493 50007 11549 50056
rect 11601 50004 11657 50056
rect 11709 50004 11765 50056
rect 3162 49976 3424 50004
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50004
rect 11554 49961 11662 49976
rect 3316 49950 11662 49961
rect 3316 49392 3327 49950
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49699 4871 49712
rect 4923 49699 4979 49712
rect 5031 49699 7247 49712
rect 7299 49699 7355 49712
rect 7407 49699 7463 49712
rect 7515 49699 7571 49712
rect 7623 49699 7679 49712
rect 7731 49699 9947 49712
rect 9999 49699 10055 49712
rect 10107 49699 11489 49712
rect 3489 49643 11489 49699
rect 3489 49630 4871 49643
rect 4923 49630 4979 49643
rect 5031 49630 7247 49643
rect 7299 49630 7355 49643
rect 7407 49630 7463 49643
rect 7515 49630 7571 49643
rect 7623 49630 7679 49643
rect 7731 49630 9947 49643
rect 9999 49630 10055 49643
rect 10107 49630 11489 49643
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 11651 49392 11662 49950
rect 3316 49381 11662 49392
rect 3316 49366 3424 49381
rect 3162 49338 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49338 11816 49366
rect 3213 49286 3269 49338
rect 3321 49286 3377 49338
rect 3429 49286 3485 49335
rect 3537 49286 3593 49335
rect 3645 49286 3701 49335
rect 3753 49286 3809 49335
rect 3861 49286 3917 49335
rect 3969 49286 4025 49335
rect 4077 49286 4133 49335
rect 4185 49286 4241 49335
rect 4293 49286 4349 49335
rect 4401 49286 4457 49335
rect 4509 49286 4565 49335
rect 4617 49286 4673 49335
rect 4725 49286 5138 49335
rect 5190 49286 5246 49335
rect 5298 49286 5354 49335
rect 5406 49286 5462 49335
rect 5514 49286 5570 49335
rect 5622 49286 5678 49335
rect 5730 49286 5786 49335
rect 5838 49286 5894 49335
rect 5946 49286 6002 49335
rect 6054 49286 6110 49335
rect 6162 49286 6218 49335
rect 6270 49286 6326 49335
rect 6378 49286 6434 49335
rect 6486 49286 6542 49335
rect 6594 49286 6650 49335
rect 6702 49286 6758 49335
rect 6810 49286 6866 49335
rect 6918 49286 6974 49335
rect 7026 49286 7082 49335
rect 7134 49286 7844 49335
rect 7896 49286 7952 49335
rect 8004 49286 8060 49335
rect 8112 49286 8168 49335
rect 8220 49286 8276 49335
rect 8328 49286 8384 49335
rect 8436 49286 8492 49335
rect 8544 49286 8600 49335
rect 8652 49286 8708 49335
rect 8760 49286 8816 49335
rect 8868 49286 8924 49335
rect 8976 49286 9032 49335
rect 9084 49286 9140 49335
rect 9192 49286 9248 49335
rect 9300 49286 9356 49335
rect 9408 49286 9464 49335
rect 9516 49286 9572 49335
rect 9624 49286 9680 49335
rect 9732 49286 9788 49335
rect 9840 49286 10253 49335
rect 10305 49286 10361 49335
rect 10413 49286 10469 49335
rect 10521 49286 10577 49335
rect 10629 49286 10685 49335
rect 10737 49286 10793 49335
rect 10845 49286 10901 49335
rect 10953 49286 11009 49335
rect 11061 49286 11117 49335
rect 11169 49286 11225 49335
rect 11277 49286 11333 49335
rect 11385 49286 11441 49335
rect 11493 49286 11549 49335
rect 11601 49286 11657 49338
rect 11709 49286 11765 49338
rect 3162 49230 11816 49286
rect 3213 49178 3269 49230
rect 3321 49227 3377 49230
rect 3429 49227 3485 49230
rect 3537 49227 3593 49230
rect 3645 49227 3701 49230
rect 3753 49227 3809 49230
rect 3861 49227 3917 49230
rect 3969 49227 4025 49230
rect 4077 49227 4133 49230
rect 4185 49227 4241 49230
rect 4293 49227 4349 49230
rect 4401 49227 4457 49230
rect 4509 49227 4565 49230
rect 4617 49227 4673 49230
rect 4725 49227 5138 49230
rect 5190 49227 5246 49230
rect 5298 49227 5354 49230
rect 5406 49227 5462 49230
rect 5514 49227 5570 49230
rect 5622 49227 5678 49230
rect 5730 49227 5786 49230
rect 5838 49227 5894 49230
rect 5946 49227 6002 49230
rect 6054 49227 6110 49230
rect 6162 49227 6218 49230
rect 6270 49227 6326 49230
rect 6378 49227 6434 49230
rect 6486 49227 6542 49230
rect 6594 49227 6650 49230
rect 6702 49227 6758 49230
rect 6810 49227 6866 49230
rect 6918 49227 6974 49230
rect 7026 49227 7082 49230
rect 7134 49227 7844 49230
rect 7896 49227 7952 49230
rect 8004 49227 8060 49230
rect 8112 49227 8168 49230
rect 8220 49227 8276 49230
rect 8328 49227 8384 49230
rect 8436 49227 8492 49230
rect 8544 49227 8600 49230
rect 8652 49227 8708 49230
rect 8760 49227 8816 49230
rect 8868 49227 8924 49230
rect 8976 49227 9032 49230
rect 9084 49227 9140 49230
rect 9192 49227 9248 49230
rect 9300 49227 9356 49230
rect 9408 49227 9464 49230
rect 9516 49227 9572 49230
rect 9624 49227 9680 49230
rect 9732 49227 9788 49230
rect 9840 49227 10253 49230
rect 10305 49227 10361 49230
rect 10413 49227 10469 49230
rect 10521 49227 10577 49230
rect 10629 49227 10685 49230
rect 10737 49227 10793 49230
rect 10845 49227 10901 49230
rect 10953 49227 11009 49230
rect 11061 49227 11117 49230
rect 11169 49227 11225 49230
rect 11277 49227 11333 49230
rect 11385 49227 11441 49230
rect 11493 49227 11549 49230
rect 11601 49227 11657 49230
rect 3321 49181 3330 49227
rect 11648 49181 11657 49227
rect 3321 49178 3377 49181
rect 3429 49178 3485 49181
rect 3537 49178 3593 49181
rect 3645 49178 3701 49181
rect 3753 49178 3809 49181
rect 3861 49178 3917 49181
rect 3969 49178 4025 49181
rect 4077 49178 4133 49181
rect 4185 49178 4241 49181
rect 4293 49178 4349 49181
rect 4401 49178 4457 49181
rect 4509 49178 4565 49181
rect 4617 49178 4673 49181
rect 4725 49178 5138 49181
rect 5190 49178 5246 49181
rect 5298 49178 5354 49181
rect 5406 49178 5462 49181
rect 5514 49178 5570 49181
rect 5622 49178 5678 49181
rect 5730 49178 5786 49181
rect 5838 49178 5894 49181
rect 5946 49178 6002 49181
rect 6054 49178 6110 49181
rect 6162 49178 6218 49181
rect 6270 49178 6326 49181
rect 6378 49178 6434 49181
rect 6486 49178 6542 49181
rect 6594 49178 6650 49181
rect 6702 49178 6758 49181
rect 6810 49178 6866 49181
rect 6918 49178 6974 49181
rect 7026 49178 7082 49181
rect 7134 49178 7844 49181
rect 7896 49178 7952 49181
rect 8004 49178 8060 49181
rect 8112 49178 8168 49181
rect 8220 49178 8276 49181
rect 8328 49178 8384 49181
rect 8436 49178 8492 49181
rect 8544 49178 8600 49181
rect 8652 49178 8708 49181
rect 8760 49178 8816 49181
rect 8868 49178 8924 49181
rect 8976 49178 9032 49181
rect 9084 49178 9140 49181
rect 9192 49178 9248 49181
rect 9300 49178 9356 49181
rect 9408 49178 9464 49181
rect 9516 49178 9572 49181
rect 9624 49178 9680 49181
rect 9732 49178 9788 49181
rect 9840 49178 10253 49181
rect 10305 49178 10361 49181
rect 10413 49178 10469 49181
rect 10521 49178 10577 49181
rect 10629 49178 10685 49181
rect 10737 49178 10793 49181
rect 10845 49178 10901 49181
rect 10953 49178 11009 49181
rect 11061 49178 11117 49181
rect 11169 49178 11225 49181
rect 11277 49178 11333 49181
rect 11385 49178 11441 49181
rect 11493 49178 11549 49181
rect 11601 49178 11657 49181
rect 11709 49178 11765 49230
rect 3162 49122 11816 49178
rect 3213 49070 3269 49122
rect 3321 49070 3377 49122
rect 3429 49073 3485 49122
rect 3537 49073 3593 49122
rect 3645 49073 3701 49122
rect 3753 49073 3809 49122
rect 3861 49073 3917 49122
rect 3969 49073 4025 49122
rect 4077 49073 4133 49122
rect 4185 49073 4241 49122
rect 4293 49073 4349 49122
rect 4401 49073 4457 49122
rect 4509 49073 4565 49122
rect 4617 49073 4673 49122
rect 4725 49073 5138 49122
rect 5190 49073 5246 49122
rect 5298 49073 5354 49122
rect 5406 49073 5462 49122
rect 5514 49073 5570 49122
rect 5622 49073 5678 49122
rect 5730 49073 5786 49122
rect 5838 49073 5894 49122
rect 5946 49073 6002 49122
rect 6054 49073 6110 49122
rect 6162 49073 6218 49122
rect 6270 49073 6326 49122
rect 6378 49073 6434 49122
rect 6486 49073 6542 49122
rect 6594 49073 6650 49122
rect 6702 49073 6758 49122
rect 6810 49073 6866 49122
rect 6918 49073 6974 49122
rect 7026 49073 7082 49122
rect 7134 49073 7844 49122
rect 7896 49073 7952 49122
rect 8004 49073 8060 49122
rect 8112 49073 8168 49122
rect 8220 49073 8276 49122
rect 8328 49073 8384 49122
rect 8436 49073 8492 49122
rect 8544 49073 8600 49122
rect 8652 49073 8708 49122
rect 8760 49073 8816 49122
rect 8868 49073 8924 49122
rect 8976 49073 9032 49122
rect 9084 49073 9140 49122
rect 9192 49073 9248 49122
rect 9300 49073 9356 49122
rect 9408 49073 9464 49122
rect 9516 49073 9572 49122
rect 9624 49073 9680 49122
rect 9732 49073 9788 49122
rect 9840 49073 10253 49122
rect 10305 49073 10361 49122
rect 10413 49073 10469 49122
rect 10521 49073 10577 49122
rect 10629 49073 10685 49122
rect 10737 49073 10793 49122
rect 10845 49073 10901 49122
rect 10953 49073 11009 49122
rect 11061 49073 11117 49122
rect 11169 49073 11225 49122
rect 11277 49073 11333 49122
rect 11385 49073 11441 49122
rect 11493 49073 11549 49122
rect 11601 49070 11657 49122
rect 11709 49070 11765 49122
rect 3162 49042 3424 49070
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49070
rect 11554 49027 11662 49042
rect 3316 49016 11662 49027
rect 3316 48458 3327 49016
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48765 4871 48778
rect 4923 48765 4979 48778
rect 5031 48765 7247 48778
rect 7299 48765 7355 48778
rect 7407 48765 7463 48778
rect 7515 48765 7571 48778
rect 7623 48765 7679 48778
rect 7731 48765 9947 48778
rect 9999 48765 10055 48778
rect 10107 48765 11489 48778
rect 3489 48709 11489 48765
rect 3489 48696 4871 48709
rect 4923 48696 4979 48709
rect 5031 48696 7247 48709
rect 7299 48696 7355 48709
rect 7407 48696 7463 48709
rect 7515 48696 7571 48709
rect 7623 48696 7679 48709
rect 7731 48696 9947 48709
rect 9999 48696 10055 48709
rect 10107 48696 11489 48709
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
rect 11651 48458 11662 49016
rect 3316 48447 11662 48458
rect 3316 48432 3424 48447
rect 3162 48427 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48427 11816 48432
rect 3105 48375 3161 48376
rect 3213 48375 3269 48427
rect 3321 48375 3377 48427
rect 3429 48375 3485 48401
rect 3537 48375 3593 48401
rect 3645 48375 3701 48401
rect 3753 48375 3809 48401
rect 3861 48375 3917 48401
rect 3969 48375 4025 48401
rect 4077 48375 4133 48401
rect 4185 48375 4241 48401
rect 4293 48375 4349 48401
rect 4401 48375 4457 48401
rect 4509 48375 4565 48401
rect 4617 48375 4673 48401
rect 4725 48375 5138 48401
rect 5190 48375 5246 48401
rect 5298 48375 5354 48401
rect 5406 48375 5462 48401
rect 5514 48375 5570 48401
rect 5622 48375 5678 48401
rect 5730 48375 5786 48401
rect 5838 48375 5894 48401
rect 5946 48375 6002 48401
rect 6054 48375 6110 48401
rect 6162 48375 6218 48401
rect 6270 48375 6326 48401
rect 6378 48375 6434 48401
rect 6486 48375 6542 48401
rect 6594 48375 6650 48401
rect 6702 48375 6758 48401
rect 6810 48375 6866 48401
rect 6918 48375 6974 48401
rect 7026 48375 7082 48401
rect 7134 48375 7844 48401
rect 7896 48375 7952 48401
rect 8004 48375 8060 48401
rect 8112 48375 8168 48401
rect 8220 48375 8276 48401
rect 8328 48375 8384 48401
rect 8436 48375 8492 48401
rect 8544 48375 8600 48401
rect 8652 48375 8708 48401
rect 8760 48375 8816 48401
rect 8868 48375 8924 48401
rect 8976 48375 9032 48401
rect 9084 48375 9140 48401
rect 9192 48375 9248 48401
rect 9300 48375 9356 48401
rect 9408 48375 9464 48401
rect 9516 48375 9572 48401
rect 9624 48375 9680 48401
rect 9732 48375 9788 48401
rect 9840 48375 10253 48401
rect 10305 48375 10361 48401
rect 10413 48375 10469 48401
rect 10521 48375 10577 48401
rect 10629 48375 10685 48401
rect 10737 48375 10793 48401
rect 10845 48375 10901 48401
rect 10953 48375 11009 48401
rect 11061 48375 11117 48401
rect 11169 48375 11225 48401
rect 11277 48375 11333 48401
rect 11385 48375 11441 48401
rect 11493 48375 11549 48401
rect 11601 48375 11657 48427
rect 11709 48375 11765 48427
rect 11862 48376 11873 51900
rect 11817 48375 11873 48376
rect 3105 48319 11873 48375
rect 3105 48293 3161 48319
rect 3213 48293 3269 48319
rect 3321 48293 3377 48319
rect 3429 48293 3485 48319
rect 3537 48293 3593 48319
rect 3645 48293 3701 48319
rect 3753 48293 3809 48319
rect 3861 48293 3917 48319
rect 3969 48293 4025 48319
rect 4077 48293 4133 48319
rect 4185 48293 4241 48319
rect 4293 48293 4349 48319
rect 4401 48293 4457 48319
rect 4509 48293 4565 48319
rect 4617 48293 4673 48319
rect 4725 48293 5138 48319
rect 5190 48293 5246 48319
rect 5298 48293 5354 48319
rect 5406 48293 5462 48319
rect 5514 48293 5570 48319
rect 5622 48293 5678 48319
rect 5730 48293 5786 48319
rect 5838 48293 5894 48319
rect 5946 48293 6002 48319
rect 6054 48293 6110 48319
rect 6162 48293 6218 48319
rect 6270 48293 6326 48319
rect 6378 48293 6434 48319
rect 6486 48293 6542 48319
rect 6594 48293 6650 48319
rect 6702 48293 6758 48319
rect 6810 48293 6866 48319
rect 6918 48293 6974 48319
rect 7026 48293 7082 48319
rect 7134 48293 7844 48319
rect 7896 48293 7952 48319
rect 8004 48293 8060 48319
rect 8112 48293 8168 48319
rect 8220 48293 8276 48319
rect 8328 48293 8384 48319
rect 8436 48293 8492 48319
rect 8544 48293 8600 48319
rect 8652 48293 8708 48319
rect 8760 48293 8816 48319
rect 8868 48293 8924 48319
rect 8976 48293 9032 48319
rect 9084 48293 9140 48319
rect 9192 48293 9248 48319
rect 9300 48293 9356 48319
rect 9408 48293 9464 48319
rect 9516 48293 9572 48319
rect 9624 48293 9680 48319
rect 9732 48293 9788 48319
rect 9840 48293 10253 48319
rect 10305 48293 10361 48319
rect 10413 48293 10469 48319
rect 10521 48293 10577 48319
rect 10629 48293 10685 48319
rect 10737 48293 10793 48319
rect 10845 48293 10901 48319
rect 10953 48293 11009 48319
rect 11061 48293 11117 48319
rect 11169 48293 11225 48319
rect 11277 48293 11333 48319
rect 11385 48293 11441 48319
rect 11493 48293 11549 48319
rect 11601 48293 11657 48319
rect 11709 48293 11765 48319
rect 11817 48293 11873 48319
rect 3105 48247 3142 48293
rect 11836 48247 11873 48293
rect 3105 48236 11873 48247
rect 12059 48022 12070 52254
rect 2908 48011 12070 48022
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12427 52611
rect 2551 47654 12427 47665
rect 12753 52611 14907 52622
rect 12753 47665 12764 52611
rect 14710 52586 14907 52611
rect 14710 52574 14968 52586
rect 14710 52522 14904 52574
rect 14956 52522 14968 52574
rect 14710 52466 14968 52522
rect 14710 52414 14904 52466
rect 14956 52414 14968 52466
rect 14710 52358 14968 52414
rect 14710 52306 14904 52358
rect 14956 52306 14968 52358
rect 14710 52250 14968 52306
rect 14710 52198 14904 52250
rect 14956 52198 14968 52250
rect 14710 52142 14968 52198
rect 14710 52090 14904 52142
rect 14956 52090 14968 52142
rect 14710 52034 14968 52090
rect 14710 51982 14904 52034
rect 14956 51982 14968 52034
rect 14710 51926 14968 51982
rect 14710 51874 14904 51926
rect 14956 51874 14968 51926
rect 14710 51818 14968 51874
rect 14710 51766 14904 51818
rect 14956 51766 14968 51818
rect 14710 51710 14968 51766
rect 14710 51658 14904 51710
rect 14956 51658 14968 51710
rect 14710 51622 14968 51658
rect 14710 51422 14721 51622
rect 14892 51602 14968 51622
rect 14892 51550 14904 51602
rect 14956 51550 14968 51602
rect 14892 51494 14968 51550
rect 14892 51442 14904 51494
rect 14956 51442 14968 51494
rect 14892 51422 14968 51442
rect 14710 51386 14968 51422
rect 14710 51334 14904 51386
rect 14956 51334 14968 51386
rect 14710 51278 14968 51334
rect 14710 51226 14904 51278
rect 14956 51226 14968 51278
rect 14710 51214 14968 51226
rect 14710 50422 14907 51214
rect 14710 49854 14721 50422
rect 14710 49386 14907 49854
rect 14710 49374 14968 49386
rect 14710 49322 14904 49374
rect 14956 49322 14968 49374
rect 14710 49266 14968 49322
rect 14710 49214 14904 49266
rect 14956 49214 14968 49266
rect 14710 49158 14968 49214
rect 14710 49106 14904 49158
rect 14956 49106 14968 49158
rect 14710 49050 14968 49106
rect 14710 48998 14904 49050
rect 14956 48998 14968 49050
rect 14710 48942 14968 48998
rect 14710 48890 14904 48942
rect 14956 48890 14968 48942
rect 14710 48854 14968 48890
rect 14710 48654 14721 48854
rect 14892 48834 14968 48854
rect 14892 48782 14904 48834
rect 14956 48782 14968 48834
rect 14892 48726 14968 48782
rect 14892 48674 14904 48726
rect 14956 48674 14968 48726
rect 14892 48654 14968 48674
rect 14710 48618 14968 48654
rect 14710 48566 14904 48618
rect 14956 48566 14968 48618
rect 14710 48510 14968 48566
rect 14710 48458 14904 48510
rect 14956 48458 14968 48510
rect 14710 48402 14968 48458
rect 14710 48350 14904 48402
rect 14956 48350 14968 48402
rect 14710 48294 14968 48350
rect 14710 48242 14904 48294
rect 14956 48242 14968 48294
rect 14710 48186 14968 48242
rect 14710 48134 14904 48186
rect 14956 48134 14968 48186
rect 14710 48078 14968 48134
rect 14710 48026 14904 48078
rect 14956 48026 14968 48078
rect 14710 48014 14968 48026
rect 14710 47665 14907 48014
rect 12753 47654 14907 47665
rect 10 46174 86 46186
rect 10 46122 22 46174
rect 74 46122 86 46174
rect 10 46066 86 46122
rect 10 46014 22 46066
rect 74 46014 86 46066
rect 10 45958 86 46014
rect 10 45906 22 45958
rect 74 45906 86 45958
rect 10 45850 86 45906
rect 10 45798 22 45850
rect 74 45798 86 45850
rect 10 45742 86 45798
rect 10 45690 22 45742
rect 74 45690 86 45742
rect 10 45634 86 45690
rect 10 45582 22 45634
rect 74 45582 86 45634
rect 10 45526 86 45582
rect 10 45474 22 45526
rect 74 45474 86 45526
rect 10 45418 86 45474
rect 10 45366 22 45418
rect 74 45366 86 45418
rect 10 45310 86 45366
rect 10 45258 22 45310
rect 74 45258 86 45310
rect 10 45202 86 45258
rect 10 45150 22 45202
rect 74 45150 86 45202
rect 10 45094 86 45150
rect 10 45042 22 45094
rect 74 45042 86 45094
rect 10 44986 86 45042
rect 10 44934 22 44986
rect 74 44934 86 44986
rect 10 44878 86 44934
rect 10 44826 22 44878
rect 74 44826 86 44878
rect 10 44814 86 44826
rect 14892 46174 14968 46186
rect 14892 46122 14904 46174
rect 14956 46122 14968 46174
rect 14892 46066 14968 46122
rect 14892 46014 14904 46066
rect 14956 46014 14968 46066
rect 14892 45958 14968 46014
rect 14892 45906 14904 45958
rect 14956 45906 14968 45958
rect 14892 45850 14968 45906
rect 14892 45798 14904 45850
rect 14956 45798 14968 45850
rect 14892 45742 14968 45798
rect 14892 45690 14904 45742
rect 14956 45690 14968 45742
rect 14892 45634 14968 45690
rect 14892 45582 14904 45634
rect 14956 45582 14968 45634
rect 14892 45526 14968 45582
rect 14892 45474 14904 45526
rect 14956 45474 14968 45526
rect 14892 45418 14968 45474
rect 14892 45366 14904 45418
rect 14956 45366 14968 45418
rect 14892 45310 14968 45366
rect 14892 45258 14904 45310
rect 14956 45258 14968 45310
rect 14892 45202 14968 45258
rect 14892 45150 14904 45202
rect 14956 45150 14968 45202
rect 14892 45094 14968 45150
rect 14892 45042 14904 45094
rect 14956 45042 14968 45094
rect 14892 44986 14968 45042
rect 14892 44934 14904 44986
rect 14956 44934 14968 44986
rect 14892 44878 14968 44934
rect 14892 44826 14904 44878
rect 14956 44826 14968 44878
rect 14892 44814 14968 44826
rect 71 42647 725 42658
rect 71 41658 268 42647
rect 257 41458 268 41658
rect 71 40458 268 41458
rect 257 40258 268 40458
rect 71 39258 268 40258
rect 257 39058 268 39258
rect 71 38186 268 39058
rect 10 38174 268 38186
rect 10 38122 22 38174
rect 74 38122 268 38174
rect 10 38066 268 38122
rect 10 38014 22 38066
rect 74 38058 268 38066
rect 74 38014 86 38058
rect 10 37958 86 38014
rect 10 37906 22 37958
rect 74 37906 86 37958
rect 10 37858 86 37906
rect 257 37858 268 38058
rect 10 37850 268 37858
rect 10 37798 22 37850
rect 74 37798 268 37850
rect 10 37742 268 37798
rect 10 37690 22 37742
rect 74 37690 268 37742
rect 10 37634 268 37690
rect 10 37582 22 37634
rect 74 37582 268 37634
rect 10 37526 268 37582
rect 10 37474 22 37526
rect 74 37474 268 37526
rect 10 37418 268 37474
rect 10 37366 22 37418
rect 74 37366 268 37418
rect 10 37310 268 37366
rect 10 37258 22 37310
rect 74 37258 268 37310
rect 10 37202 268 37258
rect 10 37150 22 37202
rect 74 37150 268 37202
rect 10 37094 268 37150
rect 10 37042 22 37094
rect 74 37042 268 37094
rect 10 36986 268 37042
rect 10 36934 22 36986
rect 74 36934 268 36986
rect 10 36878 268 36934
rect 10 36826 22 36878
rect 74 36858 268 36878
rect 74 36826 86 36858
rect 10 36814 86 36826
rect 257 36658 268 36858
rect 71 36596 268 36658
rect 10 36584 268 36596
rect 10 36532 22 36584
rect 74 36532 268 36584
rect 10 36476 268 36532
rect 10 36424 22 36476
rect 74 36424 268 36476
rect 10 36368 268 36424
rect 10 36316 22 36368
rect 74 36316 268 36368
rect 10 36260 268 36316
rect 10 36208 22 36260
rect 74 36208 268 36260
rect 10 36152 268 36208
rect 10 36100 22 36152
rect 74 36100 268 36152
rect 10 36044 268 36100
rect 10 35992 22 36044
rect 74 35992 268 36044
rect 10 35936 268 35992
rect 10 35884 22 35936
rect 74 35884 268 35936
rect 10 35828 268 35884
rect 10 35776 22 35828
rect 74 35776 268 35828
rect 10 35720 268 35776
rect 10 35668 22 35720
rect 74 35668 268 35720
rect 10 35658 268 35668
rect 10 35612 86 35658
rect 10 35560 22 35612
rect 74 35560 86 35612
rect 10 35504 86 35560
rect 10 35452 22 35504
rect 74 35458 86 35504
rect 257 35458 268 35658
rect 74 35452 268 35458
rect 10 35396 268 35452
rect 10 35344 22 35396
rect 74 35344 268 35396
rect 10 35288 268 35344
rect 10 35236 22 35288
rect 74 35236 268 35288
rect 10 35180 268 35236
rect 10 35128 22 35180
rect 74 35128 268 35180
rect 10 35072 268 35128
rect 10 35020 22 35072
rect 74 35020 268 35072
rect 10 34964 268 35020
rect 10 34912 22 34964
rect 74 34912 268 34964
rect 10 34856 268 34912
rect 10 34804 22 34856
rect 74 34804 268 34856
rect 10 34748 268 34804
rect 10 34696 22 34748
rect 74 34696 268 34748
rect 10 34640 268 34696
rect 10 34588 22 34640
rect 74 34588 268 34640
rect 10 34532 268 34588
rect 10 34480 22 34532
rect 74 34480 268 34532
rect 10 34458 268 34480
rect 10 34424 86 34458
rect 10 34372 22 34424
rect 74 34372 86 34424
rect 10 34316 86 34372
rect 10 34264 22 34316
rect 74 34264 86 34316
rect 10 34258 86 34264
rect 257 34258 268 34458
rect 10 34208 268 34258
rect 10 34156 22 34208
rect 74 34156 268 34208
rect 10 34100 268 34156
rect 10 34048 22 34100
rect 74 34048 268 34100
rect 10 33992 268 34048
rect 10 33940 22 33992
rect 74 33940 268 33992
rect 10 33884 268 33940
rect 10 33832 22 33884
rect 74 33832 268 33884
rect 10 33776 268 33832
rect 10 33724 22 33776
rect 74 33724 268 33776
rect 10 33668 268 33724
rect 10 33616 22 33668
rect 74 33616 268 33668
rect 10 33604 268 33616
rect 71 33258 268 33604
rect 257 33058 268 33258
rect 71 32058 268 33058
rect 257 31858 268 32058
rect 71 30858 268 31858
rect 257 30658 268 30858
rect 71 29658 268 30658
rect 257 29458 268 29658
rect 71 28586 268 29458
rect 10 28574 268 28586
rect 10 28522 22 28574
rect 74 28522 268 28574
rect 10 28466 268 28522
rect 10 28414 22 28466
rect 74 28458 268 28466
rect 74 28414 86 28458
rect 10 28358 86 28414
rect 10 28306 22 28358
rect 74 28306 86 28358
rect 10 28258 86 28306
rect 257 28258 268 28458
rect 10 28250 268 28258
rect 10 28198 22 28250
rect 74 28198 268 28250
rect 10 28142 268 28198
rect 10 28090 22 28142
rect 74 28090 268 28142
rect 10 28034 268 28090
rect 10 27982 22 28034
rect 74 27982 268 28034
rect 10 27926 268 27982
rect 10 27874 22 27926
rect 74 27874 268 27926
rect 10 27818 268 27874
rect 10 27766 22 27818
rect 74 27766 268 27818
rect 10 27710 268 27766
rect 10 27658 22 27710
rect 74 27658 268 27710
rect 10 27602 268 27658
rect 10 27550 22 27602
rect 74 27550 268 27602
rect 10 27494 268 27550
rect 10 27442 22 27494
rect 74 27442 268 27494
rect 10 27386 268 27442
rect 10 27334 22 27386
rect 74 27334 268 27386
rect 10 27278 268 27334
rect 10 27226 22 27278
rect 74 27258 268 27278
rect 74 27226 86 27258
rect 10 27214 86 27226
rect 257 27058 268 27258
rect 71 26058 268 27058
rect 257 25858 268 26058
rect 71 24858 268 25858
rect 257 24658 268 24858
rect 71 23658 268 24658
rect 257 23458 268 23658
rect 71 22458 268 23458
rect 257 21390 268 22458
rect 71 20390 268 21390
rect 257 20190 268 20390
rect 71 19190 268 20190
rect 257 18990 268 19190
rect 71 17990 268 18990
rect 257 17790 268 17990
rect 71 16790 268 17790
rect 257 16590 268 16790
rect 71 15590 268 16590
rect 257 15390 268 15590
rect 71 14390 268 15390
rect 257 14190 268 14390
rect 71 14186 268 14190
rect 10 14174 268 14186
rect 10 14122 22 14174
rect 74 14122 268 14174
rect 10 14066 268 14122
rect 10 14014 22 14066
rect 74 14014 268 14066
rect 10 13958 268 14014
rect 10 13906 22 13958
rect 74 13906 268 13958
rect 10 13850 268 13906
rect 10 13798 22 13850
rect 74 13798 268 13850
rect 10 13742 268 13798
rect 10 13690 22 13742
rect 74 13690 268 13742
rect 10 13634 268 13690
rect 10 13582 22 13634
rect 74 13582 268 13634
rect 10 13526 268 13582
rect 10 13474 22 13526
rect 74 13474 268 13526
rect 10 13418 268 13474
rect 10 13366 22 13418
rect 74 13366 268 13418
rect 10 13310 268 13366
rect 10 13258 22 13310
rect 74 13258 268 13310
rect 10 13202 268 13258
rect 10 13150 22 13202
rect 74 13190 268 13202
rect 74 13150 86 13190
rect 10 13094 86 13150
rect 10 13042 22 13094
rect 74 13042 86 13094
rect 10 12990 86 13042
rect 257 12990 268 13190
rect 10 12986 268 12990
rect 10 12934 22 12986
rect 74 12934 268 12986
rect 10 12878 268 12934
rect 10 12826 22 12878
rect 74 12826 268 12878
rect 10 12814 268 12826
rect 71 11990 268 12814
rect 257 11790 268 11990
rect 71 10996 268 11790
rect 10 10984 268 10996
rect 10 10932 22 10984
rect 74 10932 268 10984
rect 10 10876 268 10932
rect 10 10824 22 10876
rect 74 10824 268 10876
rect 10 10790 268 10824
rect 10 10768 86 10790
rect 10 10716 22 10768
rect 74 10716 86 10768
rect 10 10660 86 10716
rect 10 10608 22 10660
rect 74 10608 86 10660
rect 10 10590 86 10608
rect 257 10590 268 10790
rect 10 10552 268 10590
rect 10 10500 22 10552
rect 74 10500 268 10552
rect 10 10444 268 10500
rect 10 10392 22 10444
rect 74 10392 268 10444
rect 10 10336 268 10392
rect 10 10284 22 10336
rect 74 10284 268 10336
rect 10 10228 268 10284
rect 10 10176 22 10228
rect 74 10176 268 10228
rect 10 10120 268 10176
rect 10 10068 22 10120
rect 74 10068 268 10120
rect 10 10012 268 10068
rect 10 9960 22 10012
rect 74 9960 268 10012
rect 10 9904 268 9960
rect 10 9852 22 9904
rect 74 9852 268 9904
rect 10 9796 268 9852
rect 10 9744 22 9796
rect 74 9744 268 9796
rect 10 9688 268 9744
rect 10 9636 22 9688
rect 74 9636 268 9688
rect 10 9590 268 9636
rect 10 9580 86 9590
rect 10 9528 22 9580
rect 74 9528 86 9580
rect 10 9472 86 9528
rect 10 9420 22 9472
rect 74 9420 86 9472
rect 10 9390 86 9420
rect 257 9390 268 9590
rect 10 9364 268 9390
rect 10 9312 22 9364
rect 74 9312 268 9364
rect 10 9256 268 9312
rect 10 9204 22 9256
rect 74 9204 268 9256
rect 10 9148 268 9204
rect 10 9096 22 9148
rect 74 9096 268 9148
rect 10 9040 268 9096
rect 10 8988 22 9040
rect 74 8988 268 9040
rect 10 8932 268 8988
rect 10 8880 22 8932
rect 74 8880 268 8932
rect 10 8824 268 8880
rect 10 8772 22 8824
rect 74 8772 268 8824
rect 10 8716 268 8772
rect 10 8664 22 8716
rect 74 8664 268 8716
rect 10 8608 268 8664
rect 10 8556 22 8608
rect 74 8556 268 8608
rect 10 8500 268 8556
rect 10 8448 22 8500
rect 74 8448 268 8500
rect 10 8392 268 8448
rect 10 8340 22 8392
rect 74 8390 268 8392
rect 74 8340 86 8390
rect 10 8284 86 8340
rect 10 8232 22 8284
rect 74 8232 86 8284
rect 10 8190 86 8232
rect 257 8190 268 8390
rect 10 8176 268 8190
rect 10 8124 22 8176
rect 74 8124 268 8176
rect 10 8068 268 8124
rect 10 8016 22 8068
rect 74 8016 268 8068
rect 10 8004 268 8016
rect 71 7796 268 8004
rect 10 7784 268 7796
rect 10 7732 22 7784
rect 74 7732 268 7784
rect 10 7676 268 7732
rect 10 7624 22 7676
rect 74 7624 268 7676
rect 10 7568 268 7624
rect 10 7516 22 7568
rect 74 7516 268 7568
rect 10 7460 268 7516
rect 10 7408 22 7460
rect 74 7408 268 7460
rect 10 7352 268 7408
rect 10 7300 22 7352
rect 74 7300 268 7352
rect 10 7244 268 7300
rect 10 7192 22 7244
rect 74 7192 268 7244
rect 10 7190 268 7192
rect 10 7136 86 7190
rect 10 7084 22 7136
rect 74 7084 86 7136
rect 10 7028 86 7084
rect 10 6976 22 7028
rect 74 6990 86 7028
rect 257 6990 268 7190
rect 74 6976 268 6990
rect 10 6920 268 6976
rect 10 6868 22 6920
rect 74 6868 268 6920
rect 10 6812 268 6868
rect 10 6760 22 6812
rect 74 6760 268 6812
rect 10 6704 268 6760
rect 10 6652 22 6704
rect 74 6652 268 6704
rect 10 6596 268 6652
rect 10 6544 22 6596
rect 74 6544 268 6596
rect 10 6488 268 6544
rect 10 6436 22 6488
rect 74 6436 268 6488
rect 10 6380 268 6436
rect 10 6328 22 6380
rect 74 6328 268 6380
rect 10 6272 268 6328
rect 10 6220 22 6272
rect 74 6220 268 6272
rect 10 6164 268 6220
rect 10 6112 22 6164
rect 74 6112 268 6164
rect 10 6056 268 6112
rect 10 6004 22 6056
rect 74 6004 268 6056
rect 10 5990 268 6004
rect 10 5948 86 5990
rect 10 5896 22 5948
rect 74 5896 86 5948
rect 10 5840 86 5896
rect 10 5788 22 5840
rect 74 5790 86 5840
rect 257 5790 268 5990
rect 74 5788 268 5790
rect 10 5732 268 5788
rect 10 5680 22 5732
rect 74 5680 268 5732
rect 10 5624 268 5680
rect 10 5572 22 5624
rect 74 5572 268 5624
rect 10 5516 268 5572
rect 10 5464 22 5516
rect 74 5464 268 5516
rect 10 5408 268 5464
rect 10 5356 22 5408
rect 74 5356 268 5408
rect 10 5300 268 5356
rect 10 5248 22 5300
rect 74 5248 268 5300
rect 10 5192 268 5248
rect 10 5140 22 5192
rect 74 5140 268 5192
rect 10 5084 268 5140
rect 10 5032 22 5084
rect 74 5032 268 5084
rect 10 4976 268 5032
rect 10 4924 22 4976
rect 74 4924 268 4976
rect 10 4868 268 4924
rect 10 4816 22 4868
rect 74 4816 268 4868
rect 10 4804 268 4816
rect 71 4790 268 4804
rect 10 4590 86 4596
rect 257 4590 268 4790
rect 10 4584 268 4590
rect 10 4532 22 4584
rect 74 4532 268 4584
rect 10 4476 268 4532
rect 10 4424 22 4476
rect 74 4424 268 4476
rect 10 4368 268 4424
rect 10 4316 22 4368
rect 74 4316 268 4368
rect 10 4260 268 4316
rect 10 4208 22 4260
rect 74 4208 268 4260
rect 10 4152 268 4208
rect 10 4100 22 4152
rect 74 4100 268 4152
rect 10 4044 268 4100
rect 10 3992 22 4044
rect 74 3992 268 4044
rect 10 3936 268 3992
rect 10 3884 22 3936
rect 74 3884 268 3936
rect 10 3828 268 3884
rect 10 3776 22 3828
rect 74 3776 268 3828
rect 10 3720 268 3776
rect 10 3668 22 3720
rect 74 3668 268 3720
rect 10 3612 268 3668
rect 10 3560 22 3612
rect 74 3590 268 3612
rect 74 3560 86 3590
rect 10 3504 86 3560
rect 10 3452 22 3504
rect 74 3452 86 3504
rect 10 3396 86 3452
rect 10 3344 22 3396
rect 74 3390 86 3396
rect 257 3390 268 3590
rect 74 3344 268 3390
rect 10 3288 268 3344
rect 10 3236 22 3288
rect 74 3236 268 3288
rect 10 3180 268 3236
rect 10 3128 22 3180
rect 74 3128 268 3180
rect 10 3072 268 3128
rect 10 3020 22 3072
rect 74 3020 268 3072
rect 10 2964 268 3020
rect 10 2912 22 2964
rect 74 2912 268 2964
rect 10 2856 268 2912
rect 10 2804 22 2856
rect 74 2804 268 2856
rect 10 2748 268 2804
rect 10 2696 22 2748
rect 74 2696 268 2748
rect 10 2640 268 2696
rect 10 2588 22 2640
rect 74 2588 268 2640
rect 10 2532 268 2588
rect 10 2480 22 2532
rect 74 2480 268 2532
rect 10 2424 268 2480
rect 10 2372 22 2424
rect 74 2390 268 2424
rect 74 2372 86 2390
rect 10 2316 86 2372
rect 10 2264 22 2316
rect 74 2264 86 2316
rect 10 2208 86 2264
rect 10 2156 22 2208
rect 74 2190 86 2208
rect 257 2190 268 2390
rect 74 2156 268 2190
rect 10 2100 268 2156
rect 10 2048 22 2100
rect 74 2048 268 2100
rect 10 1992 268 2048
rect 10 1940 22 1992
rect 74 1940 268 1992
rect 10 1884 268 1940
rect 10 1832 22 1884
rect 74 1832 268 1884
rect 10 1776 268 1832
rect 10 1724 22 1776
rect 74 1724 268 1776
rect 10 1668 268 1724
rect 10 1616 22 1668
rect 74 1616 268 1668
rect 10 1604 268 1616
rect 71 1201 268 1604
rect 714 1201 725 42647
rect 13012 42647 14907 42658
rect 13012 27201 13023 42647
rect 13969 41658 14264 42647
rect 13969 41458 13980 41658
rect 14253 41458 14264 41658
rect 13969 40458 14264 41458
rect 13969 40258 13980 40458
rect 14253 40258 14264 40458
rect 13969 39258 14264 40258
rect 13969 39058 13980 39258
rect 14253 39058 14264 39258
rect 13969 38058 14264 39058
rect 13969 37858 13980 38058
rect 14253 37858 14264 38058
rect 13969 36858 14264 37858
rect 13969 36658 13980 36858
rect 14253 36658 14264 36858
rect 13969 35658 14264 36658
rect 13969 35458 13980 35658
rect 14253 35458 14264 35658
rect 13969 34458 14264 35458
rect 13969 34258 13980 34458
rect 14253 34258 14264 34458
rect 13969 33258 14264 34258
rect 13969 33058 13980 33258
rect 14253 33058 14264 33258
rect 13969 32058 14264 33058
rect 13969 31858 13980 32058
rect 14253 31858 14264 32058
rect 13969 30858 14264 31858
rect 13969 30658 13980 30858
rect 14253 30658 14264 30858
rect 13969 29658 14264 30658
rect 13969 29458 13980 29658
rect 14253 29458 14264 29658
rect 13969 28458 14264 29458
rect 13969 28190 13980 28458
rect 14253 28190 14264 28458
rect 13969 27201 14264 28190
rect 13012 27190 14264 27201
rect 71 1190 725 1201
rect 14253 1201 14264 27190
rect 14710 41658 14907 42647
rect 14710 41458 14721 41658
rect 14710 40458 14907 41458
rect 14710 40258 14721 40458
rect 14710 39258 14907 40258
rect 14710 39058 14721 39258
rect 14710 38186 14907 39058
rect 14710 38174 14968 38186
rect 14710 38122 14904 38174
rect 14956 38122 14968 38174
rect 14710 38066 14968 38122
rect 14710 38058 14904 38066
rect 14710 37858 14721 38058
rect 14892 38014 14904 38058
rect 14956 38014 14968 38066
rect 14892 37958 14968 38014
rect 14892 37906 14904 37958
rect 14956 37906 14968 37958
rect 14892 37858 14968 37906
rect 14710 37850 14968 37858
rect 14710 37798 14904 37850
rect 14956 37798 14968 37850
rect 14710 37742 14968 37798
rect 14710 37690 14904 37742
rect 14956 37690 14968 37742
rect 14710 37634 14968 37690
rect 14710 37582 14904 37634
rect 14956 37582 14968 37634
rect 14710 37526 14968 37582
rect 14710 37474 14904 37526
rect 14956 37474 14968 37526
rect 14710 37418 14968 37474
rect 14710 37366 14904 37418
rect 14956 37366 14968 37418
rect 14710 37310 14968 37366
rect 14710 37258 14904 37310
rect 14956 37258 14968 37310
rect 14710 37202 14968 37258
rect 14710 37150 14904 37202
rect 14956 37150 14968 37202
rect 14710 37094 14968 37150
rect 14710 37042 14904 37094
rect 14956 37042 14968 37094
rect 14710 36986 14968 37042
rect 14710 36934 14904 36986
rect 14956 36934 14968 36986
rect 14710 36878 14968 36934
rect 14710 36858 14904 36878
rect 14710 36658 14721 36858
rect 14892 36826 14904 36858
rect 14956 36826 14968 36878
rect 14892 36814 14968 36826
rect 14710 36596 14907 36658
rect 14710 36584 14968 36596
rect 14710 36532 14904 36584
rect 14956 36532 14968 36584
rect 14710 36476 14968 36532
rect 14710 36424 14904 36476
rect 14956 36424 14968 36476
rect 14710 36368 14968 36424
rect 14710 36316 14904 36368
rect 14956 36316 14968 36368
rect 14710 36260 14968 36316
rect 14710 36208 14904 36260
rect 14956 36208 14968 36260
rect 14710 36152 14968 36208
rect 14710 36100 14904 36152
rect 14956 36100 14968 36152
rect 14710 36044 14968 36100
rect 14710 35992 14904 36044
rect 14956 35992 14968 36044
rect 14710 35936 14968 35992
rect 14710 35884 14904 35936
rect 14956 35884 14968 35936
rect 14710 35828 14968 35884
rect 14710 35776 14904 35828
rect 14956 35776 14968 35828
rect 14710 35720 14968 35776
rect 14710 35668 14904 35720
rect 14956 35668 14968 35720
rect 14710 35658 14968 35668
rect 14710 35458 14721 35658
rect 14892 35612 14968 35658
rect 14892 35560 14904 35612
rect 14956 35560 14968 35612
rect 14892 35504 14968 35560
rect 14892 35458 14904 35504
rect 14710 35452 14904 35458
rect 14956 35452 14968 35504
rect 14710 35396 14968 35452
rect 14710 35344 14904 35396
rect 14956 35344 14968 35396
rect 14710 35288 14968 35344
rect 14710 35236 14904 35288
rect 14956 35236 14968 35288
rect 14710 35180 14968 35236
rect 14710 35128 14904 35180
rect 14956 35128 14968 35180
rect 14710 35072 14968 35128
rect 14710 35020 14904 35072
rect 14956 35020 14968 35072
rect 14710 34964 14968 35020
rect 14710 34912 14904 34964
rect 14956 34912 14968 34964
rect 14710 34856 14968 34912
rect 14710 34804 14904 34856
rect 14956 34804 14968 34856
rect 14710 34748 14968 34804
rect 14710 34696 14904 34748
rect 14956 34696 14968 34748
rect 14710 34640 14968 34696
rect 14710 34588 14904 34640
rect 14956 34588 14968 34640
rect 14710 34532 14968 34588
rect 14710 34480 14904 34532
rect 14956 34480 14968 34532
rect 14710 34458 14968 34480
rect 14710 34258 14721 34458
rect 14892 34424 14968 34458
rect 14892 34372 14904 34424
rect 14956 34372 14968 34424
rect 14892 34316 14968 34372
rect 14892 34264 14904 34316
rect 14956 34264 14968 34316
rect 14892 34258 14968 34264
rect 14710 34208 14968 34258
rect 14710 34156 14904 34208
rect 14956 34156 14968 34208
rect 14710 34100 14968 34156
rect 14710 34048 14904 34100
rect 14956 34048 14968 34100
rect 14710 33992 14968 34048
rect 14710 33940 14904 33992
rect 14956 33940 14968 33992
rect 14710 33884 14968 33940
rect 14710 33832 14904 33884
rect 14956 33832 14968 33884
rect 14710 33776 14968 33832
rect 14710 33724 14904 33776
rect 14956 33724 14968 33776
rect 14710 33668 14968 33724
rect 14710 33616 14904 33668
rect 14956 33616 14968 33668
rect 14710 33604 14968 33616
rect 14710 33258 14907 33604
rect 14710 33058 14721 33258
rect 14710 32058 14907 33058
rect 14710 31858 14721 32058
rect 14710 30858 14907 31858
rect 14710 30658 14721 30858
rect 14710 29658 14907 30658
rect 14710 29458 14721 29658
rect 14710 28586 14907 29458
rect 14710 28574 14968 28586
rect 14710 28522 14904 28574
rect 14956 28522 14968 28574
rect 14710 28466 14968 28522
rect 14710 28458 14904 28466
rect 14710 28258 14721 28458
rect 14892 28414 14904 28458
rect 14956 28414 14968 28466
rect 14892 28358 14968 28414
rect 14892 28306 14904 28358
rect 14956 28306 14968 28358
rect 14892 28258 14968 28306
rect 14710 28250 14968 28258
rect 14710 28198 14904 28250
rect 14956 28198 14968 28250
rect 14710 28142 14968 28198
rect 14710 28090 14904 28142
rect 14956 28090 14968 28142
rect 14710 28034 14968 28090
rect 14710 27982 14904 28034
rect 14956 27982 14968 28034
rect 14710 27926 14968 27982
rect 14710 27874 14904 27926
rect 14956 27874 14968 27926
rect 14710 27818 14968 27874
rect 14710 27766 14904 27818
rect 14956 27766 14968 27818
rect 14710 27710 14968 27766
rect 14710 27658 14904 27710
rect 14956 27658 14968 27710
rect 14710 27602 14968 27658
rect 14710 27550 14904 27602
rect 14956 27550 14968 27602
rect 14710 27494 14968 27550
rect 14710 27442 14904 27494
rect 14956 27442 14968 27494
rect 14710 27386 14968 27442
rect 14710 27334 14904 27386
rect 14956 27334 14968 27386
rect 14710 27278 14968 27334
rect 14710 27258 14904 27278
rect 14710 27058 14721 27258
rect 14892 27226 14904 27258
rect 14956 27226 14968 27278
rect 14892 27214 14968 27226
rect 14710 26058 14907 27058
rect 14710 25858 14721 26058
rect 14710 24858 14907 25858
rect 14710 24658 14721 24858
rect 14710 23658 14907 24658
rect 14710 23458 14721 23658
rect 14710 22458 14907 23458
rect 14710 21390 14721 22458
rect 14710 20390 14907 21390
rect 14710 20190 14721 20390
rect 14710 19190 14907 20190
rect 14710 18990 14721 19190
rect 14710 17990 14907 18990
rect 14710 17790 14721 17990
rect 14710 16790 14907 17790
rect 14710 16590 14721 16790
rect 14710 15590 14907 16590
rect 14710 15390 14721 15590
rect 14710 14390 14907 15390
rect 14710 14190 14721 14390
rect 14710 14186 14907 14190
rect 14710 14174 14968 14186
rect 14710 14122 14904 14174
rect 14956 14122 14968 14174
rect 14710 14066 14968 14122
rect 14710 14014 14904 14066
rect 14956 14014 14968 14066
rect 14710 13958 14968 14014
rect 14710 13906 14904 13958
rect 14956 13906 14968 13958
rect 14710 13850 14968 13906
rect 14710 13798 14904 13850
rect 14956 13798 14968 13850
rect 14710 13742 14968 13798
rect 14710 13690 14904 13742
rect 14956 13690 14968 13742
rect 14710 13634 14968 13690
rect 14710 13582 14904 13634
rect 14956 13582 14968 13634
rect 14710 13526 14968 13582
rect 14710 13474 14904 13526
rect 14956 13474 14968 13526
rect 14710 13418 14968 13474
rect 14710 13366 14904 13418
rect 14956 13366 14968 13418
rect 14710 13310 14968 13366
rect 14710 13258 14904 13310
rect 14956 13258 14968 13310
rect 14710 13202 14968 13258
rect 14710 13190 14904 13202
rect 14710 12990 14721 13190
rect 14892 13150 14904 13190
rect 14956 13150 14968 13202
rect 14892 13094 14968 13150
rect 14892 13042 14904 13094
rect 14956 13042 14968 13094
rect 14892 12990 14968 13042
rect 14710 12986 14968 12990
rect 14710 12934 14904 12986
rect 14956 12934 14968 12986
rect 14710 12878 14968 12934
rect 14710 12826 14904 12878
rect 14956 12826 14968 12878
rect 14710 12814 14968 12826
rect 14710 11990 14907 12814
rect 14710 11790 14721 11990
rect 14710 10996 14907 11790
rect 14710 10984 14968 10996
rect 14710 10932 14904 10984
rect 14956 10932 14968 10984
rect 14710 10876 14968 10932
rect 14710 10824 14904 10876
rect 14956 10824 14968 10876
rect 14710 10790 14968 10824
rect 14710 10590 14721 10790
rect 14892 10768 14968 10790
rect 14892 10716 14904 10768
rect 14956 10716 14968 10768
rect 14892 10660 14968 10716
rect 14892 10608 14904 10660
rect 14956 10608 14968 10660
rect 14892 10590 14968 10608
rect 14710 10552 14968 10590
rect 14710 10500 14904 10552
rect 14956 10500 14968 10552
rect 14710 10444 14968 10500
rect 14710 10392 14904 10444
rect 14956 10392 14968 10444
rect 14710 10336 14968 10392
rect 14710 10284 14904 10336
rect 14956 10284 14968 10336
rect 14710 10228 14968 10284
rect 14710 10176 14904 10228
rect 14956 10176 14968 10228
rect 14710 10120 14968 10176
rect 14710 10068 14904 10120
rect 14956 10068 14968 10120
rect 14710 10012 14968 10068
rect 14710 9960 14904 10012
rect 14956 9960 14968 10012
rect 14710 9904 14968 9960
rect 14710 9852 14904 9904
rect 14956 9852 14968 9904
rect 14710 9796 14968 9852
rect 14710 9744 14904 9796
rect 14956 9744 14968 9796
rect 14710 9688 14968 9744
rect 14710 9636 14904 9688
rect 14956 9636 14968 9688
rect 14710 9590 14968 9636
rect 14710 9390 14721 9590
rect 14892 9580 14968 9590
rect 14892 9528 14904 9580
rect 14956 9528 14968 9580
rect 14892 9472 14968 9528
rect 14892 9420 14904 9472
rect 14956 9420 14968 9472
rect 14892 9390 14968 9420
rect 14710 9364 14968 9390
rect 14710 9312 14904 9364
rect 14956 9312 14968 9364
rect 14710 9256 14968 9312
rect 14710 9204 14904 9256
rect 14956 9204 14968 9256
rect 14710 9148 14968 9204
rect 14710 9096 14904 9148
rect 14956 9096 14968 9148
rect 14710 9040 14968 9096
rect 14710 8988 14904 9040
rect 14956 8988 14968 9040
rect 14710 8932 14968 8988
rect 14710 8880 14904 8932
rect 14956 8880 14968 8932
rect 14710 8824 14968 8880
rect 14710 8772 14904 8824
rect 14956 8772 14968 8824
rect 14710 8716 14968 8772
rect 14710 8664 14904 8716
rect 14956 8664 14968 8716
rect 14710 8608 14968 8664
rect 14710 8556 14904 8608
rect 14956 8556 14968 8608
rect 14710 8500 14968 8556
rect 14710 8448 14904 8500
rect 14956 8448 14968 8500
rect 14710 8392 14968 8448
rect 14710 8390 14904 8392
rect 14710 8190 14721 8390
rect 14892 8340 14904 8390
rect 14956 8340 14968 8392
rect 14892 8284 14968 8340
rect 14892 8232 14904 8284
rect 14956 8232 14968 8284
rect 14892 8190 14968 8232
rect 14710 8176 14968 8190
rect 14710 8124 14904 8176
rect 14956 8124 14968 8176
rect 14710 8068 14968 8124
rect 14710 8016 14904 8068
rect 14956 8016 14968 8068
rect 14710 8004 14968 8016
rect 14710 7796 14907 8004
rect 14710 7784 14968 7796
rect 14710 7732 14904 7784
rect 14956 7732 14968 7784
rect 14710 7676 14968 7732
rect 14710 7624 14904 7676
rect 14956 7624 14968 7676
rect 14710 7568 14968 7624
rect 14710 7516 14904 7568
rect 14956 7516 14968 7568
rect 14710 7460 14968 7516
rect 14710 7408 14904 7460
rect 14956 7408 14968 7460
rect 14710 7352 14968 7408
rect 14710 7300 14904 7352
rect 14956 7300 14968 7352
rect 14710 7244 14968 7300
rect 14710 7192 14904 7244
rect 14956 7192 14968 7244
rect 14710 7190 14968 7192
rect 14710 6990 14721 7190
rect 14892 7136 14968 7190
rect 14892 7084 14904 7136
rect 14956 7084 14968 7136
rect 14892 7028 14968 7084
rect 14892 6990 14904 7028
rect 14710 6976 14904 6990
rect 14956 6976 14968 7028
rect 14710 6920 14968 6976
rect 14710 6868 14904 6920
rect 14956 6868 14968 6920
rect 14710 6812 14968 6868
rect 14710 6760 14904 6812
rect 14956 6760 14968 6812
rect 14710 6704 14968 6760
rect 14710 6652 14904 6704
rect 14956 6652 14968 6704
rect 14710 6596 14968 6652
rect 14710 6544 14904 6596
rect 14956 6544 14968 6596
rect 14710 6488 14968 6544
rect 14710 6436 14904 6488
rect 14956 6436 14968 6488
rect 14710 6380 14968 6436
rect 14710 6328 14904 6380
rect 14956 6328 14968 6380
rect 14710 6272 14968 6328
rect 14710 6220 14904 6272
rect 14956 6220 14968 6272
rect 14710 6164 14968 6220
rect 14710 6112 14904 6164
rect 14956 6112 14968 6164
rect 14710 6056 14968 6112
rect 14710 6004 14904 6056
rect 14956 6004 14968 6056
rect 14710 5990 14968 6004
rect 14710 5790 14721 5990
rect 14892 5948 14968 5990
rect 14892 5896 14904 5948
rect 14956 5896 14968 5948
rect 14892 5840 14968 5896
rect 14892 5790 14904 5840
rect 14710 5788 14904 5790
rect 14956 5788 14968 5840
rect 14710 5732 14968 5788
rect 14710 5680 14904 5732
rect 14956 5680 14968 5732
rect 14710 5624 14968 5680
rect 14710 5572 14904 5624
rect 14956 5572 14968 5624
rect 14710 5516 14968 5572
rect 14710 5464 14904 5516
rect 14956 5464 14968 5516
rect 14710 5408 14968 5464
rect 14710 5356 14904 5408
rect 14956 5356 14968 5408
rect 14710 5300 14968 5356
rect 14710 5248 14904 5300
rect 14956 5248 14968 5300
rect 14710 5192 14968 5248
rect 14710 5140 14904 5192
rect 14956 5140 14968 5192
rect 14710 5084 14968 5140
rect 14710 5032 14904 5084
rect 14956 5032 14968 5084
rect 14710 4976 14968 5032
rect 14710 4924 14904 4976
rect 14956 4924 14968 4976
rect 14710 4868 14968 4924
rect 14710 4816 14904 4868
rect 14956 4816 14968 4868
rect 14710 4804 14968 4816
rect 14710 4790 14907 4804
rect 14710 4590 14721 4790
rect 14892 4590 14968 4596
rect 14710 4584 14968 4590
rect 14710 4532 14904 4584
rect 14956 4532 14968 4584
rect 14710 4476 14968 4532
rect 14710 4424 14904 4476
rect 14956 4424 14968 4476
rect 14710 4368 14968 4424
rect 14710 4316 14904 4368
rect 14956 4316 14968 4368
rect 14710 4260 14968 4316
rect 14710 4208 14904 4260
rect 14956 4208 14968 4260
rect 14710 4152 14968 4208
rect 14710 4100 14904 4152
rect 14956 4100 14968 4152
rect 14710 4044 14968 4100
rect 14710 3992 14904 4044
rect 14956 3992 14968 4044
rect 14710 3936 14968 3992
rect 14710 3884 14904 3936
rect 14956 3884 14968 3936
rect 14710 3828 14968 3884
rect 14710 3776 14904 3828
rect 14956 3776 14968 3828
rect 14710 3720 14968 3776
rect 14710 3668 14904 3720
rect 14956 3668 14968 3720
rect 14710 3612 14968 3668
rect 14710 3590 14904 3612
rect 14710 3390 14721 3590
rect 14892 3560 14904 3590
rect 14956 3560 14968 3612
rect 14892 3504 14968 3560
rect 14892 3452 14904 3504
rect 14956 3452 14968 3504
rect 14892 3396 14968 3452
rect 14892 3390 14904 3396
rect 14710 3344 14904 3390
rect 14956 3344 14968 3396
rect 14710 3288 14968 3344
rect 14710 3236 14904 3288
rect 14956 3236 14968 3288
rect 14710 3180 14968 3236
rect 14710 3128 14904 3180
rect 14956 3128 14968 3180
rect 14710 3072 14968 3128
rect 14710 3020 14904 3072
rect 14956 3020 14968 3072
rect 14710 2964 14968 3020
rect 14710 2912 14904 2964
rect 14956 2912 14968 2964
rect 14710 2856 14968 2912
rect 14710 2804 14904 2856
rect 14956 2804 14968 2856
rect 14710 2748 14968 2804
rect 14710 2696 14904 2748
rect 14956 2696 14968 2748
rect 14710 2640 14968 2696
rect 14710 2588 14904 2640
rect 14956 2588 14968 2640
rect 14710 2532 14968 2588
rect 14710 2480 14904 2532
rect 14956 2480 14968 2532
rect 14710 2424 14968 2480
rect 14710 2390 14904 2424
rect 14710 2190 14721 2390
rect 14892 2372 14904 2390
rect 14956 2372 14968 2424
rect 14892 2316 14968 2372
rect 14892 2264 14904 2316
rect 14956 2264 14968 2316
rect 14892 2208 14968 2264
rect 14892 2190 14904 2208
rect 14710 2156 14904 2190
rect 14956 2156 14968 2208
rect 14710 2100 14968 2156
rect 14710 2048 14904 2100
rect 14956 2048 14968 2100
rect 14710 1992 14968 2048
rect 14710 1940 14904 1992
rect 14956 1940 14968 1992
rect 14710 1884 14968 1940
rect 14710 1832 14904 1884
rect 14956 1832 14968 1884
rect 14710 1776 14968 1832
rect 14710 1724 14904 1776
rect 14956 1724 14968 1776
rect 14710 1668 14968 1724
rect 14710 1616 14904 1668
rect 14956 1616 14968 1668
rect 14710 1604 14968 1616
rect 14710 1201 14907 1604
rect 14253 1190 14907 1201
rect 309 818 2113 830
rect 309 766 321 818
rect 373 766 429 818
rect 481 766 537 818
rect 589 766 645 818
rect 697 766 753 818
rect 805 766 861 818
rect 913 766 969 818
rect 1021 766 1077 818
rect 1129 766 1185 818
rect 1237 766 1293 818
rect 1345 766 1401 818
rect 1453 766 1509 818
rect 1561 766 1617 818
rect 1669 766 1725 818
rect 1777 766 1833 818
rect 1885 766 1941 818
rect 1993 766 2049 818
rect 2101 766 2113 818
rect 309 754 2113 766
rect 2864 818 4668 830
rect 2864 766 2876 818
rect 2928 766 2984 818
rect 3036 766 3092 818
rect 3144 766 3200 818
rect 3252 766 3308 818
rect 3360 766 3416 818
rect 3468 766 3524 818
rect 3576 766 3632 818
rect 3684 766 3740 818
rect 3792 766 3848 818
rect 3900 766 3956 818
rect 4008 766 4064 818
rect 4116 766 4172 818
rect 4224 766 4280 818
rect 4332 766 4388 818
rect 4440 766 4496 818
rect 4548 766 4604 818
rect 4656 766 4668 818
rect 2864 754 4668 766
rect 5234 818 7038 830
rect 5234 766 5246 818
rect 5298 766 5354 818
rect 5406 766 5462 818
rect 5514 766 5570 818
rect 5622 766 5678 818
rect 5730 766 5786 818
rect 5838 766 5894 818
rect 5946 766 6002 818
rect 6054 766 6110 818
rect 6162 766 6218 818
rect 6270 766 6326 818
rect 6378 766 6434 818
rect 6486 766 6542 818
rect 6594 766 6650 818
rect 6702 766 6758 818
rect 6810 766 6866 818
rect 6918 766 6974 818
rect 7026 766 7038 818
rect 5234 754 7038 766
rect 7940 818 9744 830
rect 7940 766 7952 818
rect 8004 766 8060 818
rect 8112 766 8168 818
rect 8220 766 8276 818
rect 8328 766 8384 818
rect 8436 766 8492 818
rect 8544 766 8600 818
rect 8652 766 8708 818
rect 8760 766 8816 818
rect 8868 766 8924 818
rect 8976 766 9032 818
rect 9084 766 9140 818
rect 9192 766 9248 818
rect 9300 766 9356 818
rect 9408 766 9464 818
rect 9516 766 9572 818
rect 9624 766 9680 818
rect 9732 766 9744 818
rect 7940 754 9744 766
rect 10310 818 12114 830
rect 10310 766 10322 818
rect 10374 766 10430 818
rect 10482 766 10538 818
rect 10590 766 10646 818
rect 10698 766 10754 818
rect 10806 766 10862 818
rect 10914 766 10970 818
rect 11022 766 11078 818
rect 11130 766 11186 818
rect 11238 766 11294 818
rect 11346 766 11402 818
rect 11454 766 11510 818
rect 11562 766 11618 818
rect 11670 766 11726 818
rect 11778 766 11834 818
rect 11886 766 11942 818
rect 11994 766 12050 818
rect 12102 766 12114 818
rect 10310 754 12114 766
rect 12865 818 14669 830
rect 12865 766 12877 818
rect 12929 766 12985 818
rect 13037 766 13093 818
rect 13145 766 13201 818
rect 13253 766 13309 818
rect 13361 766 13417 818
rect 13469 766 13525 818
rect 13577 766 13633 818
rect 13685 766 13741 818
rect 13793 766 13849 818
rect 13901 766 13957 818
rect 14009 766 14065 818
rect 14117 766 14173 818
rect 14225 766 14281 818
rect 14333 766 14389 818
rect 14441 766 14497 818
rect 14549 766 14605 818
rect 14657 766 14669 818
rect 12865 754 14669 766
<< via1 >>
rect 321 57447 373 57499
rect 429 57447 481 57499
rect 537 57447 589 57499
rect 645 57447 697 57499
rect 753 57447 805 57499
rect 861 57447 913 57499
rect 969 57447 1021 57499
rect 1077 57447 1129 57499
rect 1185 57447 1237 57499
rect 1293 57447 1345 57499
rect 1401 57447 1453 57499
rect 1509 57447 1561 57499
rect 1617 57447 1669 57499
rect 1725 57447 1777 57499
rect 1833 57447 1885 57499
rect 1941 57447 1993 57499
rect 2049 57447 2101 57499
rect 2876 57447 2928 57499
rect 2984 57447 3036 57499
rect 3092 57447 3144 57499
rect 3200 57447 3252 57499
rect 3308 57447 3360 57499
rect 3416 57447 3468 57499
rect 3524 57447 3576 57499
rect 3632 57447 3684 57499
rect 3740 57447 3792 57499
rect 3848 57447 3900 57499
rect 3956 57447 4008 57499
rect 4064 57447 4116 57499
rect 4172 57447 4224 57499
rect 4280 57447 4332 57499
rect 4388 57447 4440 57499
rect 4496 57447 4548 57499
rect 4604 57447 4656 57499
rect 5246 57447 5298 57499
rect 5354 57447 5406 57499
rect 5462 57447 5514 57499
rect 5570 57447 5622 57499
rect 5678 57447 5730 57499
rect 5786 57447 5838 57499
rect 5894 57447 5946 57499
rect 6002 57447 6054 57499
rect 6110 57447 6162 57499
rect 6218 57447 6270 57499
rect 6326 57447 6378 57499
rect 6434 57447 6486 57499
rect 6542 57447 6594 57499
rect 6650 57447 6702 57499
rect 6758 57447 6810 57499
rect 6866 57447 6918 57499
rect 6974 57447 7026 57499
rect 7952 57447 8004 57499
rect 8060 57447 8112 57499
rect 8168 57447 8220 57499
rect 8276 57447 8328 57499
rect 8384 57447 8436 57499
rect 8492 57447 8544 57499
rect 8600 57447 8652 57499
rect 8708 57447 8760 57499
rect 8816 57447 8868 57499
rect 8924 57447 8976 57499
rect 9032 57447 9084 57499
rect 9140 57447 9192 57499
rect 9248 57447 9300 57499
rect 9356 57447 9408 57499
rect 9464 57447 9516 57499
rect 9572 57447 9624 57499
rect 9680 57447 9732 57499
rect 10322 57447 10374 57499
rect 10430 57447 10482 57499
rect 10538 57447 10590 57499
rect 10646 57447 10698 57499
rect 10754 57447 10806 57499
rect 10862 57447 10914 57499
rect 10970 57447 11022 57499
rect 11078 57447 11130 57499
rect 11186 57447 11238 57499
rect 11294 57447 11346 57499
rect 11402 57447 11454 57499
rect 11510 57447 11562 57499
rect 11618 57447 11670 57499
rect 11726 57447 11778 57499
rect 11834 57447 11886 57499
rect 11942 57447 11994 57499
rect 12050 57447 12102 57499
rect 12877 57447 12929 57499
rect 12985 57447 13037 57499
rect 13093 57447 13145 57499
rect 13201 57447 13253 57499
rect 13309 57447 13361 57499
rect 13417 57447 13469 57499
rect 13525 57447 13577 57499
rect 13633 57447 13685 57499
rect 13741 57447 13793 57499
rect 13849 57447 13901 57499
rect 13957 57447 14009 57499
rect 14065 57447 14117 57499
rect 14173 57447 14225 57499
rect 14281 57447 14333 57499
rect 14389 57447 14441 57499
rect 14497 57447 14549 57499
rect 14605 57447 14657 57499
rect 22 57207 74 57259
rect 22 57099 74 57151
rect 14904 57207 14956 57259
rect 22 56991 74 57043
rect 22 56883 74 56935
rect 22 56775 74 56827
rect 22 56667 74 56719
rect 22 56559 74 56611
rect 22 56451 74 56503
rect 22 56343 74 56395
rect 22 56235 74 56287
rect 22 56127 74 56179
rect 22 56019 74 56071
rect 22 54122 74 54174
rect 22 54014 74 54066
rect 22 53906 74 53958
rect 22 53798 74 53850
rect 22 53690 74 53742
rect 22 53582 74 53634
rect 22 53474 74 53526
rect 22 53366 74 53418
rect 22 53258 74 53310
rect 22 53150 74 53202
rect 375 57052 402 57104
rect 402 57052 427 57104
rect 483 57059 510 57104
rect 510 57059 535 57104
rect 591 57059 643 57104
rect 699 57059 751 57104
rect 807 57059 859 57104
rect 915 57059 967 57104
rect 1023 57059 1075 57104
rect 1131 57059 1183 57104
rect 1239 57059 1291 57104
rect 1347 57059 1399 57104
rect 1455 57059 1507 57104
rect 1563 57059 1615 57104
rect 1671 57059 1723 57104
rect 1779 57059 1831 57104
rect 1887 57059 1939 57104
rect 1995 57059 2047 57104
rect 2768 57059 2820 57104
rect 2876 57059 2928 57104
rect 2984 57059 3036 57104
rect 3092 57059 3144 57104
rect 3200 57059 3252 57104
rect 3308 57059 3360 57104
rect 3416 57059 3468 57104
rect 3524 57059 3576 57104
rect 3632 57059 3684 57104
rect 3740 57059 3792 57104
rect 3848 57059 3900 57104
rect 3956 57059 4008 57104
rect 4064 57059 4116 57104
rect 4172 57059 4224 57104
rect 4280 57059 4332 57104
rect 4388 57059 4440 57104
rect 4496 57059 4548 57104
rect 4604 57059 4656 57104
rect 4712 57059 4764 57104
rect 5138 57059 5190 57104
rect 5246 57059 5298 57104
rect 5354 57059 5406 57104
rect 5462 57059 5514 57104
rect 5570 57059 5622 57104
rect 5678 57059 5730 57104
rect 5786 57059 5838 57104
rect 5894 57059 5946 57104
rect 6002 57059 6054 57104
rect 6110 57059 6162 57104
rect 6218 57059 6270 57104
rect 6326 57059 6378 57104
rect 6434 57059 6486 57104
rect 6542 57059 6594 57104
rect 6650 57059 6702 57104
rect 6758 57059 6810 57104
rect 6866 57059 6918 57104
rect 6974 57059 7026 57104
rect 7082 57059 7134 57104
rect 7844 57059 7896 57104
rect 7952 57059 8004 57104
rect 8060 57059 8112 57104
rect 8168 57059 8220 57104
rect 8276 57059 8328 57104
rect 8384 57059 8436 57104
rect 8492 57059 8544 57104
rect 8600 57059 8652 57104
rect 8708 57059 8760 57104
rect 8816 57059 8868 57104
rect 8924 57059 8976 57104
rect 9032 57059 9084 57104
rect 9140 57059 9192 57104
rect 9248 57059 9300 57104
rect 9356 57059 9408 57104
rect 9464 57059 9516 57104
rect 9572 57059 9624 57104
rect 9680 57059 9732 57104
rect 9788 57059 9840 57104
rect 10214 57059 10266 57104
rect 10322 57059 10374 57104
rect 10430 57059 10482 57104
rect 10538 57059 10590 57104
rect 10646 57059 10698 57104
rect 10754 57059 10806 57104
rect 10862 57059 10914 57104
rect 10970 57059 11022 57104
rect 11078 57059 11130 57104
rect 11186 57059 11238 57104
rect 11294 57059 11346 57104
rect 11402 57059 11454 57104
rect 11510 57059 11562 57104
rect 11618 57059 11670 57104
rect 11726 57059 11778 57104
rect 11834 57059 11886 57104
rect 11942 57059 11994 57104
rect 12050 57059 12102 57104
rect 12158 57059 12210 57104
rect 12931 57059 12983 57104
rect 13039 57059 13091 57104
rect 13147 57059 13199 57104
rect 13255 57059 13307 57104
rect 13363 57059 13415 57104
rect 13471 57059 13523 57104
rect 13579 57059 13631 57104
rect 13687 57059 13739 57104
rect 13795 57059 13847 57104
rect 13903 57059 13955 57104
rect 14011 57059 14063 57104
rect 14119 57059 14171 57104
rect 14227 57059 14279 57104
rect 14335 57059 14387 57104
rect 14443 57059 14468 57104
rect 14468 57059 14495 57104
rect 483 57052 535 57059
rect 591 57052 643 57059
rect 699 57052 751 57059
rect 807 57052 859 57059
rect 915 57052 967 57059
rect 1023 57052 1075 57059
rect 1131 57052 1183 57059
rect 1239 57052 1291 57059
rect 1347 57052 1399 57059
rect 1455 57052 1507 57059
rect 1563 57052 1615 57059
rect 1671 57052 1723 57059
rect 1779 57052 1831 57059
rect 1887 57052 1939 57059
rect 1995 57052 2047 57059
rect 2768 57052 2820 57059
rect 2876 57052 2928 57059
rect 2984 57052 3036 57059
rect 3092 57052 3144 57059
rect 3200 57052 3252 57059
rect 3308 57052 3360 57059
rect 3416 57052 3468 57059
rect 3524 57052 3576 57059
rect 3632 57052 3684 57059
rect 3740 57052 3792 57059
rect 3848 57052 3900 57059
rect 3956 57052 4008 57059
rect 4064 57052 4116 57059
rect 4172 57052 4224 57059
rect 4280 57052 4332 57059
rect 4388 57052 4440 57059
rect 4496 57052 4548 57059
rect 4604 57052 4656 57059
rect 4712 57052 4764 57059
rect 5138 57052 5190 57059
rect 5246 57052 5298 57059
rect 5354 57052 5406 57059
rect 5462 57052 5514 57059
rect 5570 57052 5622 57059
rect 5678 57052 5730 57059
rect 5786 57052 5838 57059
rect 5894 57052 5946 57059
rect 6002 57052 6054 57059
rect 6110 57052 6162 57059
rect 6218 57052 6270 57059
rect 6326 57052 6378 57059
rect 6434 57052 6486 57059
rect 6542 57052 6594 57059
rect 6650 57052 6702 57059
rect 6758 57052 6810 57059
rect 6866 57052 6918 57059
rect 6974 57052 7026 57059
rect 7082 57052 7134 57059
rect 7844 57052 7896 57059
rect 7952 57052 8004 57059
rect 8060 57052 8112 57059
rect 8168 57052 8220 57059
rect 8276 57052 8328 57059
rect 8384 57052 8436 57059
rect 8492 57052 8544 57059
rect 8600 57052 8652 57059
rect 8708 57052 8760 57059
rect 8816 57052 8868 57059
rect 8924 57052 8976 57059
rect 9032 57052 9084 57059
rect 9140 57052 9192 57059
rect 9248 57052 9300 57059
rect 9356 57052 9408 57059
rect 9464 57052 9516 57059
rect 9572 57052 9624 57059
rect 9680 57052 9732 57059
rect 9788 57052 9840 57059
rect 10214 57052 10266 57059
rect 10322 57052 10374 57059
rect 10430 57052 10482 57059
rect 10538 57052 10590 57059
rect 10646 57052 10698 57059
rect 10754 57052 10806 57059
rect 10862 57052 10914 57059
rect 10970 57052 11022 57059
rect 11078 57052 11130 57059
rect 11186 57052 11238 57059
rect 11294 57052 11346 57059
rect 11402 57052 11454 57059
rect 11510 57052 11562 57059
rect 11618 57052 11670 57059
rect 11726 57052 11778 57059
rect 11834 57052 11886 57059
rect 11942 57052 11994 57059
rect 12050 57052 12102 57059
rect 12158 57052 12210 57059
rect 12931 57052 12983 57059
rect 13039 57052 13091 57059
rect 13147 57052 13199 57059
rect 13255 57052 13307 57059
rect 13363 57052 13415 57059
rect 13471 57052 13523 57059
rect 13579 57052 13631 57059
rect 13687 57052 13739 57059
rect 13795 57052 13847 57059
rect 13903 57052 13955 57059
rect 14011 57052 14063 57059
rect 14119 57052 14171 57059
rect 14227 57052 14279 57059
rect 14335 57052 14387 57059
rect 14443 57052 14495 57059
rect 14551 57052 14576 57104
rect 14576 57052 14603 57104
rect 2501 56734 2553 56741
rect 2609 56734 2661 56741
rect 2501 56689 2553 56734
rect 2609 56689 2661 56734
rect 369 56591 402 56643
rect 402 56591 421 56643
rect 493 56591 545 56643
rect 617 56591 669 56643
rect 741 56618 793 56643
rect 741 56591 760 56618
rect 760 56591 793 56618
rect 369 56467 402 56519
rect 402 56467 421 56519
rect 493 56467 545 56519
rect 617 56467 669 56519
rect 741 56467 760 56519
rect 760 56467 793 56519
rect 369 56343 402 56395
rect 402 56343 421 56395
rect 493 56343 545 56395
rect 617 56343 669 56395
rect 741 56343 760 56395
rect 760 56343 793 56395
rect 369 56219 402 56271
rect 402 56219 421 56271
rect 493 56219 545 56271
rect 617 56219 669 56271
rect 741 56219 760 56271
rect 760 56219 793 56271
rect 369 56095 402 56147
rect 402 56095 421 56147
rect 493 56095 545 56147
rect 617 56095 669 56147
rect 741 56095 760 56147
rect 760 56095 793 56147
rect 369 55971 402 56023
rect 402 55971 421 56023
rect 493 55971 545 56023
rect 617 55971 669 56023
rect 741 55971 760 56023
rect 760 55971 793 56023
rect 369 55847 402 55899
rect 402 55847 421 55899
rect 493 55847 545 55899
rect 617 55847 669 55899
rect 741 55847 760 55899
rect 760 55847 793 55899
rect 369 55723 402 55775
rect 402 55723 421 55775
rect 493 55723 545 55775
rect 617 55723 669 55775
rect 741 55723 760 55775
rect 760 55723 793 55775
rect 369 55599 402 55651
rect 402 55599 421 55651
rect 493 55599 545 55651
rect 617 55599 669 55651
rect 741 55599 760 55651
rect 760 55599 793 55651
rect 369 55475 402 55527
rect 402 55475 421 55527
rect 493 55475 545 55527
rect 617 55475 669 55527
rect 741 55475 760 55527
rect 760 55475 793 55527
rect 369 55351 402 55403
rect 402 55351 421 55403
rect 493 55351 545 55403
rect 617 55351 669 55403
rect 741 55351 760 55403
rect 760 55351 793 55403
rect 369 55227 402 55279
rect 402 55227 421 55279
rect 493 55227 545 55279
rect 617 55227 669 55279
rect 741 55227 760 55279
rect 760 55227 793 55279
rect 369 55103 402 55155
rect 402 55103 421 55155
rect 493 55103 545 55155
rect 617 55103 669 55155
rect 741 55103 760 55155
rect 760 55103 793 55155
rect 369 54979 402 55031
rect 402 54979 421 55031
rect 493 54979 545 55031
rect 617 54979 669 55031
rect 741 54979 760 55031
rect 760 54979 793 55031
rect 369 54855 402 54907
rect 402 54855 421 54907
rect 493 54855 545 54907
rect 617 54855 669 54907
rect 741 54855 760 54907
rect 760 54855 793 54907
rect 369 54731 402 54783
rect 402 54731 421 54783
rect 493 54731 545 54783
rect 617 54731 669 54783
rect 741 54731 760 54783
rect 760 54731 793 54783
rect 369 54607 402 54659
rect 402 54607 421 54659
rect 493 54607 545 54659
rect 617 54607 669 54659
rect 741 54607 760 54659
rect 760 54607 793 54659
rect 369 54483 402 54535
rect 402 54483 421 54535
rect 493 54483 545 54535
rect 617 54483 669 54535
rect 741 54483 760 54535
rect 760 54483 793 54535
rect 369 54359 402 54411
rect 402 54359 421 54411
rect 493 54359 545 54411
rect 617 54359 669 54411
rect 741 54359 760 54411
rect 760 54359 793 54411
rect 369 54235 402 54287
rect 402 54235 421 54287
rect 493 54235 545 54287
rect 617 54235 669 54287
rect 741 54235 760 54287
rect 760 54235 793 54287
rect 369 54111 402 54163
rect 402 54111 421 54163
rect 493 54111 545 54163
rect 617 54111 669 54163
rect 741 54111 760 54163
rect 760 54111 793 54163
rect 369 53987 402 54039
rect 402 53987 421 54039
rect 493 53987 545 54039
rect 617 53987 669 54039
rect 741 53987 760 54039
rect 760 53987 793 54039
rect 369 53863 402 53915
rect 402 53863 421 53915
rect 493 53863 545 53915
rect 617 53863 669 53915
rect 741 53863 760 53915
rect 760 53863 793 53915
rect 369 53739 402 53791
rect 402 53739 421 53791
rect 493 53739 545 53791
rect 617 53739 669 53791
rect 741 53739 760 53791
rect 760 53739 793 53791
rect 369 53615 402 53667
rect 402 53615 421 53667
rect 493 53615 545 53667
rect 617 53615 669 53667
rect 741 53615 793 53667
rect 4871 56688 4923 56693
rect 4979 56688 5031 56693
rect 2501 53576 2553 53621
rect 2609 53576 2661 53621
rect 2501 53569 2553 53576
rect 2609 53569 2661 53576
rect 3903 56618 3955 56643
rect 3903 56591 3910 56618
rect 3910 56591 3955 56618
rect 4027 56591 4079 56643
rect 4151 56618 4203 56643
rect 4151 56591 4196 56618
rect 4196 56591 4203 56618
rect 3903 56467 3910 56519
rect 3910 56467 3955 56519
rect 4027 56467 4079 56519
rect 4151 56467 4196 56519
rect 4196 56467 4203 56519
rect 3903 56343 3910 56395
rect 3910 56343 3955 56395
rect 4027 56343 4079 56395
rect 4151 56343 4196 56395
rect 4196 56343 4203 56395
rect 3903 56219 3910 56271
rect 3910 56219 3955 56271
rect 4027 56219 4079 56271
rect 4151 56219 4196 56271
rect 4196 56219 4203 56271
rect 3903 56095 3910 56147
rect 3910 56095 3955 56147
rect 4027 56095 4079 56147
rect 4151 56095 4196 56147
rect 4196 56095 4203 56147
rect 3903 55971 3910 56023
rect 3910 55971 3955 56023
rect 4027 55971 4079 56023
rect 4151 55971 4196 56023
rect 4196 55971 4203 56023
rect 3903 55847 3910 55899
rect 3910 55847 3955 55899
rect 4027 55847 4079 55899
rect 4151 55847 4196 55899
rect 4196 55847 4203 55899
rect 3903 55723 3910 55775
rect 3910 55723 3955 55775
rect 4027 55723 4079 55775
rect 4151 55723 4196 55775
rect 4196 55723 4203 55775
rect 3903 55599 3910 55651
rect 3910 55599 3955 55651
rect 4027 55599 4079 55651
rect 4151 55599 4196 55651
rect 4196 55599 4203 55651
rect 3903 55475 3910 55527
rect 3910 55475 3955 55527
rect 4027 55475 4079 55527
rect 4151 55475 4196 55527
rect 4196 55475 4203 55527
rect 3903 55351 3910 55403
rect 3910 55351 3955 55403
rect 4027 55351 4079 55403
rect 4151 55351 4196 55403
rect 4196 55351 4203 55403
rect 3903 55227 3910 55279
rect 3910 55227 3955 55279
rect 4027 55227 4079 55279
rect 4151 55227 4196 55279
rect 4196 55227 4203 55279
rect 3903 55103 3910 55155
rect 3910 55103 3955 55155
rect 4027 55103 4079 55155
rect 4151 55103 4196 55155
rect 4196 55103 4203 55155
rect 3903 54979 3910 55031
rect 3910 54979 3955 55031
rect 4027 54979 4079 55031
rect 4151 54979 4196 55031
rect 4196 54979 4203 55031
rect 3903 54855 3910 54907
rect 3910 54855 3955 54907
rect 4027 54855 4079 54907
rect 4151 54855 4196 54907
rect 4196 54855 4203 54907
rect 3903 54731 3910 54783
rect 3910 54731 3955 54783
rect 4027 54731 4079 54783
rect 4151 54731 4196 54783
rect 4196 54731 4203 54783
rect 3903 54607 3910 54659
rect 3910 54607 3955 54659
rect 4027 54607 4079 54659
rect 4151 54607 4196 54659
rect 4196 54607 4203 54659
rect 3903 54483 3910 54535
rect 3910 54483 3955 54535
rect 4027 54483 4079 54535
rect 4151 54483 4196 54535
rect 4196 54483 4203 54535
rect 3903 54359 3910 54411
rect 3910 54359 3955 54411
rect 4027 54359 4079 54411
rect 4151 54359 4196 54411
rect 4196 54359 4203 54411
rect 3903 54235 3910 54287
rect 3910 54235 3955 54287
rect 4027 54235 4079 54287
rect 4151 54235 4196 54287
rect 4196 54235 4203 54287
rect 3903 54111 3910 54163
rect 3910 54111 3955 54163
rect 4027 54111 4079 54163
rect 4151 54111 4196 54163
rect 4196 54111 4203 54163
rect 3903 53987 3910 54039
rect 3910 53987 3955 54039
rect 4027 53987 4079 54039
rect 4151 53987 4196 54039
rect 4196 53987 4203 54039
rect 3903 53863 3910 53915
rect 3910 53863 3955 53915
rect 4027 53863 4079 53915
rect 4151 53863 4196 53915
rect 4196 53863 4203 53915
rect 3903 53739 3910 53791
rect 3910 53739 3955 53791
rect 4027 53739 4079 53791
rect 4151 53739 4196 53791
rect 4196 53739 4203 53791
rect 3903 53615 3955 53667
rect 4027 53615 4079 53667
rect 4151 53615 4203 53667
rect 369 53491 402 53543
rect 402 53491 421 53543
rect 493 53491 545 53543
rect 617 53491 669 53543
rect 741 53491 793 53543
rect 4871 56641 4923 56688
rect 4979 56641 5031 56688
rect 4871 56533 4923 56585
rect 4979 56533 5031 56585
rect 4871 56425 4923 56477
rect 4979 56425 5031 56477
rect 4871 56317 4923 56369
rect 4979 56317 5031 56369
rect 4871 56209 4923 56261
rect 4979 56209 5031 56261
rect 4871 56101 4923 56153
rect 4979 56101 5031 56153
rect 4871 55993 4923 56045
rect 4979 55993 5031 56045
rect 4871 55885 4923 55937
rect 4979 55885 5031 55937
rect 4871 55777 4923 55829
rect 4979 55777 5031 55829
rect 4871 55669 4923 55721
rect 4979 55669 5031 55721
rect 4871 55561 4923 55613
rect 4979 55561 5031 55613
rect 4871 55453 4923 55505
rect 4979 55453 5031 55505
rect 4871 55345 4923 55397
rect 4979 55345 5031 55397
rect 4871 55237 4923 55289
rect 4979 55237 5031 55289
rect 4871 55129 4923 55181
rect 4979 55129 5031 55181
rect 4871 55021 4923 55073
rect 4979 55021 5031 55073
rect 4871 54913 4923 54965
rect 4979 54913 5031 54965
rect 4871 54805 4923 54857
rect 4979 54805 5031 54857
rect 4871 54697 4923 54749
rect 4979 54697 5031 54749
rect 4871 54589 4923 54641
rect 4979 54589 5031 54641
rect 4871 54481 4923 54533
rect 4979 54481 5031 54533
rect 4871 54373 4923 54425
rect 4979 54373 5031 54425
rect 4871 54265 4923 54317
rect 4979 54265 5031 54317
rect 4871 54157 4923 54209
rect 4979 54157 5031 54209
rect 4871 54049 4923 54101
rect 4979 54049 5031 54101
rect 4871 53941 4923 53993
rect 4979 53941 5031 53993
rect 4871 53833 4923 53885
rect 4979 53833 5031 53885
rect 4871 53725 4923 53777
rect 4979 53725 5031 53777
rect 4871 53622 4923 53669
rect 4979 53622 5031 53669
rect 9947 56688 9999 56693
rect 10055 56688 10107 56693
rect 4871 53617 4923 53622
rect 4979 53617 5031 53622
rect 3903 53491 3955 53543
rect 4027 53491 4079 53543
rect 4151 53491 4203 53543
rect 9947 56641 9999 56688
rect 10055 56641 10107 56688
rect 12317 56734 12369 56741
rect 12425 56734 12477 56741
rect 12317 56689 12369 56734
rect 12425 56689 12477 56734
rect 9947 56533 9999 56585
rect 10055 56533 10107 56585
rect 9947 56425 9999 56477
rect 10055 56425 10107 56477
rect 9947 56317 9999 56369
rect 10055 56317 10107 56369
rect 9947 56209 9999 56261
rect 10055 56209 10107 56261
rect 9947 56101 9999 56153
rect 10055 56101 10107 56153
rect 9947 55993 9999 56045
rect 10055 55993 10107 56045
rect 9947 55885 9999 55937
rect 10055 55885 10107 55937
rect 9947 55777 9999 55829
rect 10055 55777 10107 55829
rect 9947 55669 9999 55721
rect 10055 55669 10107 55721
rect 9947 55561 9999 55613
rect 10055 55561 10107 55613
rect 9947 55453 9999 55505
rect 10055 55453 10107 55505
rect 9947 55345 9999 55397
rect 10055 55345 10107 55397
rect 9947 55237 9999 55289
rect 10055 55237 10107 55289
rect 9947 55129 9999 55181
rect 10055 55129 10107 55181
rect 9947 55021 9999 55073
rect 10055 55021 10107 55073
rect 9947 54913 9999 54965
rect 10055 54913 10107 54965
rect 9947 54805 9999 54857
rect 10055 54805 10107 54857
rect 9947 54697 9999 54749
rect 10055 54697 10107 54749
rect 9947 54589 9999 54641
rect 10055 54589 10107 54641
rect 9947 54481 9999 54533
rect 10055 54481 10107 54533
rect 9947 54373 9999 54425
rect 10055 54373 10107 54425
rect 9947 54265 9999 54317
rect 10055 54265 10107 54317
rect 9947 54157 9999 54209
rect 10055 54157 10107 54209
rect 9947 54049 9999 54101
rect 10055 54049 10107 54101
rect 9947 53941 9999 53993
rect 10055 53941 10107 53993
rect 9947 53833 9999 53885
rect 10055 53833 10107 53885
rect 9947 53725 9999 53777
rect 10055 53725 10107 53777
rect 9947 53622 9999 53669
rect 10055 53622 10107 53669
rect 9947 53617 9999 53622
rect 10055 53617 10107 53622
rect 10775 56618 10827 56643
rect 10775 56591 10782 56618
rect 10782 56591 10827 56618
rect 10899 56591 10951 56643
rect 11023 56618 11075 56643
rect 11023 56591 11068 56618
rect 11068 56591 11075 56618
rect 10775 56467 10782 56519
rect 10782 56467 10827 56519
rect 10899 56467 10951 56519
rect 11023 56467 11068 56519
rect 11068 56467 11075 56519
rect 10775 56343 10782 56395
rect 10782 56343 10827 56395
rect 10899 56343 10951 56395
rect 11023 56343 11068 56395
rect 11068 56343 11075 56395
rect 10775 56219 10782 56271
rect 10782 56219 10827 56271
rect 10899 56219 10951 56271
rect 11023 56219 11068 56271
rect 11068 56219 11075 56271
rect 10775 56095 10782 56147
rect 10782 56095 10827 56147
rect 10899 56095 10951 56147
rect 11023 56095 11068 56147
rect 11068 56095 11075 56147
rect 10775 55971 10782 56023
rect 10782 55971 10827 56023
rect 10899 55971 10951 56023
rect 11023 55971 11068 56023
rect 11068 55971 11075 56023
rect 10775 55847 10782 55899
rect 10782 55847 10827 55899
rect 10899 55847 10951 55899
rect 11023 55847 11068 55899
rect 11068 55847 11075 55899
rect 10775 55723 10782 55775
rect 10782 55723 10827 55775
rect 10899 55723 10951 55775
rect 11023 55723 11068 55775
rect 11068 55723 11075 55775
rect 10775 55599 10782 55651
rect 10782 55599 10827 55651
rect 10899 55599 10951 55651
rect 11023 55599 11068 55651
rect 11068 55599 11075 55651
rect 10775 55475 10782 55527
rect 10782 55475 10827 55527
rect 10899 55475 10951 55527
rect 11023 55475 11068 55527
rect 11068 55475 11075 55527
rect 10775 55351 10782 55403
rect 10782 55351 10827 55403
rect 10899 55351 10951 55403
rect 11023 55351 11068 55403
rect 11068 55351 11075 55403
rect 10775 55227 10782 55279
rect 10782 55227 10827 55279
rect 10899 55227 10951 55279
rect 11023 55227 11068 55279
rect 11068 55227 11075 55279
rect 10775 55103 10782 55155
rect 10782 55103 10827 55155
rect 10899 55103 10951 55155
rect 11023 55103 11068 55155
rect 11068 55103 11075 55155
rect 10775 54979 10782 55031
rect 10782 54979 10827 55031
rect 10899 54979 10951 55031
rect 11023 54979 11068 55031
rect 11068 54979 11075 55031
rect 10775 54855 10782 54907
rect 10782 54855 10827 54907
rect 10899 54855 10951 54907
rect 11023 54855 11068 54907
rect 11068 54855 11075 54907
rect 10775 54731 10782 54783
rect 10782 54731 10827 54783
rect 10899 54731 10951 54783
rect 11023 54731 11068 54783
rect 11068 54731 11075 54783
rect 10775 54607 10782 54659
rect 10782 54607 10827 54659
rect 10899 54607 10951 54659
rect 11023 54607 11068 54659
rect 11068 54607 11075 54659
rect 10775 54483 10782 54535
rect 10782 54483 10827 54535
rect 10899 54483 10951 54535
rect 11023 54483 11068 54535
rect 11068 54483 11075 54535
rect 10775 54359 10782 54411
rect 10782 54359 10827 54411
rect 10899 54359 10951 54411
rect 11023 54359 11068 54411
rect 11068 54359 11075 54411
rect 10775 54235 10782 54287
rect 10782 54235 10827 54287
rect 10899 54235 10951 54287
rect 11023 54235 11068 54287
rect 11068 54235 11075 54287
rect 10775 54111 10782 54163
rect 10782 54111 10827 54163
rect 10899 54111 10951 54163
rect 11023 54111 11068 54163
rect 11068 54111 11075 54163
rect 10775 53987 10782 54039
rect 10782 53987 10827 54039
rect 10899 53987 10951 54039
rect 11023 53987 11068 54039
rect 11068 53987 11075 54039
rect 10775 53863 10782 53915
rect 10782 53863 10827 53915
rect 10899 53863 10951 53915
rect 11023 53863 11068 53915
rect 11068 53863 11075 53915
rect 10775 53739 10782 53791
rect 10782 53739 10827 53791
rect 10899 53739 10951 53791
rect 11023 53739 11068 53791
rect 11068 53739 11075 53791
rect 10775 53615 10827 53667
rect 10899 53615 10951 53667
rect 11023 53615 11075 53667
rect 12317 53576 12369 53621
rect 12425 53576 12477 53621
rect 12317 53569 12369 53576
rect 12425 53569 12477 53576
rect 14185 56618 14237 56643
rect 14185 56591 14218 56618
rect 14218 56591 14237 56618
rect 14309 56591 14361 56643
rect 14433 56591 14485 56643
rect 14557 56591 14576 56643
rect 14576 56591 14609 56643
rect 14185 56467 14218 56519
rect 14218 56467 14237 56519
rect 14309 56467 14361 56519
rect 14433 56467 14485 56519
rect 14557 56467 14576 56519
rect 14576 56467 14609 56519
rect 14185 56343 14218 56395
rect 14218 56343 14237 56395
rect 14309 56343 14361 56395
rect 14433 56343 14485 56395
rect 14557 56343 14576 56395
rect 14576 56343 14609 56395
rect 14185 56219 14218 56271
rect 14218 56219 14237 56271
rect 14309 56219 14361 56271
rect 14433 56219 14485 56271
rect 14557 56219 14576 56271
rect 14576 56219 14609 56271
rect 14185 56095 14218 56147
rect 14218 56095 14237 56147
rect 14309 56095 14361 56147
rect 14433 56095 14485 56147
rect 14557 56095 14576 56147
rect 14576 56095 14609 56147
rect 14185 55971 14218 56023
rect 14218 55971 14237 56023
rect 14309 55971 14361 56023
rect 14433 55971 14485 56023
rect 14557 55971 14576 56023
rect 14576 55971 14609 56023
rect 14185 55847 14218 55899
rect 14218 55847 14237 55899
rect 14309 55847 14361 55899
rect 14433 55847 14485 55899
rect 14557 55847 14576 55899
rect 14576 55847 14609 55899
rect 14185 55723 14218 55775
rect 14218 55723 14237 55775
rect 14309 55723 14361 55775
rect 14433 55723 14485 55775
rect 14557 55723 14576 55775
rect 14576 55723 14609 55775
rect 14185 55599 14218 55651
rect 14218 55599 14237 55651
rect 14309 55599 14361 55651
rect 14433 55599 14485 55651
rect 14557 55599 14576 55651
rect 14576 55599 14609 55651
rect 14185 55475 14218 55527
rect 14218 55475 14237 55527
rect 14309 55475 14361 55527
rect 14433 55475 14485 55527
rect 14557 55475 14576 55527
rect 14576 55475 14609 55527
rect 14185 55351 14218 55403
rect 14218 55351 14237 55403
rect 14309 55351 14361 55403
rect 14433 55351 14485 55403
rect 14557 55351 14576 55403
rect 14576 55351 14609 55403
rect 14185 55227 14218 55279
rect 14218 55227 14237 55279
rect 14309 55227 14361 55279
rect 14433 55227 14485 55279
rect 14557 55227 14576 55279
rect 14576 55227 14609 55279
rect 14185 55103 14218 55155
rect 14218 55103 14237 55155
rect 14309 55103 14361 55155
rect 14433 55103 14485 55155
rect 14557 55103 14576 55155
rect 14576 55103 14609 55155
rect 14185 54979 14218 55031
rect 14218 54979 14237 55031
rect 14309 54979 14361 55031
rect 14433 54979 14485 55031
rect 14557 54979 14576 55031
rect 14576 54979 14609 55031
rect 14185 54855 14218 54907
rect 14218 54855 14237 54907
rect 14309 54855 14361 54907
rect 14433 54855 14485 54907
rect 14557 54855 14576 54907
rect 14576 54855 14609 54907
rect 14185 54731 14218 54783
rect 14218 54731 14237 54783
rect 14309 54731 14361 54783
rect 14433 54731 14485 54783
rect 14557 54731 14576 54783
rect 14576 54731 14609 54783
rect 14185 54607 14218 54659
rect 14218 54607 14237 54659
rect 14309 54607 14361 54659
rect 14433 54607 14485 54659
rect 14557 54607 14576 54659
rect 14576 54607 14609 54659
rect 14185 54483 14218 54535
rect 14218 54483 14237 54535
rect 14309 54483 14361 54535
rect 14433 54483 14485 54535
rect 14557 54483 14576 54535
rect 14576 54483 14609 54535
rect 14185 54359 14218 54411
rect 14218 54359 14237 54411
rect 14309 54359 14361 54411
rect 14433 54359 14485 54411
rect 14557 54359 14576 54411
rect 14576 54359 14609 54411
rect 14185 54235 14218 54287
rect 14218 54235 14237 54287
rect 14309 54235 14361 54287
rect 14433 54235 14485 54287
rect 14557 54235 14576 54287
rect 14576 54235 14609 54287
rect 14185 54111 14218 54163
rect 14218 54111 14237 54163
rect 14309 54111 14361 54163
rect 14433 54111 14485 54163
rect 14557 54111 14576 54163
rect 14576 54111 14609 54163
rect 14185 53987 14218 54039
rect 14218 53987 14237 54039
rect 14309 53987 14361 54039
rect 14433 53987 14485 54039
rect 14557 53987 14576 54039
rect 14576 53987 14609 54039
rect 14185 53863 14218 53915
rect 14218 53863 14237 53915
rect 14309 53863 14361 53915
rect 14433 53863 14485 53915
rect 14557 53863 14576 53915
rect 14576 53863 14609 53915
rect 14185 53739 14218 53791
rect 14218 53739 14237 53791
rect 14309 53739 14361 53791
rect 14433 53739 14485 53791
rect 14557 53739 14576 53791
rect 14576 53739 14609 53791
rect 14185 53615 14237 53667
rect 14309 53615 14361 53667
rect 14433 53615 14485 53667
rect 14557 53615 14576 53667
rect 14576 53615 14609 53667
rect 10775 53491 10827 53543
rect 10899 53491 10951 53543
rect 11023 53491 11075 53543
rect 14185 53491 14237 53543
rect 14309 53491 14361 53543
rect 14433 53491 14485 53543
rect 14557 53491 14576 53543
rect 14576 53491 14609 53543
rect 869 53431 921 53483
rect 977 53431 1029 53483
rect 1085 53431 1137 53483
rect 1193 53431 1245 53483
rect 1301 53431 1353 53483
rect 1409 53431 1461 53483
rect 1517 53431 1569 53483
rect 1625 53431 1677 53483
rect 1733 53431 1785 53483
rect 1841 53431 1893 53483
rect 1949 53431 2001 53483
rect 2057 53431 2109 53483
rect 2763 53431 2815 53483
rect 2871 53431 2923 53483
rect 2979 53431 3031 53483
rect 3087 53431 3139 53483
rect 3195 53431 3247 53483
rect 3303 53431 3355 53483
rect 3411 53431 3463 53483
rect 3519 53431 3571 53483
rect 3627 53431 3679 53483
rect 3735 53431 3787 53483
rect 5138 53431 5190 53483
rect 5246 53431 5298 53483
rect 5354 53431 5406 53483
rect 5462 53431 5514 53483
rect 5570 53431 5622 53483
rect 5678 53431 5730 53483
rect 5786 53431 5838 53483
rect 5894 53431 5946 53483
rect 6002 53431 6054 53483
rect 6110 53431 6162 53483
rect 6218 53431 6270 53483
rect 6326 53431 6378 53483
rect 6434 53431 6486 53483
rect 6542 53431 6594 53483
rect 6650 53431 6702 53483
rect 6758 53431 6810 53483
rect 6866 53431 6918 53483
rect 6974 53431 7026 53483
rect 7082 53431 7134 53483
rect 7844 53431 7896 53483
rect 7952 53431 8004 53483
rect 8060 53431 8112 53483
rect 8168 53431 8220 53483
rect 8276 53431 8328 53483
rect 8384 53431 8436 53483
rect 8492 53431 8544 53483
rect 8600 53431 8652 53483
rect 8708 53431 8760 53483
rect 8816 53431 8868 53483
rect 8924 53431 8976 53483
rect 9032 53431 9084 53483
rect 9140 53431 9192 53483
rect 9248 53431 9300 53483
rect 9356 53431 9408 53483
rect 9464 53431 9516 53483
rect 9572 53431 9624 53483
rect 9680 53431 9732 53483
rect 9788 53431 9840 53483
rect 11191 53431 11243 53483
rect 11299 53431 11351 53483
rect 11407 53431 11459 53483
rect 11515 53431 11567 53483
rect 11623 53431 11675 53483
rect 11731 53431 11783 53483
rect 11839 53431 11891 53483
rect 11947 53431 11999 53483
rect 12055 53431 12107 53483
rect 12163 53431 12215 53483
rect 12869 53431 12921 53483
rect 12977 53431 13029 53483
rect 13085 53431 13137 53483
rect 13193 53431 13245 53483
rect 13301 53431 13353 53483
rect 13409 53431 13461 53483
rect 13517 53431 13569 53483
rect 13625 53431 13677 53483
rect 13733 53431 13785 53483
rect 13841 53431 13893 53483
rect 13949 53431 14001 53483
rect 14057 53431 14109 53483
rect 369 53367 402 53419
rect 402 53367 421 53419
rect 493 53367 545 53419
rect 617 53367 669 53419
rect 741 53367 793 53419
rect 869 53323 921 53375
rect 977 53323 1029 53375
rect 1085 53323 1137 53375
rect 1193 53323 1245 53375
rect 1301 53323 1353 53375
rect 1409 53323 1461 53375
rect 1517 53323 1569 53375
rect 1625 53323 1677 53375
rect 1733 53323 1785 53375
rect 1841 53323 1893 53375
rect 1949 53323 2001 53375
rect 2057 53323 2109 53375
rect 2763 53323 2815 53375
rect 2871 53323 2923 53375
rect 2979 53323 3031 53375
rect 3087 53323 3139 53375
rect 3195 53323 3247 53375
rect 3303 53323 3355 53375
rect 3411 53323 3463 53375
rect 3519 53323 3571 53375
rect 3627 53323 3679 53375
rect 3735 53323 3787 53375
rect 3903 53367 3955 53419
rect 4027 53367 4079 53419
rect 4151 53367 4203 53419
rect 5138 53323 5190 53375
rect 5246 53323 5298 53375
rect 5354 53323 5406 53375
rect 5462 53323 5514 53375
rect 5570 53323 5622 53375
rect 5678 53323 5730 53375
rect 5786 53323 5838 53375
rect 5894 53323 5946 53375
rect 6002 53323 6054 53375
rect 6110 53323 6162 53375
rect 6218 53323 6270 53375
rect 6326 53323 6378 53375
rect 6434 53323 6486 53375
rect 6542 53323 6594 53375
rect 6650 53323 6702 53375
rect 6758 53323 6810 53375
rect 6866 53323 6918 53375
rect 6974 53323 7026 53375
rect 7082 53323 7134 53375
rect 7844 53323 7896 53375
rect 7952 53323 8004 53375
rect 8060 53323 8112 53375
rect 8168 53323 8220 53375
rect 8276 53323 8328 53375
rect 8384 53323 8436 53375
rect 8492 53323 8544 53375
rect 8600 53323 8652 53375
rect 8708 53323 8760 53375
rect 8816 53323 8868 53375
rect 8924 53323 8976 53375
rect 9032 53323 9084 53375
rect 9140 53323 9192 53375
rect 9248 53323 9300 53375
rect 9356 53323 9408 53375
rect 9464 53323 9516 53375
rect 9572 53323 9624 53375
rect 9680 53323 9732 53375
rect 9788 53323 9840 53375
rect 10775 53367 10827 53419
rect 10899 53367 10951 53419
rect 11023 53367 11075 53419
rect 11191 53323 11243 53375
rect 11299 53323 11351 53375
rect 11407 53323 11459 53375
rect 11515 53323 11567 53375
rect 11623 53323 11675 53375
rect 11731 53323 11783 53375
rect 11839 53323 11891 53375
rect 11947 53323 11999 53375
rect 12055 53323 12107 53375
rect 12163 53323 12215 53375
rect 12869 53323 12921 53375
rect 12977 53323 13029 53375
rect 13085 53323 13137 53375
rect 13193 53323 13245 53375
rect 13301 53323 13353 53375
rect 13409 53323 13461 53375
rect 13517 53323 13569 53375
rect 13625 53323 13677 53375
rect 13733 53323 13785 53375
rect 13841 53323 13893 53375
rect 13949 53323 14001 53375
rect 14057 53323 14109 53375
rect 14185 53367 14237 53419
rect 14309 53367 14361 53419
rect 14433 53367 14485 53419
rect 14557 53367 14576 53419
rect 14576 53367 14609 53419
rect 369 53243 402 53295
rect 402 53243 421 53295
rect 493 53251 545 53295
rect 617 53251 669 53295
rect 741 53251 793 53295
rect 869 53251 921 53267
rect 977 53251 1029 53267
rect 1085 53251 1137 53267
rect 1193 53251 1245 53267
rect 1301 53251 1353 53267
rect 1409 53251 1461 53267
rect 1517 53251 1569 53267
rect 1625 53251 1677 53267
rect 1733 53251 1785 53267
rect 1841 53251 1893 53267
rect 1949 53251 2001 53267
rect 2057 53251 2109 53267
rect 2763 53251 2815 53267
rect 2871 53251 2923 53267
rect 2979 53251 3031 53267
rect 3087 53251 3139 53267
rect 3195 53251 3247 53267
rect 3303 53251 3355 53267
rect 3411 53251 3463 53267
rect 3519 53251 3571 53267
rect 3627 53251 3679 53267
rect 3735 53251 3787 53267
rect 3903 53251 3955 53295
rect 4027 53251 4079 53295
rect 4151 53251 4203 53295
rect 5138 53251 5190 53267
rect 5246 53251 5298 53267
rect 5354 53251 5406 53267
rect 5462 53251 5514 53267
rect 5570 53251 5622 53267
rect 5678 53251 5730 53267
rect 5786 53251 5838 53267
rect 5894 53251 5946 53267
rect 6002 53251 6054 53267
rect 6110 53251 6162 53267
rect 6218 53251 6270 53267
rect 6326 53251 6378 53267
rect 6434 53251 6486 53267
rect 6542 53251 6594 53267
rect 6650 53251 6702 53267
rect 6758 53251 6810 53267
rect 6866 53251 6918 53267
rect 6974 53251 7026 53267
rect 7082 53251 7134 53267
rect 7844 53251 7896 53267
rect 7952 53251 8004 53267
rect 8060 53251 8112 53267
rect 8168 53251 8220 53267
rect 8276 53251 8328 53267
rect 8384 53251 8436 53267
rect 8492 53251 8544 53267
rect 8600 53251 8652 53267
rect 8708 53251 8760 53267
rect 8816 53251 8868 53267
rect 8924 53251 8976 53267
rect 9032 53251 9084 53267
rect 9140 53251 9192 53267
rect 9248 53251 9300 53267
rect 9356 53251 9408 53267
rect 9464 53251 9516 53267
rect 9572 53251 9624 53267
rect 9680 53251 9732 53267
rect 9788 53251 9840 53267
rect 10775 53251 10827 53295
rect 10899 53251 10951 53295
rect 11023 53251 11075 53295
rect 11191 53251 11243 53267
rect 11299 53251 11351 53267
rect 11407 53251 11459 53267
rect 11515 53251 11567 53267
rect 11623 53251 11675 53267
rect 11731 53251 11783 53267
rect 11839 53251 11891 53267
rect 11947 53251 11999 53267
rect 12055 53251 12107 53267
rect 12163 53251 12215 53267
rect 12869 53251 12921 53267
rect 12977 53251 13029 53267
rect 13085 53251 13137 53267
rect 13193 53251 13245 53267
rect 13301 53251 13353 53267
rect 13409 53251 13461 53267
rect 13517 53251 13569 53267
rect 13625 53251 13677 53267
rect 13733 53251 13785 53267
rect 13841 53251 13893 53267
rect 13949 53251 14001 53267
rect 14057 53251 14109 53267
rect 14185 53251 14237 53295
rect 14309 53251 14361 53295
rect 14433 53251 14485 53295
rect 493 53243 510 53251
rect 510 53243 545 53251
rect 617 53243 669 53251
rect 741 53243 793 53251
rect 869 53215 921 53251
rect 977 53215 1029 53251
rect 1085 53215 1137 53251
rect 1193 53215 1245 53251
rect 1301 53215 1353 53251
rect 1409 53215 1461 53251
rect 1517 53215 1569 53251
rect 1625 53215 1677 53251
rect 1733 53215 1785 53251
rect 1841 53215 1893 53251
rect 1949 53215 2001 53251
rect 2057 53215 2109 53251
rect 2763 53215 2815 53251
rect 2871 53215 2923 53251
rect 2979 53215 3031 53251
rect 3087 53215 3139 53251
rect 3195 53215 3247 53251
rect 3303 53215 3355 53251
rect 3411 53215 3463 53251
rect 3519 53215 3571 53251
rect 3627 53215 3679 53251
rect 3735 53215 3787 53251
rect 3903 53243 3955 53251
rect 4027 53243 4079 53251
rect 4151 53243 4203 53251
rect 5138 53215 5190 53251
rect 5246 53215 5298 53251
rect 5354 53215 5406 53251
rect 5462 53215 5514 53251
rect 5570 53215 5622 53251
rect 5678 53215 5730 53251
rect 5786 53215 5838 53251
rect 5894 53215 5946 53251
rect 6002 53215 6054 53251
rect 6110 53215 6162 53251
rect 6218 53215 6270 53251
rect 6326 53215 6378 53251
rect 6434 53215 6486 53251
rect 6542 53215 6594 53251
rect 6650 53215 6702 53251
rect 6758 53215 6810 53251
rect 6866 53215 6918 53251
rect 6974 53215 7026 53251
rect 7082 53215 7134 53251
rect 7844 53215 7896 53251
rect 7952 53215 8004 53251
rect 8060 53215 8112 53251
rect 8168 53215 8220 53251
rect 8276 53215 8328 53251
rect 8384 53215 8436 53251
rect 8492 53215 8544 53251
rect 8600 53215 8652 53251
rect 8708 53215 8760 53251
rect 8816 53215 8868 53251
rect 8924 53215 8976 53251
rect 9032 53215 9084 53251
rect 9140 53215 9192 53251
rect 9248 53215 9300 53251
rect 9356 53215 9408 53251
rect 9464 53215 9516 53251
rect 9572 53215 9624 53251
rect 9680 53215 9732 53251
rect 9788 53215 9840 53251
rect 10775 53243 10827 53251
rect 10899 53243 10951 53251
rect 11023 53243 11075 53251
rect 11191 53215 11243 53251
rect 11299 53215 11351 53251
rect 11407 53215 11459 53251
rect 11515 53215 11567 53251
rect 11623 53215 11675 53251
rect 11731 53215 11783 53251
rect 11839 53215 11891 53251
rect 11947 53215 11999 53251
rect 12055 53215 12107 53251
rect 12163 53215 12215 53251
rect 12869 53215 12921 53251
rect 12977 53215 13029 53251
rect 13085 53215 13137 53251
rect 13193 53215 13245 53251
rect 13301 53215 13353 53251
rect 13409 53215 13461 53251
rect 13517 53215 13569 53251
rect 13625 53215 13677 53251
rect 13733 53215 13785 53251
rect 13841 53215 13893 53251
rect 13949 53215 14001 53251
rect 14057 53215 14109 53251
rect 14185 53243 14237 53251
rect 14309 53243 14361 53251
rect 14433 53243 14468 53251
rect 14468 53243 14485 53251
rect 14557 53243 14576 53295
rect 14576 53243 14609 53295
rect 14904 57099 14956 57151
rect 14904 56991 14956 57043
rect 14904 56883 14956 56935
rect 14904 56775 14956 56827
rect 14904 56667 14956 56719
rect 14904 56559 14956 56611
rect 14904 56451 14956 56503
rect 14904 56343 14956 56395
rect 14904 56235 14956 56287
rect 14904 56127 14956 56179
rect 14904 56019 14956 56071
rect 14904 54122 14956 54174
rect 14904 54014 14956 54066
rect 14904 53906 14956 53958
rect 14904 53798 14956 53850
rect 14904 53690 14956 53742
rect 14904 53582 14956 53634
rect 14904 53474 14956 53526
rect 14904 53366 14956 53418
rect 14904 53258 14956 53310
rect 22 53042 74 53094
rect 22 52934 74 52986
rect 22 52826 74 52878
rect 14904 53150 14956 53202
rect 14904 53042 14956 53094
rect 14904 52934 14956 52986
rect 14904 52826 14956 52878
rect 22 52522 74 52574
rect 22 52414 74 52466
rect 22 52306 74 52358
rect 22 52198 74 52250
rect 22 52090 74 52142
rect 22 51982 74 52034
rect 22 51874 74 51926
rect 22 51766 74 51818
rect 22 51658 74 51710
rect 22 51550 74 51602
rect 22 51442 74 51494
rect 22 51334 74 51386
rect 22 51226 74 51278
rect 22 49322 74 49374
rect 22 49214 74 49266
rect 22 49106 74 49158
rect 22 48998 74 49050
rect 22 48890 74 48942
rect 22 48782 74 48834
rect 22 48674 74 48726
rect 22 48566 74 48618
rect 22 48458 74 48510
rect 22 48350 74 48402
rect 22 48242 74 48294
rect 22 48134 74 48186
rect 22 48026 74 48078
rect 2590 52542 2642 52594
rect 2590 52434 2642 52486
rect 2590 52326 2642 52378
rect 2590 52218 2642 52270
rect 4871 52520 4923 52572
rect 4979 52520 5031 52572
rect 7247 52520 7299 52572
rect 7355 52520 7407 52572
rect 7463 52520 7515 52572
rect 7571 52520 7623 52572
rect 7679 52520 7731 52572
rect 9947 52520 9999 52572
rect 10055 52520 10107 52572
rect 4871 52412 4923 52464
rect 4979 52412 5031 52464
rect 7247 52412 7299 52464
rect 7355 52412 7407 52464
rect 7463 52412 7515 52464
rect 7571 52412 7623 52464
rect 7679 52412 7731 52464
rect 9947 52412 9999 52464
rect 10055 52412 10107 52464
rect 4871 52304 4923 52356
rect 4979 52304 5031 52356
rect 7247 52304 7299 52356
rect 7355 52304 7407 52356
rect 7463 52304 7515 52356
rect 7571 52304 7623 52356
rect 7679 52304 7731 52356
rect 9947 52304 9999 52356
rect 10055 52304 10107 52356
rect 12336 52542 12388 52594
rect 12336 52434 12388 52486
rect 12336 52326 12388 52378
rect 2590 52110 2642 52162
rect 2590 52002 2642 52054
rect 2590 51894 2642 51946
rect 2590 51786 2642 51838
rect 2590 51678 2642 51730
rect 2590 51570 2642 51622
rect 2590 51462 2642 51514
rect 2590 51354 2642 51406
rect 2590 51246 2642 51298
rect 2590 51138 2642 51190
rect 2590 51030 2642 51082
rect 2590 50922 2642 50974
rect 2590 50814 2642 50866
rect 2590 50706 2642 50758
rect 2590 50598 2642 50650
rect 2590 50490 2642 50542
rect 2590 50382 2642 50434
rect 2590 50274 2642 50326
rect 2590 50166 2642 50218
rect 2590 50058 2642 50110
rect 2590 49950 2642 50002
rect 2590 49842 2642 49894
rect 2590 49734 2642 49786
rect 2590 49626 2642 49678
rect 2590 49518 2642 49570
rect 2590 49410 2642 49462
rect 2590 49302 2642 49354
rect 2590 49194 2642 49246
rect 2590 49086 2642 49138
rect 2590 48978 2642 49030
rect 2590 48870 2642 48922
rect 2590 48762 2642 48814
rect 2590 48654 2642 48706
rect 2590 48546 2642 48598
rect 2590 48438 2642 48490
rect 2590 48330 2642 48382
rect 2590 48222 2642 48274
rect 2590 48114 2642 48166
rect 2590 48006 2642 48058
rect 3161 51983 3213 52009
rect 3269 51983 3321 52009
rect 3377 51983 3429 52009
rect 3485 51983 3537 52009
rect 3593 51983 3645 52009
rect 3701 51983 3753 52009
rect 3809 51983 3861 52009
rect 3917 51983 3969 52009
rect 4025 51983 4077 52009
rect 4133 51983 4185 52009
rect 4241 51983 4293 52009
rect 4349 51983 4401 52009
rect 4457 51983 4509 52009
rect 4565 51983 4617 52009
rect 4673 51983 4725 52009
rect 5138 51983 5190 52009
rect 5246 51983 5298 52009
rect 5354 51983 5406 52009
rect 5462 51983 5514 52009
rect 5570 51983 5622 52009
rect 5678 51983 5730 52009
rect 5786 51983 5838 52009
rect 5894 51983 5946 52009
rect 6002 51983 6054 52009
rect 6110 51983 6162 52009
rect 6218 51983 6270 52009
rect 6326 51983 6378 52009
rect 6434 51983 6486 52009
rect 6542 51983 6594 52009
rect 6650 51983 6702 52009
rect 6758 51983 6810 52009
rect 6866 51983 6918 52009
rect 6974 51983 7026 52009
rect 7082 51983 7134 52009
rect 7844 51983 7896 52009
rect 7952 51983 8004 52009
rect 8060 51983 8112 52009
rect 8168 51983 8220 52009
rect 8276 51983 8328 52009
rect 8384 51983 8436 52009
rect 8492 51983 8544 52009
rect 8600 51983 8652 52009
rect 8708 51983 8760 52009
rect 8816 51983 8868 52009
rect 8924 51983 8976 52009
rect 9032 51983 9084 52009
rect 9140 51983 9192 52009
rect 9248 51983 9300 52009
rect 9356 51983 9408 52009
rect 9464 51983 9516 52009
rect 9572 51983 9624 52009
rect 9680 51983 9732 52009
rect 9788 51983 9840 52009
rect 10253 51983 10305 52009
rect 10361 51983 10413 52009
rect 10469 51983 10521 52009
rect 10577 51983 10629 52009
rect 10685 51983 10737 52009
rect 10793 51983 10845 52009
rect 10901 51983 10953 52009
rect 11009 51983 11061 52009
rect 11117 51983 11169 52009
rect 11225 51983 11277 52009
rect 11333 51983 11385 52009
rect 11441 51983 11493 52009
rect 11549 51983 11601 52009
rect 11657 51983 11709 52009
rect 11765 51983 11817 52009
rect 3161 51957 3213 51983
rect 3269 51957 3321 51983
rect 3377 51957 3429 51983
rect 3485 51957 3537 51983
rect 3593 51957 3645 51983
rect 3701 51957 3753 51983
rect 3809 51957 3861 51983
rect 3917 51957 3969 51983
rect 4025 51957 4077 51983
rect 4133 51957 4185 51983
rect 4241 51957 4293 51983
rect 4349 51957 4401 51983
rect 4457 51957 4509 51983
rect 4565 51957 4617 51983
rect 4673 51957 4725 51983
rect 5138 51957 5190 51983
rect 5246 51957 5298 51983
rect 5354 51957 5406 51983
rect 5462 51957 5514 51983
rect 5570 51957 5622 51983
rect 5678 51957 5730 51983
rect 5786 51957 5838 51983
rect 5894 51957 5946 51983
rect 6002 51957 6054 51983
rect 6110 51957 6162 51983
rect 6218 51957 6270 51983
rect 6326 51957 6378 51983
rect 6434 51957 6486 51983
rect 6542 51957 6594 51983
rect 6650 51957 6702 51983
rect 6758 51957 6810 51983
rect 6866 51957 6918 51983
rect 6974 51957 7026 51983
rect 7082 51957 7134 51983
rect 7844 51957 7896 51983
rect 7952 51957 8004 51983
rect 8060 51957 8112 51983
rect 8168 51957 8220 51983
rect 8276 51957 8328 51983
rect 8384 51957 8436 51983
rect 8492 51957 8544 51983
rect 8600 51957 8652 51983
rect 8708 51957 8760 51983
rect 8816 51957 8868 51983
rect 8924 51957 8976 51983
rect 9032 51957 9084 51983
rect 9140 51957 9192 51983
rect 9248 51957 9300 51983
rect 9356 51957 9408 51983
rect 9464 51957 9516 51983
rect 9572 51957 9624 51983
rect 9680 51957 9732 51983
rect 9788 51957 9840 51983
rect 10253 51957 10305 51983
rect 10361 51957 10413 51983
rect 10469 51957 10521 51983
rect 10577 51957 10629 51983
rect 10685 51957 10737 51983
rect 10793 51957 10845 51983
rect 10901 51957 10953 51983
rect 11009 51957 11061 51983
rect 11117 51957 11169 51983
rect 11225 51957 11277 51983
rect 11333 51957 11385 51983
rect 11441 51957 11493 51983
rect 11549 51957 11601 51983
rect 11657 51957 11709 51983
rect 11765 51957 11817 51983
rect 3161 51900 3213 51901
rect 3161 51849 3162 51900
rect 3162 51849 3213 51900
rect 3269 51849 3321 51901
rect 3377 51875 3429 51901
rect 3485 51875 3537 51901
rect 3593 51875 3645 51901
rect 3701 51875 3753 51901
rect 3809 51875 3861 51901
rect 3917 51875 3969 51901
rect 4025 51875 4077 51901
rect 4133 51875 4185 51901
rect 4241 51875 4293 51901
rect 4349 51875 4401 51901
rect 4457 51875 4509 51901
rect 4565 51875 4617 51901
rect 4673 51875 4725 51901
rect 5138 51875 5190 51901
rect 5246 51875 5298 51901
rect 5354 51875 5406 51901
rect 5462 51875 5514 51901
rect 5570 51875 5622 51901
rect 5678 51875 5730 51901
rect 5786 51875 5838 51901
rect 5894 51875 5946 51901
rect 6002 51875 6054 51901
rect 6110 51875 6162 51901
rect 6218 51875 6270 51901
rect 6326 51875 6378 51901
rect 6434 51875 6486 51901
rect 6542 51875 6594 51901
rect 6650 51875 6702 51901
rect 6758 51875 6810 51901
rect 6866 51875 6918 51901
rect 6974 51875 7026 51901
rect 7082 51875 7134 51901
rect 7844 51875 7896 51901
rect 7952 51875 8004 51901
rect 8060 51875 8112 51901
rect 8168 51875 8220 51901
rect 8276 51875 8328 51901
rect 8384 51875 8436 51901
rect 8492 51875 8544 51901
rect 8600 51875 8652 51901
rect 8708 51875 8760 51901
rect 8816 51875 8868 51901
rect 8924 51875 8976 51901
rect 9032 51875 9084 51901
rect 9140 51875 9192 51901
rect 9248 51875 9300 51901
rect 9356 51875 9408 51901
rect 9464 51875 9516 51901
rect 9572 51875 9624 51901
rect 9680 51875 9732 51901
rect 9788 51875 9840 51901
rect 10253 51875 10305 51901
rect 10361 51875 10413 51901
rect 10469 51875 10521 51901
rect 10577 51875 10629 51901
rect 10685 51875 10737 51901
rect 10793 51875 10845 51901
rect 10901 51875 10953 51901
rect 11009 51875 11061 51901
rect 11117 51875 11169 51901
rect 11225 51875 11277 51901
rect 11333 51875 11385 51901
rect 11441 51875 11493 51901
rect 11549 51875 11601 51901
rect 3377 51849 3424 51875
rect 3424 51849 3429 51875
rect 3485 51849 3537 51875
rect 3593 51849 3645 51875
rect 3701 51849 3753 51875
rect 3809 51849 3861 51875
rect 3917 51849 3969 51875
rect 4025 51849 4077 51875
rect 4133 51849 4185 51875
rect 4241 51849 4293 51875
rect 4349 51849 4401 51875
rect 4457 51849 4509 51875
rect 4565 51849 4617 51875
rect 4673 51849 4725 51875
rect 5138 51849 5190 51875
rect 5246 51849 5298 51875
rect 5354 51849 5406 51875
rect 5462 51849 5514 51875
rect 5570 51849 5622 51875
rect 5678 51849 5730 51875
rect 5786 51849 5838 51875
rect 5894 51849 5946 51875
rect 6002 51849 6054 51875
rect 6110 51849 6162 51875
rect 6218 51849 6270 51875
rect 6326 51849 6378 51875
rect 6434 51849 6486 51875
rect 6542 51849 6594 51875
rect 6650 51849 6702 51875
rect 6758 51849 6810 51875
rect 6866 51849 6918 51875
rect 6974 51849 7026 51875
rect 7082 51849 7134 51875
rect 7844 51849 7896 51875
rect 7952 51849 8004 51875
rect 8060 51849 8112 51875
rect 8168 51849 8220 51875
rect 8276 51849 8328 51875
rect 8384 51849 8436 51875
rect 8492 51849 8544 51875
rect 8600 51849 8652 51875
rect 8708 51849 8760 51875
rect 8816 51849 8868 51875
rect 8924 51849 8976 51875
rect 9032 51849 9084 51875
rect 9140 51849 9192 51875
rect 9248 51849 9300 51875
rect 9356 51849 9408 51875
rect 9464 51849 9516 51875
rect 9572 51849 9624 51875
rect 9680 51849 9732 51875
rect 9788 51849 9840 51875
rect 10253 51849 10305 51875
rect 10361 51849 10413 51875
rect 10469 51849 10521 51875
rect 10577 51849 10629 51875
rect 10685 51849 10737 51875
rect 10793 51849 10845 51875
rect 10901 51849 10953 51875
rect 11009 51849 11061 51875
rect 11117 51849 11169 51875
rect 11225 51849 11277 51875
rect 11333 51849 11385 51875
rect 11441 51849 11493 51875
rect 11549 51849 11554 51875
rect 11554 51849 11601 51875
rect 11657 51849 11709 51901
rect 11765 51900 11817 51901
rect 11765 51849 11816 51900
rect 11816 51849 11817 51900
rect 4871 51580 4923 51619
rect 4979 51580 5031 51619
rect 7247 51580 7299 51619
rect 7355 51580 7407 51619
rect 7463 51580 7515 51619
rect 7571 51580 7623 51619
rect 7679 51580 7731 51619
rect 9947 51580 9999 51619
rect 10055 51580 10107 51619
rect 4871 51567 4923 51580
rect 4979 51567 5031 51580
rect 7247 51567 7299 51580
rect 7355 51567 7407 51580
rect 7463 51567 7515 51580
rect 7571 51567 7623 51580
rect 7679 51567 7731 51580
rect 9947 51567 9999 51580
rect 10055 51567 10107 51580
rect 4871 51498 4923 51511
rect 4979 51498 5031 51511
rect 7247 51498 7299 51511
rect 7355 51498 7407 51511
rect 7463 51498 7515 51511
rect 7571 51498 7623 51511
rect 7679 51498 7731 51511
rect 9947 51498 9999 51511
rect 10055 51498 10107 51511
rect 4871 51459 4923 51498
rect 4979 51459 5031 51498
rect 7247 51459 7299 51498
rect 7355 51459 7407 51498
rect 7463 51459 7515 51498
rect 7571 51459 7623 51498
rect 7679 51459 7731 51498
rect 9947 51459 9999 51498
rect 10055 51459 10107 51498
rect 3161 51154 3162 51206
rect 3162 51154 3213 51206
rect 3269 51154 3321 51206
rect 3377 51203 3424 51206
rect 3424 51203 3429 51206
rect 3485 51203 3537 51206
rect 3593 51203 3645 51206
rect 3701 51203 3753 51206
rect 3809 51203 3861 51206
rect 3917 51203 3969 51206
rect 4025 51203 4077 51206
rect 4133 51203 4185 51206
rect 4241 51203 4293 51206
rect 4349 51203 4401 51206
rect 4457 51203 4509 51206
rect 4565 51203 4617 51206
rect 4673 51203 4725 51206
rect 5138 51203 5190 51206
rect 5246 51203 5298 51206
rect 5354 51203 5406 51206
rect 5462 51203 5514 51206
rect 5570 51203 5622 51206
rect 5678 51203 5730 51206
rect 5786 51203 5838 51206
rect 5894 51203 5946 51206
rect 6002 51203 6054 51206
rect 6110 51203 6162 51206
rect 6218 51203 6270 51206
rect 6326 51203 6378 51206
rect 6434 51203 6486 51206
rect 6542 51203 6594 51206
rect 6650 51203 6702 51206
rect 6758 51203 6810 51206
rect 6866 51203 6918 51206
rect 6974 51203 7026 51206
rect 7082 51203 7134 51206
rect 7844 51203 7896 51206
rect 7952 51203 8004 51206
rect 8060 51203 8112 51206
rect 8168 51203 8220 51206
rect 8276 51203 8328 51206
rect 8384 51203 8436 51206
rect 8492 51203 8544 51206
rect 8600 51203 8652 51206
rect 8708 51203 8760 51206
rect 8816 51203 8868 51206
rect 8924 51203 8976 51206
rect 9032 51203 9084 51206
rect 9140 51203 9192 51206
rect 9248 51203 9300 51206
rect 9356 51203 9408 51206
rect 9464 51203 9516 51206
rect 9572 51203 9624 51206
rect 9680 51203 9732 51206
rect 9788 51203 9840 51206
rect 10253 51203 10305 51206
rect 10361 51203 10413 51206
rect 10469 51203 10521 51206
rect 10577 51203 10629 51206
rect 10685 51203 10737 51206
rect 10793 51203 10845 51206
rect 10901 51203 10953 51206
rect 11009 51203 11061 51206
rect 11117 51203 11169 51206
rect 11225 51203 11277 51206
rect 11333 51203 11385 51206
rect 11441 51203 11493 51206
rect 11549 51203 11554 51206
rect 11554 51203 11601 51206
rect 3377 51154 3429 51203
rect 3485 51154 3537 51203
rect 3593 51154 3645 51203
rect 3701 51154 3753 51203
rect 3809 51154 3861 51203
rect 3917 51154 3969 51203
rect 4025 51154 4077 51203
rect 4133 51154 4185 51203
rect 4241 51154 4293 51203
rect 4349 51154 4401 51203
rect 4457 51154 4509 51203
rect 4565 51154 4617 51203
rect 4673 51154 4725 51203
rect 5138 51154 5190 51203
rect 5246 51154 5298 51203
rect 5354 51154 5406 51203
rect 5462 51154 5514 51203
rect 5570 51154 5622 51203
rect 5678 51154 5730 51203
rect 5786 51154 5838 51203
rect 5894 51154 5946 51203
rect 6002 51154 6054 51203
rect 6110 51154 6162 51203
rect 6218 51154 6270 51203
rect 6326 51154 6378 51203
rect 6434 51154 6486 51203
rect 6542 51154 6594 51203
rect 6650 51154 6702 51203
rect 6758 51154 6810 51203
rect 6866 51154 6918 51203
rect 6974 51154 7026 51203
rect 7082 51154 7134 51203
rect 7844 51154 7896 51203
rect 7952 51154 8004 51203
rect 8060 51154 8112 51203
rect 8168 51154 8220 51203
rect 8276 51154 8328 51203
rect 8384 51154 8436 51203
rect 8492 51154 8544 51203
rect 8600 51154 8652 51203
rect 8708 51154 8760 51203
rect 8816 51154 8868 51203
rect 8924 51154 8976 51203
rect 9032 51154 9084 51203
rect 9140 51154 9192 51203
rect 9248 51154 9300 51203
rect 9356 51154 9408 51203
rect 9464 51154 9516 51203
rect 9572 51154 9624 51203
rect 9680 51154 9732 51203
rect 9788 51154 9840 51203
rect 10253 51154 10305 51203
rect 10361 51154 10413 51203
rect 10469 51154 10521 51203
rect 10577 51154 10629 51203
rect 10685 51154 10737 51203
rect 10793 51154 10845 51203
rect 10901 51154 10953 51203
rect 11009 51154 11061 51203
rect 11117 51154 11169 51203
rect 11225 51154 11277 51203
rect 11333 51154 11385 51203
rect 11441 51154 11493 51203
rect 11549 51154 11601 51203
rect 11657 51154 11709 51206
rect 11765 51154 11816 51206
rect 11816 51154 11817 51206
rect 3161 51046 3162 51098
rect 3162 51046 3213 51098
rect 3269 51046 3321 51098
rect 3377 51095 3429 51098
rect 3485 51095 3537 51098
rect 3593 51095 3645 51098
rect 3701 51095 3753 51098
rect 3809 51095 3861 51098
rect 3917 51095 3969 51098
rect 4025 51095 4077 51098
rect 4133 51095 4185 51098
rect 4241 51095 4293 51098
rect 4349 51095 4401 51098
rect 4457 51095 4509 51098
rect 4565 51095 4617 51098
rect 4673 51095 4725 51098
rect 5138 51095 5190 51098
rect 5246 51095 5298 51098
rect 5354 51095 5406 51098
rect 5462 51095 5514 51098
rect 5570 51095 5622 51098
rect 5678 51095 5730 51098
rect 5786 51095 5838 51098
rect 5894 51095 5946 51098
rect 6002 51095 6054 51098
rect 6110 51095 6162 51098
rect 6218 51095 6270 51098
rect 6326 51095 6378 51098
rect 6434 51095 6486 51098
rect 6542 51095 6594 51098
rect 6650 51095 6702 51098
rect 6758 51095 6810 51098
rect 6866 51095 6918 51098
rect 6974 51095 7026 51098
rect 7082 51095 7134 51098
rect 7844 51095 7896 51098
rect 7952 51095 8004 51098
rect 8060 51095 8112 51098
rect 8168 51095 8220 51098
rect 8276 51095 8328 51098
rect 8384 51095 8436 51098
rect 8492 51095 8544 51098
rect 8600 51095 8652 51098
rect 8708 51095 8760 51098
rect 8816 51095 8868 51098
rect 8924 51095 8976 51098
rect 9032 51095 9084 51098
rect 9140 51095 9192 51098
rect 9248 51095 9300 51098
rect 9356 51095 9408 51098
rect 9464 51095 9516 51098
rect 9572 51095 9624 51098
rect 9680 51095 9732 51098
rect 9788 51095 9840 51098
rect 10253 51095 10305 51098
rect 10361 51095 10413 51098
rect 10469 51095 10521 51098
rect 10577 51095 10629 51098
rect 10685 51095 10737 51098
rect 10793 51095 10845 51098
rect 10901 51095 10953 51098
rect 11009 51095 11061 51098
rect 11117 51095 11169 51098
rect 11225 51095 11277 51098
rect 11333 51095 11385 51098
rect 11441 51095 11493 51098
rect 11549 51095 11601 51098
rect 3377 51049 3429 51095
rect 3485 51049 3537 51095
rect 3593 51049 3645 51095
rect 3701 51049 3753 51095
rect 3809 51049 3861 51095
rect 3917 51049 3969 51095
rect 4025 51049 4077 51095
rect 4133 51049 4185 51095
rect 4241 51049 4293 51095
rect 4349 51049 4401 51095
rect 4457 51049 4509 51095
rect 4565 51049 4617 51095
rect 4673 51049 4725 51095
rect 5138 51049 5190 51095
rect 5246 51049 5298 51095
rect 5354 51049 5406 51095
rect 5462 51049 5514 51095
rect 5570 51049 5622 51095
rect 5678 51049 5730 51095
rect 5786 51049 5838 51095
rect 5894 51049 5946 51095
rect 6002 51049 6054 51095
rect 6110 51049 6162 51095
rect 6218 51049 6270 51095
rect 6326 51049 6378 51095
rect 6434 51049 6486 51095
rect 6542 51049 6594 51095
rect 6650 51049 6702 51095
rect 6758 51049 6810 51095
rect 6866 51049 6918 51095
rect 6974 51049 7026 51095
rect 7082 51049 7134 51095
rect 7844 51049 7896 51095
rect 7952 51049 8004 51095
rect 8060 51049 8112 51095
rect 8168 51049 8220 51095
rect 8276 51049 8328 51095
rect 8384 51049 8436 51095
rect 8492 51049 8544 51095
rect 8600 51049 8652 51095
rect 8708 51049 8760 51095
rect 8816 51049 8868 51095
rect 8924 51049 8976 51095
rect 9032 51049 9084 51095
rect 9140 51049 9192 51095
rect 9248 51049 9300 51095
rect 9356 51049 9408 51095
rect 9464 51049 9516 51095
rect 9572 51049 9624 51095
rect 9680 51049 9732 51095
rect 9788 51049 9840 51095
rect 10253 51049 10305 51095
rect 10361 51049 10413 51095
rect 10469 51049 10521 51095
rect 10577 51049 10629 51095
rect 10685 51049 10737 51095
rect 10793 51049 10845 51095
rect 10901 51049 10953 51095
rect 11009 51049 11061 51095
rect 11117 51049 11169 51095
rect 11225 51049 11277 51095
rect 11333 51049 11385 51095
rect 11441 51049 11493 51095
rect 11549 51049 11601 51095
rect 3377 51046 3429 51049
rect 3485 51046 3537 51049
rect 3593 51046 3645 51049
rect 3701 51046 3753 51049
rect 3809 51046 3861 51049
rect 3917 51046 3969 51049
rect 4025 51046 4077 51049
rect 4133 51046 4185 51049
rect 4241 51046 4293 51049
rect 4349 51046 4401 51049
rect 4457 51046 4509 51049
rect 4565 51046 4617 51049
rect 4673 51046 4725 51049
rect 5138 51046 5190 51049
rect 5246 51046 5298 51049
rect 5354 51046 5406 51049
rect 5462 51046 5514 51049
rect 5570 51046 5622 51049
rect 5678 51046 5730 51049
rect 5786 51046 5838 51049
rect 5894 51046 5946 51049
rect 6002 51046 6054 51049
rect 6110 51046 6162 51049
rect 6218 51046 6270 51049
rect 6326 51046 6378 51049
rect 6434 51046 6486 51049
rect 6542 51046 6594 51049
rect 6650 51046 6702 51049
rect 6758 51046 6810 51049
rect 6866 51046 6918 51049
rect 6974 51046 7026 51049
rect 7082 51046 7134 51049
rect 7844 51046 7896 51049
rect 7952 51046 8004 51049
rect 8060 51046 8112 51049
rect 8168 51046 8220 51049
rect 8276 51046 8328 51049
rect 8384 51046 8436 51049
rect 8492 51046 8544 51049
rect 8600 51046 8652 51049
rect 8708 51046 8760 51049
rect 8816 51046 8868 51049
rect 8924 51046 8976 51049
rect 9032 51046 9084 51049
rect 9140 51046 9192 51049
rect 9248 51046 9300 51049
rect 9356 51046 9408 51049
rect 9464 51046 9516 51049
rect 9572 51046 9624 51049
rect 9680 51046 9732 51049
rect 9788 51046 9840 51049
rect 10253 51046 10305 51049
rect 10361 51046 10413 51049
rect 10469 51046 10521 51049
rect 10577 51046 10629 51049
rect 10685 51046 10737 51049
rect 10793 51046 10845 51049
rect 10901 51046 10953 51049
rect 11009 51046 11061 51049
rect 11117 51046 11169 51049
rect 11225 51046 11277 51049
rect 11333 51046 11385 51049
rect 11441 51046 11493 51049
rect 11549 51046 11601 51049
rect 11657 51046 11709 51098
rect 11765 51046 11816 51098
rect 11816 51046 11817 51098
rect 3161 50938 3162 50990
rect 3162 50938 3213 50990
rect 3269 50938 3321 50990
rect 3377 50941 3429 50990
rect 3485 50941 3537 50990
rect 3593 50941 3645 50990
rect 3701 50941 3753 50990
rect 3809 50941 3861 50990
rect 3917 50941 3969 50990
rect 4025 50941 4077 50990
rect 4133 50941 4185 50990
rect 4241 50941 4293 50990
rect 4349 50941 4401 50990
rect 4457 50941 4509 50990
rect 4565 50941 4617 50990
rect 4673 50941 4725 50990
rect 5138 50941 5190 50990
rect 5246 50941 5298 50990
rect 5354 50941 5406 50990
rect 5462 50941 5514 50990
rect 5570 50941 5622 50990
rect 5678 50941 5730 50990
rect 5786 50941 5838 50990
rect 5894 50941 5946 50990
rect 6002 50941 6054 50990
rect 6110 50941 6162 50990
rect 6218 50941 6270 50990
rect 6326 50941 6378 50990
rect 6434 50941 6486 50990
rect 6542 50941 6594 50990
rect 6650 50941 6702 50990
rect 6758 50941 6810 50990
rect 6866 50941 6918 50990
rect 6974 50941 7026 50990
rect 7082 50941 7134 50990
rect 7844 50941 7896 50990
rect 7952 50941 8004 50990
rect 8060 50941 8112 50990
rect 8168 50941 8220 50990
rect 8276 50941 8328 50990
rect 8384 50941 8436 50990
rect 8492 50941 8544 50990
rect 8600 50941 8652 50990
rect 8708 50941 8760 50990
rect 8816 50941 8868 50990
rect 8924 50941 8976 50990
rect 9032 50941 9084 50990
rect 9140 50941 9192 50990
rect 9248 50941 9300 50990
rect 9356 50941 9408 50990
rect 9464 50941 9516 50990
rect 9572 50941 9624 50990
rect 9680 50941 9732 50990
rect 9788 50941 9840 50990
rect 10253 50941 10305 50990
rect 10361 50941 10413 50990
rect 10469 50941 10521 50990
rect 10577 50941 10629 50990
rect 10685 50941 10737 50990
rect 10793 50941 10845 50990
rect 10901 50941 10953 50990
rect 11009 50941 11061 50990
rect 11117 50941 11169 50990
rect 11225 50941 11277 50990
rect 11333 50941 11385 50990
rect 11441 50941 11493 50990
rect 11549 50941 11601 50990
rect 3377 50938 3424 50941
rect 3424 50938 3429 50941
rect 3485 50938 3537 50941
rect 3593 50938 3645 50941
rect 3701 50938 3753 50941
rect 3809 50938 3861 50941
rect 3917 50938 3969 50941
rect 4025 50938 4077 50941
rect 4133 50938 4185 50941
rect 4241 50938 4293 50941
rect 4349 50938 4401 50941
rect 4457 50938 4509 50941
rect 4565 50938 4617 50941
rect 4673 50938 4725 50941
rect 5138 50938 5190 50941
rect 5246 50938 5298 50941
rect 5354 50938 5406 50941
rect 5462 50938 5514 50941
rect 5570 50938 5622 50941
rect 5678 50938 5730 50941
rect 5786 50938 5838 50941
rect 5894 50938 5946 50941
rect 6002 50938 6054 50941
rect 6110 50938 6162 50941
rect 6218 50938 6270 50941
rect 6326 50938 6378 50941
rect 6434 50938 6486 50941
rect 6542 50938 6594 50941
rect 6650 50938 6702 50941
rect 6758 50938 6810 50941
rect 6866 50938 6918 50941
rect 6974 50938 7026 50941
rect 7082 50938 7134 50941
rect 7844 50938 7896 50941
rect 7952 50938 8004 50941
rect 8060 50938 8112 50941
rect 8168 50938 8220 50941
rect 8276 50938 8328 50941
rect 8384 50938 8436 50941
rect 8492 50938 8544 50941
rect 8600 50938 8652 50941
rect 8708 50938 8760 50941
rect 8816 50938 8868 50941
rect 8924 50938 8976 50941
rect 9032 50938 9084 50941
rect 9140 50938 9192 50941
rect 9248 50938 9300 50941
rect 9356 50938 9408 50941
rect 9464 50938 9516 50941
rect 9572 50938 9624 50941
rect 9680 50938 9732 50941
rect 9788 50938 9840 50941
rect 10253 50938 10305 50941
rect 10361 50938 10413 50941
rect 10469 50938 10521 50941
rect 10577 50938 10629 50941
rect 10685 50938 10737 50941
rect 10793 50938 10845 50941
rect 10901 50938 10953 50941
rect 11009 50938 11061 50941
rect 11117 50938 11169 50941
rect 11225 50938 11277 50941
rect 11333 50938 11385 50941
rect 11441 50938 11493 50941
rect 11549 50938 11554 50941
rect 11554 50938 11601 50941
rect 11657 50938 11709 50990
rect 11765 50938 11816 50990
rect 11816 50938 11817 50990
rect 4871 50646 4923 50685
rect 4979 50646 5031 50685
rect 7247 50646 7299 50685
rect 7355 50646 7407 50685
rect 7463 50646 7515 50685
rect 7571 50646 7623 50685
rect 7679 50646 7731 50685
rect 9947 50646 9999 50685
rect 10055 50646 10107 50685
rect 4871 50633 4923 50646
rect 4979 50633 5031 50646
rect 7247 50633 7299 50646
rect 7355 50633 7407 50646
rect 7463 50633 7515 50646
rect 7571 50633 7623 50646
rect 7679 50633 7731 50646
rect 9947 50633 9999 50646
rect 10055 50633 10107 50646
rect 4871 50564 4923 50577
rect 4979 50564 5031 50577
rect 7247 50564 7299 50577
rect 7355 50564 7407 50577
rect 7463 50564 7515 50577
rect 7571 50564 7623 50577
rect 7679 50564 7731 50577
rect 9947 50564 9999 50577
rect 10055 50564 10107 50577
rect 4871 50525 4923 50564
rect 4979 50525 5031 50564
rect 7247 50525 7299 50564
rect 7355 50525 7407 50564
rect 7463 50525 7515 50564
rect 7571 50525 7623 50564
rect 7679 50525 7731 50564
rect 9947 50525 9999 50564
rect 10055 50525 10107 50564
rect 3161 50220 3162 50272
rect 3162 50220 3213 50272
rect 3269 50220 3321 50272
rect 3377 50269 3424 50272
rect 3424 50269 3429 50272
rect 3485 50269 3537 50272
rect 3593 50269 3645 50272
rect 3701 50269 3753 50272
rect 3809 50269 3861 50272
rect 3917 50269 3969 50272
rect 4025 50269 4077 50272
rect 4133 50269 4185 50272
rect 4241 50269 4293 50272
rect 4349 50269 4401 50272
rect 4457 50269 4509 50272
rect 4565 50269 4617 50272
rect 4673 50269 4725 50272
rect 5138 50269 5190 50272
rect 5246 50269 5298 50272
rect 5354 50269 5406 50272
rect 5462 50269 5514 50272
rect 5570 50269 5622 50272
rect 5678 50269 5730 50272
rect 5786 50269 5838 50272
rect 5894 50269 5946 50272
rect 6002 50269 6054 50272
rect 6110 50269 6162 50272
rect 6218 50269 6270 50272
rect 6326 50269 6378 50272
rect 6434 50269 6486 50272
rect 6542 50269 6594 50272
rect 6650 50269 6702 50272
rect 6758 50269 6810 50272
rect 6866 50269 6918 50272
rect 6974 50269 7026 50272
rect 7082 50269 7134 50272
rect 7844 50269 7896 50272
rect 7952 50269 8004 50272
rect 8060 50269 8112 50272
rect 8168 50269 8220 50272
rect 8276 50269 8328 50272
rect 8384 50269 8436 50272
rect 8492 50269 8544 50272
rect 8600 50269 8652 50272
rect 8708 50269 8760 50272
rect 8816 50269 8868 50272
rect 8924 50269 8976 50272
rect 9032 50269 9084 50272
rect 9140 50269 9192 50272
rect 9248 50269 9300 50272
rect 9356 50269 9408 50272
rect 9464 50269 9516 50272
rect 9572 50269 9624 50272
rect 9680 50269 9732 50272
rect 9788 50269 9840 50272
rect 10253 50269 10305 50272
rect 10361 50269 10413 50272
rect 10469 50269 10521 50272
rect 10577 50269 10629 50272
rect 10685 50269 10737 50272
rect 10793 50269 10845 50272
rect 10901 50269 10953 50272
rect 11009 50269 11061 50272
rect 11117 50269 11169 50272
rect 11225 50269 11277 50272
rect 11333 50269 11385 50272
rect 11441 50269 11493 50272
rect 11549 50269 11554 50272
rect 11554 50269 11601 50272
rect 3377 50220 3429 50269
rect 3485 50220 3537 50269
rect 3593 50220 3645 50269
rect 3701 50220 3753 50269
rect 3809 50220 3861 50269
rect 3917 50220 3969 50269
rect 4025 50220 4077 50269
rect 4133 50220 4185 50269
rect 4241 50220 4293 50269
rect 4349 50220 4401 50269
rect 4457 50220 4509 50269
rect 4565 50220 4617 50269
rect 4673 50220 4725 50269
rect 5138 50220 5190 50269
rect 5246 50220 5298 50269
rect 5354 50220 5406 50269
rect 5462 50220 5514 50269
rect 5570 50220 5622 50269
rect 5678 50220 5730 50269
rect 5786 50220 5838 50269
rect 5894 50220 5946 50269
rect 6002 50220 6054 50269
rect 6110 50220 6162 50269
rect 6218 50220 6270 50269
rect 6326 50220 6378 50269
rect 6434 50220 6486 50269
rect 6542 50220 6594 50269
rect 6650 50220 6702 50269
rect 6758 50220 6810 50269
rect 6866 50220 6918 50269
rect 6974 50220 7026 50269
rect 7082 50220 7134 50269
rect 7844 50220 7896 50269
rect 7952 50220 8004 50269
rect 8060 50220 8112 50269
rect 8168 50220 8220 50269
rect 8276 50220 8328 50269
rect 8384 50220 8436 50269
rect 8492 50220 8544 50269
rect 8600 50220 8652 50269
rect 8708 50220 8760 50269
rect 8816 50220 8868 50269
rect 8924 50220 8976 50269
rect 9032 50220 9084 50269
rect 9140 50220 9192 50269
rect 9248 50220 9300 50269
rect 9356 50220 9408 50269
rect 9464 50220 9516 50269
rect 9572 50220 9624 50269
rect 9680 50220 9732 50269
rect 9788 50220 9840 50269
rect 10253 50220 10305 50269
rect 10361 50220 10413 50269
rect 10469 50220 10521 50269
rect 10577 50220 10629 50269
rect 10685 50220 10737 50269
rect 10793 50220 10845 50269
rect 10901 50220 10953 50269
rect 11009 50220 11061 50269
rect 11117 50220 11169 50269
rect 11225 50220 11277 50269
rect 11333 50220 11385 50269
rect 11441 50220 11493 50269
rect 11549 50220 11601 50269
rect 11657 50220 11709 50272
rect 11765 50220 11816 50272
rect 11816 50220 11817 50272
rect 3161 50112 3162 50164
rect 3162 50112 3213 50164
rect 3269 50112 3321 50164
rect 3377 50161 3429 50164
rect 3485 50161 3537 50164
rect 3593 50161 3645 50164
rect 3701 50161 3753 50164
rect 3809 50161 3861 50164
rect 3917 50161 3969 50164
rect 4025 50161 4077 50164
rect 4133 50161 4185 50164
rect 4241 50161 4293 50164
rect 4349 50161 4401 50164
rect 4457 50161 4509 50164
rect 4565 50161 4617 50164
rect 4673 50161 4725 50164
rect 5138 50161 5190 50164
rect 5246 50161 5298 50164
rect 5354 50161 5406 50164
rect 5462 50161 5514 50164
rect 5570 50161 5622 50164
rect 5678 50161 5730 50164
rect 5786 50161 5838 50164
rect 5894 50161 5946 50164
rect 6002 50161 6054 50164
rect 6110 50161 6162 50164
rect 6218 50161 6270 50164
rect 6326 50161 6378 50164
rect 6434 50161 6486 50164
rect 6542 50161 6594 50164
rect 6650 50161 6702 50164
rect 6758 50161 6810 50164
rect 6866 50161 6918 50164
rect 6974 50161 7026 50164
rect 7082 50161 7134 50164
rect 7844 50161 7896 50164
rect 7952 50161 8004 50164
rect 8060 50161 8112 50164
rect 8168 50161 8220 50164
rect 8276 50161 8328 50164
rect 8384 50161 8436 50164
rect 8492 50161 8544 50164
rect 8600 50161 8652 50164
rect 8708 50161 8760 50164
rect 8816 50161 8868 50164
rect 8924 50161 8976 50164
rect 9032 50161 9084 50164
rect 9140 50161 9192 50164
rect 9248 50161 9300 50164
rect 9356 50161 9408 50164
rect 9464 50161 9516 50164
rect 9572 50161 9624 50164
rect 9680 50161 9732 50164
rect 9788 50161 9840 50164
rect 10253 50161 10305 50164
rect 10361 50161 10413 50164
rect 10469 50161 10521 50164
rect 10577 50161 10629 50164
rect 10685 50161 10737 50164
rect 10793 50161 10845 50164
rect 10901 50161 10953 50164
rect 11009 50161 11061 50164
rect 11117 50161 11169 50164
rect 11225 50161 11277 50164
rect 11333 50161 11385 50164
rect 11441 50161 11493 50164
rect 11549 50161 11601 50164
rect 3377 50115 3429 50161
rect 3485 50115 3537 50161
rect 3593 50115 3645 50161
rect 3701 50115 3753 50161
rect 3809 50115 3861 50161
rect 3917 50115 3969 50161
rect 4025 50115 4077 50161
rect 4133 50115 4185 50161
rect 4241 50115 4293 50161
rect 4349 50115 4401 50161
rect 4457 50115 4509 50161
rect 4565 50115 4617 50161
rect 4673 50115 4725 50161
rect 5138 50115 5190 50161
rect 5246 50115 5298 50161
rect 5354 50115 5406 50161
rect 5462 50115 5514 50161
rect 5570 50115 5622 50161
rect 5678 50115 5730 50161
rect 5786 50115 5838 50161
rect 5894 50115 5946 50161
rect 6002 50115 6054 50161
rect 6110 50115 6162 50161
rect 6218 50115 6270 50161
rect 6326 50115 6378 50161
rect 6434 50115 6486 50161
rect 6542 50115 6594 50161
rect 6650 50115 6702 50161
rect 6758 50115 6810 50161
rect 6866 50115 6918 50161
rect 6974 50115 7026 50161
rect 7082 50115 7134 50161
rect 7844 50115 7896 50161
rect 7952 50115 8004 50161
rect 8060 50115 8112 50161
rect 8168 50115 8220 50161
rect 8276 50115 8328 50161
rect 8384 50115 8436 50161
rect 8492 50115 8544 50161
rect 8600 50115 8652 50161
rect 8708 50115 8760 50161
rect 8816 50115 8868 50161
rect 8924 50115 8976 50161
rect 9032 50115 9084 50161
rect 9140 50115 9192 50161
rect 9248 50115 9300 50161
rect 9356 50115 9408 50161
rect 9464 50115 9516 50161
rect 9572 50115 9624 50161
rect 9680 50115 9732 50161
rect 9788 50115 9840 50161
rect 10253 50115 10305 50161
rect 10361 50115 10413 50161
rect 10469 50115 10521 50161
rect 10577 50115 10629 50161
rect 10685 50115 10737 50161
rect 10793 50115 10845 50161
rect 10901 50115 10953 50161
rect 11009 50115 11061 50161
rect 11117 50115 11169 50161
rect 11225 50115 11277 50161
rect 11333 50115 11385 50161
rect 11441 50115 11493 50161
rect 11549 50115 11601 50161
rect 3377 50112 3429 50115
rect 3485 50112 3537 50115
rect 3593 50112 3645 50115
rect 3701 50112 3753 50115
rect 3809 50112 3861 50115
rect 3917 50112 3969 50115
rect 4025 50112 4077 50115
rect 4133 50112 4185 50115
rect 4241 50112 4293 50115
rect 4349 50112 4401 50115
rect 4457 50112 4509 50115
rect 4565 50112 4617 50115
rect 4673 50112 4725 50115
rect 5138 50112 5190 50115
rect 5246 50112 5298 50115
rect 5354 50112 5406 50115
rect 5462 50112 5514 50115
rect 5570 50112 5622 50115
rect 5678 50112 5730 50115
rect 5786 50112 5838 50115
rect 5894 50112 5946 50115
rect 6002 50112 6054 50115
rect 6110 50112 6162 50115
rect 6218 50112 6270 50115
rect 6326 50112 6378 50115
rect 6434 50112 6486 50115
rect 6542 50112 6594 50115
rect 6650 50112 6702 50115
rect 6758 50112 6810 50115
rect 6866 50112 6918 50115
rect 6974 50112 7026 50115
rect 7082 50112 7134 50115
rect 7844 50112 7896 50115
rect 7952 50112 8004 50115
rect 8060 50112 8112 50115
rect 8168 50112 8220 50115
rect 8276 50112 8328 50115
rect 8384 50112 8436 50115
rect 8492 50112 8544 50115
rect 8600 50112 8652 50115
rect 8708 50112 8760 50115
rect 8816 50112 8868 50115
rect 8924 50112 8976 50115
rect 9032 50112 9084 50115
rect 9140 50112 9192 50115
rect 9248 50112 9300 50115
rect 9356 50112 9408 50115
rect 9464 50112 9516 50115
rect 9572 50112 9624 50115
rect 9680 50112 9732 50115
rect 9788 50112 9840 50115
rect 10253 50112 10305 50115
rect 10361 50112 10413 50115
rect 10469 50112 10521 50115
rect 10577 50112 10629 50115
rect 10685 50112 10737 50115
rect 10793 50112 10845 50115
rect 10901 50112 10953 50115
rect 11009 50112 11061 50115
rect 11117 50112 11169 50115
rect 11225 50112 11277 50115
rect 11333 50112 11385 50115
rect 11441 50112 11493 50115
rect 11549 50112 11601 50115
rect 11657 50112 11709 50164
rect 11765 50112 11816 50164
rect 11816 50112 11817 50164
rect 3161 50004 3162 50056
rect 3162 50004 3213 50056
rect 3269 50004 3321 50056
rect 3377 50007 3429 50056
rect 3485 50007 3537 50056
rect 3593 50007 3645 50056
rect 3701 50007 3753 50056
rect 3809 50007 3861 50056
rect 3917 50007 3969 50056
rect 4025 50007 4077 50056
rect 4133 50007 4185 50056
rect 4241 50007 4293 50056
rect 4349 50007 4401 50056
rect 4457 50007 4509 50056
rect 4565 50007 4617 50056
rect 4673 50007 4725 50056
rect 5138 50007 5190 50056
rect 5246 50007 5298 50056
rect 5354 50007 5406 50056
rect 5462 50007 5514 50056
rect 5570 50007 5622 50056
rect 5678 50007 5730 50056
rect 5786 50007 5838 50056
rect 5894 50007 5946 50056
rect 6002 50007 6054 50056
rect 6110 50007 6162 50056
rect 6218 50007 6270 50056
rect 6326 50007 6378 50056
rect 6434 50007 6486 50056
rect 6542 50007 6594 50056
rect 6650 50007 6702 50056
rect 6758 50007 6810 50056
rect 6866 50007 6918 50056
rect 6974 50007 7026 50056
rect 7082 50007 7134 50056
rect 7844 50007 7896 50056
rect 7952 50007 8004 50056
rect 8060 50007 8112 50056
rect 8168 50007 8220 50056
rect 8276 50007 8328 50056
rect 8384 50007 8436 50056
rect 8492 50007 8544 50056
rect 8600 50007 8652 50056
rect 8708 50007 8760 50056
rect 8816 50007 8868 50056
rect 8924 50007 8976 50056
rect 9032 50007 9084 50056
rect 9140 50007 9192 50056
rect 9248 50007 9300 50056
rect 9356 50007 9408 50056
rect 9464 50007 9516 50056
rect 9572 50007 9624 50056
rect 9680 50007 9732 50056
rect 9788 50007 9840 50056
rect 10253 50007 10305 50056
rect 10361 50007 10413 50056
rect 10469 50007 10521 50056
rect 10577 50007 10629 50056
rect 10685 50007 10737 50056
rect 10793 50007 10845 50056
rect 10901 50007 10953 50056
rect 11009 50007 11061 50056
rect 11117 50007 11169 50056
rect 11225 50007 11277 50056
rect 11333 50007 11385 50056
rect 11441 50007 11493 50056
rect 11549 50007 11601 50056
rect 3377 50004 3424 50007
rect 3424 50004 3429 50007
rect 3485 50004 3537 50007
rect 3593 50004 3645 50007
rect 3701 50004 3753 50007
rect 3809 50004 3861 50007
rect 3917 50004 3969 50007
rect 4025 50004 4077 50007
rect 4133 50004 4185 50007
rect 4241 50004 4293 50007
rect 4349 50004 4401 50007
rect 4457 50004 4509 50007
rect 4565 50004 4617 50007
rect 4673 50004 4725 50007
rect 5138 50004 5190 50007
rect 5246 50004 5298 50007
rect 5354 50004 5406 50007
rect 5462 50004 5514 50007
rect 5570 50004 5622 50007
rect 5678 50004 5730 50007
rect 5786 50004 5838 50007
rect 5894 50004 5946 50007
rect 6002 50004 6054 50007
rect 6110 50004 6162 50007
rect 6218 50004 6270 50007
rect 6326 50004 6378 50007
rect 6434 50004 6486 50007
rect 6542 50004 6594 50007
rect 6650 50004 6702 50007
rect 6758 50004 6810 50007
rect 6866 50004 6918 50007
rect 6974 50004 7026 50007
rect 7082 50004 7134 50007
rect 7844 50004 7896 50007
rect 7952 50004 8004 50007
rect 8060 50004 8112 50007
rect 8168 50004 8220 50007
rect 8276 50004 8328 50007
rect 8384 50004 8436 50007
rect 8492 50004 8544 50007
rect 8600 50004 8652 50007
rect 8708 50004 8760 50007
rect 8816 50004 8868 50007
rect 8924 50004 8976 50007
rect 9032 50004 9084 50007
rect 9140 50004 9192 50007
rect 9248 50004 9300 50007
rect 9356 50004 9408 50007
rect 9464 50004 9516 50007
rect 9572 50004 9624 50007
rect 9680 50004 9732 50007
rect 9788 50004 9840 50007
rect 10253 50004 10305 50007
rect 10361 50004 10413 50007
rect 10469 50004 10521 50007
rect 10577 50004 10629 50007
rect 10685 50004 10737 50007
rect 10793 50004 10845 50007
rect 10901 50004 10953 50007
rect 11009 50004 11061 50007
rect 11117 50004 11169 50007
rect 11225 50004 11277 50007
rect 11333 50004 11385 50007
rect 11441 50004 11493 50007
rect 11549 50004 11554 50007
rect 11554 50004 11601 50007
rect 11657 50004 11709 50056
rect 11765 50004 11816 50056
rect 11816 50004 11817 50056
rect 4871 49712 4923 49751
rect 4979 49712 5031 49751
rect 7247 49712 7299 49751
rect 7355 49712 7407 49751
rect 7463 49712 7515 49751
rect 7571 49712 7623 49751
rect 7679 49712 7731 49751
rect 9947 49712 9999 49751
rect 10055 49712 10107 49751
rect 4871 49699 4923 49712
rect 4979 49699 5031 49712
rect 7247 49699 7299 49712
rect 7355 49699 7407 49712
rect 7463 49699 7515 49712
rect 7571 49699 7623 49712
rect 7679 49699 7731 49712
rect 9947 49699 9999 49712
rect 10055 49699 10107 49712
rect 4871 49630 4923 49643
rect 4979 49630 5031 49643
rect 7247 49630 7299 49643
rect 7355 49630 7407 49643
rect 7463 49630 7515 49643
rect 7571 49630 7623 49643
rect 7679 49630 7731 49643
rect 9947 49630 9999 49643
rect 10055 49630 10107 49643
rect 4871 49591 4923 49630
rect 4979 49591 5031 49630
rect 7247 49591 7299 49630
rect 7355 49591 7407 49630
rect 7463 49591 7515 49630
rect 7571 49591 7623 49630
rect 7679 49591 7731 49630
rect 9947 49591 9999 49630
rect 10055 49591 10107 49630
rect 3161 49286 3162 49338
rect 3162 49286 3213 49338
rect 3269 49286 3321 49338
rect 3377 49335 3424 49338
rect 3424 49335 3429 49338
rect 3485 49335 3537 49338
rect 3593 49335 3645 49338
rect 3701 49335 3753 49338
rect 3809 49335 3861 49338
rect 3917 49335 3969 49338
rect 4025 49335 4077 49338
rect 4133 49335 4185 49338
rect 4241 49335 4293 49338
rect 4349 49335 4401 49338
rect 4457 49335 4509 49338
rect 4565 49335 4617 49338
rect 4673 49335 4725 49338
rect 5138 49335 5190 49338
rect 5246 49335 5298 49338
rect 5354 49335 5406 49338
rect 5462 49335 5514 49338
rect 5570 49335 5622 49338
rect 5678 49335 5730 49338
rect 5786 49335 5838 49338
rect 5894 49335 5946 49338
rect 6002 49335 6054 49338
rect 6110 49335 6162 49338
rect 6218 49335 6270 49338
rect 6326 49335 6378 49338
rect 6434 49335 6486 49338
rect 6542 49335 6594 49338
rect 6650 49335 6702 49338
rect 6758 49335 6810 49338
rect 6866 49335 6918 49338
rect 6974 49335 7026 49338
rect 7082 49335 7134 49338
rect 7844 49335 7896 49338
rect 7952 49335 8004 49338
rect 8060 49335 8112 49338
rect 8168 49335 8220 49338
rect 8276 49335 8328 49338
rect 8384 49335 8436 49338
rect 8492 49335 8544 49338
rect 8600 49335 8652 49338
rect 8708 49335 8760 49338
rect 8816 49335 8868 49338
rect 8924 49335 8976 49338
rect 9032 49335 9084 49338
rect 9140 49335 9192 49338
rect 9248 49335 9300 49338
rect 9356 49335 9408 49338
rect 9464 49335 9516 49338
rect 9572 49335 9624 49338
rect 9680 49335 9732 49338
rect 9788 49335 9840 49338
rect 10253 49335 10305 49338
rect 10361 49335 10413 49338
rect 10469 49335 10521 49338
rect 10577 49335 10629 49338
rect 10685 49335 10737 49338
rect 10793 49335 10845 49338
rect 10901 49335 10953 49338
rect 11009 49335 11061 49338
rect 11117 49335 11169 49338
rect 11225 49335 11277 49338
rect 11333 49335 11385 49338
rect 11441 49335 11493 49338
rect 11549 49335 11554 49338
rect 11554 49335 11601 49338
rect 3377 49286 3429 49335
rect 3485 49286 3537 49335
rect 3593 49286 3645 49335
rect 3701 49286 3753 49335
rect 3809 49286 3861 49335
rect 3917 49286 3969 49335
rect 4025 49286 4077 49335
rect 4133 49286 4185 49335
rect 4241 49286 4293 49335
rect 4349 49286 4401 49335
rect 4457 49286 4509 49335
rect 4565 49286 4617 49335
rect 4673 49286 4725 49335
rect 5138 49286 5190 49335
rect 5246 49286 5298 49335
rect 5354 49286 5406 49335
rect 5462 49286 5514 49335
rect 5570 49286 5622 49335
rect 5678 49286 5730 49335
rect 5786 49286 5838 49335
rect 5894 49286 5946 49335
rect 6002 49286 6054 49335
rect 6110 49286 6162 49335
rect 6218 49286 6270 49335
rect 6326 49286 6378 49335
rect 6434 49286 6486 49335
rect 6542 49286 6594 49335
rect 6650 49286 6702 49335
rect 6758 49286 6810 49335
rect 6866 49286 6918 49335
rect 6974 49286 7026 49335
rect 7082 49286 7134 49335
rect 7844 49286 7896 49335
rect 7952 49286 8004 49335
rect 8060 49286 8112 49335
rect 8168 49286 8220 49335
rect 8276 49286 8328 49335
rect 8384 49286 8436 49335
rect 8492 49286 8544 49335
rect 8600 49286 8652 49335
rect 8708 49286 8760 49335
rect 8816 49286 8868 49335
rect 8924 49286 8976 49335
rect 9032 49286 9084 49335
rect 9140 49286 9192 49335
rect 9248 49286 9300 49335
rect 9356 49286 9408 49335
rect 9464 49286 9516 49335
rect 9572 49286 9624 49335
rect 9680 49286 9732 49335
rect 9788 49286 9840 49335
rect 10253 49286 10305 49335
rect 10361 49286 10413 49335
rect 10469 49286 10521 49335
rect 10577 49286 10629 49335
rect 10685 49286 10737 49335
rect 10793 49286 10845 49335
rect 10901 49286 10953 49335
rect 11009 49286 11061 49335
rect 11117 49286 11169 49335
rect 11225 49286 11277 49335
rect 11333 49286 11385 49335
rect 11441 49286 11493 49335
rect 11549 49286 11601 49335
rect 11657 49286 11709 49338
rect 11765 49286 11816 49338
rect 11816 49286 11817 49338
rect 3161 49178 3162 49230
rect 3162 49178 3213 49230
rect 3269 49178 3321 49230
rect 3377 49227 3429 49230
rect 3485 49227 3537 49230
rect 3593 49227 3645 49230
rect 3701 49227 3753 49230
rect 3809 49227 3861 49230
rect 3917 49227 3969 49230
rect 4025 49227 4077 49230
rect 4133 49227 4185 49230
rect 4241 49227 4293 49230
rect 4349 49227 4401 49230
rect 4457 49227 4509 49230
rect 4565 49227 4617 49230
rect 4673 49227 4725 49230
rect 5138 49227 5190 49230
rect 5246 49227 5298 49230
rect 5354 49227 5406 49230
rect 5462 49227 5514 49230
rect 5570 49227 5622 49230
rect 5678 49227 5730 49230
rect 5786 49227 5838 49230
rect 5894 49227 5946 49230
rect 6002 49227 6054 49230
rect 6110 49227 6162 49230
rect 6218 49227 6270 49230
rect 6326 49227 6378 49230
rect 6434 49227 6486 49230
rect 6542 49227 6594 49230
rect 6650 49227 6702 49230
rect 6758 49227 6810 49230
rect 6866 49227 6918 49230
rect 6974 49227 7026 49230
rect 7082 49227 7134 49230
rect 7844 49227 7896 49230
rect 7952 49227 8004 49230
rect 8060 49227 8112 49230
rect 8168 49227 8220 49230
rect 8276 49227 8328 49230
rect 8384 49227 8436 49230
rect 8492 49227 8544 49230
rect 8600 49227 8652 49230
rect 8708 49227 8760 49230
rect 8816 49227 8868 49230
rect 8924 49227 8976 49230
rect 9032 49227 9084 49230
rect 9140 49227 9192 49230
rect 9248 49227 9300 49230
rect 9356 49227 9408 49230
rect 9464 49227 9516 49230
rect 9572 49227 9624 49230
rect 9680 49227 9732 49230
rect 9788 49227 9840 49230
rect 10253 49227 10305 49230
rect 10361 49227 10413 49230
rect 10469 49227 10521 49230
rect 10577 49227 10629 49230
rect 10685 49227 10737 49230
rect 10793 49227 10845 49230
rect 10901 49227 10953 49230
rect 11009 49227 11061 49230
rect 11117 49227 11169 49230
rect 11225 49227 11277 49230
rect 11333 49227 11385 49230
rect 11441 49227 11493 49230
rect 11549 49227 11601 49230
rect 3377 49181 3429 49227
rect 3485 49181 3537 49227
rect 3593 49181 3645 49227
rect 3701 49181 3753 49227
rect 3809 49181 3861 49227
rect 3917 49181 3969 49227
rect 4025 49181 4077 49227
rect 4133 49181 4185 49227
rect 4241 49181 4293 49227
rect 4349 49181 4401 49227
rect 4457 49181 4509 49227
rect 4565 49181 4617 49227
rect 4673 49181 4725 49227
rect 5138 49181 5190 49227
rect 5246 49181 5298 49227
rect 5354 49181 5406 49227
rect 5462 49181 5514 49227
rect 5570 49181 5622 49227
rect 5678 49181 5730 49227
rect 5786 49181 5838 49227
rect 5894 49181 5946 49227
rect 6002 49181 6054 49227
rect 6110 49181 6162 49227
rect 6218 49181 6270 49227
rect 6326 49181 6378 49227
rect 6434 49181 6486 49227
rect 6542 49181 6594 49227
rect 6650 49181 6702 49227
rect 6758 49181 6810 49227
rect 6866 49181 6918 49227
rect 6974 49181 7026 49227
rect 7082 49181 7134 49227
rect 7844 49181 7896 49227
rect 7952 49181 8004 49227
rect 8060 49181 8112 49227
rect 8168 49181 8220 49227
rect 8276 49181 8328 49227
rect 8384 49181 8436 49227
rect 8492 49181 8544 49227
rect 8600 49181 8652 49227
rect 8708 49181 8760 49227
rect 8816 49181 8868 49227
rect 8924 49181 8976 49227
rect 9032 49181 9084 49227
rect 9140 49181 9192 49227
rect 9248 49181 9300 49227
rect 9356 49181 9408 49227
rect 9464 49181 9516 49227
rect 9572 49181 9624 49227
rect 9680 49181 9732 49227
rect 9788 49181 9840 49227
rect 10253 49181 10305 49227
rect 10361 49181 10413 49227
rect 10469 49181 10521 49227
rect 10577 49181 10629 49227
rect 10685 49181 10737 49227
rect 10793 49181 10845 49227
rect 10901 49181 10953 49227
rect 11009 49181 11061 49227
rect 11117 49181 11169 49227
rect 11225 49181 11277 49227
rect 11333 49181 11385 49227
rect 11441 49181 11493 49227
rect 11549 49181 11601 49227
rect 3377 49178 3429 49181
rect 3485 49178 3537 49181
rect 3593 49178 3645 49181
rect 3701 49178 3753 49181
rect 3809 49178 3861 49181
rect 3917 49178 3969 49181
rect 4025 49178 4077 49181
rect 4133 49178 4185 49181
rect 4241 49178 4293 49181
rect 4349 49178 4401 49181
rect 4457 49178 4509 49181
rect 4565 49178 4617 49181
rect 4673 49178 4725 49181
rect 5138 49178 5190 49181
rect 5246 49178 5298 49181
rect 5354 49178 5406 49181
rect 5462 49178 5514 49181
rect 5570 49178 5622 49181
rect 5678 49178 5730 49181
rect 5786 49178 5838 49181
rect 5894 49178 5946 49181
rect 6002 49178 6054 49181
rect 6110 49178 6162 49181
rect 6218 49178 6270 49181
rect 6326 49178 6378 49181
rect 6434 49178 6486 49181
rect 6542 49178 6594 49181
rect 6650 49178 6702 49181
rect 6758 49178 6810 49181
rect 6866 49178 6918 49181
rect 6974 49178 7026 49181
rect 7082 49178 7134 49181
rect 7844 49178 7896 49181
rect 7952 49178 8004 49181
rect 8060 49178 8112 49181
rect 8168 49178 8220 49181
rect 8276 49178 8328 49181
rect 8384 49178 8436 49181
rect 8492 49178 8544 49181
rect 8600 49178 8652 49181
rect 8708 49178 8760 49181
rect 8816 49178 8868 49181
rect 8924 49178 8976 49181
rect 9032 49178 9084 49181
rect 9140 49178 9192 49181
rect 9248 49178 9300 49181
rect 9356 49178 9408 49181
rect 9464 49178 9516 49181
rect 9572 49178 9624 49181
rect 9680 49178 9732 49181
rect 9788 49178 9840 49181
rect 10253 49178 10305 49181
rect 10361 49178 10413 49181
rect 10469 49178 10521 49181
rect 10577 49178 10629 49181
rect 10685 49178 10737 49181
rect 10793 49178 10845 49181
rect 10901 49178 10953 49181
rect 11009 49178 11061 49181
rect 11117 49178 11169 49181
rect 11225 49178 11277 49181
rect 11333 49178 11385 49181
rect 11441 49178 11493 49181
rect 11549 49178 11601 49181
rect 11657 49178 11709 49230
rect 11765 49178 11816 49230
rect 11816 49178 11817 49230
rect 3161 49070 3162 49122
rect 3162 49070 3213 49122
rect 3269 49070 3321 49122
rect 3377 49073 3429 49122
rect 3485 49073 3537 49122
rect 3593 49073 3645 49122
rect 3701 49073 3753 49122
rect 3809 49073 3861 49122
rect 3917 49073 3969 49122
rect 4025 49073 4077 49122
rect 4133 49073 4185 49122
rect 4241 49073 4293 49122
rect 4349 49073 4401 49122
rect 4457 49073 4509 49122
rect 4565 49073 4617 49122
rect 4673 49073 4725 49122
rect 5138 49073 5190 49122
rect 5246 49073 5298 49122
rect 5354 49073 5406 49122
rect 5462 49073 5514 49122
rect 5570 49073 5622 49122
rect 5678 49073 5730 49122
rect 5786 49073 5838 49122
rect 5894 49073 5946 49122
rect 6002 49073 6054 49122
rect 6110 49073 6162 49122
rect 6218 49073 6270 49122
rect 6326 49073 6378 49122
rect 6434 49073 6486 49122
rect 6542 49073 6594 49122
rect 6650 49073 6702 49122
rect 6758 49073 6810 49122
rect 6866 49073 6918 49122
rect 6974 49073 7026 49122
rect 7082 49073 7134 49122
rect 7844 49073 7896 49122
rect 7952 49073 8004 49122
rect 8060 49073 8112 49122
rect 8168 49073 8220 49122
rect 8276 49073 8328 49122
rect 8384 49073 8436 49122
rect 8492 49073 8544 49122
rect 8600 49073 8652 49122
rect 8708 49073 8760 49122
rect 8816 49073 8868 49122
rect 8924 49073 8976 49122
rect 9032 49073 9084 49122
rect 9140 49073 9192 49122
rect 9248 49073 9300 49122
rect 9356 49073 9408 49122
rect 9464 49073 9516 49122
rect 9572 49073 9624 49122
rect 9680 49073 9732 49122
rect 9788 49073 9840 49122
rect 10253 49073 10305 49122
rect 10361 49073 10413 49122
rect 10469 49073 10521 49122
rect 10577 49073 10629 49122
rect 10685 49073 10737 49122
rect 10793 49073 10845 49122
rect 10901 49073 10953 49122
rect 11009 49073 11061 49122
rect 11117 49073 11169 49122
rect 11225 49073 11277 49122
rect 11333 49073 11385 49122
rect 11441 49073 11493 49122
rect 11549 49073 11601 49122
rect 3377 49070 3424 49073
rect 3424 49070 3429 49073
rect 3485 49070 3537 49073
rect 3593 49070 3645 49073
rect 3701 49070 3753 49073
rect 3809 49070 3861 49073
rect 3917 49070 3969 49073
rect 4025 49070 4077 49073
rect 4133 49070 4185 49073
rect 4241 49070 4293 49073
rect 4349 49070 4401 49073
rect 4457 49070 4509 49073
rect 4565 49070 4617 49073
rect 4673 49070 4725 49073
rect 5138 49070 5190 49073
rect 5246 49070 5298 49073
rect 5354 49070 5406 49073
rect 5462 49070 5514 49073
rect 5570 49070 5622 49073
rect 5678 49070 5730 49073
rect 5786 49070 5838 49073
rect 5894 49070 5946 49073
rect 6002 49070 6054 49073
rect 6110 49070 6162 49073
rect 6218 49070 6270 49073
rect 6326 49070 6378 49073
rect 6434 49070 6486 49073
rect 6542 49070 6594 49073
rect 6650 49070 6702 49073
rect 6758 49070 6810 49073
rect 6866 49070 6918 49073
rect 6974 49070 7026 49073
rect 7082 49070 7134 49073
rect 7844 49070 7896 49073
rect 7952 49070 8004 49073
rect 8060 49070 8112 49073
rect 8168 49070 8220 49073
rect 8276 49070 8328 49073
rect 8384 49070 8436 49073
rect 8492 49070 8544 49073
rect 8600 49070 8652 49073
rect 8708 49070 8760 49073
rect 8816 49070 8868 49073
rect 8924 49070 8976 49073
rect 9032 49070 9084 49073
rect 9140 49070 9192 49073
rect 9248 49070 9300 49073
rect 9356 49070 9408 49073
rect 9464 49070 9516 49073
rect 9572 49070 9624 49073
rect 9680 49070 9732 49073
rect 9788 49070 9840 49073
rect 10253 49070 10305 49073
rect 10361 49070 10413 49073
rect 10469 49070 10521 49073
rect 10577 49070 10629 49073
rect 10685 49070 10737 49073
rect 10793 49070 10845 49073
rect 10901 49070 10953 49073
rect 11009 49070 11061 49073
rect 11117 49070 11169 49073
rect 11225 49070 11277 49073
rect 11333 49070 11385 49073
rect 11441 49070 11493 49073
rect 11549 49070 11554 49073
rect 11554 49070 11601 49073
rect 11657 49070 11709 49122
rect 11765 49070 11816 49122
rect 11816 49070 11817 49122
rect 4871 48778 4923 48817
rect 4979 48778 5031 48817
rect 7247 48778 7299 48817
rect 7355 48778 7407 48817
rect 7463 48778 7515 48817
rect 7571 48778 7623 48817
rect 7679 48778 7731 48817
rect 9947 48778 9999 48817
rect 10055 48778 10107 48817
rect 4871 48765 4923 48778
rect 4979 48765 5031 48778
rect 7247 48765 7299 48778
rect 7355 48765 7407 48778
rect 7463 48765 7515 48778
rect 7571 48765 7623 48778
rect 7679 48765 7731 48778
rect 9947 48765 9999 48778
rect 10055 48765 10107 48778
rect 4871 48696 4923 48709
rect 4979 48696 5031 48709
rect 7247 48696 7299 48709
rect 7355 48696 7407 48709
rect 7463 48696 7515 48709
rect 7571 48696 7623 48709
rect 7679 48696 7731 48709
rect 9947 48696 9999 48709
rect 10055 48696 10107 48709
rect 4871 48657 4923 48696
rect 4979 48657 5031 48696
rect 7247 48657 7299 48696
rect 7355 48657 7407 48696
rect 7463 48657 7515 48696
rect 7571 48657 7623 48696
rect 7679 48657 7731 48696
rect 9947 48657 9999 48696
rect 10055 48657 10107 48696
rect 3161 48376 3162 48427
rect 3162 48376 3213 48427
rect 3161 48375 3213 48376
rect 3269 48375 3321 48427
rect 3377 48401 3424 48427
rect 3424 48401 3429 48427
rect 3485 48401 3537 48427
rect 3593 48401 3645 48427
rect 3701 48401 3753 48427
rect 3809 48401 3861 48427
rect 3917 48401 3969 48427
rect 4025 48401 4077 48427
rect 4133 48401 4185 48427
rect 4241 48401 4293 48427
rect 4349 48401 4401 48427
rect 4457 48401 4509 48427
rect 4565 48401 4617 48427
rect 4673 48401 4725 48427
rect 5138 48401 5190 48427
rect 5246 48401 5298 48427
rect 5354 48401 5406 48427
rect 5462 48401 5514 48427
rect 5570 48401 5622 48427
rect 5678 48401 5730 48427
rect 5786 48401 5838 48427
rect 5894 48401 5946 48427
rect 6002 48401 6054 48427
rect 6110 48401 6162 48427
rect 6218 48401 6270 48427
rect 6326 48401 6378 48427
rect 6434 48401 6486 48427
rect 6542 48401 6594 48427
rect 6650 48401 6702 48427
rect 6758 48401 6810 48427
rect 6866 48401 6918 48427
rect 6974 48401 7026 48427
rect 7082 48401 7134 48427
rect 7844 48401 7896 48427
rect 7952 48401 8004 48427
rect 8060 48401 8112 48427
rect 8168 48401 8220 48427
rect 8276 48401 8328 48427
rect 8384 48401 8436 48427
rect 8492 48401 8544 48427
rect 8600 48401 8652 48427
rect 8708 48401 8760 48427
rect 8816 48401 8868 48427
rect 8924 48401 8976 48427
rect 9032 48401 9084 48427
rect 9140 48401 9192 48427
rect 9248 48401 9300 48427
rect 9356 48401 9408 48427
rect 9464 48401 9516 48427
rect 9572 48401 9624 48427
rect 9680 48401 9732 48427
rect 9788 48401 9840 48427
rect 10253 48401 10305 48427
rect 10361 48401 10413 48427
rect 10469 48401 10521 48427
rect 10577 48401 10629 48427
rect 10685 48401 10737 48427
rect 10793 48401 10845 48427
rect 10901 48401 10953 48427
rect 11009 48401 11061 48427
rect 11117 48401 11169 48427
rect 11225 48401 11277 48427
rect 11333 48401 11385 48427
rect 11441 48401 11493 48427
rect 11549 48401 11554 48427
rect 11554 48401 11601 48427
rect 3377 48375 3429 48401
rect 3485 48375 3537 48401
rect 3593 48375 3645 48401
rect 3701 48375 3753 48401
rect 3809 48375 3861 48401
rect 3917 48375 3969 48401
rect 4025 48375 4077 48401
rect 4133 48375 4185 48401
rect 4241 48375 4293 48401
rect 4349 48375 4401 48401
rect 4457 48375 4509 48401
rect 4565 48375 4617 48401
rect 4673 48375 4725 48401
rect 5138 48375 5190 48401
rect 5246 48375 5298 48401
rect 5354 48375 5406 48401
rect 5462 48375 5514 48401
rect 5570 48375 5622 48401
rect 5678 48375 5730 48401
rect 5786 48375 5838 48401
rect 5894 48375 5946 48401
rect 6002 48375 6054 48401
rect 6110 48375 6162 48401
rect 6218 48375 6270 48401
rect 6326 48375 6378 48401
rect 6434 48375 6486 48401
rect 6542 48375 6594 48401
rect 6650 48375 6702 48401
rect 6758 48375 6810 48401
rect 6866 48375 6918 48401
rect 6974 48375 7026 48401
rect 7082 48375 7134 48401
rect 7844 48375 7896 48401
rect 7952 48375 8004 48401
rect 8060 48375 8112 48401
rect 8168 48375 8220 48401
rect 8276 48375 8328 48401
rect 8384 48375 8436 48401
rect 8492 48375 8544 48401
rect 8600 48375 8652 48401
rect 8708 48375 8760 48401
rect 8816 48375 8868 48401
rect 8924 48375 8976 48401
rect 9032 48375 9084 48401
rect 9140 48375 9192 48401
rect 9248 48375 9300 48401
rect 9356 48375 9408 48401
rect 9464 48375 9516 48401
rect 9572 48375 9624 48401
rect 9680 48375 9732 48401
rect 9788 48375 9840 48401
rect 10253 48375 10305 48401
rect 10361 48375 10413 48401
rect 10469 48375 10521 48401
rect 10577 48375 10629 48401
rect 10685 48375 10737 48401
rect 10793 48375 10845 48401
rect 10901 48375 10953 48401
rect 11009 48375 11061 48401
rect 11117 48375 11169 48401
rect 11225 48375 11277 48401
rect 11333 48375 11385 48401
rect 11441 48375 11493 48401
rect 11549 48375 11601 48401
rect 11657 48375 11709 48427
rect 11765 48376 11816 48427
rect 11816 48376 11817 48427
rect 11765 48375 11817 48376
rect 3161 48293 3213 48319
rect 3269 48293 3321 48319
rect 3377 48293 3429 48319
rect 3485 48293 3537 48319
rect 3593 48293 3645 48319
rect 3701 48293 3753 48319
rect 3809 48293 3861 48319
rect 3917 48293 3969 48319
rect 4025 48293 4077 48319
rect 4133 48293 4185 48319
rect 4241 48293 4293 48319
rect 4349 48293 4401 48319
rect 4457 48293 4509 48319
rect 4565 48293 4617 48319
rect 4673 48293 4725 48319
rect 5138 48293 5190 48319
rect 5246 48293 5298 48319
rect 5354 48293 5406 48319
rect 5462 48293 5514 48319
rect 5570 48293 5622 48319
rect 5678 48293 5730 48319
rect 5786 48293 5838 48319
rect 5894 48293 5946 48319
rect 6002 48293 6054 48319
rect 6110 48293 6162 48319
rect 6218 48293 6270 48319
rect 6326 48293 6378 48319
rect 6434 48293 6486 48319
rect 6542 48293 6594 48319
rect 6650 48293 6702 48319
rect 6758 48293 6810 48319
rect 6866 48293 6918 48319
rect 6974 48293 7026 48319
rect 7082 48293 7134 48319
rect 7844 48293 7896 48319
rect 7952 48293 8004 48319
rect 8060 48293 8112 48319
rect 8168 48293 8220 48319
rect 8276 48293 8328 48319
rect 8384 48293 8436 48319
rect 8492 48293 8544 48319
rect 8600 48293 8652 48319
rect 8708 48293 8760 48319
rect 8816 48293 8868 48319
rect 8924 48293 8976 48319
rect 9032 48293 9084 48319
rect 9140 48293 9192 48319
rect 9248 48293 9300 48319
rect 9356 48293 9408 48319
rect 9464 48293 9516 48319
rect 9572 48293 9624 48319
rect 9680 48293 9732 48319
rect 9788 48293 9840 48319
rect 10253 48293 10305 48319
rect 10361 48293 10413 48319
rect 10469 48293 10521 48319
rect 10577 48293 10629 48319
rect 10685 48293 10737 48319
rect 10793 48293 10845 48319
rect 10901 48293 10953 48319
rect 11009 48293 11061 48319
rect 11117 48293 11169 48319
rect 11225 48293 11277 48319
rect 11333 48293 11385 48319
rect 11441 48293 11493 48319
rect 11549 48293 11601 48319
rect 11657 48293 11709 48319
rect 11765 48293 11817 48319
rect 3161 48267 3213 48293
rect 3269 48267 3321 48293
rect 3377 48267 3429 48293
rect 3485 48267 3537 48293
rect 3593 48267 3645 48293
rect 3701 48267 3753 48293
rect 3809 48267 3861 48293
rect 3917 48267 3969 48293
rect 4025 48267 4077 48293
rect 4133 48267 4185 48293
rect 4241 48267 4293 48293
rect 4349 48267 4401 48293
rect 4457 48267 4509 48293
rect 4565 48267 4617 48293
rect 4673 48267 4725 48293
rect 5138 48267 5190 48293
rect 5246 48267 5298 48293
rect 5354 48267 5406 48293
rect 5462 48267 5514 48293
rect 5570 48267 5622 48293
rect 5678 48267 5730 48293
rect 5786 48267 5838 48293
rect 5894 48267 5946 48293
rect 6002 48267 6054 48293
rect 6110 48267 6162 48293
rect 6218 48267 6270 48293
rect 6326 48267 6378 48293
rect 6434 48267 6486 48293
rect 6542 48267 6594 48293
rect 6650 48267 6702 48293
rect 6758 48267 6810 48293
rect 6866 48267 6918 48293
rect 6974 48267 7026 48293
rect 7082 48267 7134 48293
rect 7844 48267 7896 48293
rect 7952 48267 8004 48293
rect 8060 48267 8112 48293
rect 8168 48267 8220 48293
rect 8276 48267 8328 48293
rect 8384 48267 8436 48293
rect 8492 48267 8544 48293
rect 8600 48267 8652 48293
rect 8708 48267 8760 48293
rect 8816 48267 8868 48293
rect 8924 48267 8976 48293
rect 9032 48267 9084 48293
rect 9140 48267 9192 48293
rect 9248 48267 9300 48293
rect 9356 48267 9408 48293
rect 9464 48267 9516 48293
rect 9572 48267 9624 48293
rect 9680 48267 9732 48293
rect 9788 48267 9840 48293
rect 10253 48267 10305 48293
rect 10361 48267 10413 48293
rect 10469 48267 10521 48293
rect 10577 48267 10629 48293
rect 10685 48267 10737 48293
rect 10793 48267 10845 48293
rect 10901 48267 10953 48293
rect 11009 48267 11061 48293
rect 11117 48267 11169 48293
rect 11225 48267 11277 48293
rect 11333 48267 11385 48293
rect 11441 48267 11493 48293
rect 11549 48267 11601 48293
rect 11657 48267 11709 48293
rect 11765 48267 11817 48293
rect 12336 52218 12388 52270
rect 12336 52110 12388 52162
rect 12336 52002 12388 52054
rect 12336 51894 12388 51946
rect 12336 51786 12388 51838
rect 12336 51678 12388 51730
rect 12336 51570 12388 51622
rect 12336 51462 12388 51514
rect 12336 51354 12388 51406
rect 12336 51246 12388 51298
rect 12336 51138 12388 51190
rect 12336 51030 12388 51082
rect 12336 50922 12388 50974
rect 12336 50814 12388 50866
rect 12336 50706 12388 50758
rect 12336 50598 12388 50650
rect 12336 50490 12388 50542
rect 12336 50382 12388 50434
rect 12336 50274 12388 50326
rect 12336 50166 12388 50218
rect 12336 50058 12388 50110
rect 12336 49950 12388 50002
rect 12336 49842 12388 49894
rect 12336 49734 12388 49786
rect 12336 49626 12388 49678
rect 12336 49518 12388 49570
rect 12336 49410 12388 49462
rect 12336 49302 12388 49354
rect 12336 49194 12388 49246
rect 12336 49086 12388 49138
rect 12336 48978 12388 49030
rect 12336 48870 12388 48922
rect 12336 48762 12388 48814
rect 12336 48654 12388 48706
rect 12336 48546 12388 48598
rect 12336 48438 12388 48490
rect 12336 48330 12388 48382
rect 12336 48222 12388 48274
rect 12336 48114 12388 48166
rect 2590 47898 2642 47950
rect 2590 47790 2642 47842
rect 2590 47682 2642 47734
rect 4871 47920 4923 47972
rect 4979 47920 5031 47972
rect 7247 47920 7299 47972
rect 7355 47920 7407 47972
rect 7463 47920 7515 47972
rect 7571 47920 7623 47972
rect 7679 47920 7731 47972
rect 9947 47920 9999 47972
rect 10055 47920 10107 47972
rect 4871 47812 4923 47864
rect 4979 47812 5031 47864
rect 7247 47812 7299 47864
rect 7355 47812 7407 47864
rect 7463 47812 7515 47864
rect 7571 47812 7623 47864
rect 7679 47812 7731 47864
rect 9947 47812 9999 47864
rect 10055 47812 10107 47864
rect 4871 47704 4923 47756
rect 4979 47704 5031 47756
rect 7247 47704 7299 47756
rect 7355 47704 7407 47756
rect 7463 47704 7515 47756
rect 7571 47704 7623 47756
rect 7679 47704 7731 47756
rect 9947 47704 9999 47756
rect 10055 47704 10107 47756
rect 12336 48006 12388 48058
rect 12336 47898 12388 47950
rect 12336 47790 12388 47842
rect 12336 47682 12388 47734
rect 14904 52522 14956 52574
rect 14904 52414 14956 52466
rect 14904 52306 14956 52358
rect 14904 52198 14956 52250
rect 14904 52090 14956 52142
rect 14904 51982 14956 52034
rect 14904 51874 14956 51926
rect 14904 51766 14956 51818
rect 14904 51658 14956 51710
rect 14904 51550 14956 51602
rect 14904 51442 14956 51494
rect 14904 51334 14956 51386
rect 14904 51226 14956 51278
rect 14904 49322 14956 49374
rect 14904 49214 14956 49266
rect 14904 49106 14956 49158
rect 14904 48998 14956 49050
rect 14904 48890 14956 48942
rect 14904 48782 14956 48834
rect 14904 48674 14956 48726
rect 14904 48566 14956 48618
rect 14904 48458 14956 48510
rect 14904 48350 14956 48402
rect 14904 48242 14956 48294
rect 14904 48134 14956 48186
rect 14904 48026 14956 48078
rect 22 46122 74 46174
rect 22 46014 74 46066
rect 22 45906 74 45958
rect 22 45798 74 45850
rect 22 45690 74 45742
rect 22 45582 74 45634
rect 22 45474 74 45526
rect 22 45366 74 45418
rect 22 45258 74 45310
rect 22 45150 74 45202
rect 22 45042 74 45094
rect 22 44934 74 44986
rect 22 44826 74 44878
rect 14904 46122 14956 46174
rect 14904 46014 14956 46066
rect 14904 45906 14956 45958
rect 14904 45798 14956 45850
rect 14904 45690 14956 45742
rect 14904 45582 14956 45634
rect 14904 45474 14956 45526
rect 14904 45366 14956 45418
rect 14904 45258 14956 45310
rect 14904 45150 14956 45202
rect 14904 45042 14956 45094
rect 14904 44934 14956 44986
rect 14904 44826 14956 44878
rect 22 38122 74 38174
rect 22 38014 74 38066
rect 22 37906 74 37958
rect 22 37798 74 37850
rect 22 37690 74 37742
rect 22 37582 74 37634
rect 22 37474 74 37526
rect 22 37366 74 37418
rect 22 37258 74 37310
rect 22 37150 74 37202
rect 22 37042 74 37094
rect 22 36934 74 36986
rect 22 36826 74 36878
rect 22 36532 74 36584
rect 22 36424 74 36476
rect 22 36316 74 36368
rect 22 36208 74 36260
rect 22 36100 74 36152
rect 22 35992 74 36044
rect 22 35884 74 35936
rect 22 35776 74 35828
rect 22 35668 74 35720
rect 22 35560 74 35612
rect 22 35452 74 35504
rect 22 35344 74 35396
rect 22 35236 74 35288
rect 22 35128 74 35180
rect 22 35020 74 35072
rect 22 34912 74 34964
rect 22 34804 74 34856
rect 22 34696 74 34748
rect 22 34588 74 34640
rect 22 34480 74 34532
rect 22 34372 74 34424
rect 22 34264 74 34316
rect 22 34156 74 34208
rect 22 34048 74 34100
rect 22 33940 74 33992
rect 22 33832 74 33884
rect 22 33724 74 33776
rect 22 33616 74 33668
rect 22 28522 74 28574
rect 22 28414 74 28466
rect 22 28306 74 28358
rect 22 28198 74 28250
rect 22 28090 74 28142
rect 22 27982 74 28034
rect 22 27874 74 27926
rect 22 27766 74 27818
rect 22 27658 74 27710
rect 22 27550 74 27602
rect 22 27442 74 27494
rect 22 27334 74 27386
rect 22 27226 74 27278
rect 22 14122 74 14174
rect 22 14014 74 14066
rect 22 13906 74 13958
rect 22 13798 74 13850
rect 22 13690 74 13742
rect 22 13582 74 13634
rect 22 13474 74 13526
rect 22 13366 74 13418
rect 22 13258 74 13310
rect 22 13150 74 13202
rect 22 13042 74 13094
rect 22 12934 74 12986
rect 22 12826 74 12878
rect 22 10932 74 10984
rect 22 10824 74 10876
rect 22 10716 74 10768
rect 22 10608 74 10660
rect 22 10500 74 10552
rect 22 10392 74 10444
rect 22 10284 74 10336
rect 22 10176 74 10228
rect 22 10068 74 10120
rect 22 9960 74 10012
rect 22 9852 74 9904
rect 22 9744 74 9796
rect 22 9636 74 9688
rect 22 9528 74 9580
rect 22 9420 74 9472
rect 22 9312 74 9364
rect 22 9204 74 9256
rect 22 9096 74 9148
rect 22 8988 74 9040
rect 22 8880 74 8932
rect 22 8772 74 8824
rect 22 8664 74 8716
rect 22 8556 74 8608
rect 22 8448 74 8500
rect 22 8340 74 8392
rect 22 8232 74 8284
rect 22 8124 74 8176
rect 22 8016 74 8068
rect 22 7732 74 7784
rect 22 7624 74 7676
rect 22 7516 74 7568
rect 22 7408 74 7460
rect 22 7300 74 7352
rect 22 7192 74 7244
rect 22 7084 74 7136
rect 22 6976 74 7028
rect 22 6868 74 6920
rect 22 6760 74 6812
rect 22 6652 74 6704
rect 22 6544 74 6596
rect 22 6436 74 6488
rect 22 6328 74 6380
rect 22 6220 74 6272
rect 22 6112 74 6164
rect 22 6004 74 6056
rect 22 5896 74 5948
rect 22 5788 74 5840
rect 22 5680 74 5732
rect 22 5572 74 5624
rect 22 5464 74 5516
rect 22 5356 74 5408
rect 22 5248 74 5300
rect 22 5140 74 5192
rect 22 5032 74 5084
rect 22 4924 74 4976
rect 22 4816 74 4868
rect 22 4532 74 4584
rect 22 4424 74 4476
rect 22 4316 74 4368
rect 22 4208 74 4260
rect 22 4100 74 4152
rect 22 3992 74 4044
rect 22 3884 74 3936
rect 22 3776 74 3828
rect 22 3668 74 3720
rect 22 3560 74 3612
rect 22 3452 74 3504
rect 22 3344 74 3396
rect 22 3236 74 3288
rect 22 3128 74 3180
rect 22 3020 74 3072
rect 22 2912 74 2964
rect 22 2804 74 2856
rect 22 2696 74 2748
rect 22 2588 74 2640
rect 22 2480 74 2532
rect 22 2372 74 2424
rect 22 2264 74 2316
rect 22 2156 74 2208
rect 22 2048 74 2100
rect 22 1940 74 1992
rect 22 1832 74 1884
rect 22 1724 74 1776
rect 22 1616 74 1668
rect 14904 38122 14956 38174
rect 14904 38014 14956 38066
rect 14904 37906 14956 37958
rect 14904 37798 14956 37850
rect 14904 37690 14956 37742
rect 14904 37582 14956 37634
rect 14904 37474 14956 37526
rect 14904 37366 14956 37418
rect 14904 37258 14956 37310
rect 14904 37150 14956 37202
rect 14904 37042 14956 37094
rect 14904 36934 14956 36986
rect 14904 36826 14956 36878
rect 14904 36532 14956 36584
rect 14904 36424 14956 36476
rect 14904 36316 14956 36368
rect 14904 36208 14956 36260
rect 14904 36100 14956 36152
rect 14904 35992 14956 36044
rect 14904 35884 14956 35936
rect 14904 35776 14956 35828
rect 14904 35668 14956 35720
rect 14904 35560 14956 35612
rect 14904 35452 14956 35504
rect 14904 35344 14956 35396
rect 14904 35236 14956 35288
rect 14904 35128 14956 35180
rect 14904 35020 14956 35072
rect 14904 34912 14956 34964
rect 14904 34804 14956 34856
rect 14904 34696 14956 34748
rect 14904 34588 14956 34640
rect 14904 34480 14956 34532
rect 14904 34372 14956 34424
rect 14904 34264 14956 34316
rect 14904 34156 14956 34208
rect 14904 34048 14956 34100
rect 14904 33940 14956 33992
rect 14904 33832 14956 33884
rect 14904 33724 14956 33776
rect 14904 33616 14956 33668
rect 14904 28522 14956 28574
rect 14904 28414 14956 28466
rect 14904 28306 14956 28358
rect 14904 28198 14956 28250
rect 14904 28090 14956 28142
rect 14904 27982 14956 28034
rect 14904 27874 14956 27926
rect 14904 27766 14956 27818
rect 14904 27658 14956 27710
rect 14904 27550 14956 27602
rect 14904 27442 14956 27494
rect 14904 27334 14956 27386
rect 14904 27226 14956 27278
rect 14904 14122 14956 14174
rect 14904 14014 14956 14066
rect 14904 13906 14956 13958
rect 14904 13798 14956 13850
rect 14904 13690 14956 13742
rect 14904 13582 14956 13634
rect 14904 13474 14956 13526
rect 14904 13366 14956 13418
rect 14904 13258 14956 13310
rect 14904 13150 14956 13202
rect 14904 13042 14956 13094
rect 14904 12934 14956 12986
rect 14904 12826 14956 12878
rect 14904 10932 14956 10984
rect 14904 10824 14956 10876
rect 14904 10716 14956 10768
rect 14904 10608 14956 10660
rect 14904 10500 14956 10552
rect 14904 10392 14956 10444
rect 14904 10284 14956 10336
rect 14904 10176 14956 10228
rect 14904 10068 14956 10120
rect 14904 9960 14956 10012
rect 14904 9852 14956 9904
rect 14904 9744 14956 9796
rect 14904 9636 14956 9688
rect 14904 9528 14956 9580
rect 14904 9420 14956 9472
rect 14904 9312 14956 9364
rect 14904 9204 14956 9256
rect 14904 9096 14956 9148
rect 14904 8988 14956 9040
rect 14904 8880 14956 8932
rect 14904 8772 14956 8824
rect 14904 8664 14956 8716
rect 14904 8556 14956 8608
rect 14904 8448 14956 8500
rect 14904 8340 14956 8392
rect 14904 8232 14956 8284
rect 14904 8124 14956 8176
rect 14904 8016 14956 8068
rect 14904 7732 14956 7784
rect 14904 7624 14956 7676
rect 14904 7516 14956 7568
rect 14904 7408 14956 7460
rect 14904 7300 14956 7352
rect 14904 7192 14956 7244
rect 14904 7084 14956 7136
rect 14904 6976 14956 7028
rect 14904 6868 14956 6920
rect 14904 6760 14956 6812
rect 14904 6652 14956 6704
rect 14904 6544 14956 6596
rect 14904 6436 14956 6488
rect 14904 6328 14956 6380
rect 14904 6220 14956 6272
rect 14904 6112 14956 6164
rect 14904 6004 14956 6056
rect 14904 5896 14956 5948
rect 14904 5788 14956 5840
rect 14904 5680 14956 5732
rect 14904 5572 14956 5624
rect 14904 5464 14956 5516
rect 14904 5356 14956 5408
rect 14904 5248 14956 5300
rect 14904 5140 14956 5192
rect 14904 5032 14956 5084
rect 14904 4924 14956 4976
rect 14904 4816 14956 4868
rect 14904 4532 14956 4584
rect 14904 4424 14956 4476
rect 14904 4316 14956 4368
rect 14904 4208 14956 4260
rect 14904 4100 14956 4152
rect 14904 3992 14956 4044
rect 14904 3884 14956 3936
rect 14904 3776 14956 3828
rect 14904 3668 14956 3720
rect 14904 3560 14956 3612
rect 14904 3452 14956 3504
rect 14904 3344 14956 3396
rect 14904 3236 14956 3288
rect 14904 3128 14956 3180
rect 14904 3020 14956 3072
rect 14904 2912 14956 2964
rect 14904 2804 14956 2856
rect 14904 2696 14956 2748
rect 14904 2588 14956 2640
rect 14904 2480 14956 2532
rect 14904 2372 14956 2424
rect 14904 2264 14956 2316
rect 14904 2156 14956 2208
rect 14904 2048 14956 2100
rect 14904 1940 14956 1992
rect 14904 1832 14956 1884
rect 14904 1724 14956 1776
rect 14904 1616 14956 1668
rect 321 766 373 818
rect 429 766 481 818
rect 537 766 589 818
rect 645 766 697 818
rect 753 766 805 818
rect 861 766 913 818
rect 969 766 1021 818
rect 1077 766 1129 818
rect 1185 766 1237 818
rect 1293 766 1345 818
rect 1401 766 1453 818
rect 1509 766 1561 818
rect 1617 766 1669 818
rect 1725 766 1777 818
rect 1833 766 1885 818
rect 1941 766 1993 818
rect 2049 766 2101 818
rect 2876 766 2928 818
rect 2984 766 3036 818
rect 3092 766 3144 818
rect 3200 766 3252 818
rect 3308 766 3360 818
rect 3416 766 3468 818
rect 3524 766 3576 818
rect 3632 766 3684 818
rect 3740 766 3792 818
rect 3848 766 3900 818
rect 3956 766 4008 818
rect 4064 766 4116 818
rect 4172 766 4224 818
rect 4280 766 4332 818
rect 4388 766 4440 818
rect 4496 766 4548 818
rect 4604 766 4656 818
rect 5246 766 5298 818
rect 5354 766 5406 818
rect 5462 766 5514 818
rect 5570 766 5622 818
rect 5678 766 5730 818
rect 5786 766 5838 818
rect 5894 766 5946 818
rect 6002 766 6054 818
rect 6110 766 6162 818
rect 6218 766 6270 818
rect 6326 766 6378 818
rect 6434 766 6486 818
rect 6542 766 6594 818
rect 6650 766 6702 818
rect 6758 766 6810 818
rect 6866 766 6918 818
rect 6974 766 7026 818
rect 7952 766 8004 818
rect 8060 766 8112 818
rect 8168 766 8220 818
rect 8276 766 8328 818
rect 8384 766 8436 818
rect 8492 766 8544 818
rect 8600 766 8652 818
rect 8708 766 8760 818
rect 8816 766 8868 818
rect 8924 766 8976 818
rect 9032 766 9084 818
rect 9140 766 9192 818
rect 9248 766 9300 818
rect 9356 766 9408 818
rect 9464 766 9516 818
rect 9572 766 9624 818
rect 9680 766 9732 818
rect 10322 766 10374 818
rect 10430 766 10482 818
rect 10538 766 10590 818
rect 10646 766 10698 818
rect 10754 766 10806 818
rect 10862 766 10914 818
rect 10970 766 11022 818
rect 11078 766 11130 818
rect 11186 766 11238 818
rect 11294 766 11346 818
rect 11402 766 11454 818
rect 11510 766 11562 818
rect 11618 766 11670 818
rect 11726 766 11778 818
rect 11834 766 11886 818
rect 11942 766 11994 818
rect 12050 766 12102 818
rect 12877 766 12929 818
rect 12985 766 13037 818
rect 13093 766 13145 818
rect 13201 766 13253 818
rect 13309 766 13361 818
rect 13417 766 13469 818
rect 13525 766 13577 818
rect 13633 766 13685 818
rect 13741 766 13793 818
rect 13849 766 13901 818
rect 13957 766 14009 818
rect 14065 766 14117 818
rect 14173 766 14225 818
rect 14281 766 14333 818
rect 14389 766 14441 818
rect 14497 766 14549 818
rect 14605 766 14657 818
<< metal2 >>
rect 261 57499 2161 57600
rect 261 57447 321 57499
rect 373 57447 429 57499
rect 481 57447 537 57499
rect 589 57447 645 57499
rect 697 57447 753 57499
rect 805 57447 861 57499
rect 913 57447 969 57499
rect 1021 57447 1077 57499
rect 1129 57447 1185 57499
rect 1237 57447 1293 57499
rect 1345 57447 1401 57499
rect 1453 57447 1509 57499
rect 1561 57447 1617 57499
rect 1669 57447 1725 57499
rect 1777 57447 1833 57499
rect 1885 57447 1941 57499
rect 1993 57447 2049 57499
rect 2101 57447 2161 57499
rect -11 57261 86 57271
rect -11 56017 20 57261
rect 76 56017 86 57261
rect -11 56007 86 56017
rect 261 57225 2161 57447
rect 2741 57499 4791 57600
rect 2741 57447 2876 57499
rect 2928 57447 2984 57499
rect 3036 57447 3092 57499
rect 3144 57447 3200 57499
rect 3252 57447 3308 57499
rect 3360 57447 3416 57499
rect 3468 57447 3524 57499
rect 3576 57447 3632 57499
rect 3684 57447 3740 57499
rect 3792 57447 3848 57499
rect 3900 57447 3956 57499
rect 4008 57447 4064 57499
rect 4116 57447 4172 57499
rect 4224 57447 4280 57499
rect 4332 57447 4388 57499
rect 4440 57447 4496 57499
rect 4548 57447 4604 57499
rect 4656 57447 4791 57499
rect 261 57169 315 57225
rect 371 57169 439 57225
rect 495 57169 563 57225
rect 619 57169 687 57225
rect 743 57169 811 57225
rect 867 57169 935 57225
rect 991 57169 1059 57225
rect 1115 57169 1183 57225
rect 1239 57169 1307 57225
rect 1363 57169 1431 57225
rect 1487 57169 1555 57225
rect 1611 57169 1679 57225
rect 1735 57169 1803 57225
rect 1859 57169 1927 57225
rect 1983 57169 2051 57225
rect 2107 57169 2161 57225
rect 261 57104 2161 57169
rect 261 57101 375 57104
rect 261 57045 315 57101
rect 371 57052 375 57101
rect 427 57101 483 57104
rect 535 57101 591 57104
rect 643 57101 699 57104
rect 427 57052 439 57101
rect 535 57052 563 57101
rect 643 57052 687 57101
rect 751 57052 807 57104
rect 859 57101 915 57104
rect 967 57101 1023 57104
rect 1075 57101 1131 57104
rect 867 57052 915 57101
rect 991 57052 1023 57101
rect 1115 57052 1131 57101
rect 1183 57101 1239 57104
rect 371 57045 439 57052
rect 495 57045 563 57052
rect 619 57045 687 57052
rect 743 57045 811 57052
rect 867 57045 935 57052
rect 991 57045 1059 57052
rect 1115 57045 1183 57052
rect 1291 57101 1347 57104
rect 1399 57101 1455 57104
rect 1507 57101 1563 57104
rect 1291 57052 1307 57101
rect 1399 57052 1431 57101
rect 1507 57052 1555 57101
rect 1615 57052 1671 57104
rect 1723 57101 1779 57104
rect 1831 57101 1887 57104
rect 1939 57101 1995 57104
rect 1735 57052 1779 57101
rect 1859 57052 1887 57101
rect 1983 57052 1995 57101
rect 2047 57101 2161 57104
rect 2047 57052 2051 57101
rect 1239 57045 1307 57052
rect 1363 57045 1431 57052
rect 1487 57045 1555 57052
rect 1611 57045 1679 57052
rect 1735 57045 1803 57052
rect 1859 57045 1927 57052
rect 1983 57045 2051 57052
rect 2107 57045 2161 57101
rect 261 56977 2161 57045
rect 261 56921 315 56977
rect 371 56921 439 56977
rect 495 56921 563 56977
rect 619 56921 687 56977
rect 743 56921 811 56977
rect 867 56921 935 56977
rect 991 56921 1059 56977
rect 1115 56921 1183 56977
rect 1239 56921 1307 56977
rect 1363 56921 1431 56977
rect 1487 56921 1555 56977
rect 1611 56921 1679 56977
rect 1735 56921 1803 56977
rect 1859 56921 1927 56977
rect 1983 56921 2051 56977
rect 2107 56921 2161 56977
rect 261 56853 2161 56921
rect 261 56797 315 56853
rect 371 56797 439 56853
rect 495 56797 563 56853
rect 619 56797 687 56853
rect 743 56797 811 56853
rect 867 56797 935 56853
rect 991 56797 1059 56853
rect 1115 56797 1183 56853
rect 1239 56797 1307 56853
rect 1363 56797 1431 56853
rect 1487 56797 1555 56853
rect 1611 56797 1679 56853
rect 1735 56797 1803 56853
rect 1859 56797 1927 56853
rect 1983 56797 2051 56853
rect 2107 56797 2161 56853
rect 261 56729 2161 56797
rect 261 56673 315 56729
rect 371 56673 439 56729
rect 495 56673 563 56729
rect 619 56673 687 56729
rect 743 56673 811 56729
rect 867 56673 935 56729
rect 991 56673 1059 56729
rect 1115 56673 1183 56729
rect 1239 56673 1307 56729
rect 1363 56673 1431 56729
rect 1487 56673 1555 56729
rect 1611 56673 1679 56729
rect 1735 56673 1803 56729
rect 1859 56673 1927 56729
rect 1983 56673 2051 56729
rect 2107 56673 2161 56729
rect 261 56643 2161 56673
rect 261 56605 369 56643
rect 421 56605 493 56643
rect 545 56605 617 56643
rect 669 56605 741 56643
rect 793 56605 2161 56643
rect 261 56549 315 56605
rect 421 56591 439 56605
rect 545 56591 563 56605
rect 669 56591 687 56605
rect 793 56591 811 56605
rect 371 56549 439 56591
rect 495 56549 563 56591
rect 619 56549 687 56591
rect 743 56549 811 56591
rect 867 56549 935 56605
rect 991 56549 1059 56605
rect 1115 56549 1183 56605
rect 1239 56549 1307 56605
rect 1363 56549 1431 56605
rect 1487 56549 1555 56605
rect 1611 56549 1679 56605
rect 1735 56549 1803 56605
rect 1859 56549 1927 56605
rect 1983 56549 2051 56605
rect 2107 56549 2161 56605
rect 261 56519 2161 56549
rect 261 56481 369 56519
rect 421 56481 493 56519
rect 545 56481 617 56519
rect 669 56481 741 56519
rect 793 56481 2161 56519
rect 261 56425 315 56481
rect 421 56467 439 56481
rect 545 56467 563 56481
rect 669 56467 687 56481
rect 793 56467 811 56481
rect 371 56425 439 56467
rect 495 56425 563 56467
rect 619 56425 687 56467
rect 743 56425 811 56467
rect 867 56425 935 56481
rect 991 56425 1059 56481
rect 1115 56425 1183 56481
rect 1239 56425 1307 56481
rect 1363 56425 1431 56481
rect 1487 56425 1555 56481
rect 1611 56425 1679 56481
rect 1735 56425 1803 56481
rect 1859 56425 1927 56481
rect 1983 56425 2051 56481
rect 2107 56425 2161 56481
rect 261 56395 2161 56425
rect 261 56357 369 56395
rect 421 56357 493 56395
rect 545 56357 617 56395
rect 669 56357 741 56395
rect 793 56357 2161 56395
rect 261 56301 315 56357
rect 421 56343 439 56357
rect 545 56343 563 56357
rect 669 56343 687 56357
rect 793 56343 811 56357
rect 371 56301 439 56343
rect 495 56301 563 56343
rect 619 56301 687 56343
rect 743 56301 811 56343
rect 867 56301 935 56357
rect 991 56301 1059 56357
rect 1115 56301 1183 56357
rect 1239 56301 1307 56357
rect 1363 56301 1431 56357
rect 1487 56301 1555 56357
rect 1611 56301 1679 56357
rect 1735 56301 1803 56357
rect 1859 56301 1927 56357
rect 1983 56301 2051 56357
rect 2107 56301 2161 56357
rect 261 56271 2161 56301
rect 261 56233 369 56271
rect 421 56233 493 56271
rect 545 56233 617 56271
rect 669 56233 741 56271
rect 793 56233 2161 56271
rect 261 56177 315 56233
rect 421 56219 439 56233
rect 545 56219 563 56233
rect 669 56219 687 56233
rect 793 56219 811 56233
rect 371 56177 439 56219
rect 495 56177 563 56219
rect 619 56177 687 56219
rect 743 56177 811 56219
rect 867 56177 935 56233
rect 991 56177 1059 56233
rect 1115 56177 1183 56233
rect 1239 56177 1307 56233
rect 1363 56177 1431 56233
rect 1487 56177 1555 56233
rect 1611 56177 1679 56233
rect 1735 56177 1803 56233
rect 1859 56177 1927 56233
rect 1983 56177 2051 56233
rect 2107 56177 2161 56233
rect 261 56147 2161 56177
rect 261 56109 369 56147
rect 421 56109 493 56147
rect 545 56109 617 56147
rect 669 56109 741 56147
rect 793 56109 2161 56147
rect 261 56053 315 56109
rect 421 56095 439 56109
rect 545 56095 563 56109
rect 669 56095 687 56109
rect 793 56095 811 56109
rect 371 56053 439 56095
rect 495 56053 563 56095
rect 619 56053 687 56095
rect 743 56053 811 56095
rect 867 56053 935 56109
rect 991 56053 1059 56109
rect 1115 56053 1183 56109
rect 1239 56053 1307 56109
rect 1363 56053 1431 56109
rect 1487 56053 1555 56109
rect 1611 56053 1679 56109
rect 1735 56053 1803 56109
rect 1859 56053 1927 56109
rect 1983 56053 2051 56109
rect 2107 56053 2161 56109
rect 261 56023 2161 56053
rect 261 55971 369 56023
rect 421 55971 493 56023
rect 545 55971 617 56023
rect 669 55971 741 56023
rect 793 55971 2161 56023
rect 261 55899 2161 55971
rect 261 55847 369 55899
rect 421 55847 493 55899
rect 545 55847 617 55899
rect 669 55847 741 55899
rect 793 55847 2161 55899
rect 261 55775 2161 55847
rect 261 55723 369 55775
rect 421 55723 493 55775
rect 545 55723 617 55775
rect 669 55723 741 55775
rect 793 55723 2161 55775
rect 261 55651 2161 55723
rect 261 55599 369 55651
rect 421 55599 493 55651
rect 545 55599 617 55651
rect 669 55599 741 55651
rect 793 55599 2161 55651
rect 261 55527 2161 55599
rect 261 55475 369 55527
rect 421 55475 493 55527
rect 545 55475 617 55527
rect 669 55475 741 55527
rect 793 55475 2161 55527
rect 261 55403 2161 55475
rect 261 55351 369 55403
rect 421 55351 493 55403
rect 545 55351 617 55403
rect 669 55351 741 55403
rect 793 55351 2161 55403
rect 261 55279 2161 55351
rect 261 55227 369 55279
rect 421 55227 493 55279
rect 545 55227 617 55279
rect 669 55227 741 55279
rect 793 55227 2161 55279
rect 261 55155 2161 55227
rect 261 55103 369 55155
rect 421 55103 493 55155
rect 545 55103 617 55155
rect 669 55103 741 55155
rect 793 55103 2161 55155
rect 261 55031 2161 55103
rect 261 54979 369 55031
rect 421 54979 493 55031
rect 545 54979 617 55031
rect 669 54979 741 55031
rect 793 54979 2161 55031
rect 261 54907 2161 54979
rect 261 54855 369 54907
rect 421 54855 493 54907
rect 545 54855 617 54907
rect 669 54855 741 54907
rect 793 54855 2161 54907
rect 261 54783 2161 54855
rect 261 54731 369 54783
rect 421 54731 493 54783
rect 545 54731 617 54783
rect 669 54731 741 54783
rect 793 54731 2161 54783
rect 261 54659 2161 54731
rect 261 54607 369 54659
rect 421 54607 493 54659
rect 545 54607 617 54659
rect 669 54607 741 54659
rect 793 54607 2161 54659
rect 261 54535 2161 54607
rect 261 54483 369 54535
rect 421 54483 493 54535
rect 545 54483 617 54535
rect 669 54483 741 54535
rect 793 54483 2161 54535
rect 261 54411 2161 54483
rect 261 54359 369 54411
rect 421 54359 493 54411
rect 545 54359 617 54411
rect 669 54359 741 54411
rect 793 54359 2161 54411
rect 261 54287 2161 54359
rect 261 54235 369 54287
rect 421 54235 493 54287
rect 545 54235 617 54287
rect 669 54235 741 54287
rect 793 54235 2161 54287
rect -11 54176 86 54186
rect -11 52824 20 54176
rect 76 52824 86 54176
rect -11 52814 86 52824
rect 261 54163 2161 54235
rect 261 54148 369 54163
rect 421 54148 493 54163
rect 545 54148 617 54163
rect 669 54148 741 54163
rect 793 54148 2161 54163
rect 261 54092 315 54148
rect 421 54111 439 54148
rect 545 54111 563 54148
rect 669 54111 687 54148
rect 793 54111 811 54148
rect 371 54092 439 54111
rect 495 54092 563 54111
rect 619 54092 687 54111
rect 743 54092 811 54111
rect 867 54092 935 54148
rect 991 54092 1059 54148
rect 1115 54092 1183 54148
rect 1239 54092 1307 54148
rect 1363 54092 1431 54148
rect 1487 54092 1555 54148
rect 1611 54092 1679 54148
rect 1735 54092 1803 54148
rect 1859 54092 1927 54148
rect 1983 54092 2051 54148
rect 2107 54092 2161 54148
rect 261 54039 2161 54092
rect 261 54024 369 54039
rect 421 54024 493 54039
rect 545 54024 617 54039
rect 669 54024 741 54039
rect 793 54024 2161 54039
rect 261 53968 315 54024
rect 421 53987 439 54024
rect 545 53987 563 54024
rect 669 53987 687 54024
rect 793 53987 811 54024
rect 371 53968 439 53987
rect 495 53968 563 53987
rect 619 53968 687 53987
rect 743 53968 811 53987
rect 867 53968 935 54024
rect 991 53968 1059 54024
rect 1115 53968 1183 54024
rect 1239 53968 1307 54024
rect 1363 53968 1431 54024
rect 1487 53968 1555 54024
rect 1611 53968 1679 54024
rect 1735 53968 1803 54024
rect 1859 53968 1927 54024
rect 1983 53968 2051 54024
rect 2107 53968 2161 54024
rect 261 53915 2161 53968
rect 261 53900 369 53915
rect 421 53900 493 53915
rect 545 53900 617 53915
rect 669 53900 741 53915
rect 793 53900 2161 53915
rect 261 53844 315 53900
rect 421 53863 439 53900
rect 545 53863 563 53900
rect 669 53863 687 53900
rect 793 53863 811 53900
rect 371 53844 439 53863
rect 495 53844 563 53863
rect 619 53844 687 53863
rect 743 53844 811 53863
rect 867 53844 935 53900
rect 991 53844 1059 53900
rect 1115 53844 1183 53900
rect 1239 53844 1307 53900
rect 1363 53844 1431 53900
rect 1487 53844 1555 53900
rect 1611 53844 1679 53900
rect 1735 53844 1803 53900
rect 1859 53844 1927 53900
rect 1983 53844 2051 53900
rect 2107 53844 2161 53900
rect 261 53791 2161 53844
rect 261 53776 369 53791
rect 421 53776 493 53791
rect 545 53776 617 53791
rect 669 53776 741 53791
rect 793 53776 2161 53791
rect 261 53720 315 53776
rect 421 53739 439 53776
rect 545 53739 563 53776
rect 669 53739 687 53776
rect 793 53739 811 53776
rect 371 53720 439 53739
rect 495 53720 563 53739
rect 619 53720 687 53739
rect 743 53720 811 53739
rect 867 53720 935 53776
rect 991 53720 1059 53776
rect 1115 53720 1183 53776
rect 1239 53720 1307 53776
rect 1363 53720 1431 53776
rect 1487 53720 1555 53776
rect 1611 53720 1679 53776
rect 1735 53720 1803 53776
rect 1859 53720 1927 53776
rect 1983 53720 2051 53776
rect 2107 53720 2161 53776
rect 261 53667 2161 53720
rect 261 53652 369 53667
rect 421 53652 493 53667
rect 545 53652 617 53667
rect 669 53652 741 53667
rect 793 53652 2161 53667
rect 261 53596 315 53652
rect 421 53615 439 53652
rect 545 53615 563 53652
rect 669 53615 687 53652
rect 793 53615 811 53652
rect 371 53596 439 53615
rect 495 53596 563 53615
rect 619 53596 687 53615
rect 743 53596 811 53615
rect 867 53596 935 53652
rect 991 53596 1059 53652
rect 1115 53596 1183 53652
rect 1239 53596 1307 53652
rect 1363 53596 1431 53652
rect 1487 53596 1555 53652
rect 1611 53596 1679 53652
rect 1735 53596 1803 53652
rect 1859 53596 1927 53652
rect 1983 53596 2051 53652
rect 2107 53596 2161 53652
rect 261 53543 2161 53596
rect 261 53528 369 53543
rect 421 53528 493 53543
rect 545 53528 617 53543
rect 669 53528 741 53543
rect 793 53528 2161 53543
rect 261 53472 315 53528
rect 421 53491 439 53528
rect 545 53491 563 53528
rect 669 53491 687 53528
rect 793 53491 811 53528
rect 371 53472 439 53491
rect 495 53472 563 53491
rect 619 53472 687 53491
rect 743 53472 811 53491
rect 867 53483 935 53528
rect 991 53483 1059 53528
rect 1115 53483 1183 53528
rect 1239 53483 1307 53528
rect 1363 53483 1431 53528
rect 1487 53483 1555 53528
rect 1611 53483 1679 53528
rect 1735 53483 1803 53528
rect 1859 53483 1927 53528
rect 1983 53483 2051 53528
rect 2107 53483 2161 53528
rect 867 53472 869 53483
rect 261 53431 869 53472
rect 921 53472 935 53483
rect 1029 53472 1059 53483
rect 1137 53472 1183 53483
rect 921 53431 977 53472
rect 1029 53431 1085 53472
rect 1137 53431 1193 53472
rect 1245 53431 1301 53483
rect 1363 53472 1409 53483
rect 1487 53472 1517 53483
rect 1611 53472 1625 53483
rect 1353 53431 1409 53472
rect 1461 53431 1517 53472
rect 1569 53431 1625 53472
rect 1677 53472 1679 53483
rect 1785 53472 1803 53483
rect 1893 53472 1927 53483
rect 2001 53472 2051 53483
rect 1677 53431 1733 53472
rect 1785 53431 1841 53472
rect 1893 53431 1949 53472
rect 2001 53431 2057 53472
rect 2109 53431 2161 53483
rect 261 53419 2161 53431
rect 261 53404 369 53419
rect 421 53404 493 53419
rect 545 53404 617 53419
rect 669 53404 741 53419
rect 793 53404 2161 53419
rect 261 53348 315 53404
rect 421 53367 439 53404
rect 545 53367 563 53404
rect 669 53367 687 53404
rect 793 53367 811 53404
rect 371 53348 439 53367
rect 495 53348 563 53367
rect 619 53348 687 53367
rect 743 53348 811 53367
rect 867 53375 935 53404
rect 991 53375 1059 53404
rect 1115 53375 1183 53404
rect 1239 53375 1307 53404
rect 1363 53375 1431 53404
rect 1487 53375 1555 53404
rect 1611 53375 1679 53404
rect 1735 53375 1803 53404
rect 1859 53375 1927 53404
rect 1983 53375 2051 53404
rect 2107 53375 2161 53404
rect 867 53348 869 53375
rect 261 53323 869 53348
rect 921 53348 935 53375
rect 1029 53348 1059 53375
rect 1137 53348 1183 53375
rect 921 53323 977 53348
rect 1029 53323 1085 53348
rect 1137 53323 1193 53348
rect 1245 53323 1301 53375
rect 1363 53348 1409 53375
rect 1487 53348 1517 53375
rect 1611 53348 1625 53375
rect 1353 53323 1409 53348
rect 1461 53323 1517 53348
rect 1569 53323 1625 53348
rect 1677 53348 1679 53375
rect 1785 53348 1803 53375
rect 1893 53348 1927 53375
rect 2001 53348 2051 53375
rect 1677 53323 1733 53348
rect 1785 53323 1841 53348
rect 1893 53323 1949 53348
rect 2001 53323 2057 53348
rect 2109 53323 2161 53375
rect 261 53295 2161 53323
rect 261 53280 369 53295
rect 421 53280 493 53295
rect 545 53280 617 53295
rect 669 53280 741 53295
rect 793 53280 2161 53295
rect 261 53224 315 53280
rect 421 53243 439 53280
rect 545 53243 563 53280
rect 669 53243 687 53280
rect 793 53243 811 53280
rect 371 53224 439 53243
rect 495 53224 563 53243
rect 619 53224 687 53243
rect 743 53224 811 53243
rect 867 53267 935 53280
rect 991 53267 1059 53280
rect 1115 53267 1183 53280
rect 1239 53267 1307 53280
rect 1363 53267 1431 53280
rect 1487 53267 1555 53280
rect 1611 53267 1679 53280
rect 1735 53267 1803 53280
rect 1859 53267 1927 53280
rect 1983 53267 2051 53280
rect 2107 53267 2161 53280
rect 867 53224 869 53267
rect 261 53215 869 53224
rect 921 53224 935 53267
rect 1029 53224 1059 53267
rect 1137 53224 1183 53267
rect 921 53215 977 53224
rect 1029 53215 1085 53224
rect 1137 53215 1193 53224
rect 1245 53215 1301 53267
rect 1363 53224 1409 53267
rect 1487 53224 1517 53267
rect 1611 53224 1625 53267
rect 1353 53215 1409 53224
rect 1461 53215 1517 53224
rect 1569 53215 1625 53224
rect 1677 53224 1679 53267
rect 1785 53224 1803 53267
rect 1893 53224 1927 53267
rect 2001 53224 2051 53267
rect 1677 53215 1733 53224
rect 1785 53215 1841 53224
rect 1893 53215 1949 53224
rect 2001 53215 2057 53224
rect 2109 53215 2161 53267
rect 261 53156 2161 53215
rect 261 53100 315 53156
rect 371 53100 439 53156
rect 495 53100 563 53156
rect 619 53100 687 53156
rect 743 53100 811 53156
rect 867 53100 935 53156
rect 991 53100 1059 53156
rect 1115 53100 1183 53156
rect 1239 53100 1307 53156
rect 1363 53100 1431 53156
rect 1487 53100 1555 53156
rect 1611 53100 1679 53156
rect 1735 53100 1803 53156
rect 1859 53100 1927 53156
rect 1983 53100 2051 53156
rect 2107 53100 2161 53156
rect 261 53032 2161 53100
rect 261 52976 315 53032
rect 371 52976 439 53032
rect 495 52976 563 53032
rect 619 52976 687 53032
rect 743 52976 811 53032
rect 867 52976 935 53032
rect 991 52976 1059 53032
rect 1115 52976 1183 53032
rect 1239 52976 1307 53032
rect 1363 52976 1431 53032
rect 1487 52976 1555 53032
rect 1611 52976 1679 53032
rect 1735 52976 1803 53032
rect 1859 52976 1927 53032
rect 1983 52976 2051 53032
rect 2107 52976 2161 53032
rect 261 52908 2161 52976
rect 261 52852 315 52908
rect 371 52852 439 52908
rect 495 52852 563 52908
rect 619 52852 687 52908
rect 743 52852 811 52908
rect 867 52852 935 52908
rect 991 52852 1059 52908
rect 1115 52852 1183 52908
rect 1239 52852 1307 52908
rect 1363 52852 1431 52908
rect 1487 52852 1555 52908
rect 1611 52852 1679 52908
rect 1735 52852 1803 52908
rect 1859 52852 1927 52908
rect 1983 52852 2051 52908
rect 2107 52852 2161 52908
rect -11 52576 86 52600
rect -11 51224 20 52576
rect 76 51224 86 52576
rect -11 51200 86 51224
rect 261 52548 2161 52852
rect 261 52492 315 52548
rect 371 52492 439 52548
rect 495 52492 563 52548
rect 619 52492 687 52548
rect 743 52492 811 52548
rect 867 52492 935 52548
rect 991 52492 1059 52548
rect 1115 52492 1183 52548
rect 1239 52492 1307 52548
rect 1363 52492 1431 52548
rect 1487 52492 1555 52548
rect 1611 52492 1679 52548
rect 1735 52492 1803 52548
rect 1859 52492 1927 52548
rect 1983 52492 2051 52548
rect 2107 52492 2161 52548
rect 261 52424 2161 52492
rect 261 52368 315 52424
rect 371 52368 439 52424
rect 495 52368 563 52424
rect 619 52368 687 52424
rect 743 52368 811 52424
rect 867 52368 935 52424
rect 991 52368 1059 52424
rect 1115 52368 1183 52424
rect 1239 52368 1307 52424
rect 1363 52368 1431 52424
rect 1487 52368 1555 52424
rect 1611 52368 1679 52424
rect 1735 52368 1803 52424
rect 1859 52368 1927 52424
rect 1983 52368 2051 52424
rect 2107 52368 2161 52424
rect 261 52300 2161 52368
rect 261 52244 315 52300
rect 371 52244 439 52300
rect 495 52244 563 52300
rect 619 52244 687 52300
rect 743 52244 811 52300
rect 867 52244 935 52300
rect 991 52244 1059 52300
rect 1115 52244 1183 52300
rect 1239 52244 1307 52300
rect 1363 52244 1431 52300
rect 1487 52244 1555 52300
rect 1611 52244 1679 52300
rect 1735 52244 1803 52300
rect 1859 52244 1927 52300
rect 1983 52244 2051 52300
rect 2107 52244 2161 52300
rect 261 52176 2161 52244
rect 261 52120 315 52176
rect 371 52120 439 52176
rect 495 52120 563 52176
rect 619 52120 687 52176
rect 743 52120 811 52176
rect 867 52120 935 52176
rect 991 52120 1059 52176
rect 1115 52120 1183 52176
rect 1239 52120 1307 52176
rect 1363 52120 1431 52176
rect 1487 52120 1555 52176
rect 1611 52120 1679 52176
rect 1735 52120 1803 52176
rect 1859 52120 1927 52176
rect 1983 52120 2051 52176
rect 2107 52120 2161 52176
rect 261 52052 2161 52120
rect 261 51996 315 52052
rect 371 51996 439 52052
rect 495 51996 563 52052
rect 619 51996 687 52052
rect 743 51996 811 52052
rect 867 51996 935 52052
rect 991 51996 1059 52052
rect 1115 51996 1183 52052
rect 1239 51996 1307 52052
rect 1363 51996 1431 52052
rect 1487 51996 1555 52052
rect 1611 51996 1679 52052
rect 1735 51996 1803 52052
rect 1859 51996 1927 52052
rect 1983 51996 2051 52052
rect 2107 51996 2161 52052
rect 261 51928 2161 51996
rect 261 51872 315 51928
rect 371 51872 439 51928
rect 495 51872 563 51928
rect 619 51872 687 51928
rect 743 51872 811 51928
rect 867 51872 935 51928
rect 991 51872 1059 51928
rect 1115 51872 1183 51928
rect 1239 51872 1307 51928
rect 1363 51872 1431 51928
rect 1487 51872 1555 51928
rect 1611 51872 1679 51928
rect 1735 51872 1803 51928
rect 1859 51872 1927 51928
rect 1983 51872 2051 51928
rect 2107 51872 2161 51928
rect 261 51804 2161 51872
rect 261 51748 315 51804
rect 371 51748 439 51804
rect 495 51748 563 51804
rect 619 51748 687 51804
rect 743 51748 811 51804
rect 867 51748 935 51804
rect 991 51748 1059 51804
rect 1115 51748 1183 51804
rect 1239 51748 1307 51804
rect 1363 51748 1431 51804
rect 1487 51748 1555 51804
rect 1611 51748 1679 51804
rect 1735 51748 1803 51804
rect 1859 51748 1927 51804
rect 1983 51748 2051 51804
rect 2107 51748 2161 51804
rect 261 51680 2161 51748
rect 261 51624 315 51680
rect 371 51624 439 51680
rect 495 51624 563 51680
rect 619 51624 687 51680
rect 743 51624 811 51680
rect 867 51624 935 51680
rect 991 51624 1059 51680
rect 1115 51624 1183 51680
rect 1239 51624 1307 51680
rect 1363 51624 1431 51680
rect 1487 51624 1555 51680
rect 1611 51624 1679 51680
rect 1735 51624 1803 51680
rect 1859 51624 1927 51680
rect 1983 51624 2051 51680
rect 2107 51624 2161 51680
rect 261 51556 2161 51624
rect 261 51500 315 51556
rect 371 51500 439 51556
rect 495 51500 563 51556
rect 619 51500 687 51556
rect 743 51500 811 51556
rect 867 51500 935 51556
rect 991 51500 1059 51556
rect 1115 51500 1183 51556
rect 1239 51500 1307 51556
rect 1363 51500 1431 51556
rect 1487 51500 1555 51556
rect 1611 51500 1679 51556
rect 1735 51500 1803 51556
rect 1859 51500 1927 51556
rect 1983 51500 2051 51556
rect 2107 51500 2161 51556
rect 261 51432 2161 51500
rect 261 51376 315 51432
rect 371 51376 439 51432
rect 495 51376 563 51432
rect 619 51376 687 51432
rect 743 51376 811 51432
rect 867 51376 935 51432
rect 991 51376 1059 51432
rect 1115 51376 1183 51432
rect 1239 51376 1307 51432
rect 1363 51376 1431 51432
rect 1487 51376 1555 51432
rect 1611 51376 1679 51432
rect 1735 51376 1803 51432
rect 1859 51376 1927 51432
rect 1983 51376 2051 51432
rect 2107 51376 2161 51432
rect 261 51308 2161 51376
rect 261 51252 315 51308
rect 371 51252 439 51308
rect 495 51252 563 51308
rect 619 51252 687 51308
rect 743 51252 811 51308
rect 867 51252 935 51308
rect 991 51252 1059 51308
rect 1115 51252 1183 51308
rect 1239 51252 1307 51308
rect 1363 51252 1431 51308
rect 1487 51252 1555 51308
rect 1611 51252 1679 51308
rect 1735 51252 1803 51308
rect 1859 51252 1927 51308
rect 1983 51252 2051 51308
rect 2107 51252 2161 51308
rect -11 49376 86 49386
rect -11 48024 20 49376
rect 76 48024 86 49376
rect -11 48014 86 48024
rect 261 49348 2161 51252
rect 2481 56741 2681 57278
rect 2481 56689 2501 56741
rect 2553 56689 2609 56741
rect 2661 56689 2681 56741
rect 2481 55748 2681 56689
rect 2481 55692 2491 55748
rect 2547 55692 2615 55748
rect 2671 55692 2681 55748
rect 2481 55624 2681 55692
rect 2481 55568 2491 55624
rect 2547 55568 2615 55624
rect 2671 55568 2681 55624
rect 2481 55500 2681 55568
rect 2481 55444 2491 55500
rect 2547 55444 2615 55500
rect 2671 55444 2681 55500
rect 2481 55376 2681 55444
rect 2481 55320 2491 55376
rect 2547 55320 2615 55376
rect 2671 55320 2681 55376
rect 2481 55252 2681 55320
rect 2481 55196 2491 55252
rect 2547 55196 2615 55252
rect 2671 55196 2681 55252
rect 2481 55128 2681 55196
rect 2481 55072 2491 55128
rect 2547 55072 2615 55128
rect 2671 55072 2681 55128
rect 2481 55004 2681 55072
rect 2481 54948 2491 55004
rect 2547 54948 2615 55004
rect 2671 54948 2681 55004
rect 2481 54880 2681 54948
rect 2481 54824 2491 54880
rect 2547 54824 2615 54880
rect 2671 54824 2681 54880
rect 2481 54756 2681 54824
rect 2481 54700 2491 54756
rect 2547 54700 2615 54756
rect 2671 54700 2681 54756
rect 2481 54632 2681 54700
rect 2481 54576 2491 54632
rect 2547 54576 2615 54632
rect 2671 54576 2681 54632
rect 2481 54508 2681 54576
rect 2481 54452 2491 54508
rect 2547 54452 2615 54508
rect 2671 54452 2681 54508
rect 2481 53621 2681 54452
rect 2481 53569 2501 53621
rect 2553 53569 2609 53621
rect 2661 53569 2681 53621
rect 2481 52594 2681 53569
rect 2481 52542 2590 52594
rect 2642 52542 2681 52594
rect 2481 52486 2681 52542
rect 2481 52434 2590 52486
rect 2642 52434 2681 52486
rect 2481 52378 2681 52434
rect 2481 52326 2590 52378
rect 2642 52326 2681 52378
rect 2481 52270 2681 52326
rect 2481 52218 2590 52270
rect 2642 52218 2681 52270
rect 2481 52162 2681 52218
rect 2481 52110 2590 52162
rect 2642 52110 2681 52162
rect 2481 52054 2681 52110
rect 2481 52002 2590 52054
rect 2642 52002 2681 52054
rect 2481 51946 2681 52002
rect 2481 51894 2590 51946
rect 2642 51894 2681 51946
rect 2481 51838 2681 51894
rect 2481 51786 2590 51838
rect 2642 51786 2681 51838
rect 2481 51730 2681 51786
rect 2481 51678 2590 51730
rect 2642 51678 2681 51730
rect 2481 51622 2681 51678
rect 2481 51570 2590 51622
rect 2642 51570 2681 51622
rect 2481 51514 2681 51570
rect 2481 51462 2590 51514
rect 2642 51462 2681 51514
rect 2481 51406 2681 51462
rect 2481 51354 2590 51406
rect 2642 51354 2681 51406
rect 2481 51298 2681 51354
rect 2481 51246 2590 51298
rect 2642 51246 2681 51298
rect 2481 51190 2681 51246
rect 2481 51138 2590 51190
rect 2642 51138 2681 51190
rect 2481 51082 2681 51138
rect 2481 51030 2590 51082
rect 2642 51030 2681 51082
rect 261 49292 315 49348
rect 371 49292 439 49348
rect 495 49292 563 49348
rect 619 49292 687 49348
rect 743 49292 811 49348
rect 867 49292 935 49348
rect 991 49292 1059 49348
rect 1115 49292 1183 49348
rect 1239 49292 1307 49348
rect 1363 49292 1431 49348
rect 1487 49292 1555 49348
rect 1611 49292 1679 49348
rect 1735 49292 1803 49348
rect 1859 49292 1927 49348
rect 1983 49292 2051 49348
rect 2107 49292 2161 49348
rect 261 49224 2161 49292
rect 261 49168 315 49224
rect 371 49168 439 49224
rect 495 49168 563 49224
rect 619 49168 687 49224
rect 743 49168 811 49224
rect 867 49168 935 49224
rect 991 49168 1059 49224
rect 1115 49168 1183 49224
rect 1239 49168 1307 49224
rect 1363 49168 1431 49224
rect 1487 49168 1555 49224
rect 1611 49168 1679 49224
rect 1735 49168 1803 49224
rect 1859 49168 1927 49224
rect 1983 49168 2051 49224
rect 2107 49168 2161 49224
rect 261 49100 2161 49168
rect 261 49044 315 49100
rect 371 49044 439 49100
rect 495 49044 563 49100
rect 619 49044 687 49100
rect 743 49044 811 49100
rect 867 49044 935 49100
rect 991 49044 1059 49100
rect 1115 49044 1183 49100
rect 1239 49044 1307 49100
rect 1363 49044 1431 49100
rect 1487 49044 1555 49100
rect 1611 49044 1679 49100
rect 1735 49044 1803 49100
rect 1859 49044 1927 49100
rect 1983 49044 2051 49100
rect 2107 49044 2161 49100
rect 261 48976 2161 49044
rect 261 48920 315 48976
rect 371 48920 439 48976
rect 495 48920 563 48976
rect 619 48920 687 48976
rect 743 48920 811 48976
rect 867 48920 935 48976
rect 991 48920 1059 48976
rect 1115 48920 1183 48976
rect 1239 48920 1307 48976
rect 1363 48920 1431 48976
rect 1487 48920 1555 48976
rect 1611 48920 1679 48976
rect 1735 48920 1803 48976
rect 1859 48920 1927 48976
rect 1983 48920 2051 48976
rect 2107 48920 2161 48976
rect 261 48852 2161 48920
rect 261 48796 315 48852
rect 371 48796 439 48852
rect 495 48796 563 48852
rect 619 48796 687 48852
rect 743 48796 811 48852
rect 867 48796 935 48852
rect 991 48796 1059 48852
rect 1115 48796 1183 48852
rect 1239 48796 1307 48852
rect 1363 48796 1431 48852
rect 1487 48796 1555 48852
rect 1611 48796 1679 48852
rect 1735 48796 1803 48852
rect 1859 48796 1927 48852
rect 1983 48796 2051 48852
rect 2107 48796 2161 48852
rect 261 48728 2161 48796
rect 261 48672 315 48728
rect 371 48672 439 48728
rect 495 48672 563 48728
rect 619 48672 687 48728
rect 743 48672 811 48728
rect 867 48672 935 48728
rect 991 48672 1059 48728
rect 1115 48672 1183 48728
rect 1239 48672 1307 48728
rect 1363 48672 1431 48728
rect 1487 48672 1555 48728
rect 1611 48672 1679 48728
rect 1735 48672 1803 48728
rect 1859 48672 1927 48728
rect 1983 48672 2051 48728
rect 2107 48672 2161 48728
rect 261 48604 2161 48672
rect 261 48548 315 48604
rect 371 48548 439 48604
rect 495 48548 563 48604
rect 619 48548 687 48604
rect 743 48548 811 48604
rect 867 48548 935 48604
rect 991 48548 1059 48604
rect 1115 48548 1183 48604
rect 1239 48548 1307 48604
rect 1363 48548 1431 48604
rect 1487 48548 1555 48604
rect 1611 48548 1679 48604
rect 1735 48548 1803 48604
rect 1859 48548 1927 48604
rect 1983 48548 2051 48604
rect 2107 48548 2161 48604
rect 261 48480 2161 48548
rect 261 48424 315 48480
rect 371 48424 439 48480
rect 495 48424 563 48480
rect 619 48424 687 48480
rect 743 48424 811 48480
rect 867 48424 935 48480
rect 991 48424 1059 48480
rect 1115 48424 1183 48480
rect 1239 48424 1307 48480
rect 1363 48424 1431 48480
rect 1487 48424 1555 48480
rect 1611 48424 1679 48480
rect 1735 48424 1803 48480
rect 1859 48424 1927 48480
rect 1983 48424 2051 48480
rect 2107 48424 2161 48480
rect 261 48356 2161 48424
rect 261 48300 315 48356
rect 371 48300 439 48356
rect 495 48300 563 48356
rect 619 48300 687 48356
rect 743 48300 811 48356
rect 867 48300 935 48356
rect 991 48300 1059 48356
rect 1115 48300 1183 48356
rect 1239 48300 1307 48356
rect 1363 48300 1431 48356
rect 1487 48300 1555 48356
rect 1611 48300 1679 48356
rect 1735 48300 1803 48356
rect 1859 48300 1927 48356
rect 1983 48300 2051 48356
rect 2107 48300 2161 48356
rect 261 48232 2161 48300
rect 261 48176 315 48232
rect 371 48176 439 48232
rect 495 48176 563 48232
rect 619 48176 687 48232
rect 743 48176 811 48232
rect 867 48176 935 48232
rect 991 48176 1059 48232
rect 1115 48176 1183 48232
rect 1239 48176 1307 48232
rect 1363 48176 1431 48232
rect 1487 48176 1555 48232
rect 1611 48176 1679 48232
rect 1735 48176 1803 48232
rect 1859 48176 1927 48232
rect 1983 48176 2051 48232
rect 2107 48176 2161 48232
rect 261 48108 2161 48176
rect 261 48052 315 48108
rect 371 48052 439 48108
rect 495 48052 563 48108
rect 619 48052 687 48108
rect 743 48052 811 48108
rect 867 48052 935 48108
rect 991 48052 1059 48108
rect 1115 48052 1183 48108
rect 1239 48052 1307 48108
rect 1363 48052 1431 48108
rect 1487 48052 1555 48108
rect 1611 48052 1679 48108
rect 1735 48052 1803 48108
rect 1859 48052 1927 48108
rect 1983 48052 2051 48108
rect 2107 48052 2161 48108
rect 261 47163 2161 48052
rect 2292 50926 2368 51000
rect 2292 50870 2302 50926
rect 2358 50870 2368 50926
rect 2292 50794 2368 50870
rect 2292 50738 2302 50794
rect 2358 50738 2368 50794
rect 2292 50662 2368 50738
rect 2292 50606 2302 50662
rect 2358 50606 2368 50662
rect 2292 50530 2368 50606
rect 2292 50474 2302 50530
rect 2358 50474 2368 50530
rect 2292 50398 2368 50474
rect 2292 50342 2302 50398
rect 2358 50342 2368 50398
rect 2292 50266 2368 50342
rect 2292 50210 2302 50266
rect 2358 50210 2368 50266
rect 2292 50134 2368 50210
rect 2292 50078 2302 50134
rect 2358 50078 2368 50134
rect 2292 50002 2368 50078
rect 2292 49946 2302 50002
rect 2358 49946 2368 50002
rect 2292 49870 2368 49946
rect 2292 49814 2302 49870
rect 2358 49814 2368 49870
rect 2292 49738 2368 49814
rect 2292 49682 2302 49738
rect 2358 49682 2368 49738
rect -11 46176 86 46186
rect -11 44824 20 46176
rect 76 44824 86 46176
rect 305 46148 2117 46158
rect 305 46092 315 46148
rect 371 46092 439 46148
rect 495 46092 563 46148
rect 619 46092 687 46148
rect 743 46092 811 46148
rect 867 46092 935 46148
rect 991 46092 1059 46148
rect 1115 46092 1183 46148
rect 1239 46092 1307 46148
rect 1363 46092 1431 46148
rect 1487 46092 1555 46148
rect 1611 46092 1679 46148
rect 1735 46092 1803 46148
rect 1859 46092 1927 46148
rect 1983 46092 2051 46148
rect 2107 46092 2117 46148
rect 305 46024 2117 46092
rect 305 45968 315 46024
rect 371 45968 439 46024
rect 495 45968 563 46024
rect 619 45968 687 46024
rect 743 45968 811 46024
rect 867 45968 935 46024
rect 991 45968 1059 46024
rect 1115 45968 1183 46024
rect 1239 45968 1307 46024
rect 1363 45968 1431 46024
rect 1487 45968 1555 46024
rect 1611 45968 1679 46024
rect 1735 45968 1803 46024
rect 1859 45968 1927 46024
rect 1983 45968 2051 46024
rect 2107 45968 2117 46024
rect 305 45900 2117 45968
rect 305 45844 315 45900
rect 371 45844 439 45900
rect 495 45844 563 45900
rect 619 45844 687 45900
rect 743 45844 811 45900
rect 867 45844 935 45900
rect 991 45844 1059 45900
rect 1115 45844 1183 45900
rect 1239 45844 1307 45900
rect 1363 45844 1431 45900
rect 1487 45844 1555 45900
rect 1611 45844 1679 45900
rect 1735 45844 1803 45900
rect 1859 45844 1927 45900
rect 1983 45844 2051 45900
rect 2107 45844 2117 45900
rect 305 45776 2117 45844
rect 305 45720 315 45776
rect 371 45720 439 45776
rect 495 45720 563 45776
rect 619 45720 687 45776
rect 743 45720 811 45776
rect 867 45720 935 45776
rect 991 45720 1059 45776
rect 1115 45720 1183 45776
rect 1239 45720 1307 45776
rect 1363 45720 1431 45776
rect 1487 45720 1555 45776
rect 1611 45720 1679 45776
rect 1735 45720 1803 45776
rect 1859 45720 1927 45776
rect 1983 45720 2051 45776
rect 2107 45720 2117 45776
rect 305 45652 2117 45720
rect 305 45596 315 45652
rect 371 45596 439 45652
rect 495 45596 563 45652
rect 619 45596 687 45652
rect 743 45596 811 45652
rect 867 45596 935 45652
rect 991 45596 1059 45652
rect 1115 45596 1183 45652
rect 1239 45596 1307 45652
rect 1363 45596 1431 45652
rect 1487 45596 1555 45652
rect 1611 45596 1679 45652
rect 1735 45596 1803 45652
rect 1859 45596 1927 45652
rect 1983 45596 2051 45652
rect 2107 45596 2117 45652
rect 305 45528 2117 45596
rect 305 45472 315 45528
rect 371 45472 439 45528
rect 495 45472 563 45528
rect 619 45472 687 45528
rect 743 45472 811 45528
rect 867 45472 935 45528
rect 991 45472 1059 45528
rect 1115 45472 1183 45528
rect 1239 45472 1307 45528
rect 1363 45472 1431 45528
rect 1487 45472 1555 45528
rect 1611 45472 1679 45528
rect 1735 45472 1803 45528
rect 1859 45472 1927 45528
rect 1983 45472 2051 45528
rect 2107 45472 2117 45528
rect 305 45404 2117 45472
rect 305 45348 315 45404
rect 371 45348 439 45404
rect 495 45348 563 45404
rect 619 45348 687 45404
rect 743 45348 811 45404
rect 867 45348 935 45404
rect 991 45348 1059 45404
rect 1115 45348 1183 45404
rect 1239 45348 1307 45404
rect 1363 45348 1431 45404
rect 1487 45348 1555 45404
rect 1611 45348 1679 45404
rect 1735 45348 1803 45404
rect 1859 45348 1927 45404
rect 1983 45348 2051 45404
rect 2107 45348 2117 45404
rect 305 45280 2117 45348
rect 305 45224 315 45280
rect 371 45224 439 45280
rect 495 45224 563 45280
rect 619 45224 687 45280
rect 743 45224 811 45280
rect 867 45224 935 45280
rect 991 45224 1059 45280
rect 1115 45224 1183 45280
rect 1239 45224 1307 45280
rect 1363 45224 1431 45280
rect 1487 45224 1555 45280
rect 1611 45224 1679 45280
rect 1735 45224 1803 45280
rect 1859 45224 1927 45280
rect 1983 45224 2051 45280
rect 2107 45224 2117 45280
rect 305 45156 2117 45224
rect 305 45100 315 45156
rect 371 45100 439 45156
rect 495 45100 563 45156
rect 619 45100 687 45156
rect 743 45100 811 45156
rect 867 45100 935 45156
rect 991 45100 1059 45156
rect 1115 45100 1183 45156
rect 1239 45100 1307 45156
rect 1363 45100 1431 45156
rect 1487 45100 1555 45156
rect 1611 45100 1679 45156
rect 1735 45100 1803 45156
rect 1859 45100 1927 45156
rect 1983 45100 2051 45156
rect 2107 45100 2117 45156
rect 305 45032 2117 45100
rect 305 44976 315 45032
rect 371 44976 439 45032
rect 495 44976 563 45032
rect 619 44976 687 45032
rect 743 44976 811 45032
rect 867 44976 935 45032
rect 991 44976 1059 45032
rect 1115 44976 1183 45032
rect 1239 44976 1307 45032
rect 1363 44976 1431 45032
rect 1487 44976 1555 45032
rect 1611 44976 1679 45032
rect 1735 44976 1803 45032
rect 1859 44976 1927 45032
rect 1983 44976 2051 45032
rect 2107 44976 2117 45032
rect 305 44908 2117 44976
rect 305 44852 315 44908
rect 371 44852 439 44908
rect 495 44852 563 44908
rect 619 44852 687 44908
rect 743 44852 811 44908
rect 867 44852 935 44908
rect 991 44852 1059 44908
rect 1115 44852 1183 44908
rect 1239 44852 1307 44908
rect 1363 44852 1431 44908
rect 1487 44852 1555 44908
rect 1611 44852 1679 44908
rect 1735 44852 1803 44908
rect 1859 44852 1927 44908
rect 1983 44852 2051 44908
rect 2107 44852 2117 44908
rect 305 44842 2117 44852
rect -11 44814 86 44824
rect 2292 39727 2368 49682
rect 2481 50974 2681 51030
rect 2481 50922 2590 50974
rect 2642 50922 2681 50974
rect 2481 50866 2681 50922
rect 2481 50814 2590 50866
rect 2642 50814 2681 50866
rect 2481 50758 2681 50814
rect 2481 50706 2590 50758
rect 2642 50706 2681 50758
rect 2481 50650 2681 50706
rect 2481 50598 2590 50650
rect 2642 50598 2681 50650
rect 2481 50542 2681 50598
rect 2481 50490 2590 50542
rect 2642 50490 2681 50542
rect 2481 50434 2681 50490
rect 2481 50382 2590 50434
rect 2642 50382 2681 50434
rect 2481 50326 2681 50382
rect 2481 50274 2590 50326
rect 2642 50274 2681 50326
rect 2481 50218 2681 50274
rect 2481 50166 2590 50218
rect 2642 50166 2681 50218
rect 2481 50110 2681 50166
rect 2481 50058 2590 50110
rect 2642 50058 2681 50110
rect 2481 50002 2681 50058
rect 2481 49950 2590 50002
rect 2642 49950 2681 50002
rect 2481 49894 2681 49950
rect 2481 49842 2590 49894
rect 2642 49842 2681 49894
rect 2481 49786 2681 49842
rect 2481 49734 2590 49786
rect 2642 49734 2681 49786
rect 2481 49678 2681 49734
rect 2481 49626 2590 49678
rect 2642 49626 2681 49678
rect 2481 49570 2681 49626
rect 2481 49518 2590 49570
rect 2642 49518 2681 49570
rect 2481 49462 2681 49518
rect 2481 49410 2590 49462
rect 2642 49410 2681 49462
rect 2481 49354 2681 49410
rect 2481 49302 2590 49354
rect 2642 49302 2681 49354
rect 2481 49246 2681 49302
rect 2481 49194 2590 49246
rect 2642 49194 2681 49246
rect 2481 49138 2681 49194
rect 2481 49086 2590 49138
rect 2642 49086 2681 49138
rect 2481 49030 2681 49086
rect 2481 48978 2590 49030
rect 2642 48978 2681 49030
rect 2481 48922 2681 48978
rect 2481 48870 2590 48922
rect 2642 48870 2681 48922
rect 2481 48814 2681 48870
rect 2481 48762 2590 48814
rect 2642 48762 2681 48814
rect 2481 48706 2681 48762
rect 2481 48654 2590 48706
rect 2642 48654 2681 48706
rect 2481 48598 2681 48654
rect 2481 48546 2590 48598
rect 2642 48546 2681 48598
rect 2481 48490 2681 48546
rect 2481 48438 2590 48490
rect 2642 48438 2681 48490
rect 2481 48382 2681 48438
rect 2481 48330 2590 48382
rect 2642 48330 2681 48382
rect 2481 48274 2681 48330
rect 2481 48222 2590 48274
rect 2642 48222 2681 48274
rect 2481 48166 2681 48222
rect 2481 48114 2590 48166
rect 2642 48114 2681 48166
rect 2481 48058 2681 48114
rect 2481 48006 2590 48058
rect 2642 48006 2681 48058
rect 2481 47950 2681 48006
rect 2481 47898 2590 47950
rect 2642 47898 2681 47950
rect 2481 47842 2681 47898
rect 2481 47790 2590 47842
rect 2642 47790 2681 47842
rect 2481 47748 2681 47790
rect 2481 47692 2491 47748
rect 2547 47734 2615 47748
rect 2547 47692 2590 47734
rect 2671 47692 2681 47748
rect 2481 47682 2590 47692
rect 2642 47682 2681 47692
rect 2481 47624 2681 47682
rect 2481 47568 2491 47624
rect 2547 47568 2615 47624
rect 2671 47568 2681 47624
rect 2481 47500 2681 47568
rect 2481 47444 2491 47500
rect 2547 47444 2615 47500
rect 2671 47444 2681 47500
rect 2481 47376 2681 47444
rect 2481 47320 2491 47376
rect 2547 47320 2615 47376
rect 2671 47320 2681 47376
rect 2481 47252 2681 47320
rect 2481 47196 2491 47252
rect 2547 47196 2615 47252
rect 2671 47196 2681 47252
rect 2481 47128 2681 47196
rect 2741 57225 4791 57447
rect 5111 57499 7161 57600
rect 5111 57447 5246 57499
rect 5298 57447 5354 57499
rect 5406 57447 5462 57499
rect 5514 57447 5570 57499
rect 5622 57447 5678 57499
rect 5730 57447 5786 57499
rect 5838 57447 5894 57499
rect 5946 57447 6002 57499
rect 6054 57447 6110 57499
rect 6162 57447 6218 57499
rect 6270 57447 6326 57499
rect 6378 57447 6434 57499
rect 6486 57447 6542 57499
rect 6594 57447 6650 57499
rect 6702 57447 6758 57499
rect 6810 57447 6866 57499
rect 6918 57447 6974 57499
rect 7026 57447 7161 57499
rect 2741 57169 2808 57225
rect 2864 57169 2932 57225
rect 2988 57169 3056 57225
rect 3112 57169 3180 57225
rect 3236 57169 3304 57225
rect 3360 57169 3428 57225
rect 3484 57169 3552 57225
rect 3608 57169 3676 57225
rect 3732 57169 3800 57225
rect 3856 57169 3924 57225
rect 3980 57169 4048 57225
rect 4104 57169 4172 57225
rect 4228 57169 4296 57225
rect 4352 57169 4420 57225
rect 4476 57169 4544 57225
rect 4600 57169 4668 57225
rect 4724 57169 4791 57225
rect 2741 57104 4791 57169
rect 2741 57052 2768 57104
rect 2820 57101 2876 57104
rect 2864 57052 2876 57101
rect 2928 57101 2984 57104
rect 3036 57101 3092 57104
rect 3144 57101 3200 57104
rect 3252 57101 3308 57104
rect 2928 57052 2932 57101
rect 3036 57052 3056 57101
rect 3144 57052 3180 57101
rect 3252 57052 3304 57101
rect 3360 57052 3416 57104
rect 3468 57101 3524 57104
rect 3576 57101 3632 57104
rect 3684 57101 3740 57104
rect 3484 57052 3524 57101
rect 3608 57052 3632 57101
rect 3732 57052 3740 57101
rect 3792 57101 3848 57104
rect 3900 57101 3956 57104
rect 4008 57101 4064 57104
rect 3792 57052 3800 57101
rect 3900 57052 3924 57101
rect 4008 57052 4048 57101
rect 4116 57052 4172 57104
rect 4224 57101 4280 57104
rect 4332 57101 4388 57104
rect 4440 57101 4496 57104
rect 4548 57101 4604 57104
rect 4228 57052 4280 57101
rect 4352 57052 4388 57101
rect 4476 57052 4496 57101
rect 4600 57052 4604 57101
rect 4656 57101 4712 57104
rect 4656 57052 4668 57101
rect 4764 57052 4791 57104
rect 2741 57045 2808 57052
rect 2864 57045 2932 57052
rect 2988 57045 3056 57052
rect 3112 57045 3180 57052
rect 3236 57045 3304 57052
rect 3360 57045 3428 57052
rect 3484 57045 3552 57052
rect 3608 57045 3676 57052
rect 3732 57045 3800 57052
rect 3856 57045 3924 57052
rect 3980 57045 4048 57052
rect 4104 57045 4172 57052
rect 4228 57045 4296 57052
rect 4352 57045 4420 57052
rect 4476 57045 4544 57052
rect 4600 57045 4668 57052
rect 4724 57045 4791 57052
rect 2741 56977 4791 57045
rect 2741 56921 2808 56977
rect 2864 56921 2932 56977
rect 2988 56921 3056 56977
rect 3112 56921 3180 56977
rect 3236 56921 3304 56977
rect 3360 56921 3428 56977
rect 3484 56921 3552 56977
rect 3608 56921 3676 56977
rect 3732 56921 3800 56977
rect 3856 56921 3924 56977
rect 3980 56921 4048 56977
rect 4104 56921 4172 56977
rect 4228 56921 4296 56977
rect 4352 56921 4420 56977
rect 4476 56921 4544 56977
rect 4600 56921 4668 56977
rect 4724 56921 4791 56977
rect 2741 56853 4791 56921
rect 2741 56797 2808 56853
rect 2864 56797 2932 56853
rect 2988 56797 3056 56853
rect 3112 56797 3180 56853
rect 3236 56797 3304 56853
rect 3360 56797 3428 56853
rect 3484 56797 3552 56853
rect 3608 56797 3676 56853
rect 3732 56797 3800 56853
rect 3856 56797 3924 56853
rect 3980 56797 4048 56853
rect 4104 56797 4172 56853
rect 4228 56797 4296 56853
rect 4352 56797 4420 56853
rect 4476 56797 4544 56853
rect 4600 56797 4668 56853
rect 4724 56797 4791 56853
rect 2741 56729 4791 56797
rect 2741 56673 2808 56729
rect 2864 56673 2932 56729
rect 2988 56673 3056 56729
rect 3112 56673 3180 56729
rect 3236 56673 3304 56729
rect 3360 56673 3428 56729
rect 3484 56673 3552 56729
rect 3608 56673 3676 56729
rect 3732 56673 3800 56729
rect 3856 56673 3924 56729
rect 3980 56673 4048 56729
rect 4104 56673 4172 56729
rect 4228 56673 4296 56729
rect 4352 56673 4420 56729
rect 4476 56673 4544 56729
rect 4600 56673 4668 56729
rect 4724 56673 4791 56729
rect 2741 56643 4791 56673
rect 2741 56605 3903 56643
rect 3955 56605 4027 56643
rect 4079 56605 4151 56643
rect 4203 56605 4791 56643
rect 2741 56549 2808 56605
rect 2864 56549 2932 56605
rect 2988 56549 3056 56605
rect 3112 56549 3180 56605
rect 3236 56549 3304 56605
rect 3360 56549 3428 56605
rect 3484 56549 3552 56605
rect 3608 56549 3676 56605
rect 3732 56549 3800 56605
rect 3856 56591 3903 56605
rect 3980 56591 4027 56605
rect 4104 56591 4151 56605
rect 3856 56549 3924 56591
rect 3980 56549 4048 56591
rect 4104 56549 4172 56591
rect 4228 56549 4296 56605
rect 4352 56549 4420 56605
rect 4476 56549 4544 56605
rect 4600 56549 4668 56605
rect 4724 56549 4791 56605
rect 2741 56519 4791 56549
rect 2741 56481 3903 56519
rect 3955 56481 4027 56519
rect 4079 56481 4151 56519
rect 4203 56481 4791 56519
rect 2741 56425 2808 56481
rect 2864 56425 2932 56481
rect 2988 56425 3056 56481
rect 3112 56425 3180 56481
rect 3236 56425 3304 56481
rect 3360 56425 3428 56481
rect 3484 56425 3552 56481
rect 3608 56425 3676 56481
rect 3732 56425 3800 56481
rect 3856 56467 3903 56481
rect 3980 56467 4027 56481
rect 4104 56467 4151 56481
rect 3856 56425 3924 56467
rect 3980 56425 4048 56467
rect 4104 56425 4172 56467
rect 4228 56425 4296 56481
rect 4352 56425 4420 56481
rect 4476 56425 4544 56481
rect 4600 56425 4668 56481
rect 4724 56425 4791 56481
rect 2741 56395 4791 56425
rect 2741 56357 3903 56395
rect 3955 56357 4027 56395
rect 4079 56357 4151 56395
rect 4203 56357 4791 56395
rect 2741 56301 2808 56357
rect 2864 56301 2932 56357
rect 2988 56301 3056 56357
rect 3112 56301 3180 56357
rect 3236 56301 3304 56357
rect 3360 56301 3428 56357
rect 3484 56301 3552 56357
rect 3608 56301 3676 56357
rect 3732 56301 3800 56357
rect 3856 56343 3903 56357
rect 3980 56343 4027 56357
rect 4104 56343 4151 56357
rect 3856 56301 3924 56343
rect 3980 56301 4048 56343
rect 4104 56301 4172 56343
rect 4228 56301 4296 56357
rect 4352 56301 4420 56357
rect 4476 56301 4544 56357
rect 4600 56301 4668 56357
rect 4724 56301 4791 56357
rect 2741 56271 4791 56301
rect 2741 56233 3903 56271
rect 3955 56233 4027 56271
rect 4079 56233 4151 56271
rect 4203 56233 4791 56271
rect 2741 56177 2808 56233
rect 2864 56177 2932 56233
rect 2988 56177 3056 56233
rect 3112 56177 3180 56233
rect 3236 56177 3304 56233
rect 3360 56177 3428 56233
rect 3484 56177 3552 56233
rect 3608 56177 3676 56233
rect 3732 56177 3800 56233
rect 3856 56219 3903 56233
rect 3980 56219 4027 56233
rect 4104 56219 4151 56233
rect 3856 56177 3924 56219
rect 3980 56177 4048 56219
rect 4104 56177 4172 56219
rect 4228 56177 4296 56233
rect 4352 56177 4420 56233
rect 4476 56177 4544 56233
rect 4600 56177 4668 56233
rect 4724 56177 4791 56233
rect 2741 56147 4791 56177
rect 2741 56109 3903 56147
rect 3955 56109 4027 56147
rect 4079 56109 4151 56147
rect 4203 56109 4791 56147
rect 2741 56053 2808 56109
rect 2864 56053 2932 56109
rect 2988 56053 3056 56109
rect 3112 56053 3180 56109
rect 3236 56053 3304 56109
rect 3360 56053 3428 56109
rect 3484 56053 3552 56109
rect 3608 56053 3676 56109
rect 3732 56053 3800 56109
rect 3856 56095 3903 56109
rect 3980 56095 4027 56109
rect 4104 56095 4151 56109
rect 3856 56053 3924 56095
rect 3980 56053 4048 56095
rect 4104 56053 4172 56095
rect 4228 56053 4296 56109
rect 4352 56053 4420 56109
rect 4476 56053 4544 56109
rect 4600 56053 4668 56109
rect 4724 56053 4791 56109
rect 2741 56023 4791 56053
rect 2741 55971 3903 56023
rect 3955 55971 4027 56023
rect 4079 55971 4151 56023
rect 4203 55971 4791 56023
rect 2741 55899 4791 55971
rect 2741 55847 3903 55899
rect 3955 55847 4027 55899
rect 4079 55847 4151 55899
rect 4203 55847 4791 55899
rect 2741 55775 4791 55847
rect 2741 55723 3903 55775
rect 3955 55723 4027 55775
rect 4079 55723 4151 55775
rect 4203 55723 4791 55775
rect 2741 55651 4791 55723
rect 2741 55599 3903 55651
rect 3955 55599 4027 55651
rect 4079 55599 4151 55651
rect 4203 55599 4791 55651
rect 2741 55527 4791 55599
rect 2741 55475 3903 55527
rect 3955 55475 4027 55527
rect 4079 55475 4151 55527
rect 4203 55475 4791 55527
rect 2741 55403 4791 55475
rect 2741 55351 3903 55403
rect 3955 55351 4027 55403
rect 4079 55351 4151 55403
rect 4203 55351 4791 55403
rect 2741 55279 4791 55351
rect 2741 55227 3903 55279
rect 3955 55227 4027 55279
rect 4079 55227 4151 55279
rect 4203 55227 4791 55279
rect 2741 55155 4791 55227
rect 2741 55103 3903 55155
rect 3955 55103 4027 55155
rect 4079 55103 4151 55155
rect 4203 55103 4791 55155
rect 2741 55031 4791 55103
rect 2741 54979 3903 55031
rect 3955 54979 4027 55031
rect 4079 54979 4151 55031
rect 4203 54979 4791 55031
rect 2741 54907 4791 54979
rect 2741 54855 3903 54907
rect 3955 54855 4027 54907
rect 4079 54855 4151 54907
rect 4203 54855 4791 54907
rect 2741 54783 4791 54855
rect 2741 54731 3903 54783
rect 3955 54731 4027 54783
rect 4079 54731 4151 54783
rect 4203 54731 4791 54783
rect 2741 54659 4791 54731
rect 2741 54607 3903 54659
rect 3955 54607 4027 54659
rect 4079 54607 4151 54659
rect 4203 54607 4791 54659
rect 2741 54535 4791 54607
rect 2741 54483 3903 54535
rect 3955 54483 4027 54535
rect 4079 54483 4151 54535
rect 4203 54483 4791 54535
rect 2741 54411 4791 54483
rect 2741 54359 3903 54411
rect 3955 54359 4027 54411
rect 4079 54359 4151 54411
rect 4203 54359 4791 54411
rect 2741 54287 4791 54359
rect 2741 54235 3903 54287
rect 3955 54235 4027 54287
rect 4079 54235 4151 54287
rect 4203 54235 4791 54287
rect 2741 54163 4791 54235
rect 2741 54148 3903 54163
rect 3955 54148 4027 54163
rect 4079 54148 4151 54163
rect 4203 54148 4791 54163
rect 2741 54092 2808 54148
rect 2864 54092 2932 54148
rect 2988 54092 3056 54148
rect 3112 54092 3180 54148
rect 3236 54092 3304 54148
rect 3360 54092 3428 54148
rect 3484 54092 3552 54148
rect 3608 54092 3676 54148
rect 3732 54092 3800 54148
rect 3856 54111 3903 54148
rect 3980 54111 4027 54148
rect 4104 54111 4151 54148
rect 3856 54092 3924 54111
rect 3980 54092 4048 54111
rect 4104 54092 4172 54111
rect 4228 54092 4296 54148
rect 4352 54092 4420 54148
rect 4476 54092 4544 54148
rect 4600 54092 4668 54148
rect 4724 54092 4791 54148
rect 2741 54039 4791 54092
rect 2741 54024 3903 54039
rect 3955 54024 4027 54039
rect 4079 54024 4151 54039
rect 4203 54024 4791 54039
rect 2741 53968 2808 54024
rect 2864 53968 2932 54024
rect 2988 53968 3056 54024
rect 3112 53968 3180 54024
rect 3236 53968 3304 54024
rect 3360 53968 3428 54024
rect 3484 53968 3552 54024
rect 3608 53968 3676 54024
rect 3732 53968 3800 54024
rect 3856 53987 3903 54024
rect 3980 53987 4027 54024
rect 4104 53987 4151 54024
rect 3856 53968 3924 53987
rect 3980 53968 4048 53987
rect 4104 53968 4172 53987
rect 4228 53968 4296 54024
rect 4352 53968 4420 54024
rect 4476 53968 4544 54024
rect 4600 53968 4668 54024
rect 4724 53968 4791 54024
rect 2741 53915 4791 53968
rect 2741 53900 3903 53915
rect 3955 53900 4027 53915
rect 4079 53900 4151 53915
rect 4203 53900 4791 53915
rect 2741 53844 2808 53900
rect 2864 53844 2932 53900
rect 2988 53844 3056 53900
rect 3112 53844 3180 53900
rect 3236 53844 3304 53900
rect 3360 53844 3428 53900
rect 3484 53844 3552 53900
rect 3608 53844 3676 53900
rect 3732 53844 3800 53900
rect 3856 53863 3903 53900
rect 3980 53863 4027 53900
rect 4104 53863 4151 53900
rect 3856 53844 3924 53863
rect 3980 53844 4048 53863
rect 4104 53844 4172 53863
rect 4228 53844 4296 53900
rect 4352 53844 4420 53900
rect 4476 53844 4544 53900
rect 4600 53844 4668 53900
rect 4724 53844 4791 53900
rect 2741 53791 4791 53844
rect 2741 53776 3903 53791
rect 3955 53776 4027 53791
rect 4079 53776 4151 53791
rect 4203 53776 4791 53791
rect 2741 53720 2808 53776
rect 2864 53720 2932 53776
rect 2988 53720 3056 53776
rect 3112 53720 3180 53776
rect 3236 53720 3304 53776
rect 3360 53720 3428 53776
rect 3484 53720 3552 53776
rect 3608 53720 3676 53776
rect 3732 53720 3800 53776
rect 3856 53739 3903 53776
rect 3980 53739 4027 53776
rect 4104 53739 4151 53776
rect 3856 53720 3924 53739
rect 3980 53720 4048 53739
rect 4104 53720 4172 53739
rect 4228 53720 4296 53776
rect 4352 53720 4420 53776
rect 4476 53720 4544 53776
rect 4600 53720 4668 53776
rect 4724 53720 4791 53776
rect 2741 53667 4791 53720
rect 2741 53652 3903 53667
rect 3955 53652 4027 53667
rect 4079 53652 4151 53667
rect 4203 53652 4791 53667
rect 2741 53596 2808 53652
rect 2864 53596 2932 53652
rect 2988 53596 3056 53652
rect 3112 53596 3180 53652
rect 3236 53596 3304 53652
rect 3360 53596 3428 53652
rect 3484 53596 3552 53652
rect 3608 53596 3676 53652
rect 3732 53596 3800 53652
rect 3856 53615 3903 53652
rect 3980 53615 4027 53652
rect 4104 53615 4151 53652
rect 3856 53596 3924 53615
rect 3980 53596 4048 53615
rect 4104 53596 4172 53615
rect 4228 53596 4296 53652
rect 4352 53596 4420 53652
rect 4476 53596 4544 53652
rect 4600 53596 4668 53652
rect 4724 53596 4791 53652
rect 2741 53543 4791 53596
rect 2741 53528 3903 53543
rect 3955 53528 4027 53543
rect 4079 53528 4151 53543
rect 4203 53528 4791 53543
rect 2741 53483 2808 53528
rect 2864 53483 2932 53528
rect 2988 53483 3056 53528
rect 3112 53483 3180 53528
rect 3236 53483 3304 53528
rect 3360 53483 3428 53528
rect 3484 53483 3552 53528
rect 3608 53483 3676 53528
rect 3732 53483 3800 53528
rect 2741 53431 2763 53483
rect 2864 53472 2871 53483
rect 2815 53431 2871 53472
rect 2923 53472 2932 53483
rect 3031 53472 3056 53483
rect 3139 53472 3180 53483
rect 2923 53431 2979 53472
rect 3031 53431 3087 53472
rect 3139 53431 3195 53472
rect 3247 53431 3303 53483
rect 3360 53472 3411 53483
rect 3484 53472 3519 53483
rect 3608 53472 3627 53483
rect 3732 53472 3735 53483
rect 3355 53431 3411 53472
rect 3463 53431 3519 53472
rect 3571 53431 3627 53472
rect 3679 53431 3735 53472
rect 3787 53472 3800 53483
rect 3856 53491 3903 53528
rect 3980 53491 4027 53528
rect 4104 53491 4151 53528
rect 3856 53472 3924 53491
rect 3980 53472 4048 53491
rect 4104 53472 4172 53491
rect 4228 53472 4296 53528
rect 4352 53472 4420 53528
rect 4476 53472 4544 53528
rect 4600 53472 4668 53528
rect 4724 53472 4791 53528
rect 3787 53431 4791 53472
rect 2741 53419 4791 53431
rect 2741 53404 3903 53419
rect 3955 53404 4027 53419
rect 4079 53404 4151 53419
rect 4203 53404 4791 53419
rect 2741 53375 2808 53404
rect 2864 53375 2932 53404
rect 2988 53375 3056 53404
rect 3112 53375 3180 53404
rect 3236 53375 3304 53404
rect 3360 53375 3428 53404
rect 3484 53375 3552 53404
rect 3608 53375 3676 53404
rect 3732 53375 3800 53404
rect 2741 53323 2763 53375
rect 2864 53348 2871 53375
rect 2815 53323 2871 53348
rect 2923 53348 2932 53375
rect 3031 53348 3056 53375
rect 3139 53348 3180 53375
rect 2923 53323 2979 53348
rect 3031 53323 3087 53348
rect 3139 53323 3195 53348
rect 3247 53323 3303 53375
rect 3360 53348 3411 53375
rect 3484 53348 3519 53375
rect 3608 53348 3627 53375
rect 3732 53348 3735 53375
rect 3355 53323 3411 53348
rect 3463 53323 3519 53348
rect 3571 53323 3627 53348
rect 3679 53323 3735 53348
rect 3787 53348 3800 53375
rect 3856 53367 3903 53404
rect 3980 53367 4027 53404
rect 4104 53367 4151 53404
rect 3856 53348 3924 53367
rect 3980 53348 4048 53367
rect 4104 53348 4172 53367
rect 4228 53348 4296 53404
rect 4352 53348 4420 53404
rect 4476 53348 4544 53404
rect 4600 53348 4668 53404
rect 4724 53348 4791 53404
rect 3787 53323 4791 53348
rect 2741 53295 4791 53323
rect 2741 53280 3903 53295
rect 3955 53280 4027 53295
rect 4079 53280 4151 53295
rect 4203 53280 4791 53295
rect 2741 53267 2808 53280
rect 2864 53267 2932 53280
rect 2988 53267 3056 53280
rect 3112 53267 3180 53280
rect 3236 53267 3304 53280
rect 3360 53267 3428 53280
rect 3484 53267 3552 53280
rect 3608 53267 3676 53280
rect 3732 53267 3800 53280
rect 2741 53215 2763 53267
rect 2864 53224 2871 53267
rect 2815 53215 2871 53224
rect 2923 53224 2932 53267
rect 3031 53224 3056 53267
rect 3139 53224 3180 53267
rect 2923 53215 2979 53224
rect 3031 53215 3087 53224
rect 3139 53215 3195 53224
rect 3247 53215 3303 53267
rect 3360 53224 3411 53267
rect 3484 53224 3519 53267
rect 3608 53224 3627 53267
rect 3732 53224 3735 53267
rect 3355 53215 3411 53224
rect 3463 53215 3519 53224
rect 3571 53215 3627 53224
rect 3679 53215 3735 53224
rect 3787 53224 3800 53267
rect 3856 53243 3903 53280
rect 3980 53243 4027 53280
rect 4104 53243 4151 53280
rect 3856 53224 3924 53243
rect 3980 53224 4048 53243
rect 4104 53224 4172 53243
rect 4228 53224 4296 53280
rect 4352 53224 4420 53280
rect 4476 53224 4544 53280
rect 4600 53224 4668 53280
rect 4724 53224 4791 53280
rect 3787 53215 4791 53224
rect 2741 53156 4791 53215
rect 2741 53100 2808 53156
rect 2864 53100 2932 53156
rect 2988 53100 3056 53156
rect 3112 53100 3180 53156
rect 3236 53100 3304 53156
rect 3360 53100 3428 53156
rect 3484 53100 3552 53156
rect 3608 53100 3676 53156
rect 3732 53100 3800 53156
rect 3856 53100 3924 53156
rect 3980 53100 4048 53156
rect 4104 53100 4172 53156
rect 4228 53100 4296 53156
rect 4352 53100 4420 53156
rect 4476 53100 4544 53156
rect 4600 53100 4668 53156
rect 4724 53100 4791 53156
rect 2741 53032 4791 53100
rect 2741 52976 2808 53032
rect 2864 52976 2932 53032
rect 2988 52976 3056 53032
rect 3112 52976 3180 53032
rect 3236 52976 3304 53032
rect 3360 52976 3428 53032
rect 3484 52976 3552 53032
rect 3608 52976 3676 53032
rect 3732 52976 3800 53032
rect 3856 52976 3924 53032
rect 3980 52976 4048 53032
rect 4104 52976 4172 53032
rect 4228 52976 4296 53032
rect 4352 52976 4420 53032
rect 4476 52976 4544 53032
rect 4600 52976 4668 53032
rect 4724 52976 4791 53032
rect 2741 52908 4791 52976
rect 2741 52852 2808 52908
rect 2864 52852 2932 52908
rect 2988 52852 3056 52908
rect 3112 52852 3180 52908
rect 3236 52852 3304 52908
rect 3360 52852 3428 52908
rect 3484 52852 3552 52908
rect 3608 52852 3676 52908
rect 3732 52852 3800 52908
rect 3856 52852 3924 52908
rect 3980 52852 4048 52908
rect 4104 52852 4172 52908
rect 4228 52852 4296 52908
rect 4352 52852 4420 52908
rect 4476 52852 4544 52908
rect 4600 52852 4668 52908
rect 4724 52852 4791 52908
rect 2741 52548 4791 52852
rect 2741 52492 2808 52548
rect 2864 52492 2932 52548
rect 2988 52492 3056 52548
rect 3112 52492 3180 52548
rect 3236 52492 3304 52548
rect 3360 52492 3428 52548
rect 3484 52492 3552 52548
rect 3608 52492 3676 52548
rect 3732 52492 3800 52548
rect 3856 52492 3924 52548
rect 3980 52492 4048 52548
rect 4104 52492 4172 52548
rect 4228 52492 4296 52548
rect 4352 52492 4420 52548
rect 4476 52492 4544 52548
rect 4600 52492 4668 52548
rect 4724 52492 4791 52548
rect 2741 52424 4791 52492
rect 2741 52368 2808 52424
rect 2864 52368 2932 52424
rect 2988 52368 3056 52424
rect 3112 52368 3180 52424
rect 3236 52368 3304 52424
rect 3360 52368 3428 52424
rect 3484 52368 3552 52424
rect 3608 52368 3676 52424
rect 3732 52368 3800 52424
rect 3856 52368 3924 52424
rect 3980 52368 4048 52424
rect 4104 52368 4172 52424
rect 4228 52368 4296 52424
rect 4352 52368 4420 52424
rect 4476 52368 4544 52424
rect 4600 52368 4668 52424
rect 4724 52368 4791 52424
rect 2741 52300 4791 52368
rect 2741 52244 2808 52300
rect 2864 52244 2932 52300
rect 2988 52244 3056 52300
rect 3112 52244 3180 52300
rect 3236 52244 3304 52300
rect 3360 52244 3428 52300
rect 3484 52244 3552 52300
rect 3608 52244 3676 52300
rect 3732 52244 3800 52300
rect 3856 52244 3924 52300
rect 3980 52244 4048 52300
rect 4104 52244 4172 52300
rect 4228 52244 4296 52300
rect 4352 52244 4420 52300
rect 4476 52244 4544 52300
rect 4600 52244 4668 52300
rect 4724 52244 4791 52300
rect 2741 52176 4791 52244
rect 2741 52120 2808 52176
rect 2864 52120 2932 52176
rect 2988 52120 3056 52176
rect 3112 52120 3180 52176
rect 3236 52120 3304 52176
rect 3360 52120 3428 52176
rect 3484 52120 3552 52176
rect 3608 52120 3676 52176
rect 3732 52120 3800 52176
rect 3856 52120 3924 52176
rect 3980 52120 4048 52176
rect 4104 52120 4172 52176
rect 4228 52120 4296 52176
rect 4352 52120 4420 52176
rect 4476 52120 4544 52176
rect 4600 52120 4668 52176
rect 4724 52120 4791 52176
rect 2741 52052 4791 52120
rect 2741 51996 2808 52052
rect 2864 51996 2932 52052
rect 2988 51996 3056 52052
rect 3112 52009 3180 52052
rect 3236 52009 3304 52052
rect 3360 52009 3428 52052
rect 3484 52009 3552 52052
rect 3608 52009 3676 52052
rect 3732 52009 3800 52052
rect 3856 52009 3924 52052
rect 3980 52009 4048 52052
rect 4104 52009 4172 52052
rect 4228 52009 4296 52052
rect 4352 52009 4420 52052
rect 4476 52009 4544 52052
rect 4600 52009 4668 52052
rect 4724 52009 4791 52052
rect 3112 51996 3161 52009
rect 3236 51996 3269 52009
rect 3360 51996 3377 52009
rect 3484 51996 3485 52009
rect 2741 51957 3161 51996
rect 3213 51957 3269 51996
rect 3321 51957 3377 51996
rect 3429 51957 3485 51996
rect 3537 51996 3552 52009
rect 3645 51996 3676 52009
rect 3753 51996 3800 52009
rect 3537 51957 3593 51996
rect 3645 51957 3701 51996
rect 3753 51957 3809 51996
rect 3861 51957 3917 52009
rect 3980 51996 4025 52009
rect 4104 51996 4133 52009
rect 4228 51996 4241 52009
rect 3969 51957 4025 51996
rect 4077 51957 4133 51996
rect 4185 51957 4241 51996
rect 4293 51996 4296 52009
rect 4401 51996 4420 52009
rect 4509 51996 4544 52009
rect 4617 51996 4668 52009
rect 4293 51957 4349 51996
rect 4401 51957 4457 51996
rect 4509 51957 4565 51996
rect 4617 51957 4673 51996
rect 4725 51957 4791 52009
rect 2741 51928 4791 51957
rect 2741 51872 2808 51928
rect 2864 51872 2932 51928
rect 2988 51872 3056 51928
rect 3112 51901 3180 51928
rect 3236 51901 3304 51928
rect 3360 51901 3428 51928
rect 3484 51901 3552 51928
rect 3608 51901 3676 51928
rect 3732 51901 3800 51928
rect 3856 51901 3924 51928
rect 3980 51901 4048 51928
rect 4104 51901 4172 51928
rect 4228 51901 4296 51928
rect 4352 51901 4420 51928
rect 4476 51901 4544 51928
rect 4600 51901 4668 51928
rect 4724 51901 4791 51928
rect 3112 51872 3161 51901
rect 3236 51872 3269 51901
rect 3360 51872 3377 51901
rect 3484 51872 3485 51901
rect 2741 51849 3161 51872
rect 3213 51849 3269 51872
rect 3321 51849 3377 51872
rect 3429 51849 3485 51872
rect 3537 51872 3552 51901
rect 3645 51872 3676 51901
rect 3753 51872 3800 51901
rect 3537 51849 3593 51872
rect 3645 51849 3701 51872
rect 3753 51849 3809 51872
rect 3861 51849 3917 51901
rect 3980 51872 4025 51901
rect 4104 51872 4133 51901
rect 4228 51872 4241 51901
rect 3969 51849 4025 51872
rect 4077 51849 4133 51872
rect 4185 51849 4241 51872
rect 4293 51872 4296 51901
rect 4401 51872 4420 51901
rect 4509 51872 4544 51901
rect 4617 51872 4668 51901
rect 4293 51849 4349 51872
rect 4401 51849 4457 51872
rect 4509 51849 4565 51872
rect 4617 51849 4673 51872
rect 4725 51849 4791 51901
rect 2741 51804 4791 51849
rect 2741 51748 2808 51804
rect 2864 51748 2932 51804
rect 2988 51748 3056 51804
rect 3112 51748 3180 51804
rect 3236 51748 3304 51804
rect 3360 51748 3428 51804
rect 3484 51748 3552 51804
rect 3608 51748 3676 51804
rect 3732 51748 3800 51804
rect 3856 51748 3924 51804
rect 3980 51748 4048 51804
rect 4104 51748 4172 51804
rect 4228 51748 4296 51804
rect 4352 51748 4420 51804
rect 4476 51748 4544 51804
rect 4600 51748 4668 51804
rect 4724 51748 4791 51804
rect 2741 51680 4791 51748
rect 2741 51624 2808 51680
rect 2864 51624 2932 51680
rect 2988 51624 3056 51680
rect 3112 51624 3180 51680
rect 3236 51624 3304 51680
rect 3360 51624 3428 51680
rect 3484 51624 3552 51680
rect 3608 51624 3676 51680
rect 3732 51624 3800 51680
rect 3856 51624 3924 51680
rect 3980 51624 4048 51680
rect 4104 51624 4172 51680
rect 4228 51624 4296 51680
rect 4352 51624 4420 51680
rect 4476 51624 4544 51680
rect 4600 51624 4668 51680
rect 4724 51624 4791 51680
rect 2741 51556 4791 51624
rect 2741 51500 2808 51556
rect 2864 51500 2932 51556
rect 2988 51500 3056 51556
rect 3112 51500 3180 51556
rect 3236 51500 3304 51556
rect 3360 51500 3428 51556
rect 3484 51500 3552 51556
rect 3608 51500 3676 51556
rect 3732 51500 3800 51556
rect 3856 51500 3924 51556
rect 3980 51500 4048 51556
rect 4104 51500 4172 51556
rect 4228 51500 4296 51556
rect 4352 51500 4420 51556
rect 4476 51500 4544 51556
rect 4600 51500 4668 51556
rect 4724 51500 4791 51556
rect 2741 51432 4791 51500
rect 2741 51376 2808 51432
rect 2864 51376 2932 51432
rect 2988 51376 3056 51432
rect 3112 51376 3180 51432
rect 3236 51376 3304 51432
rect 3360 51376 3428 51432
rect 3484 51376 3552 51432
rect 3608 51376 3676 51432
rect 3732 51376 3800 51432
rect 3856 51376 3924 51432
rect 3980 51376 4048 51432
rect 4104 51376 4172 51432
rect 4228 51376 4296 51432
rect 4352 51376 4420 51432
rect 4476 51376 4544 51432
rect 4600 51376 4668 51432
rect 4724 51376 4791 51432
rect 2741 51308 4791 51376
rect 2741 51252 2808 51308
rect 2864 51252 2932 51308
rect 2988 51252 3056 51308
rect 3112 51252 3180 51308
rect 3236 51252 3304 51308
rect 3360 51252 3428 51308
rect 3484 51252 3552 51308
rect 3608 51252 3676 51308
rect 3732 51252 3800 51308
rect 3856 51252 3924 51308
rect 3980 51252 4048 51308
rect 4104 51252 4172 51308
rect 4228 51252 4296 51308
rect 4352 51252 4420 51308
rect 4476 51252 4544 51308
rect 4600 51252 4668 51308
rect 4724 51252 4791 51308
rect 2741 51206 4791 51252
rect 2741 51154 3161 51206
rect 3213 51154 3269 51206
rect 3321 51154 3377 51206
rect 3429 51154 3485 51206
rect 3537 51154 3593 51206
rect 3645 51154 3701 51206
rect 3753 51154 3809 51206
rect 3861 51154 3917 51206
rect 3969 51154 4025 51206
rect 4077 51154 4133 51206
rect 4185 51154 4241 51206
rect 4293 51154 4349 51206
rect 4401 51154 4457 51206
rect 4509 51154 4565 51206
rect 4617 51154 4673 51206
rect 4725 51154 4791 51206
rect 2741 51098 4791 51154
rect 2741 51046 3161 51098
rect 3213 51046 3269 51098
rect 3321 51046 3377 51098
rect 3429 51046 3485 51098
rect 3537 51046 3593 51098
rect 3645 51046 3701 51098
rect 3753 51046 3809 51098
rect 3861 51046 3917 51098
rect 3969 51046 4025 51098
rect 4077 51046 4133 51098
rect 4185 51046 4241 51098
rect 4293 51046 4349 51098
rect 4401 51046 4457 51098
rect 4509 51046 4565 51098
rect 4617 51046 4673 51098
rect 4725 51046 4791 51098
rect 2741 50990 4791 51046
rect 2741 50938 3161 50990
rect 3213 50938 3269 50990
rect 3321 50938 3377 50990
rect 3429 50938 3485 50990
rect 3537 50938 3593 50990
rect 3645 50938 3701 50990
rect 3753 50938 3809 50990
rect 3861 50938 3917 50990
rect 3969 50938 4025 50990
rect 4077 50938 4133 50990
rect 4185 50938 4241 50990
rect 4293 50938 4349 50990
rect 4401 50938 4457 50990
rect 4509 50938 4565 50990
rect 4617 50938 4673 50990
rect 4725 50938 4791 50990
rect 2741 50272 4791 50938
rect 2741 50220 3161 50272
rect 3213 50220 3269 50272
rect 3321 50220 3377 50272
rect 3429 50220 3485 50272
rect 3537 50220 3593 50272
rect 3645 50220 3701 50272
rect 3753 50220 3809 50272
rect 3861 50220 3917 50272
rect 3969 50220 4025 50272
rect 4077 50220 4133 50272
rect 4185 50220 4241 50272
rect 4293 50220 4349 50272
rect 4401 50220 4457 50272
rect 4509 50220 4565 50272
rect 4617 50220 4673 50272
rect 4725 50220 4791 50272
rect 2741 50164 4791 50220
rect 2741 50112 3161 50164
rect 3213 50112 3269 50164
rect 3321 50112 3377 50164
rect 3429 50112 3485 50164
rect 3537 50112 3593 50164
rect 3645 50112 3701 50164
rect 3753 50112 3809 50164
rect 3861 50112 3917 50164
rect 3969 50112 4025 50164
rect 4077 50112 4133 50164
rect 4185 50112 4241 50164
rect 4293 50112 4349 50164
rect 4401 50112 4457 50164
rect 4509 50112 4565 50164
rect 4617 50112 4673 50164
rect 4725 50112 4791 50164
rect 2741 50056 4791 50112
rect 2741 50004 3161 50056
rect 3213 50004 3269 50056
rect 3321 50004 3377 50056
rect 3429 50004 3485 50056
rect 3537 50004 3593 50056
rect 3645 50004 3701 50056
rect 3753 50004 3809 50056
rect 3861 50004 3917 50056
rect 3969 50004 4025 50056
rect 4077 50004 4133 50056
rect 4185 50004 4241 50056
rect 4293 50004 4349 50056
rect 4401 50004 4457 50056
rect 4509 50004 4565 50056
rect 4617 50004 4673 50056
rect 4725 50004 4791 50056
rect 2741 49348 4791 50004
rect 2741 49292 2808 49348
rect 2864 49292 2932 49348
rect 2988 49292 3056 49348
rect 3112 49338 3180 49348
rect 3236 49338 3304 49348
rect 3360 49338 3428 49348
rect 3484 49338 3552 49348
rect 3608 49338 3676 49348
rect 3732 49338 3800 49348
rect 3856 49338 3924 49348
rect 3980 49338 4048 49348
rect 4104 49338 4172 49348
rect 4228 49338 4296 49348
rect 4352 49338 4420 49348
rect 4476 49338 4544 49348
rect 4600 49338 4668 49348
rect 4724 49338 4791 49348
rect 3112 49292 3161 49338
rect 3236 49292 3269 49338
rect 3360 49292 3377 49338
rect 3484 49292 3485 49338
rect 2741 49286 3161 49292
rect 3213 49286 3269 49292
rect 3321 49286 3377 49292
rect 3429 49286 3485 49292
rect 3537 49292 3552 49338
rect 3645 49292 3676 49338
rect 3753 49292 3800 49338
rect 3537 49286 3593 49292
rect 3645 49286 3701 49292
rect 3753 49286 3809 49292
rect 3861 49286 3917 49338
rect 3980 49292 4025 49338
rect 4104 49292 4133 49338
rect 4228 49292 4241 49338
rect 3969 49286 4025 49292
rect 4077 49286 4133 49292
rect 4185 49286 4241 49292
rect 4293 49292 4296 49338
rect 4401 49292 4420 49338
rect 4509 49292 4544 49338
rect 4617 49292 4668 49338
rect 4293 49286 4349 49292
rect 4401 49286 4457 49292
rect 4509 49286 4565 49292
rect 4617 49286 4673 49292
rect 4725 49286 4791 49338
rect 2741 49230 4791 49286
rect 2741 49224 3161 49230
rect 3213 49224 3269 49230
rect 3321 49224 3377 49230
rect 3429 49224 3485 49230
rect 2741 49168 2808 49224
rect 2864 49168 2932 49224
rect 2988 49168 3056 49224
rect 3112 49178 3161 49224
rect 3236 49178 3269 49224
rect 3360 49178 3377 49224
rect 3484 49178 3485 49224
rect 3537 49224 3593 49230
rect 3645 49224 3701 49230
rect 3753 49224 3809 49230
rect 3537 49178 3552 49224
rect 3645 49178 3676 49224
rect 3753 49178 3800 49224
rect 3861 49178 3917 49230
rect 3969 49224 4025 49230
rect 4077 49224 4133 49230
rect 4185 49224 4241 49230
rect 3980 49178 4025 49224
rect 4104 49178 4133 49224
rect 4228 49178 4241 49224
rect 4293 49224 4349 49230
rect 4401 49224 4457 49230
rect 4509 49224 4565 49230
rect 4617 49224 4673 49230
rect 4293 49178 4296 49224
rect 4401 49178 4420 49224
rect 4509 49178 4544 49224
rect 4617 49178 4668 49224
rect 4725 49178 4791 49230
rect 3112 49168 3180 49178
rect 3236 49168 3304 49178
rect 3360 49168 3428 49178
rect 3484 49168 3552 49178
rect 3608 49168 3676 49178
rect 3732 49168 3800 49178
rect 3856 49168 3924 49178
rect 3980 49168 4048 49178
rect 4104 49168 4172 49178
rect 4228 49168 4296 49178
rect 4352 49168 4420 49178
rect 4476 49168 4544 49178
rect 4600 49168 4668 49178
rect 4724 49168 4791 49178
rect 2741 49122 4791 49168
rect 2741 49100 3161 49122
rect 3213 49100 3269 49122
rect 3321 49100 3377 49122
rect 3429 49100 3485 49122
rect 2741 49044 2808 49100
rect 2864 49044 2932 49100
rect 2988 49044 3056 49100
rect 3112 49070 3161 49100
rect 3236 49070 3269 49100
rect 3360 49070 3377 49100
rect 3484 49070 3485 49100
rect 3537 49100 3593 49122
rect 3645 49100 3701 49122
rect 3753 49100 3809 49122
rect 3537 49070 3552 49100
rect 3645 49070 3676 49100
rect 3753 49070 3800 49100
rect 3861 49070 3917 49122
rect 3969 49100 4025 49122
rect 4077 49100 4133 49122
rect 4185 49100 4241 49122
rect 3980 49070 4025 49100
rect 4104 49070 4133 49100
rect 4228 49070 4241 49100
rect 4293 49100 4349 49122
rect 4401 49100 4457 49122
rect 4509 49100 4565 49122
rect 4617 49100 4673 49122
rect 4293 49070 4296 49100
rect 4401 49070 4420 49100
rect 4509 49070 4544 49100
rect 4617 49070 4668 49100
rect 4725 49070 4791 49122
rect 3112 49044 3180 49070
rect 3236 49044 3304 49070
rect 3360 49044 3428 49070
rect 3484 49044 3552 49070
rect 3608 49044 3676 49070
rect 3732 49044 3800 49070
rect 3856 49044 3924 49070
rect 3980 49044 4048 49070
rect 4104 49044 4172 49070
rect 4228 49044 4296 49070
rect 4352 49044 4420 49070
rect 4476 49044 4544 49070
rect 4600 49044 4668 49070
rect 4724 49044 4791 49070
rect 2741 48976 4791 49044
rect 2741 48920 2808 48976
rect 2864 48920 2932 48976
rect 2988 48920 3056 48976
rect 3112 48920 3180 48976
rect 3236 48920 3304 48976
rect 3360 48920 3428 48976
rect 3484 48920 3552 48976
rect 3608 48920 3676 48976
rect 3732 48920 3800 48976
rect 3856 48920 3924 48976
rect 3980 48920 4048 48976
rect 4104 48920 4172 48976
rect 4228 48920 4296 48976
rect 4352 48920 4420 48976
rect 4476 48920 4544 48976
rect 4600 48920 4668 48976
rect 4724 48920 4791 48976
rect 2741 48852 4791 48920
rect 2741 48796 2808 48852
rect 2864 48796 2932 48852
rect 2988 48796 3056 48852
rect 3112 48796 3180 48852
rect 3236 48796 3304 48852
rect 3360 48796 3428 48852
rect 3484 48796 3552 48852
rect 3608 48796 3676 48852
rect 3732 48796 3800 48852
rect 3856 48796 3924 48852
rect 3980 48796 4048 48852
rect 4104 48796 4172 48852
rect 4228 48796 4296 48852
rect 4352 48796 4420 48852
rect 4476 48796 4544 48852
rect 4600 48796 4668 48852
rect 4724 48796 4791 48852
rect 2741 48728 4791 48796
rect 2741 48672 2808 48728
rect 2864 48672 2932 48728
rect 2988 48672 3056 48728
rect 3112 48672 3180 48728
rect 3236 48672 3304 48728
rect 3360 48672 3428 48728
rect 3484 48672 3552 48728
rect 3608 48672 3676 48728
rect 3732 48672 3800 48728
rect 3856 48672 3924 48728
rect 3980 48672 4048 48728
rect 4104 48672 4172 48728
rect 4228 48672 4296 48728
rect 4352 48672 4420 48728
rect 4476 48672 4544 48728
rect 4600 48672 4668 48728
rect 4724 48672 4791 48728
rect 2741 48604 4791 48672
rect 2741 48548 2808 48604
rect 2864 48548 2932 48604
rect 2988 48548 3056 48604
rect 3112 48548 3180 48604
rect 3236 48548 3304 48604
rect 3360 48548 3428 48604
rect 3484 48548 3552 48604
rect 3608 48548 3676 48604
rect 3732 48548 3800 48604
rect 3856 48548 3924 48604
rect 3980 48548 4048 48604
rect 4104 48548 4172 48604
rect 4228 48548 4296 48604
rect 4352 48548 4420 48604
rect 4476 48548 4544 48604
rect 4600 48548 4668 48604
rect 4724 48548 4791 48604
rect 2741 48480 4791 48548
rect 2741 48424 2808 48480
rect 2864 48424 2932 48480
rect 2988 48424 3056 48480
rect 3112 48427 3180 48480
rect 3236 48427 3304 48480
rect 3360 48427 3428 48480
rect 3484 48427 3552 48480
rect 3608 48427 3676 48480
rect 3732 48427 3800 48480
rect 3856 48427 3924 48480
rect 3980 48427 4048 48480
rect 4104 48427 4172 48480
rect 4228 48427 4296 48480
rect 4352 48427 4420 48480
rect 4476 48427 4544 48480
rect 4600 48427 4668 48480
rect 4724 48427 4791 48480
rect 3112 48424 3161 48427
rect 3236 48424 3269 48427
rect 3360 48424 3377 48427
rect 3484 48424 3485 48427
rect 2741 48375 3161 48424
rect 3213 48375 3269 48424
rect 3321 48375 3377 48424
rect 3429 48375 3485 48424
rect 3537 48424 3552 48427
rect 3645 48424 3676 48427
rect 3753 48424 3800 48427
rect 3537 48375 3593 48424
rect 3645 48375 3701 48424
rect 3753 48375 3809 48424
rect 3861 48375 3917 48427
rect 3980 48424 4025 48427
rect 4104 48424 4133 48427
rect 4228 48424 4241 48427
rect 3969 48375 4025 48424
rect 4077 48375 4133 48424
rect 4185 48375 4241 48424
rect 4293 48424 4296 48427
rect 4401 48424 4420 48427
rect 4509 48424 4544 48427
rect 4617 48424 4668 48427
rect 4293 48375 4349 48424
rect 4401 48375 4457 48424
rect 4509 48375 4565 48424
rect 4617 48375 4673 48424
rect 4725 48375 4791 48427
rect 2741 48356 4791 48375
rect 2741 48300 2808 48356
rect 2864 48300 2932 48356
rect 2988 48300 3056 48356
rect 3112 48319 3180 48356
rect 3236 48319 3304 48356
rect 3360 48319 3428 48356
rect 3484 48319 3552 48356
rect 3608 48319 3676 48356
rect 3732 48319 3800 48356
rect 3856 48319 3924 48356
rect 3980 48319 4048 48356
rect 4104 48319 4172 48356
rect 4228 48319 4296 48356
rect 4352 48319 4420 48356
rect 4476 48319 4544 48356
rect 4600 48319 4668 48356
rect 4724 48319 4791 48356
rect 3112 48300 3161 48319
rect 3236 48300 3269 48319
rect 3360 48300 3377 48319
rect 3484 48300 3485 48319
rect 2741 48267 3161 48300
rect 3213 48267 3269 48300
rect 3321 48267 3377 48300
rect 3429 48267 3485 48300
rect 3537 48300 3552 48319
rect 3645 48300 3676 48319
rect 3753 48300 3800 48319
rect 3537 48267 3593 48300
rect 3645 48267 3701 48300
rect 3753 48267 3809 48300
rect 3861 48267 3917 48319
rect 3980 48300 4025 48319
rect 4104 48300 4133 48319
rect 4228 48300 4241 48319
rect 3969 48267 4025 48300
rect 4077 48267 4133 48300
rect 4185 48267 4241 48300
rect 4293 48300 4296 48319
rect 4401 48300 4420 48319
rect 4509 48300 4544 48319
rect 4617 48300 4668 48319
rect 4293 48267 4349 48300
rect 4401 48267 4457 48300
rect 4509 48267 4565 48300
rect 4617 48267 4673 48300
rect 4725 48267 4791 48319
rect 2741 48232 4791 48267
rect 2741 48176 2808 48232
rect 2864 48176 2932 48232
rect 2988 48176 3056 48232
rect 3112 48176 3180 48232
rect 3236 48176 3304 48232
rect 3360 48176 3428 48232
rect 3484 48176 3552 48232
rect 3608 48176 3676 48232
rect 3732 48176 3800 48232
rect 3856 48176 3924 48232
rect 3980 48176 4048 48232
rect 4104 48176 4172 48232
rect 4228 48176 4296 48232
rect 4352 48176 4420 48232
rect 4476 48176 4544 48232
rect 4600 48176 4668 48232
rect 4724 48176 4791 48232
rect 2741 48108 4791 48176
rect 2741 48052 2808 48108
rect 2864 48052 2932 48108
rect 2988 48052 3056 48108
rect 3112 48052 3180 48108
rect 3236 48052 3304 48108
rect 3360 48052 3428 48108
rect 3484 48052 3552 48108
rect 3608 48052 3676 48108
rect 3732 48052 3800 48108
rect 3856 48052 3924 48108
rect 3980 48052 4048 48108
rect 4104 48052 4172 48108
rect 4228 48052 4296 48108
rect 4352 48052 4420 48108
rect 4476 48052 4544 48108
rect 4600 48052 4668 48108
rect 4724 48052 4791 48108
rect 2741 47163 4791 48052
rect 4851 56693 5051 57278
rect 4851 56641 4871 56693
rect 4923 56641 4979 56693
rect 5031 56641 5051 56693
rect 4851 56585 5051 56641
rect 4851 56533 4871 56585
rect 4923 56533 4979 56585
rect 5031 56533 5051 56585
rect 4851 56477 5051 56533
rect 4851 56425 4871 56477
rect 4923 56425 4979 56477
rect 5031 56425 5051 56477
rect 4851 56369 5051 56425
rect 4851 56317 4871 56369
rect 4923 56317 4979 56369
rect 5031 56317 5051 56369
rect 4851 56261 5051 56317
rect 4851 56209 4871 56261
rect 4923 56209 4979 56261
rect 5031 56209 5051 56261
rect 4851 56153 5051 56209
rect 4851 56101 4871 56153
rect 4923 56101 4979 56153
rect 5031 56101 5051 56153
rect 4851 56045 5051 56101
rect 4851 55993 4871 56045
rect 4923 55993 4979 56045
rect 5031 55993 5051 56045
rect 4851 55937 5051 55993
rect 4851 55885 4871 55937
rect 4923 55885 4979 55937
rect 5031 55885 5051 55937
rect 4851 55829 5051 55885
rect 4851 55777 4871 55829
rect 4923 55777 4979 55829
rect 5031 55777 5051 55829
rect 4851 55748 5051 55777
rect 4851 55692 4861 55748
rect 4917 55721 4985 55748
rect 4851 55669 4871 55692
rect 4923 55669 4979 55721
rect 5041 55692 5051 55748
rect 5031 55669 5051 55692
rect 4851 55624 5051 55669
rect 4851 55568 4861 55624
rect 4917 55613 4985 55624
rect 4851 55561 4871 55568
rect 4923 55561 4979 55613
rect 5041 55568 5051 55624
rect 5031 55561 5051 55568
rect 4851 55505 5051 55561
rect 4851 55500 4871 55505
rect 4851 55444 4861 55500
rect 4923 55453 4979 55505
rect 5031 55500 5051 55505
rect 4917 55444 4985 55453
rect 5041 55444 5051 55500
rect 4851 55397 5051 55444
rect 4851 55376 4871 55397
rect 4851 55320 4861 55376
rect 4923 55345 4979 55397
rect 5031 55376 5051 55397
rect 4917 55320 4985 55345
rect 5041 55320 5051 55376
rect 4851 55289 5051 55320
rect 4851 55252 4871 55289
rect 4851 55196 4861 55252
rect 4923 55237 4979 55289
rect 5031 55252 5051 55289
rect 4917 55196 4985 55237
rect 5041 55196 5051 55252
rect 4851 55181 5051 55196
rect 4851 55129 4871 55181
rect 4923 55129 4979 55181
rect 5031 55129 5051 55181
rect 4851 55128 5051 55129
rect 4851 55072 4861 55128
rect 4917 55073 4985 55128
rect 4851 55021 4871 55072
rect 4923 55021 4979 55073
rect 5041 55072 5051 55128
rect 5031 55021 5051 55072
rect 4851 55004 5051 55021
rect 4851 54948 4861 55004
rect 4917 54965 4985 55004
rect 4851 54913 4871 54948
rect 4923 54913 4979 54965
rect 5041 54948 5051 55004
rect 5031 54913 5051 54948
rect 4851 54880 5051 54913
rect 4851 54824 4861 54880
rect 4917 54857 4985 54880
rect 4851 54805 4871 54824
rect 4923 54805 4979 54857
rect 5041 54824 5051 54880
rect 5031 54805 5051 54824
rect 4851 54756 5051 54805
rect 4851 54700 4861 54756
rect 4917 54749 4985 54756
rect 4851 54697 4871 54700
rect 4923 54697 4979 54749
rect 5041 54700 5051 54756
rect 5031 54697 5051 54700
rect 4851 54641 5051 54697
rect 4851 54632 4871 54641
rect 4851 54576 4861 54632
rect 4923 54589 4979 54641
rect 5031 54632 5051 54641
rect 4917 54576 4985 54589
rect 5041 54576 5051 54632
rect 4851 54533 5051 54576
rect 4851 54508 4871 54533
rect 4851 54452 4861 54508
rect 4923 54481 4979 54533
rect 5031 54508 5051 54533
rect 4917 54452 4985 54481
rect 5041 54452 5051 54508
rect 4851 54425 5051 54452
rect 4851 54373 4871 54425
rect 4923 54373 4979 54425
rect 5031 54373 5051 54425
rect 4851 54317 5051 54373
rect 4851 54265 4871 54317
rect 4923 54265 4979 54317
rect 5031 54265 5051 54317
rect 4851 54209 5051 54265
rect 4851 54157 4871 54209
rect 4923 54157 4979 54209
rect 5031 54157 5051 54209
rect 4851 54101 5051 54157
rect 4851 54049 4871 54101
rect 4923 54049 4979 54101
rect 5031 54049 5051 54101
rect 4851 53993 5051 54049
rect 4851 53941 4871 53993
rect 4923 53941 4979 53993
rect 5031 53941 5051 53993
rect 4851 53885 5051 53941
rect 4851 53833 4871 53885
rect 4923 53833 4979 53885
rect 5031 53833 5051 53885
rect 4851 53777 5051 53833
rect 4851 53725 4871 53777
rect 4923 53725 4979 53777
rect 5031 53725 5051 53777
rect 4851 53669 5051 53725
rect 4851 53617 4871 53669
rect 4923 53617 4979 53669
rect 5031 53617 5051 53669
rect 4851 52572 5051 53617
rect 4851 52520 4871 52572
rect 4923 52520 4979 52572
rect 5031 52520 5051 52572
rect 4851 52464 5051 52520
rect 4851 52412 4871 52464
rect 4923 52412 4979 52464
rect 5031 52412 5051 52464
rect 4851 52356 5051 52412
rect 4851 52304 4871 52356
rect 4923 52304 4979 52356
rect 5031 52304 5051 52356
rect 4851 51619 5051 52304
rect 4851 51567 4871 51619
rect 4923 51567 4979 51619
rect 5031 51567 5051 51619
rect 4851 51511 5051 51567
rect 4851 51459 4871 51511
rect 4923 51459 4979 51511
rect 5031 51459 5051 51511
rect 4851 50685 5051 51459
rect 4851 50633 4871 50685
rect 4923 50633 4979 50685
rect 5031 50633 5051 50685
rect 4851 50577 5051 50633
rect 4851 50525 4871 50577
rect 4923 50525 4979 50577
rect 5031 50525 5051 50577
rect 4851 49751 5051 50525
rect 4851 49699 4871 49751
rect 4923 49699 4979 49751
rect 5031 49699 5051 49751
rect 4851 49643 5051 49699
rect 4851 49591 4871 49643
rect 4923 49591 4979 49643
rect 5031 49591 5051 49643
rect 4851 48817 5051 49591
rect 4851 48765 4871 48817
rect 4923 48765 4979 48817
rect 5031 48765 5051 48817
rect 4851 48709 5051 48765
rect 4851 48657 4871 48709
rect 4923 48657 4979 48709
rect 5031 48657 5051 48709
rect 4851 47972 5051 48657
rect 4851 47920 4871 47972
rect 4923 47920 4979 47972
rect 5031 47920 5051 47972
rect 4851 47864 5051 47920
rect 4851 47812 4871 47864
rect 4923 47812 4979 47864
rect 5031 47812 5051 47864
rect 4851 47756 5051 47812
rect 4851 47748 4871 47756
rect 4851 47692 4861 47748
rect 4923 47704 4979 47756
rect 5031 47748 5051 47756
rect 4917 47692 4985 47704
rect 5041 47692 5051 47748
rect 4851 47624 5051 47692
rect 4851 47568 4861 47624
rect 4917 47568 4985 47624
rect 5041 47568 5051 47624
rect 4851 47500 5051 47568
rect 4851 47444 4861 47500
rect 4917 47444 4985 47500
rect 5041 47444 5051 47500
rect 4851 47376 5051 47444
rect 4851 47320 4861 47376
rect 4917 47320 4985 47376
rect 5041 47320 5051 47376
rect 4851 47252 5051 47320
rect 4851 47196 4861 47252
rect 4917 47196 4985 47252
rect 5041 47196 5051 47252
rect 2481 47072 2491 47128
rect 2547 47072 2615 47128
rect 2671 47072 2681 47128
rect 2481 47004 2681 47072
rect 2481 46948 2491 47004
rect 2547 46948 2615 47004
rect 2671 46948 2681 47004
rect 2481 46880 2681 46948
rect 2481 46824 2491 46880
rect 2547 46824 2615 46880
rect 2671 46824 2681 46880
rect 2481 46756 2681 46824
rect 2481 46700 2491 46756
rect 2547 46700 2615 46756
rect 2671 46700 2681 46756
rect 2481 46632 2681 46700
rect 2481 46576 2491 46632
rect 2547 46576 2615 46632
rect 2671 46576 2681 46632
rect 2481 46508 2681 46576
rect 2481 46452 2491 46508
rect 2547 46452 2615 46508
rect 2671 46452 2681 46508
rect 2481 46442 2681 46452
rect 4851 47128 5051 47196
rect 5111 57225 7161 57447
rect 7817 57499 9867 57600
rect 7817 57447 7952 57499
rect 8004 57447 8060 57499
rect 8112 57447 8168 57499
rect 8220 57447 8276 57499
rect 8328 57447 8384 57499
rect 8436 57447 8492 57499
rect 8544 57447 8600 57499
rect 8652 57447 8708 57499
rect 8760 57447 8816 57499
rect 8868 57447 8924 57499
rect 8976 57447 9032 57499
rect 9084 57447 9140 57499
rect 9192 57447 9248 57499
rect 9300 57447 9356 57499
rect 9408 57447 9464 57499
rect 9516 57447 9572 57499
rect 9624 57447 9680 57499
rect 9732 57447 9867 57499
rect 5111 57169 5178 57225
rect 5234 57169 5302 57225
rect 5358 57169 5426 57225
rect 5482 57169 5550 57225
rect 5606 57169 5674 57225
rect 5730 57169 5798 57225
rect 5854 57169 5922 57225
rect 5978 57169 6046 57225
rect 6102 57169 6170 57225
rect 6226 57169 6294 57225
rect 6350 57169 6418 57225
rect 6474 57169 6542 57225
rect 6598 57169 6666 57225
rect 6722 57169 6790 57225
rect 6846 57169 6914 57225
rect 6970 57169 7038 57225
rect 7094 57169 7161 57225
rect 5111 57104 7161 57169
rect 5111 57052 5138 57104
rect 5190 57101 5246 57104
rect 5234 57052 5246 57101
rect 5298 57101 5354 57104
rect 5406 57101 5462 57104
rect 5514 57101 5570 57104
rect 5622 57101 5678 57104
rect 5298 57052 5302 57101
rect 5406 57052 5426 57101
rect 5514 57052 5550 57101
rect 5622 57052 5674 57101
rect 5730 57052 5786 57104
rect 5838 57101 5894 57104
rect 5946 57101 6002 57104
rect 6054 57101 6110 57104
rect 5854 57052 5894 57101
rect 5978 57052 6002 57101
rect 6102 57052 6110 57101
rect 6162 57101 6218 57104
rect 6270 57101 6326 57104
rect 6378 57101 6434 57104
rect 6162 57052 6170 57101
rect 6270 57052 6294 57101
rect 6378 57052 6418 57101
rect 6486 57052 6542 57104
rect 6594 57101 6650 57104
rect 6702 57101 6758 57104
rect 6810 57101 6866 57104
rect 6918 57101 6974 57104
rect 6598 57052 6650 57101
rect 6722 57052 6758 57101
rect 6846 57052 6866 57101
rect 6970 57052 6974 57101
rect 7026 57101 7082 57104
rect 7026 57052 7038 57101
rect 7134 57052 7161 57104
rect 5111 57045 5178 57052
rect 5234 57045 5302 57052
rect 5358 57045 5426 57052
rect 5482 57045 5550 57052
rect 5606 57045 5674 57052
rect 5730 57045 5798 57052
rect 5854 57045 5922 57052
rect 5978 57045 6046 57052
rect 6102 57045 6170 57052
rect 6226 57045 6294 57052
rect 6350 57045 6418 57052
rect 6474 57045 6542 57052
rect 6598 57045 6666 57052
rect 6722 57045 6790 57052
rect 6846 57045 6914 57052
rect 6970 57045 7038 57052
rect 7094 57045 7161 57052
rect 5111 56977 7161 57045
rect 5111 56921 5178 56977
rect 5234 56921 5302 56977
rect 5358 56921 5426 56977
rect 5482 56921 5550 56977
rect 5606 56921 5674 56977
rect 5730 56921 5798 56977
rect 5854 56921 5922 56977
rect 5978 56921 6046 56977
rect 6102 56921 6170 56977
rect 6226 56921 6294 56977
rect 6350 56921 6418 56977
rect 6474 56921 6542 56977
rect 6598 56921 6666 56977
rect 6722 56921 6790 56977
rect 6846 56921 6914 56977
rect 6970 56921 7038 56977
rect 7094 56921 7161 56977
rect 5111 56853 7161 56921
rect 5111 56797 5178 56853
rect 5234 56797 5302 56853
rect 5358 56797 5426 56853
rect 5482 56797 5550 56853
rect 5606 56797 5674 56853
rect 5730 56797 5798 56853
rect 5854 56797 5922 56853
rect 5978 56797 6046 56853
rect 6102 56797 6170 56853
rect 6226 56797 6294 56853
rect 6350 56797 6418 56853
rect 6474 56797 6542 56853
rect 6598 56797 6666 56853
rect 6722 56797 6790 56853
rect 6846 56797 6914 56853
rect 6970 56797 7038 56853
rect 7094 56797 7161 56853
rect 5111 56729 7161 56797
rect 5111 56673 5178 56729
rect 5234 56673 5302 56729
rect 5358 56673 5426 56729
rect 5482 56673 5550 56729
rect 5606 56673 5674 56729
rect 5730 56673 5798 56729
rect 5854 56673 5922 56729
rect 5978 56673 6046 56729
rect 6102 56673 6170 56729
rect 6226 56673 6294 56729
rect 6350 56673 6418 56729
rect 6474 56673 6542 56729
rect 6598 56673 6666 56729
rect 6722 56673 6790 56729
rect 6846 56673 6914 56729
rect 6970 56673 7038 56729
rect 7094 56673 7161 56729
rect 5111 56605 7161 56673
rect 5111 56549 5178 56605
rect 5234 56549 5302 56605
rect 5358 56549 5426 56605
rect 5482 56549 5550 56605
rect 5606 56549 5674 56605
rect 5730 56549 5798 56605
rect 5854 56549 5922 56605
rect 5978 56549 6046 56605
rect 6102 56549 6170 56605
rect 6226 56549 6294 56605
rect 6350 56549 6418 56605
rect 6474 56549 6542 56605
rect 6598 56549 6666 56605
rect 6722 56549 6790 56605
rect 6846 56549 6914 56605
rect 6970 56549 7038 56605
rect 7094 56549 7161 56605
rect 5111 56481 7161 56549
rect 5111 56425 5178 56481
rect 5234 56425 5302 56481
rect 5358 56425 5426 56481
rect 5482 56425 5550 56481
rect 5606 56425 5674 56481
rect 5730 56425 5798 56481
rect 5854 56425 5922 56481
rect 5978 56425 6046 56481
rect 6102 56425 6170 56481
rect 6226 56425 6294 56481
rect 6350 56425 6418 56481
rect 6474 56425 6542 56481
rect 6598 56425 6666 56481
rect 6722 56425 6790 56481
rect 6846 56425 6914 56481
rect 6970 56425 7038 56481
rect 7094 56425 7161 56481
rect 5111 56357 7161 56425
rect 5111 56301 5178 56357
rect 5234 56301 5302 56357
rect 5358 56301 5426 56357
rect 5482 56301 5550 56357
rect 5606 56301 5674 56357
rect 5730 56301 5798 56357
rect 5854 56301 5922 56357
rect 5978 56301 6046 56357
rect 6102 56301 6170 56357
rect 6226 56301 6294 56357
rect 6350 56301 6418 56357
rect 6474 56301 6542 56357
rect 6598 56301 6666 56357
rect 6722 56301 6790 56357
rect 6846 56301 6914 56357
rect 6970 56301 7038 56357
rect 7094 56301 7161 56357
rect 5111 56233 7161 56301
rect 5111 56177 5178 56233
rect 5234 56177 5302 56233
rect 5358 56177 5426 56233
rect 5482 56177 5550 56233
rect 5606 56177 5674 56233
rect 5730 56177 5798 56233
rect 5854 56177 5922 56233
rect 5978 56177 6046 56233
rect 6102 56177 6170 56233
rect 6226 56177 6294 56233
rect 6350 56177 6418 56233
rect 6474 56177 6542 56233
rect 6598 56177 6666 56233
rect 6722 56177 6790 56233
rect 6846 56177 6914 56233
rect 6970 56177 7038 56233
rect 7094 56177 7161 56233
rect 5111 56109 7161 56177
rect 5111 56053 5178 56109
rect 5234 56053 5302 56109
rect 5358 56053 5426 56109
rect 5482 56053 5550 56109
rect 5606 56053 5674 56109
rect 5730 56053 5798 56109
rect 5854 56053 5922 56109
rect 5978 56053 6046 56109
rect 6102 56053 6170 56109
rect 6226 56053 6294 56109
rect 6350 56053 6418 56109
rect 6474 56053 6542 56109
rect 6598 56053 6666 56109
rect 6722 56053 6790 56109
rect 6846 56053 6914 56109
rect 6970 56053 7038 56109
rect 7094 56053 7161 56109
rect 5111 54148 7161 56053
rect 5111 54092 5178 54148
rect 5234 54092 5302 54148
rect 5358 54092 5426 54148
rect 5482 54092 5550 54148
rect 5606 54092 5674 54148
rect 5730 54092 5798 54148
rect 5854 54092 5922 54148
rect 5978 54092 6046 54148
rect 6102 54092 6170 54148
rect 6226 54092 6294 54148
rect 6350 54092 6418 54148
rect 6474 54092 6542 54148
rect 6598 54092 6666 54148
rect 6722 54092 6790 54148
rect 6846 54092 6914 54148
rect 6970 54092 7038 54148
rect 7094 54092 7161 54148
rect 5111 54024 7161 54092
rect 5111 53968 5178 54024
rect 5234 53968 5302 54024
rect 5358 53968 5426 54024
rect 5482 53968 5550 54024
rect 5606 53968 5674 54024
rect 5730 53968 5798 54024
rect 5854 53968 5922 54024
rect 5978 53968 6046 54024
rect 6102 53968 6170 54024
rect 6226 53968 6294 54024
rect 6350 53968 6418 54024
rect 6474 53968 6542 54024
rect 6598 53968 6666 54024
rect 6722 53968 6790 54024
rect 6846 53968 6914 54024
rect 6970 53968 7038 54024
rect 7094 53968 7161 54024
rect 5111 53900 7161 53968
rect 5111 53844 5178 53900
rect 5234 53844 5302 53900
rect 5358 53844 5426 53900
rect 5482 53844 5550 53900
rect 5606 53844 5674 53900
rect 5730 53844 5798 53900
rect 5854 53844 5922 53900
rect 5978 53844 6046 53900
rect 6102 53844 6170 53900
rect 6226 53844 6294 53900
rect 6350 53844 6418 53900
rect 6474 53844 6542 53900
rect 6598 53844 6666 53900
rect 6722 53844 6790 53900
rect 6846 53844 6914 53900
rect 6970 53844 7038 53900
rect 7094 53844 7161 53900
rect 5111 53776 7161 53844
rect 5111 53720 5178 53776
rect 5234 53720 5302 53776
rect 5358 53720 5426 53776
rect 5482 53720 5550 53776
rect 5606 53720 5674 53776
rect 5730 53720 5798 53776
rect 5854 53720 5922 53776
rect 5978 53720 6046 53776
rect 6102 53720 6170 53776
rect 6226 53720 6294 53776
rect 6350 53720 6418 53776
rect 6474 53720 6542 53776
rect 6598 53720 6666 53776
rect 6722 53720 6790 53776
rect 6846 53720 6914 53776
rect 6970 53720 7038 53776
rect 7094 53720 7161 53776
rect 5111 53652 7161 53720
rect 5111 53596 5178 53652
rect 5234 53596 5302 53652
rect 5358 53596 5426 53652
rect 5482 53596 5550 53652
rect 5606 53596 5674 53652
rect 5730 53596 5798 53652
rect 5854 53596 5922 53652
rect 5978 53596 6046 53652
rect 6102 53596 6170 53652
rect 6226 53596 6294 53652
rect 6350 53596 6418 53652
rect 6474 53596 6542 53652
rect 6598 53596 6666 53652
rect 6722 53596 6790 53652
rect 6846 53596 6914 53652
rect 6970 53596 7038 53652
rect 7094 53596 7161 53652
rect 5111 53528 7161 53596
rect 5111 53483 5178 53528
rect 5234 53483 5302 53528
rect 5358 53483 5426 53528
rect 5482 53483 5550 53528
rect 5606 53483 5674 53528
rect 5730 53483 5798 53528
rect 5854 53483 5922 53528
rect 5978 53483 6046 53528
rect 6102 53483 6170 53528
rect 6226 53483 6294 53528
rect 6350 53483 6418 53528
rect 6474 53483 6542 53528
rect 6598 53483 6666 53528
rect 6722 53483 6790 53528
rect 6846 53483 6914 53528
rect 6970 53483 7038 53528
rect 7094 53483 7161 53528
rect 5111 53431 5138 53483
rect 5234 53472 5246 53483
rect 5190 53431 5246 53472
rect 5298 53472 5302 53483
rect 5406 53472 5426 53483
rect 5514 53472 5550 53483
rect 5622 53472 5674 53483
rect 5298 53431 5354 53472
rect 5406 53431 5462 53472
rect 5514 53431 5570 53472
rect 5622 53431 5678 53472
rect 5730 53431 5786 53483
rect 5854 53472 5894 53483
rect 5978 53472 6002 53483
rect 6102 53472 6110 53483
rect 5838 53431 5894 53472
rect 5946 53431 6002 53472
rect 6054 53431 6110 53472
rect 6162 53472 6170 53483
rect 6270 53472 6294 53483
rect 6378 53472 6418 53483
rect 6162 53431 6218 53472
rect 6270 53431 6326 53472
rect 6378 53431 6434 53472
rect 6486 53431 6542 53483
rect 6598 53472 6650 53483
rect 6722 53472 6758 53483
rect 6846 53472 6866 53483
rect 6970 53472 6974 53483
rect 6594 53431 6650 53472
rect 6702 53431 6758 53472
rect 6810 53431 6866 53472
rect 6918 53431 6974 53472
rect 7026 53472 7038 53483
rect 7026 53431 7082 53472
rect 7134 53431 7161 53483
rect 5111 53404 7161 53431
rect 5111 53375 5178 53404
rect 5234 53375 5302 53404
rect 5358 53375 5426 53404
rect 5482 53375 5550 53404
rect 5606 53375 5674 53404
rect 5730 53375 5798 53404
rect 5854 53375 5922 53404
rect 5978 53375 6046 53404
rect 6102 53375 6170 53404
rect 6226 53375 6294 53404
rect 6350 53375 6418 53404
rect 6474 53375 6542 53404
rect 6598 53375 6666 53404
rect 6722 53375 6790 53404
rect 6846 53375 6914 53404
rect 6970 53375 7038 53404
rect 7094 53375 7161 53404
rect 5111 53323 5138 53375
rect 5234 53348 5246 53375
rect 5190 53323 5246 53348
rect 5298 53348 5302 53375
rect 5406 53348 5426 53375
rect 5514 53348 5550 53375
rect 5622 53348 5674 53375
rect 5298 53323 5354 53348
rect 5406 53323 5462 53348
rect 5514 53323 5570 53348
rect 5622 53323 5678 53348
rect 5730 53323 5786 53375
rect 5854 53348 5894 53375
rect 5978 53348 6002 53375
rect 6102 53348 6110 53375
rect 5838 53323 5894 53348
rect 5946 53323 6002 53348
rect 6054 53323 6110 53348
rect 6162 53348 6170 53375
rect 6270 53348 6294 53375
rect 6378 53348 6418 53375
rect 6162 53323 6218 53348
rect 6270 53323 6326 53348
rect 6378 53323 6434 53348
rect 6486 53323 6542 53375
rect 6598 53348 6650 53375
rect 6722 53348 6758 53375
rect 6846 53348 6866 53375
rect 6970 53348 6974 53375
rect 6594 53323 6650 53348
rect 6702 53323 6758 53348
rect 6810 53323 6866 53348
rect 6918 53323 6974 53348
rect 7026 53348 7038 53375
rect 7026 53323 7082 53348
rect 7134 53323 7161 53375
rect 5111 53280 7161 53323
rect 5111 53267 5178 53280
rect 5234 53267 5302 53280
rect 5358 53267 5426 53280
rect 5482 53267 5550 53280
rect 5606 53267 5674 53280
rect 5730 53267 5798 53280
rect 5854 53267 5922 53280
rect 5978 53267 6046 53280
rect 6102 53267 6170 53280
rect 6226 53267 6294 53280
rect 6350 53267 6418 53280
rect 6474 53267 6542 53280
rect 6598 53267 6666 53280
rect 6722 53267 6790 53280
rect 6846 53267 6914 53280
rect 6970 53267 7038 53280
rect 7094 53267 7161 53280
rect 5111 53215 5138 53267
rect 5234 53224 5246 53267
rect 5190 53215 5246 53224
rect 5298 53224 5302 53267
rect 5406 53224 5426 53267
rect 5514 53224 5550 53267
rect 5622 53224 5674 53267
rect 5298 53215 5354 53224
rect 5406 53215 5462 53224
rect 5514 53215 5570 53224
rect 5622 53215 5678 53224
rect 5730 53215 5786 53267
rect 5854 53224 5894 53267
rect 5978 53224 6002 53267
rect 6102 53224 6110 53267
rect 5838 53215 5894 53224
rect 5946 53215 6002 53224
rect 6054 53215 6110 53224
rect 6162 53224 6170 53267
rect 6270 53224 6294 53267
rect 6378 53224 6418 53267
rect 6162 53215 6218 53224
rect 6270 53215 6326 53224
rect 6378 53215 6434 53224
rect 6486 53215 6542 53267
rect 6598 53224 6650 53267
rect 6722 53224 6758 53267
rect 6846 53224 6866 53267
rect 6970 53224 6974 53267
rect 6594 53215 6650 53224
rect 6702 53215 6758 53224
rect 6810 53215 6866 53224
rect 6918 53215 6974 53224
rect 7026 53224 7038 53267
rect 7026 53215 7082 53224
rect 7134 53215 7161 53267
rect 5111 53156 7161 53215
rect 5111 53100 5178 53156
rect 5234 53100 5302 53156
rect 5358 53100 5426 53156
rect 5482 53100 5550 53156
rect 5606 53100 5674 53156
rect 5730 53100 5798 53156
rect 5854 53100 5922 53156
rect 5978 53100 6046 53156
rect 6102 53100 6170 53156
rect 6226 53100 6294 53156
rect 6350 53100 6418 53156
rect 6474 53100 6542 53156
rect 6598 53100 6666 53156
rect 6722 53100 6790 53156
rect 6846 53100 6914 53156
rect 6970 53100 7038 53156
rect 7094 53100 7161 53156
rect 5111 53032 7161 53100
rect 5111 52976 5178 53032
rect 5234 52976 5302 53032
rect 5358 52976 5426 53032
rect 5482 52976 5550 53032
rect 5606 52976 5674 53032
rect 5730 52976 5798 53032
rect 5854 52976 5922 53032
rect 5978 52976 6046 53032
rect 6102 52976 6170 53032
rect 6226 52976 6294 53032
rect 6350 52976 6418 53032
rect 6474 52976 6542 53032
rect 6598 52976 6666 53032
rect 6722 52976 6790 53032
rect 6846 52976 6914 53032
rect 6970 52976 7038 53032
rect 7094 52976 7161 53032
rect 5111 52908 7161 52976
rect 5111 52852 5178 52908
rect 5234 52852 5302 52908
rect 5358 52852 5426 52908
rect 5482 52852 5550 52908
rect 5606 52852 5674 52908
rect 5730 52852 5798 52908
rect 5854 52852 5922 52908
rect 5978 52852 6046 52908
rect 6102 52852 6170 52908
rect 6226 52852 6294 52908
rect 6350 52852 6418 52908
rect 6474 52852 6542 52908
rect 6598 52852 6666 52908
rect 6722 52852 6790 52908
rect 6846 52852 6914 52908
rect 6970 52852 7038 52908
rect 7094 52852 7161 52908
rect 5111 52548 7161 52852
rect 5111 52492 5178 52548
rect 5234 52492 5302 52548
rect 5358 52492 5426 52548
rect 5482 52492 5550 52548
rect 5606 52492 5674 52548
rect 5730 52492 5798 52548
rect 5854 52492 5922 52548
rect 5978 52492 6046 52548
rect 6102 52492 6170 52548
rect 6226 52492 6294 52548
rect 6350 52492 6418 52548
rect 6474 52492 6542 52548
rect 6598 52492 6666 52548
rect 6722 52492 6790 52548
rect 6846 52492 6914 52548
rect 6970 52492 7038 52548
rect 7094 52492 7161 52548
rect 5111 52424 7161 52492
rect 5111 52368 5178 52424
rect 5234 52368 5302 52424
rect 5358 52368 5426 52424
rect 5482 52368 5550 52424
rect 5606 52368 5674 52424
rect 5730 52368 5798 52424
rect 5854 52368 5922 52424
rect 5978 52368 6046 52424
rect 6102 52368 6170 52424
rect 6226 52368 6294 52424
rect 6350 52368 6418 52424
rect 6474 52368 6542 52424
rect 6598 52368 6666 52424
rect 6722 52368 6790 52424
rect 6846 52368 6914 52424
rect 6970 52368 7038 52424
rect 7094 52368 7161 52424
rect 5111 52300 7161 52368
rect 5111 52244 5178 52300
rect 5234 52244 5302 52300
rect 5358 52244 5426 52300
rect 5482 52244 5550 52300
rect 5606 52244 5674 52300
rect 5730 52244 5798 52300
rect 5854 52244 5922 52300
rect 5978 52244 6046 52300
rect 6102 52244 6170 52300
rect 6226 52244 6294 52300
rect 6350 52244 6418 52300
rect 6474 52244 6542 52300
rect 6598 52244 6666 52300
rect 6722 52244 6790 52300
rect 6846 52244 6914 52300
rect 6970 52244 7038 52300
rect 7094 52244 7161 52300
rect 5111 52176 7161 52244
rect 5111 52120 5178 52176
rect 5234 52120 5302 52176
rect 5358 52120 5426 52176
rect 5482 52120 5550 52176
rect 5606 52120 5674 52176
rect 5730 52120 5798 52176
rect 5854 52120 5922 52176
rect 5978 52120 6046 52176
rect 6102 52120 6170 52176
rect 6226 52120 6294 52176
rect 6350 52120 6418 52176
rect 6474 52120 6542 52176
rect 6598 52120 6666 52176
rect 6722 52120 6790 52176
rect 6846 52120 6914 52176
rect 6970 52120 7038 52176
rect 7094 52120 7161 52176
rect 5111 52052 7161 52120
rect 5111 52009 5178 52052
rect 5234 52009 5302 52052
rect 5358 52009 5426 52052
rect 5482 52009 5550 52052
rect 5606 52009 5674 52052
rect 5730 52009 5798 52052
rect 5854 52009 5922 52052
rect 5978 52009 6046 52052
rect 6102 52009 6170 52052
rect 6226 52009 6294 52052
rect 6350 52009 6418 52052
rect 6474 52009 6542 52052
rect 6598 52009 6666 52052
rect 6722 52009 6790 52052
rect 6846 52009 6914 52052
rect 6970 52009 7038 52052
rect 7094 52009 7161 52052
rect 5111 51957 5138 52009
rect 5234 51996 5246 52009
rect 5190 51957 5246 51996
rect 5298 51996 5302 52009
rect 5406 51996 5426 52009
rect 5514 51996 5550 52009
rect 5622 51996 5674 52009
rect 5298 51957 5354 51996
rect 5406 51957 5462 51996
rect 5514 51957 5570 51996
rect 5622 51957 5678 51996
rect 5730 51957 5786 52009
rect 5854 51996 5894 52009
rect 5978 51996 6002 52009
rect 6102 51996 6110 52009
rect 5838 51957 5894 51996
rect 5946 51957 6002 51996
rect 6054 51957 6110 51996
rect 6162 51996 6170 52009
rect 6270 51996 6294 52009
rect 6378 51996 6418 52009
rect 6162 51957 6218 51996
rect 6270 51957 6326 51996
rect 6378 51957 6434 51996
rect 6486 51957 6542 52009
rect 6598 51996 6650 52009
rect 6722 51996 6758 52009
rect 6846 51996 6866 52009
rect 6970 51996 6974 52009
rect 6594 51957 6650 51996
rect 6702 51957 6758 51996
rect 6810 51957 6866 51996
rect 6918 51957 6974 51996
rect 7026 51996 7038 52009
rect 7026 51957 7082 51996
rect 7134 51957 7161 52009
rect 5111 51928 7161 51957
rect 5111 51901 5178 51928
rect 5234 51901 5302 51928
rect 5358 51901 5426 51928
rect 5482 51901 5550 51928
rect 5606 51901 5674 51928
rect 5730 51901 5798 51928
rect 5854 51901 5922 51928
rect 5978 51901 6046 51928
rect 6102 51901 6170 51928
rect 6226 51901 6294 51928
rect 6350 51901 6418 51928
rect 6474 51901 6542 51928
rect 6598 51901 6666 51928
rect 6722 51901 6790 51928
rect 6846 51901 6914 51928
rect 6970 51901 7038 51928
rect 7094 51901 7161 51928
rect 5111 51849 5138 51901
rect 5234 51872 5246 51901
rect 5190 51849 5246 51872
rect 5298 51872 5302 51901
rect 5406 51872 5426 51901
rect 5514 51872 5550 51901
rect 5622 51872 5674 51901
rect 5298 51849 5354 51872
rect 5406 51849 5462 51872
rect 5514 51849 5570 51872
rect 5622 51849 5678 51872
rect 5730 51849 5786 51901
rect 5854 51872 5894 51901
rect 5978 51872 6002 51901
rect 6102 51872 6110 51901
rect 5838 51849 5894 51872
rect 5946 51849 6002 51872
rect 6054 51849 6110 51872
rect 6162 51872 6170 51901
rect 6270 51872 6294 51901
rect 6378 51872 6418 51901
rect 6162 51849 6218 51872
rect 6270 51849 6326 51872
rect 6378 51849 6434 51872
rect 6486 51849 6542 51901
rect 6598 51872 6650 51901
rect 6722 51872 6758 51901
rect 6846 51872 6866 51901
rect 6970 51872 6974 51901
rect 6594 51849 6650 51872
rect 6702 51849 6758 51872
rect 6810 51849 6866 51872
rect 6918 51849 6974 51872
rect 7026 51872 7038 51901
rect 7026 51849 7082 51872
rect 7134 51849 7161 51901
rect 5111 51804 7161 51849
rect 5111 51748 5178 51804
rect 5234 51748 5302 51804
rect 5358 51748 5426 51804
rect 5482 51748 5550 51804
rect 5606 51748 5674 51804
rect 5730 51748 5798 51804
rect 5854 51748 5922 51804
rect 5978 51748 6046 51804
rect 6102 51748 6170 51804
rect 6226 51748 6294 51804
rect 6350 51748 6418 51804
rect 6474 51748 6542 51804
rect 6598 51748 6666 51804
rect 6722 51748 6790 51804
rect 6846 51748 6914 51804
rect 6970 51748 7038 51804
rect 7094 51748 7161 51804
rect 5111 51680 7161 51748
rect 5111 51624 5178 51680
rect 5234 51624 5302 51680
rect 5358 51624 5426 51680
rect 5482 51624 5550 51680
rect 5606 51624 5674 51680
rect 5730 51624 5798 51680
rect 5854 51624 5922 51680
rect 5978 51624 6046 51680
rect 6102 51624 6170 51680
rect 6226 51624 6294 51680
rect 6350 51624 6418 51680
rect 6474 51624 6542 51680
rect 6598 51624 6666 51680
rect 6722 51624 6790 51680
rect 6846 51624 6914 51680
rect 6970 51624 7038 51680
rect 7094 51624 7161 51680
rect 5111 51556 7161 51624
rect 5111 51500 5178 51556
rect 5234 51500 5302 51556
rect 5358 51500 5426 51556
rect 5482 51500 5550 51556
rect 5606 51500 5674 51556
rect 5730 51500 5798 51556
rect 5854 51500 5922 51556
rect 5978 51500 6046 51556
rect 6102 51500 6170 51556
rect 6226 51500 6294 51556
rect 6350 51500 6418 51556
rect 6474 51500 6542 51556
rect 6598 51500 6666 51556
rect 6722 51500 6790 51556
rect 6846 51500 6914 51556
rect 6970 51500 7038 51556
rect 7094 51500 7161 51556
rect 5111 51432 7161 51500
rect 5111 51376 5178 51432
rect 5234 51376 5302 51432
rect 5358 51376 5426 51432
rect 5482 51376 5550 51432
rect 5606 51376 5674 51432
rect 5730 51376 5798 51432
rect 5854 51376 5922 51432
rect 5978 51376 6046 51432
rect 6102 51376 6170 51432
rect 6226 51376 6294 51432
rect 6350 51376 6418 51432
rect 6474 51376 6542 51432
rect 6598 51376 6666 51432
rect 6722 51376 6790 51432
rect 6846 51376 6914 51432
rect 6970 51376 7038 51432
rect 7094 51376 7161 51432
rect 5111 51308 7161 51376
rect 5111 51252 5178 51308
rect 5234 51252 5302 51308
rect 5358 51252 5426 51308
rect 5482 51252 5550 51308
rect 5606 51252 5674 51308
rect 5730 51252 5798 51308
rect 5854 51252 5922 51308
rect 5978 51252 6046 51308
rect 6102 51252 6170 51308
rect 6226 51252 6294 51308
rect 6350 51252 6418 51308
rect 6474 51252 6542 51308
rect 6598 51252 6666 51308
rect 6722 51252 6790 51308
rect 6846 51252 6914 51308
rect 6970 51252 7038 51308
rect 7094 51252 7161 51308
rect 5111 51206 7161 51252
rect 5111 51154 5138 51206
rect 5190 51154 5246 51206
rect 5298 51154 5354 51206
rect 5406 51154 5462 51206
rect 5514 51154 5570 51206
rect 5622 51154 5678 51206
rect 5730 51154 5786 51206
rect 5838 51154 5894 51206
rect 5946 51154 6002 51206
rect 6054 51154 6110 51206
rect 6162 51154 6218 51206
rect 6270 51154 6326 51206
rect 6378 51154 6434 51206
rect 6486 51154 6542 51206
rect 6594 51154 6650 51206
rect 6702 51154 6758 51206
rect 6810 51154 6866 51206
rect 6918 51154 6974 51206
rect 7026 51154 7082 51206
rect 7134 51154 7161 51206
rect 5111 51098 7161 51154
rect 5111 51046 5138 51098
rect 5190 51046 5246 51098
rect 5298 51046 5354 51098
rect 5406 51046 5462 51098
rect 5514 51046 5570 51098
rect 5622 51046 5678 51098
rect 5730 51046 5786 51098
rect 5838 51046 5894 51098
rect 5946 51046 6002 51098
rect 6054 51046 6110 51098
rect 6162 51046 6218 51098
rect 6270 51046 6326 51098
rect 6378 51046 6434 51098
rect 6486 51046 6542 51098
rect 6594 51046 6650 51098
rect 6702 51046 6758 51098
rect 6810 51046 6866 51098
rect 6918 51046 6974 51098
rect 7026 51046 7082 51098
rect 7134 51046 7161 51098
rect 5111 50990 7161 51046
rect 5111 50938 5138 50990
rect 5190 50938 5246 50990
rect 5298 50938 5354 50990
rect 5406 50938 5462 50990
rect 5514 50938 5570 50990
rect 5622 50938 5678 50990
rect 5730 50938 5786 50990
rect 5838 50938 5894 50990
rect 5946 50938 6002 50990
rect 6054 50938 6110 50990
rect 6162 50938 6218 50990
rect 6270 50938 6326 50990
rect 6378 50938 6434 50990
rect 6486 50938 6542 50990
rect 6594 50938 6650 50990
rect 6702 50938 6758 50990
rect 6810 50938 6866 50990
rect 6918 50938 6974 50990
rect 7026 50938 7082 50990
rect 7134 50938 7161 50990
rect 5111 50272 7161 50938
rect 5111 50220 5138 50272
rect 5190 50220 5246 50272
rect 5298 50220 5354 50272
rect 5406 50220 5462 50272
rect 5514 50220 5570 50272
rect 5622 50220 5678 50272
rect 5730 50220 5786 50272
rect 5838 50220 5894 50272
rect 5946 50220 6002 50272
rect 6054 50220 6110 50272
rect 6162 50220 6218 50272
rect 6270 50220 6326 50272
rect 6378 50220 6434 50272
rect 6486 50220 6542 50272
rect 6594 50220 6650 50272
rect 6702 50220 6758 50272
rect 6810 50220 6866 50272
rect 6918 50220 6974 50272
rect 7026 50220 7082 50272
rect 7134 50220 7161 50272
rect 5111 50164 7161 50220
rect 5111 50112 5138 50164
rect 5190 50112 5246 50164
rect 5298 50112 5354 50164
rect 5406 50112 5462 50164
rect 5514 50112 5570 50164
rect 5622 50112 5678 50164
rect 5730 50112 5786 50164
rect 5838 50112 5894 50164
rect 5946 50112 6002 50164
rect 6054 50112 6110 50164
rect 6162 50112 6218 50164
rect 6270 50112 6326 50164
rect 6378 50112 6434 50164
rect 6486 50112 6542 50164
rect 6594 50112 6650 50164
rect 6702 50112 6758 50164
rect 6810 50112 6866 50164
rect 6918 50112 6974 50164
rect 7026 50112 7082 50164
rect 7134 50112 7161 50164
rect 5111 50056 7161 50112
rect 5111 50004 5138 50056
rect 5190 50004 5246 50056
rect 5298 50004 5354 50056
rect 5406 50004 5462 50056
rect 5514 50004 5570 50056
rect 5622 50004 5678 50056
rect 5730 50004 5786 50056
rect 5838 50004 5894 50056
rect 5946 50004 6002 50056
rect 6054 50004 6110 50056
rect 6162 50004 6218 50056
rect 6270 50004 6326 50056
rect 6378 50004 6434 50056
rect 6486 50004 6542 50056
rect 6594 50004 6650 50056
rect 6702 50004 6758 50056
rect 6810 50004 6866 50056
rect 6918 50004 6974 50056
rect 7026 50004 7082 50056
rect 7134 50004 7161 50056
rect 5111 49348 7161 50004
rect 5111 49338 5178 49348
rect 5234 49338 5302 49348
rect 5358 49338 5426 49348
rect 5482 49338 5550 49348
rect 5606 49338 5674 49348
rect 5730 49338 5798 49348
rect 5854 49338 5922 49348
rect 5978 49338 6046 49348
rect 6102 49338 6170 49348
rect 6226 49338 6294 49348
rect 6350 49338 6418 49348
rect 6474 49338 6542 49348
rect 6598 49338 6666 49348
rect 6722 49338 6790 49348
rect 6846 49338 6914 49348
rect 6970 49338 7038 49348
rect 7094 49338 7161 49348
rect 5111 49286 5138 49338
rect 5234 49292 5246 49338
rect 5190 49286 5246 49292
rect 5298 49292 5302 49338
rect 5406 49292 5426 49338
rect 5514 49292 5550 49338
rect 5622 49292 5674 49338
rect 5298 49286 5354 49292
rect 5406 49286 5462 49292
rect 5514 49286 5570 49292
rect 5622 49286 5678 49292
rect 5730 49286 5786 49338
rect 5854 49292 5894 49338
rect 5978 49292 6002 49338
rect 6102 49292 6110 49338
rect 5838 49286 5894 49292
rect 5946 49286 6002 49292
rect 6054 49286 6110 49292
rect 6162 49292 6170 49338
rect 6270 49292 6294 49338
rect 6378 49292 6418 49338
rect 6162 49286 6218 49292
rect 6270 49286 6326 49292
rect 6378 49286 6434 49292
rect 6486 49286 6542 49338
rect 6598 49292 6650 49338
rect 6722 49292 6758 49338
rect 6846 49292 6866 49338
rect 6970 49292 6974 49338
rect 6594 49286 6650 49292
rect 6702 49286 6758 49292
rect 6810 49286 6866 49292
rect 6918 49286 6974 49292
rect 7026 49292 7038 49338
rect 7026 49286 7082 49292
rect 7134 49286 7161 49338
rect 5111 49230 7161 49286
rect 5111 49178 5138 49230
rect 5190 49224 5246 49230
rect 5234 49178 5246 49224
rect 5298 49224 5354 49230
rect 5406 49224 5462 49230
rect 5514 49224 5570 49230
rect 5622 49224 5678 49230
rect 5298 49178 5302 49224
rect 5406 49178 5426 49224
rect 5514 49178 5550 49224
rect 5622 49178 5674 49224
rect 5730 49178 5786 49230
rect 5838 49224 5894 49230
rect 5946 49224 6002 49230
rect 6054 49224 6110 49230
rect 5854 49178 5894 49224
rect 5978 49178 6002 49224
rect 6102 49178 6110 49224
rect 6162 49224 6218 49230
rect 6270 49224 6326 49230
rect 6378 49224 6434 49230
rect 6162 49178 6170 49224
rect 6270 49178 6294 49224
rect 6378 49178 6418 49224
rect 6486 49178 6542 49230
rect 6594 49224 6650 49230
rect 6702 49224 6758 49230
rect 6810 49224 6866 49230
rect 6918 49224 6974 49230
rect 6598 49178 6650 49224
rect 6722 49178 6758 49224
rect 6846 49178 6866 49224
rect 6970 49178 6974 49224
rect 7026 49224 7082 49230
rect 7026 49178 7038 49224
rect 7134 49178 7161 49230
rect 5111 49168 5178 49178
rect 5234 49168 5302 49178
rect 5358 49168 5426 49178
rect 5482 49168 5550 49178
rect 5606 49168 5674 49178
rect 5730 49168 5798 49178
rect 5854 49168 5922 49178
rect 5978 49168 6046 49178
rect 6102 49168 6170 49178
rect 6226 49168 6294 49178
rect 6350 49168 6418 49178
rect 6474 49168 6542 49178
rect 6598 49168 6666 49178
rect 6722 49168 6790 49178
rect 6846 49168 6914 49178
rect 6970 49168 7038 49178
rect 7094 49168 7161 49178
rect 5111 49122 7161 49168
rect 5111 49070 5138 49122
rect 5190 49100 5246 49122
rect 5234 49070 5246 49100
rect 5298 49100 5354 49122
rect 5406 49100 5462 49122
rect 5514 49100 5570 49122
rect 5622 49100 5678 49122
rect 5298 49070 5302 49100
rect 5406 49070 5426 49100
rect 5514 49070 5550 49100
rect 5622 49070 5674 49100
rect 5730 49070 5786 49122
rect 5838 49100 5894 49122
rect 5946 49100 6002 49122
rect 6054 49100 6110 49122
rect 5854 49070 5894 49100
rect 5978 49070 6002 49100
rect 6102 49070 6110 49100
rect 6162 49100 6218 49122
rect 6270 49100 6326 49122
rect 6378 49100 6434 49122
rect 6162 49070 6170 49100
rect 6270 49070 6294 49100
rect 6378 49070 6418 49100
rect 6486 49070 6542 49122
rect 6594 49100 6650 49122
rect 6702 49100 6758 49122
rect 6810 49100 6866 49122
rect 6918 49100 6974 49122
rect 6598 49070 6650 49100
rect 6722 49070 6758 49100
rect 6846 49070 6866 49100
rect 6970 49070 6974 49100
rect 7026 49100 7082 49122
rect 7026 49070 7038 49100
rect 7134 49070 7161 49122
rect 5111 49044 5178 49070
rect 5234 49044 5302 49070
rect 5358 49044 5426 49070
rect 5482 49044 5550 49070
rect 5606 49044 5674 49070
rect 5730 49044 5798 49070
rect 5854 49044 5922 49070
rect 5978 49044 6046 49070
rect 6102 49044 6170 49070
rect 6226 49044 6294 49070
rect 6350 49044 6418 49070
rect 6474 49044 6542 49070
rect 6598 49044 6666 49070
rect 6722 49044 6790 49070
rect 6846 49044 6914 49070
rect 6970 49044 7038 49070
rect 7094 49044 7161 49070
rect 5111 48976 7161 49044
rect 5111 48920 5178 48976
rect 5234 48920 5302 48976
rect 5358 48920 5426 48976
rect 5482 48920 5550 48976
rect 5606 48920 5674 48976
rect 5730 48920 5798 48976
rect 5854 48920 5922 48976
rect 5978 48920 6046 48976
rect 6102 48920 6170 48976
rect 6226 48920 6294 48976
rect 6350 48920 6418 48976
rect 6474 48920 6542 48976
rect 6598 48920 6666 48976
rect 6722 48920 6790 48976
rect 6846 48920 6914 48976
rect 6970 48920 7038 48976
rect 7094 48920 7161 48976
rect 5111 48852 7161 48920
rect 5111 48796 5178 48852
rect 5234 48796 5302 48852
rect 5358 48796 5426 48852
rect 5482 48796 5550 48852
rect 5606 48796 5674 48852
rect 5730 48796 5798 48852
rect 5854 48796 5922 48852
rect 5978 48796 6046 48852
rect 6102 48796 6170 48852
rect 6226 48796 6294 48852
rect 6350 48796 6418 48852
rect 6474 48796 6542 48852
rect 6598 48796 6666 48852
rect 6722 48796 6790 48852
rect 6846 48796 6914 48852
rect 6970 48796 7038 48852
rect 7094 48796 7161 48852
rect 5111 48728 7161 48796
rect 5111 48672 5178 48728
rect 5234 48672 5302 48728
rect 5358 48672 5426 48728
rect 5482 48672 5550 48728
rect 5606 48672 5674 48728
rect 5730 48672 5798 48728
rect 5854 48672 5922 48728
rect 5978 48672 6046 48728
rect 6102 48672 6170 48728
rect 6226 48672 6294 48728
rect 6350 48672 6418 48728
rect 6474 48672 6542 48728
rect 6598 48672 6666 48728
rect 6722 48672 6790 48728
rect 6846 48672 6914 48728
rect 6970 48672 7038 48728
rect 7094 48672 7161 48728
rect 5111 48604 7161 48672
rect 5111 48548 5178 48604
rect 5234 48548 5302 48604
rect 5358 48548 5426 48604
rect 5482 48548 5550 48604
rect 5606 48548 5674 48604
rect 5730 48548 5798 48604
rect 5854 48548 5922 48604
rect 5978 48548 6046 48604
rect 6102 48548 6170 48604
rect 6226 48548 6294 48604
rect 6350 48548 6418 48604
rect 6474 48548 6542 48604
rect 6598 48548 6666 48604
rect 6722 48548 6790 48604
rect 6846 48548 6914 48604
rect 6970 48548 7038 48604
rect 7094 48548 7161 48604
rect 5111 48480 7161 48548
rect 5111 48427 5178 48480
rect 5234 48427 5302 48480
rect 5358 48427 5426 48480
rect 5482 48427 5550 48480
rect 5606 48427 5674 48480
rect 5730 48427 5798 48480
rect 5854 48427 5922 48480
rect 5978 48427 6046 48480
rect 6102 48427 6170 48480
rect 6226 48427 6294 48480
rect 6350 48427 6418 48480
rect 6474 48427 6542 48480
rect 6598 48427 6666 48480
rect 6722 48427 6790 48480
rect 6846 48427 6914 48480
rect 6970 48427 7038 48480
rect 7094 48427 7161 48480
rect 5111 48375 5138 48427
rect 5234 48424 5246 48427
rect 5190 48375 5246 48424
rect 5298 48424 5302 48427
rect 5406 48424 5426 48427
rect 5514 48424 5550 48427
rect 5622 48424 5674 48427
rect 5298 48375 5354 48424
rect 5406 48375 5462 48424
rect 5514 48375 5570 48424
rect 5622 48375 5678 48424
rect 5730 48375 5786 48427
rect 5854 48424 5894 48427
rect 5978 48424 6002 48427
rect 6102 48424 6110 48427
rect 5838 48375 5894 48424
rect 5946 48375 6002 48424
rect 6054 48375 6110 48424
rect 6162 48424 6170 48427
rect 6270 48424 6294 48427
rect 6378 48424 6418 48427
rect 6162 48375 6218 48424
rect 6270 48375 6326 48424
rect 6378 48375 6434 48424
rect 6486 48375 6542 48427
rect 6598 48424 6650 48427
rect 6722 48424 6758 48427
rect 6846 48424 6866 48427
rect 6970 48424 6974 48427
rect 6594 48375 6650 48424
rect 6702 48375 6758 48424
rect 6810 48375 6866 48424
rect 6918 48375 6974 48424
rect 7026 48424 7038 48427
rect 7026 48375 7082 48424
rect 7134 48375 7161 48427
rect 5111 48356 7161 48375
rect 5111 48319 5178 48356
rect 5234 48319 5302 48356
rect 5358 48319 5426 48356
rect 5482 48319 5550 48356
rect 5606 48319 5674 48356
rect 5730 48319 5798 48356
rect 5854 48319 5922 48356
rect 5978 48319 6046 48356
rect 6102 48319 6170 48356
rect 6226 48319 6294 48356
rect 6350 48319 6418 48356
rect 6474 48319 6542 48356
rect 6598 48319 6666 48356
rect 6722 48319 6790 48356
rect 6846 48319 6914 48356
rect 6970 48319 7038 48356
rect 7094 48319 7161 48356
rect 5111 48267 5138 48319
rect 5234 48300 5246 48319
rect 5190 48267 5246 48300
rect 5298 48300 5302 48319
rect 5406 48300 5426 48319
rect 5514 48300 5550 48319
rect 5622 48300 5674 48319
rect 5298 48267 5354 48300
rect 5406 48267 5462 48300
rect 5514 48267 5570 48300
rect 5622 48267 5678 48300
rect 5730 48267 5786 48319
rect 5854 48300 5894 48319
rect 5978 48300 6002 48319
rect 6102 48300 6110 48319
rect 5838 48267 5894 48300
rect 5946 48267 6002 48300
rect 6054 48267 6110 48300
rect 6162 48300 6170 48319
rect 6270 48300 6294 48319
rect 6378 48300 6418 48319
rect 6162 48267 6218 48300
rect 6270 48267 6326 48300
rect 6378 48267 6434 48300
rect 6486 48267 6542 48319
rect 6598 48300 6650 48319
rect 6722 48300 6758 48319
rect 6846 48300 6866 48319
rect 6970 48300 6974 48319
rect 6594 48267 6650 48300
rect 6702 48267 6758 48300
rect 6810 48267 6866 48300
rect 6918 48267 6974 48300
rect 7026 48300 7038 48319
rect 7026 48267 7082 48300
rect 7134 48267 7161 48319
rect 5111 48232 7161 48267
rect 5111 48176 5178 48232
rect 5234 48176 5302 48232
rect 5358 48176 5426 48232
rect 5482 48176 5550 48232
rect 5606 48176 5674 48232
rect 5730 48176 5798 48232
rect 5854 48176 5922 48232
rect 5978 48176 6046 48232
rect 6102 48176 6170 48232
rect 6226 48176 6294 48232
rect 6350 48176 6418 48232
rect 6474 48176 6542 48232
rect 6598 48176 6666 48232
rect 6722 48176 6790 48232
rect 6846 48176 6914 48232
rect 6970 48176 7038 48232
rect 7094 48176 7161 48232
rect 5111 48108 7161 48176
rect 5111 48052 5178 48108
rect 5234 48052 5302 48108
rect 5358 48052 5426 48108
rect 5482 48052 5550 48108
rect 5606 48052 5674 48108
rect 5730 48052 5798 48108
rect 5854 48052 5922 48108
rect 5978 48052 6046 48108
rect 6102 48052 6170 48108
rect 6226 48052 6294 48108
rect 6350 48052 6418 48108
rect 6474 48052 6542 48108
rect 6598 48052 6666 48108
rect 6722 48052 6790 48108
rect 6846 48052 6914 48108
rect 6970 48052 7038 48108
rect 7094 48052 7161 48108
rect 5111 47163 7161 48052
rect 7221 55748 7757 57278
rect 7221 55692 7275 55748
rect 7331 55692 7399 55748
rect 7455 55692 7523 55748
rect 7579 55692 7647 55748
rect 7703 55692 7757 55748
rect 7221 55624 7757 55692
rect 7221 55568 7275 55624
rect 7331 55568 7399 55624
rect 7455 55568 7523 55624
rect 7579 55568 7647 55624
rect 7703 55568 7757 55624
rect 7221 55500 7757 55568
rect 7221 55444 7275 55500
rect 7331 55444 7399 55500
rect 7455 55444 7523 55500
rect 7579 55444 7647 55500
rect 7703 55444 7757 55500
rect 7221 55376 7757 55444
rect 7221 55320 7275 55376
rect 7331 55320 7399 55376
rect 7455 55320 7523 55376
rect 7579 55320 7647 55376
rect 7703 55320 7757 55376
rect 7221 55252 7757 55320
rect 7221 55196 7275 55252
rect 7331 55196 7399 55252
rect 7455 55196 7523 55252
rect 7579 55196 7647 55252
rect 7703 55196 7757 55252
rect 7221 55128 7757 55196
rect 7221 55072 7275 55128
rect 7331 55072 7399 55128
rect 7455 55072 7523 55128
rect 7579 55072 7647 55128
rect 7703 55072 7757 55128
rect 7221 55004 7757 55072
rect 7221 54948 7275 55004
rect 7331 54948 7399 55004
rect 7455 54948 7523 55004
rect 7579 54948 7647 55004
rect 7703 54948 7757 55004
rect 7221 54880 7757 54948
rect 7221 54824 7275 54880
rect 7331 54824 7399 54880
rect 7455 54824 7523 54880
rect 7579 54824 7647 54880
rect 7703 54824 7757 54880
rect 7221 54756 7757 54824
rect 7221 54700 7275 54756
rect 7331 54700 7399 54756
rect 7455 54700 7523 54756
rect 7579 54700 7647 54756
rect 7703 54700 7757 54756
rect 7221 54632 7757 54700
rect 7221 54576 7275 54632
rect 7331 54576 7399 54632
rect 7455 54576 7523 54632
rect 7579 54576 7647 54632
rect 7703 54576 7757 54632
rect 7221 54508 7757 54576
rect 7221 54452 7275 54508
rect 7331 54452 7399 54508
rect 7455 54452 7523 54508
rect 7579 54452 7647 54508
rect 7703 54452 7757 54508
rect 7221 52572 7757 54452
rect 7221 52520 7247 52572
rect 7299 52520 7355 52572
rect 7407 52520 7463 52572
rect 7515 52520 7571 52572
rect 7623 52520 7679 52572
rect 7731 52520 7757 52572
rect 7221 52464 7757 52520
rect 7221 52412 7247 52464
rect 7299 52412 7355 52464
rect 7407 52412 7463 52464
rect 7515 52412 7571 52464
rect 7623 52412 7679 52464
rect 7731 52412 7757 52464
rect 7221 52356 7757 52412
rect 7221 52304 7247 52356
rect 7299 52304 7355 52356
rect 7407 52304 7463 52356
rect 7515 52304 7571 52356
rect 7623 52304 7679 52356
rect 7731 52304 7757 52356
rect 7221 51619 7757 52304
rect 7221 51567 7247 51619
rect 7299 51567 7355 51619
rect 7407 51567 7463 51619
rect 7515 51567 7571 51619
rect 7623 51567 7679 51619
rect 7731 51567 7757 51619
rect 7221 51511 7757 51567
rect 7221 51459 7247 51511
rect 7299 51459 7355 51511
rect 7407 51459 7463 51511
rect 7515 51459 7571 51511
rect 7623 51459 7679 51511
rect 7731 51459 7757 51511
rect 7221 50685 7757 51459
rect 7221 50633 7247 50685
rect 7299 50633 7355 50685
rect 7407 50633 7463 50685
rect 7515 50633 7571 50685
rect 7623 50633 7679 50685
rect 7731 50633 7757 50685
rect 7221 50577 7757 50633
rect 7221 50525 7247 50577
rect 7299 50525 7355 50577
rect 7407 50525 7463 50577
rect 7515 50525 7571 50577
rect 7623 50525 7679 50577
rect 7731 50525 7757 50577
rect 7221 49751 7757 50525
rect 7221 49699 7247 49751
rect 7299 49699 7355 49751
rect 7407 49699 7463 49751
rect 7515 49699 7571 49751
rect 7623 49699 7679 49751
rect 7731 49699 7757 49751
rect 7221 49643 7757 49699
rect 7221 49591 7247 49643
rect 7299 49591 7355 49643
rect 7407 49591 7463 49643
rect 7515 49591 7571 49643
rect 7623 49591 7679 49643
rect 7731 49591 7757 49643
rect 7221 48817 7757 49591
rect 7221 48765 7247 48817
rect 7299 48765 7355 48817
rect 7407 48765 7463 48817
rect 7515 48765 7571 48817
rect 7623 48765 7679 48817
rect 7731 48765 7757 48817
rect 7221 48709 7757 48765
rect 7221 48657 7247 48709
rect 7299 48657 7355 48709
rect 7407 48657 7463 48709
rect 7515 48657 7571 48709
rect 7623 48657 7679 48709
rect 7731 48657 7757 48709
rect 7221 47972 7757 48657
rect 7221 47920 7247 47972
rect 7299 47920 7355 47972
rect 7407 47920 7463 47972
rect 7515 47920 7571 47972
rect 7623 47920 7679 47972
rect 7731 47920 7757 47972
rect 7221 47864 7757 47920
rect 7221 47812 7247 47864
rect 7299 47812 7355 47864
rect 7407 47812 7463 47864
rect 7515 47812 7571 47864
rect 7623 47812 7679 47864
rect 7731 47812 7757 47864
rect 7221 47756 7757 47812
rect 7221 47704 7247 47756
rect 7299 47748 7355 47756
rect 7407 47748 7463 47756
rect 7331 47704 7355 47748
rect 7455 47704 7463 47748
rect 7515 47748 7571 47756
rect 7623 47748 7679 47756
rect 7515 47704 7523 47748
rect 7623 47704 7647 47748
rect 7731 47704 7757 47756
rect 7221 47692 7275 47704
rect 7331 47692 7399 47704
rect 7455 47692 7523 47704
rect 7579 47692 7647 47704
rect 7703 47692 7757 47704
rect 7221 47624 7757 47692
rect 7221 47568 7275 47624
rect 7331 47568 7399 47624
rect 7455 47568 7523 47624
rect 7579 47568 7647 47624
rect 7703 47568 7757 47624
rect 7221 47500 7757 47568
rect 7221 47444 7275 47500
rect 7331 47444 7399 47500
rect 7455 47444 7523 47500
rect 7579 47444 7647 47500
rect 7703 47444 7757 47500
rect 7221 47376 7757 47444
rect 7221 47320 7275 47376
rect 7331 47320 7399 47376
rect 7455 47320 7523 47376
rect 7579 47320 7647 47376
rect 7703 47320 7757 47376
rect 7221 47252 7757 47320
rect 7221 47196 7275 47252
rect 7331 47196 7399 47252
rect 7455 47196 7523 47252
rect 7579 47196 7647 47252
rect 7703 47196 7757 47252
rect 7221 47163 7757 47196
rect 7817 57225 9867 57447
rect 10187 57499 12237 57600
rect 10187 57447 10322 57499
rect 10374 57447 10430 57499
rect 10482 57447 10538 57499
rect 10590 57447 10646 57499
rect 10698 57447 10754 57499
rect 10806 57447 10862 57499
rect 10914 57447 10970 57499
rect 11022 57447 11078 57499
rect 11130 57447 11186 57499
rect 11238 57447 11294 57499
rect 11346 57447 11402 57499
rect 11454 57447 11510 57499
rect 11562 57447 11618 57499
rect 11670 57447 11726 57499
rect 11778 57447 11834 57499
rect 11886 57447 11942 57499
rect 11994 57447 12050 57499
rect 12102 57447 12237 57499
rect 7817 57169 7884 57225
rect 7940 57169 8008 57225
rect 8064 57169 8132 57225
rect 8188 57169 8256 57225
rect 8312 57169 8380 57225
rect 8436 57169 8504 57225
rect 8560 57169 8628 57225
rect 8684 57169 8752 57225
rect 8808 57169 8876 57225
rect 8932 57169 9000 57225
rect 9056 57169 9124 57225
rect 9180 57169 9248 57225
rect 9304 57169 9372 57225
rect 9428 57169 9496 57225
rect 9552 57169 9620 57225
rect 9676 57169 9744 57225
rect 9800 57169 9867 57225
rect 7817 57104 9867 57169
rect 7817 57052 7844 57104
rect 7896 57101 7952 57104
rect 7940 57052 7952 57101
rect 8004 57101 8060 57104
rect 8112 57101 8168 57104
rect 8220 57101 8276 57104
rect 8328 57101 8384 57104
rect 8004 57052 8008 57101
rect 8112 57052 8132 57101
rect 8220 57052 8256 57101
rect 8328 57052 8380 57101
rect 8436 57052 8492 57104
rect 8544 57101 8600 57104
rect 8652 57101 8708 57104
rect 8760 57101 8816 57104
rect 8560 57052 8600 57101
rect 8684 57052 8708 57101
rect 8808 57052 8816 57101
rect 8868 57101 8924 57104
rect 8976 57101 9032 57104
rect 9084 57101 9140 57104
rect 8868 57052 8876 57101
rect 8976 57052 9000 57101
rect 9084 57052 9124 57101
rect 9192 57052 9248 57104
rect 9300 57101 9356 57104
rect 9408 57101 9464 57104
rect 9516 57101 9572 57104
rect 9624 57101 9680 57104
rect 9304 57052 9356 57101
rect 9428 57052 9464 57101
rect 9552 57052 9572 57101
rect 9676 57052 9680 57101
rect 9732 57101 9788 57104
rect 9732 57052 9744 57101
rect 9840 57052 9867 57104
rect 7817 57045 7884 57052
rect 7940 57045 8008 57052
rect 8064 57045 8132 57052
rect 8188 57045 8256 57052
rect 8312 57045 8380 57052
rect 8436 57045 8504 57052
rect 8560 57045 8628 57052
rect 8684 57045 8752 57052
rect 8808 57045 8876 57052
rect 8932 57045 9000 57052
rect 9056 57045 9124 57052
rect 9180 57045 9248 57052
rect 9304 57045 9372 57052
rect 9428 57045 9496 57052
rect 9552 57045 9620 57052
rect 9676 57045 9744 57052
rect 9800 57045 9867 57052
rect 7817 56977 9867 57045
rect 7817 56921 7884 56977
rect 7940 56921 8008 56977
rect 8064 56921 8132 56977
rect 8188 56921 8256 56977
rect 8312 56921 8380 56977
rect 8436 56921 8504 56977
rect 8560 56921 8628 56977
rect 8684 56921 8752 56977
rect 8808 56921 8876 56977
rect 8932 56921 9000 56977
rect 9056 56921 9124 56977
rect 9180 56921 9248 56977
rect 9304 56921 9372 56977
rect 9428 56921 9496 56977
rect 9552 56921 9620 56977
rect 9676 56921 9744 56977
rect 9800 56921 9867 56977
rect 7817 56853 9867 56921
rect 7817 56797 7884 56853
rect 7940 56797 8008 56853
rect 8064 56797 8132 56853
rect 8188 56797 8256 56853
rect 8312 56797 8380 56853
rect 8436 56797 8504 56853
rect 8560 56797 8628 56853
rect 8684 56797 8752 56853
rect 8808 56797 8876 56853
rect 8932 56797 9000 56853
rect 9056 56797 9124 56853
rect 9180 56797 9248 56853
rect 9304 56797 9372 56853
rect 9428 56797 9496 56853
rect 9552 56797 9620 56853
rect 9676 56797 9744 56853
rect 9800 56797 9867 56853
rect 7817 56729 9867 56797
rect 7817 56673 7884 56729
rect 7940 56673 8008 56729
rect 8064 56673 8132 56729
rect 8188 56673 8256 56729
rect 8312 56673 8380 56729
rect 8436 56673 8504 56729
rect 8560 56673 8628 56729
rect 8684 56673 8752 56729
rect 8808 56673 8876 56729
rect 8932 56673 9000 56729
rect 9056 56673 9124 56729
rect 9180 56673 9248 56729
rect 9304 56673 9372 56729
rect 9428 56673 9496 56729
rect 9552 56673 9620 56729
rect 9676 56673 9744 56729
rect 9800 56673 9867 56729
rect 7817 56605 9867 56673
rect 7817 56549 7884 56605
rect 7940 56549 8008 56605
rect 8064 56549 8132 56605
rect 8188 56549 8256 56605
rect 8312 56549 8380 56605
rect 8436 56549 8504 56605
rect 8560 56549 8628 56605
rect 8684 56549 8752 56605
rect 8808 56549 8876 56605
rect 8932 56549 9000 56605
rect 9056 56549 9124 56605
rect 9180 56549 9248 56605
rect 9304 56549 9372 56605
rect 9428 56549 9496 56605
rect 9552 56549 9620 56605
rect 9676 56549 9744 56605
rect 9800 56549 9867 56605
rect 7817 56481 9867 56549
rect 7817 56425 7884 56481
rect 7940 56425 8008 56481
rect 8064 56425 8132 56481
rect 8188 56425 8256 56481
rect 8312 56425 8380 56481
rect 8436 56425 8504 56481
rect 8560 56425 8628 56481
rect 8684 56425 8752 56481
rect 8808 56425 8876 56481
rect 8932 56425 9000 56481
rect 9056 56425 9124 56481
rect 9180 56425 9248 56481
rect 9304 56425 9372 56481
rect 9428 56425 9496 56481
rect 9552 56425 9620 56481
rect 9676 56425 9744 56481
rect 9800 56425 9867 56481
rect 7817 56357 9867 56425
rect 7817 56301 7884 56357
rect 7940 56301 8008 56357
rect 8064 56301 8132 56357
rect 8188 56301 8256 56357
rect 8312 56301 8380 56357
rect 8436 56301 8504 56357
rect 8560 56301 8628 56357
rect 8684 56301 8752 56357
rect 8808 56301 8876 56357
rect 8932 56301 9000 56357
rect 9056 56301 9124 56357
rect 9180 56301 9248 56357
rect 9304 56301 9372 56357
rect 9428 56301 9496 56357
rect 9552 56301 9620 56357
rect 9676 56301 9744 56357
rect 9800 56301 9867 56357
rect 7817 56233 9867 56301
rect 7817 56177 7884 56233
rect 7940 56177 8008 56233
rect 8064 56177 8132 56233
rect 8188 56177 8256 56233
rect 8312 56177 8380 56233
rect 8436 56177 8504 56233
rect 8560 56177 8628 56233
rect 8684 56177 8752 56233
rect 8808 56177 8876 56233
rect 8932 56177 9000 56233
rect 9056 56177 9124 56233
rect 9180 56177 9248 56233
rect 9304 56177 9372 56233
rect 9428 56177 9496 56233
rect 9552 56177 9620 56233
rect 9676 56177 9744 56233
rect 9800 56177 9867 56233
rect 7817 56109 9867 56177
rect 7817 56053 7884 56109
rect 7940 56053 8008 56109
rect 8064 56053 8132 56109
rect 8188 56053 8256 56109
rect 8312 56053 8380 56109
rect 8436 56053 8504 56109
rect 8560 56053 8628 56109
rect 8684 56053 8752 56109
rect 8808 56053 8876 56109
rect 8932 56053 9000 56109
rect 9056 56053 9124 56109
rect 9180 56053 9248 56109
rect 9304 56053 9372 56109
rect 9428 56053 9496 56109
rect 9552 56053 9620 56109
rect 9676 56053 9744 56109
rect 9800 56053 9867 56109
rect 7817 54148 9867 56053
rect 7817 54092 7884 54148
rect 7940 54092 8008 54148
rect 8064 54092 8132 54148
rect 8188 54092 8256 54148
rect 8312 54092 8380 54148
rect 8436 54092 8504 54148
rect 8560 54092 8628 54148
rect 8684 54092 8752 54148
rect 8808 54092 8876 54148
rect 8932 54092 9000 54148
rect 9056 54092 9124 54148
rect 9180 54092 9248 54148
rect 9304 54092 9372 54148
rect 9428 54092 9496 54148
rect 9552 54092 9620 54148
rect 9676 54092 9744 54148
rect 9800 54092 9867 54148
rect 7817 54024 9867 54092
rect 7817 53968 7884 54024
rect 7940 53968 8008 54024
rect 8064 53968 8132 54024
rect 8188 53968 8256 54024
rect 8312 53968 8380 54024
rect 8436 53968 8504 54024
rect 8560 53968 8628 54024
rect 8684 53968 8752 54024
rect 8808 53968 8876 54024
rect 8932 53968 9000 54024
rect 9056 53968 9124 54024
rect 9180 53968 9248 54024
rect 9304 53968 9372 54024
rect 9428 53968 9496 54024
rect 9552 53968 9620 54024
rect 9676 53968 9744 54024
rect 9800 53968 9867 54024
rect 7817 53900 9867 53968
rect 7817 53844 7884 53900
rect 7940 53844 8008 53900
rect 8064 53844 8132 53900
rect 8188 53844 8256 53900
rect 8312 53844 8380 53900
rect 8436 53844 8504 53900
rect 8560 53844 8628 53900
rect 8684 53844 8752 53900
rect 8808 53844 8876 53900
rect 8932 53844 9000 53900
rect 9056 53844 9124 53900
rect 9180 53844 9248 53900
rect 9304 53844 9372 53900
rect 9428 53844 9496 53900
rect 9552 53844 9620 53900
rect 9676 53844 9744 53900
rect 9800 53844 9867 53900
rect 7817 53776 9867 53844
rect 7817 53720 7884 53776
rect 7940 53720 8008 53776
rect 8064 53720 8132 53776
rect 8188 53720 8256 53776
rect 8312 53720 8380 53776
rect 8436 53720 8504 53776
rect 8560 53720 8628 53776
rect 8684 53720 8752 53776
rect 8808 53720 8876 53776
rect 8932 53720 9000 53776
rect 9056 53720 9124 53776
rect 9180 53720 9248 53776
rect 9304 53720 9372 53776
rect 9428 53720 9496 53776
rect 9552 53720 9620 53776
rect 9676 53720 9744 53776
rect 9800 53720 9867 53776
rect 7817 53652 9867 53720
rect 7817 53596 7884 53652
rect 7940 53596 8008 53652
rect 8064 53596 8132 53652
rect 8188 53596 8256 53652
rect 8312 53596 8380 53652
rect 8436 53596 8504 53652
rect 8560 53596 8628 53652
rect 8684 53596 8752 53652
rect 8808 53596 8876 53652
rect 8932 53596 9000 53652
rect 9056 53596 9124 53652
rect 9180 53596 9248 53652
rect 9304 53596 9372 53652
rect 9428 53596 9496 53652
rect 9552 53596 9620 53652
rect 9676 53596 9744 53652
rect 9800 53596 9867 53652
rect 7817 53528 9867 53596
rect 7817 53483 7884 53528
rect 7940 53483 8008 53528
rect 8064 53483 8132 53528
rect 8188 53483 8256 53528
rect 8312 53483 8380 53528
rect 8436 53483 8504 53528
rect 8560 53483 8628 53528
rect 8684 53483 8752 53528
rect 8808 53483 8876 53528
rect 8932 53483 9000 53528
rect 9056 53483 9124 53528
rect 9180 53483 9248 53528
rect 9304 53483 9372 53528
rect 9428 53483 9496 53528
rect 9552 53483 9620 53528
rect 9676 53483 9744 53528
rect 9800 53483 9867 53528
rect 7817 53431 7844 53483
rect 7940 53472 7952 53483
rect 7896 53431 7952 53472
rect 8004 53472 8008 53483
rect 8112 53472 8132 53483
rect 8220 53472 8256 53483
rect 8328 53472 8380 53483
rect 8004 53431 8060 53472
rect 8112 53431 8168 53472
rect 8220 53431 8276 53472
rect 8328 53431 8384 53472
rect 8436 53431 8492 53483
rect 8560 53472 8600 53483
rect 8684 53472 8708 53483
rect 8808 53472 8816 53483
rect 8544 53431 8600 53472
rect 8652 53431 8708 53472
rect 8760 53431 8816 53472
rect 8868 53472 8876 53483
rect 8976 53472 9000 53483
rect 9084 53472 9124 53483
rect 8868 53431 8924 53472
rect 8976 53431 9032 53472
rect 9084 53431 9140 53472
rect 9192 53431 9248 53483
rect 9304 53472 9356 53483
rect 9428 53472 9464 53483
rect 9552 53472 9572 53483
rect 9676 53472 9680 53483
rect 9300 53431 9356 53472
rect 9408 53431 9464 53472
rect 9516 53431 9572 53472
rect 9624 53431 9680 53472
rect 9732 53472 9744 53483
rect 9732 53431 9788 53472
rect 9840 53431 9867 53483
rect 7817 53404 9867 53431
rect 7817 53375 7884 53404
rect 7940 53375 8008 53404
rect 8064 53375 8132 53404
rect 8188 53375 8256 53404
rect 8312 53375 8380 53404
rect 8436 53375 8504 53404
rect 8560 53375 8628 53404
rect 8684 53375 8752 53404
rect 8808 53375 8876 53404
rect 8932 53375 9000 53404
rect 9056 53375 9124 53404
rect 9180 53375 9248 53404
rect 9304 53375 9372 53404
rect 9428 53375 9496 53404
rect 9552 53375 9620 53404
rect 9676 53375 9744 53404
rect 9800 53375 9867 53404
rect 7817 53323 7844 53375
rect 7940 53348 7952 53375
rect 7896 53323 7952 53348
rect 8004 53348 8008 53375
rect 8112 53348 8132 53375
rect 8220 53348 8256 53375
rect 8328 53348 8380 53375
rect 8004 53323 8060 53348
rect 8112 53323 8168 53348
rect 8220 53323 8276 53348
rect 8328 53323 8384 53348
rect 8436 53323 8492 53375
rect 8560 53348 8600 53375
rect 8684 53348 8708 53375
rect 8808 53348 8816 53375
rect 8544 53323 8600 53348
rect 8652 53323 8708 53348
rect 8760 53323 8816 53348
rect 8868 53348 8876 53375
rect 8976 53348 9000 53375
rect 9084 53348 9124 53375
rect 8868 53323 8924 53348
rect 8976 53323 9032 53348
rect 9084 53323 9140 53348
rect 9192 53323 9248 53375
rect 9304 53348 9356 53375
rect 9428 53348 9464 53375
rect 9552 53348 9572 53375
rect 9676 53348 9680 53375
rect 9300 53323 9356 53348
rect 9408 53323 9464 53348
rect 9516 53323 9572 53348
rect 9624 53323 9680 53348
rect 9732 53348 9744 53375
rect 9732 53323 9788 53348
rect 9840 53323 9867 53375
rect 7817 53280 9867 53323
rect 7817 53267 7884 53280
rect 7940 53267 8008 53280
rect 8064 53267 8132 53280
rect 8188 53267 8256 53280
rect 8312 53267 8380 53280
rect 8436 53267 8504 53280
rect 8560 53267 8628 53280
rect 8684 53267 8752 53280
rect 8808 53267 8876 53280
rect 8932 53267 9000 53280
rect 9056 53267 9124 53280
rect 9180 53267 9248 53280
rect 9304 53267 9372 53280
rect 9428 53267 9496 53280
rect 9552 53267 9620 53280
rect 9676 53267 9744 53280
rect 9800 53267 9867 53280
rect 7817 53215 7844 53267
rect 7940 53224 7952 53267
rect 7896 53215 7952 53224
rect 8004 53224 8008 53267
rect 8112 53224 8132 53267
rect 8220 53224 8256 53267
rect 8328 53224 8380 53267
rect 8004 53215 8060 53224
rect 8112 53215 8168 53224
rect 8220 53215 8276 53224
rect 8328 53215 8384 53224
rect 8436 53215 8492 53267
rect 8560 53224 8600 53267
rect 8684 53224 8708 53267
rect 8808 53224 8816 53267
rect 8544 53215 8600 53224
rect 8652 53215 8708 53224
rect 8760 53215 8816 53224
rect 8868 53224 8876 53267
rect 8976 53224 9000 53267
rect 9084 53224 9124 53267
rect 8868 53215 8924 53224
rect 8976 53215 9032 53224
rect 9084 53215 9140 53224
rect 9192 53215 9248 53267
rect 9304 53224 9356 53267
rect 9428 53224 9464 53267
rect 9552 53224 9572 53267
rect 9676 53224 9680 53267
rect 9300 53215 9356 53224
rect 9408 53215 9464 53224
rect 9516 53215 9572 53224
rect 9624 53215 9680 53224
rect 9732 53224 9744 53267
rect 9732 53215 9788 53224
rect 9840 53215 9867 53267
rect 7817 53156 9867 53215
rect 7817 53100 7884 53156
rect 7940 53100 8008 53156
rect 8064 53100 8132 53156
rect 8188 53100 8256 53156
rect 8312 53100 8380 53156
rect 8436 53100 8504 53156
rect 8560 53100 8628 53156
rect 8684 53100 8752 53156
rect 8808 53100 8876 53156
rect 8932 53100 9000 53156
rect 9056 53100 9124 53156
rect 9180 53100 9248 53156
rect 9304 53100 9372 53156
rect 9428 53100 9496 53156
rect 9552 53100 9620 53156
rect 9676 53100 9744 53156
rect 9800 53100 9867 53156
rect 7817 53032 9867 53100
rect 7817 52976 7884 53032
rect 7940 52976 8008 53032
rect 8064 52976 8132 53032
rect 8188 52976 8256 53032
rect 8312 52976 8380 53032
rect 8436 52976 8504 53032
rect 8560 52976 8628 53032
rect 8684 52976 8752 53032
rect 8808 52976 8876 53032
rect 8932 52976 9000 53032
rect 9056 52976 9124 53032
rect 9180 52976 9248 53032
rect 9304 52976 9372 53032
rect 9428 52976 9496 53032
rect 9552 52976 9620 53032
rect 9676 52976 9744 53032
rect 9800 52976 9867 53032
rect 7817 52908 9867 52976
rect 7817 52852 7884 52908
rect 7940 52852 8008 52908
rect 8064 52852 8132 52908
rect 8188 52852 8256 52908
rect 8312 52852 8380 52908
rect 8436 52852 8504 52908
rect 8560 52852 8628 52908
rect 8684 52852 8752 52908
rect 8808 52852 8876 52908
rect 8932 52852 9000 52908
rect 9056 52852 9124 52908
rect 9180 52852 9248 52908
rect 9304 52852 9372 52908
rect 9428 52852 9496 52908
rect 9552 52852 9620 52908
rect 9676 52852 9744 52908
rect 9800 52852 9867 52908
rect 7817 52548 9867 52852
rect 7817 52492 7884 52548
rect 7940 52492 8008 52548
rect 8064 52492 8132 52548
rect 8188 52492 8256 52548
rect 8312 52492 8380 52548
rect 8436 52492 8504 52548
rect 8560 52492 8628 52548
rect 8684 52492 8752 52548
rect 8808 52492 8876 52548
rect 8932 52492 9000 52548
rect 9056 52492 9124 52548
rect 9180 52492 9248 52548
rect 9304 52492 9372 52548
rect 9428 52492 9496 52548
rect 9552 52492 9620 52548
rect 9676 52492 9744 52548
rect 9800 52492 9867 52548
rect 7817 52424 9867 52492
rect 7817 52368 7884 52424
rect 7940 52368 8008 52424
rect 8064 52368 8132 52424
rect 8188 52368 8256 52424
rect 8312 52368 8380 52424
rect 8436 52368 8504 52424
rect 8560 52368 8628 52424
rect 8684 52368 8752 52424
rect 8808 52368 8876 52424
rect 8932 52368 9000 52424
rect 9056 52368 9124 52424
rect 9180 52368 9248 52424
rect 9304 52368 9372 52424
rect 9428 52368 9496 52424
rect 9552 52368 9620 52424
rect 9676 52368 9744 52424
rect 9800 52368 9867 52424
rect 7817 52300 9867 52368
rect 7817 52244 7884 52300
rect 7940 52244 8008 52300
rect 8064 52244 8132 52300
rect 8188 52244 8256 52300
rect 8312 52244 8380 52300
rect 8436 52244 8504 52300
rect 8560 52244 8628 52300
rect 8684 52244 8752 52300
rect 8808 52244 8876 52300
rect 8932 52244 9000 52300
rect 9056 52244 9124 52300
rect 9180 52244 9248 52300
rect 9304 52244 9372 52300
rect 9428 52244 9496 52300
rect 9552 52244 9620 52300
rect 9676 52244 9744 52300
rect 9800 52244 9867 52300
rect 7817 52176 9867 52244
rect 7817 52120 7884 52176
rect 7940 52120 8008 52176
rect 8064 52120 8132 52176
rect 8188 52120 8256 52176
rect 8312 52120 8380 52176
rect 8436 52120 8504 52176
rect 8560 52120 8628 52176
rect 8684 52120 8752 52176
rect 8808 52120 8876 52176
rect 8932 52120 9000 52176
rect 9056 52120 9124 52176
rect 9180 52120 9248 52176
rect 9304 52120 9372 52176
rect 9428 52120 9496 52176
rect 9552 52120 9620 52176
rect 9676 52120 9744 52176
rect 9800 52120 9867 52176
rect 7817 52052 9867 52120
rect 7817 52009 7884 52052
rect 7940 52009 8008 52052
rect 8064 52009 8132 52052
rect 8188 52009 8256 52052
rect 8312 52009 8380 52052
rect 8436 52009 8504 52052
rect 8560 52009 8628 52052
rect 8684 52009 8752 52052
rect 8808 52009 8876 52052
rect 8932 52009 9000 52052
rect 9056 52009 9124 52052
rect 9180 52009 9248 52052
rect 9304 52009 9372 52052
rect 9428 52009 9496 52052
rect 9552 52009 9620 52052
rect 9676 52009 9744 52052
rect 9800 52009 9867 52052
rect 7817 51957 7844 52009
rect 7940 51996 7952 52009
rect 7896 51957 7952 51996
rect 8004 51996 8008 52009
rect 8112 51996 8132 52009
rect 8220 51996 8256 52009
rect 8328 51996 8380 52009
rect 8004 51957 8060 51996
rect 8112 51957 8168 51996
rect 8220 51957 8276 51996
rect 8328 51957 8384 51996
rect 8436 51957 8492 52009
rect 8560 51996 8600 52009
rect 8684 51996 8708 52009
rect 8808 51996 8816 52009
rect 8544 51957 8600 51996
rect 8652 51957 8708 51996
rect 8760 51957 8816 51996
rect 8868 51996 8876 52009
rect 8976 51996 9000 52009
rect 9084 51996 9124 52009
rect 8868 51957 8924 51996
rect 8976 51957 9032 51996
rect 9084 51957 9140 51996
rect 9192 51957 9248 52009
rect 9304 51996 9356 52009
rect 9428 51996 9464 52009
rect 9552 51996 9572 52009
rect 9676 51996 9680 52009
rect 9300 51957 9356 51996
rect 9408 51957 9464 51996
rect 9516 51957 9572 51996
rect 9624 51957 9680 51996
rect 9732 51996 9744 52009
rect 9732 51957 9788 51996
rect 9840 51957 9867 52009
rect 7817 51928 9867 51957
rect 7817 51901 7884 51928
rect 7940 51901 8008 51928
rect 8064 51901 8132 51928
rect 8188 51901 8256 51928
rect 8312 51901 8380 51928
rect 8436 51901 8504 51928
rect 8560 51901 8628 51928
rect 8684 51901 8752 51928
rect 8808 51901 8876 51928
rect 8932 51901 9000 51928
rect 9056 51901 9124 51928
rect 9180 51901 9248 51928
rect 9304 51901 9372 51928
rect 9428 51901 9496 51928
rect 9552 51901 9620 51928
rect 9676 51901 9744 51928
rect 9800 51901 9867 51928
rect 7817 51849 7844 51901
rect 7940 51872 7952 51901
rect 7896 51849 7952 51872
rect 8004 51872 8008 51901
rect 8112 51872 8132 51901
rect 8220 51872 8256 51901
rect 8328 51872 8380 51901
rect 8004 51849 8060 51872
rect 8112 51849 8168 51872
rect 8220 51849 8276 51872
rect 8328 51849 8384 51872
rect 8436 51849 8492 51901
rect 8560 51872 8600 51901
rect 8684 51872 8708 51901
rect 8808 51872 8816 51901
rect 8544 51849 8600 51872
rect 8652 51849 8708 51872
rect 8760 51849 8816 51872
rect 8868 51872 8876 51901
rect 8976 51872 9000 51901
rect 9084 51872 9124 51901
rect 8868 51849 8924 51872
rect 8976 51849 9032 51872
rect 9084 51849 9140 51872
rect 9192 51849 9248 51901
rect 9304 51872 9356 51901
rect 9428 51872 9464 51901
rect 9552 51872 9572 51901
rect 9676 51872 9680 51901
rect 9300 51849 9356 51872
rect 9408 51849 9464 51872
rect 9516 51849 9572 51872
rect 9624 51849 9680 51872
rect 9732 51872 9744 51901
rect 9732 51849 9788 51872
rect 9840 51849 9867 51901
rect 7817 51804 9867 51849
rect 7817 51748 7884 51804
rect 7940 51748 8008 51804
rect 8064 51748 8132 51804
rect 8188 51748 8256 51804
rect 8312 51748 8380 51804
rect 8436 51748 8504 51804
rect 8560 51748 8628 51804
rect 8684 51748 8752 51804
rect 8808 51748 8876 51804
rect 8932 51748 9000 51804
rect 9056 51748 9124 51804
rect 9180 51748 9248 51804
rect 9304 51748 9372 51804
rect 9428 51748 9496 51804
rect 9552 51748 9620 51804
rect 9676 51748 9744 51804
rect 9800 51748 9867 51804
rect 7817 51680 9867 51748
rect 7817 51624 7884 51680
rect 7940 51624 8008 51680
rect 8064 51624 8132 51680
rect 8188 51624 8256 51680
rect 8312 51624 8380 51680
rect 8436 51624 8504 51680
rect 8560 51624 8628 51680
rect 8684 51624 8752 51680
rect 8808 51624 8876 51680
rect 8932 51624 9000 51680
rect 9056 51624 9124 51680
rect 9180 51624 9248 51680
rect 9304 51624 9372 51680
rect 9428 51624 9496 51680
rect 9552 51624 9620 51680
rect 9676 51624 9744 51680
rect 9800 51624 9867 51680
rect 7817 51556 9867 51624
rect 7817 51500 7884 51556
rect 7940 51500 8008 51556
rect 8064 51500 8132 51556
rect 8188 51500 8256 51556
rect 8312 51500 8380 51556
rect 8436 51500 8504 51556
rect 8560 51500 8628 51556
rect 8684 51500 8752 51556
rect 8808 51500 8876 51556
rect 8932 51500 9000 51556
rect 9056 51500 9124 51556
rect 9180 51500 9248 51556
rect 9304 51500 9372 51556
rect 9428 51500 9496 51556
rect 9552 51500 9620 51556
rect 9676 51500 9744 51556
rect 9800 51500 9867 51556
rect 7817 51432 9867 51500
rect 7817 51376 7884 51432
rect 7940 51376 8008 51432
rect 8064 51376 8132 51432
rect 8188 51376 8256 51432
rect 8312 51376 8380 51432
rect 8436 51376 8504 51432
rect 8560 51376 8628 51432
rect 8684 51376 8752 51432
rect 8808 51376 8876 51432
rect 8932 51376 9000 51432
rect 9056 51376 9124 51432
rect 9180 51376 9248 51432
rect 9304 51376 9372 51432
rect 9428 51376 9496 51432
rect 9552 51376 9620 51432
rect 9676 51376 9744 51432
rect 9800 51376 9867 51432
rect 7817 51308 9867 51376
rect 7817 51252 7884 51308
rect 7940 51252 8008 51308
rect 8064 51252 8132 51308
rect 8188 51252 8256 51308
rect 8312 51252 8380 51308
rect 8436 51252 8504 51308
rect 8560 51252 8628 51308
rect 8684 51252 8752 51308
rect 8808 51252 8876 51308
rect 8932 51252 9000 51308
rect 9056 51252 9124 51308
rect 9180 51252 9248 51308
rect 9304 51252 9372 51308
rect 9428 51252 9496 51308
rect 9552 51252 9620 51308
rect 9676 51252 9744 51308
rect 9800 51252 9867 51308
rect 7817 51206 9867 51252
rect 7817 51154 7844 51206
rect 7896 51154 7952 51206
rect 8004 51154 8060 51206
rect 8112 51154 8168 51206
rect 8220 51154 8276 51206
rect 8328 51154 8384 51206
rect 8436 51154 8492 51206
rect 8544 51154 8600 51206
rect 8652 51154 8708 51206
rect 8760 51154 8816 51206
rect 8868 51154 8924 51206
rect 8976 51154 9032 51206
rect 9084 51154 9140 51206
rect 9192 51154 9248 51206
rect 9300 51154 9356 51206
rect 9408 51154 9464 51206
rect 9516 51154 9572 51206
rect 9624 51154 9680 51206
rect 9732 51154 9788 51206
rect 9840 51154 9867 51206
rect 7817 51098 9867 51154
rect 7817 51046 7844 51098
rect 7896 51046 7952 51098
rect 8004 51046 8060 51098
rect 8112 51046 8168 51098
rect 8220 51046 8276 51098
rect 8328 51046 8384 51098
rect 8436 51046 8492 51098
rect 8544 51046 8600 51098
rect 8652 51046 8708 51098
rect 8760 51046 8816 51098
rect 8868 51046 8924 51098
rect 8976 51046 9032 51098
rect 9084 51046 9140 51098
rect 9192 51046 9248 51098
rect 9300 51046 9356 51098
rect 9408 51046 9464 51098
rect 9516 51046 9572 51098
rect 9624 51046 9680 51098
rect 9732 51046 9788 51098
rect 9840 51046 9867 51098
rect 7817 50990 9867 51046
rect 7817 50938 7844 50990
rect 7896 50938 7952 50990
rect 8004 50938 8060 50990
rect 8112 50938 8168 50990
rect 8220 50938 8276 50990
rect 8328 50938 8384 50990
rect 8436 50938 8492 50990
rect 8544 50938 8600 50990
rect 8652 50938 8708 50990
rect 8760 50938 8816 50990
rect 8868 50938 8924 50990
rect 8976 50938 9032 50990
rect 9084 50938 9140 50990
rect 9192 50938 9248 50990
rect 9300 50938 9356 50990
rect 9408 50938 9464 50990
rect 9516 50938 9572 50990
rect 9624 50938 9680 50990
rect 9732 50938 9788 50990
rect 9840 50938 9867 50990
rect 7817 50272 9867 50938
rect 7817 50220 7844 50272
rect 7896 50220 7952 50272
rect 8004 50220 8060 50272
rect 8112 50220 8168 50272
rect 8220 50220 8276 50272
rect 8328 50220 8384 50272
rect 8436 50220 8492 50272
rect 8544 50220 8600 50272
rect 8652 50220 8708 50272
rect 8760 50220 8816 50272
rect 8868 50220 8924 50272
rect 8976 50220 9032 50272
rect 9084 50220 9140 50272
rect 9192 50220 9248 50272
rect 9300 50220 9356 50272
rect 9408 50220 9464 50272
rect 9516 50220 9572 50272
rect 9624 50220 9680 50272
rect 9732 50220 9788 50272
rect 9840 50220 9867 50272
rect 7817 50164 9867 50220
rect 7817 50112 7844 50164
rect 7896 50112 7952 50164
rect 8004 50112 8060 50164
rect 8112 50112 8168 50164
rect 8220 50112 8276 50164
rect 8328 50112 8384 50164
rect 8436 50112 8492 50164
rect 8544 50112 8600 50164
rect 8652 50112 8708 50164
rect 8760 50112 8816 50164
rect 8868 50112 8924 50164
rect 8976 50112 9032 50164
rect 9084 50112 9140 50164
rect 9192 50112 9248 50164
rect 9300 50112 9356 50164
rect 9408 50112 9464 50164
rect 9516 50112 9572 50164
rect 9624 50112 9680 50164
rect 9732 50112 9788 50164
rect 9840 50112 9867 50164
rect 7817 50056 9867 50112
rect 7817 50004 7844 50056
rect 7896 50004 7952 50056
rect 8004 50004 8060 50056
rect 8112 50004 8168 50056
rect 8220 50004 8276 50056
rect 8328 50004 8384 50056
rect 8436 50004 8492 50056
rect 8544 50004 8600 50056
rect 8652 50004 8708 50056
rect 8760 50004 8816 50056
rect 8868 50004 8924 50056
rect 8976 50004 9032 50056
rect 9084 50004 9140 50056
rect 9192 50004 9248 50056
rect 9300 50004 9356 50056
rect 9408 50004 9464 50056
rect 9516 50004 9572 50056
rect 9624 50004 9680 50056
rect 9732 50004 9788 50056
rect 9840 50004 9867 50056
rect 7817 49348 9867 50004
rect 7817 49338 7884 49348
rect 7940 49338 8008 49348
rect 8064 49338 8132 49348
rect 8188 49338 8256 49348
rect 8312 49338 8380 49348
rect 8436 49338 8504 49348
rect 8560 49338 8628 49348
rect 8684 49338 8752 49348
rect 8808 49338 8876 49348
rect 8932 49338 9000 49348
rect 9056 49338 9124 49348
rect 9180 49338 9248 49348
rect 9304 49338 9372 49348
rect 9428 49338 9496 49348
rect 9552 49338 9620 49348
rect 9676 49338 9744 49348
rect 9800 49338 9867 49348
rect 7817 49286 7844 49338
rect 7940 49292 7952 49338
rect 7896 49286 7952 49292
rect 8004 49292 8008 49338
rect 8112 49292 8132 49338
rect 8220 49292 8256 49338
rect 8328 49292 8380 49338
rect 8004 49286 8060 49292
rect 8112 49286 8168 49292
rect 8220 49286 8276 49292
rect 8328 49286 8384 49292
rect 8436 49286 8492 49338
rect 8560 49292 8600 49338
rect 8684 49292 8708 49338
rect 8808 49292 8816 49338
rect 8544 49286 8600 49292
rect 8652 49286 8708 49292
rect 8760 49286 8816 49292
rect 8868 49292 8876 49338
rect 8976 49292 9000 49338
rect 9084 49292 9124 49338
rect 8868 49286 8924 49292
rect 8976 49286 9032 49292
rect 9084 49286 9140 49292
rect 9192 49286 9248 49338
rect 9304 49292 9356 49338
rect 9428 49292 9464 49338
rect 9552 49292 9572 49338
rect 9676 49292 9680 49338
rect 9300 49286 9356 49292
rect 9408 49286 9464 49292
rect 9516 49286 9572 49292
rect 9624 49286 9680 49292
rect 9732 49292 9744 49338
rect 9732 49286 9788 49292
rect 9840 49286 9867 49338
rect 7817 49230 9867 49286
rect 7817 49178 7844 49230
rect 7896 49224 7952 49230
rect 7940 49178 7952 49224
rect 8004 49224 8060 49230
rect 8112 49224 8168 49230
rect 8220 49224 8276 49230
rect 8328 49224 8384 49230
rect 8004 49178 8008 49224
rect 8112 49178 8132 49224
rect 8220 49178 8256 49224
rect 8328 49178 8380 49224
rect 8436 49178 8492 49230
rect 8544 49224 8600 49230
rect 8652 49224 8708 49230
rect 8760 49224 8816 49230
rect 8560 49178 8600 49224
rect 8684 49178 8708 49224
rect 8808 49178 8816 49224
rect 8868 49224 8924 49230
rect 8976 49224 9032 49230
rect 9084 49224 9140 49230
rect 8868 49178 8876 49224
rect 8976 49178 9000 49224
rect 9084 49178 9124 49224
rect 9192 49178 9248 49230
rect 9300 49224 9356 49230
rect 9408 49224 9464 49230
rect 9516 49224 9572 49230
rect 9624 49224 9680 49230
rect 9304 49178 9356 49224
rect 9428 49178 9464 49224
rect 9552 49178 9572 49224
rect 9676 49178 9680 49224
rect 9732 49224 9788 49230
rect 9732 49178 9744 49224
rect 9840 49178 9867 49230
rect 7817 49168 7884 49178
rect 7940 49168 8008 49178
rect 8064 49168 8132 49178
rect 8188 49168 8256 49178
rect 8312 49168 8380 49178
rect 8436 49168 8504 49178
rect 8560 49168 8628 49178
rect 8684 49168 8752 49178
rect 8808 49168 8876 49178
rect 8932 49168 9000 49178
rect 9056 49168 9124 49178
rect 9180 49168 9248 49178
rect 9304 49168 9372 49178
rect 9428 49168 9496 49178
rect 9552 49168 9620 49178
rect 9676 49168 9744 49178
rect 9800 49168 9867 49178
rect 7817 49122 9867 49168
rect 7817 49070 7844 49122
rect 7896 49100 7952 49122
rect 7940 49070 7952 49100
rect 8004 49100 8060 49122
rect 8112 49100 8168 49122
rect 8220 49100 8276 49122
rect 8328 49100 8384 49122
rect 8004 49070 8008 49100
rect 8112 49070 8132 49100
rect 8220 49070 8256 49100
rect 8328 49070 8380 49100
rect 8436 49070 8492 49122
rect 8544 49100 8600 49122
rect 8652 49100 8708 49122
rect 8760 49100 8816 49122
rect 8560 49070 8600 49100
rect 8684 49070 8708 49100
rect 8808 49070 8816 49100
rect 8868 49100 8924 49122
rect 8976 49100 9032 49122
rect 9084 49100 9140 49122
rect 8868 49070 8876 49100
rect 8976 49070 9000 49100
rect 9084 49070 9124 49100
rect 9192 49070 9248 49122
rect 9300 49100 9356 49122
rect 9408 49100 9464 49122
rect 9516 49100 9572 49122
rect 9624 49100 9680 49122
rect 9304 49070 9356 49100
rect 9428 49070 9464 49100
rect 9552 49070 9572 49100
rect 9676 49070 9680 49100
rect 9732 49100 9788 49122
rect 9732 49070 9744 49100
rect 9840 49070 9867 49122
rect 7817 49044 7884 49070
rect 7940 49044 8008 49070
rect 8064 49044 8132 49070
rect 8188 49044 8256 49070
rect 8312 49044 8380 49070
rect 8436 49044 8504 49070
rect 8560 49044 8628 49070
rect 8684 49044 8752 49070
rect 8808 49044 8876 49070
rect 8932 49044 9000 49070
rect 9056 49044 9124 49070
rect 9180 49044 9248 49070
rect 9304 49044 9372 49070
rect 9428 49044 9496 49070
rect 9552 49044 9620 49070
rect 9676 49044 9744 49070
rect 9800 49044 9867 49070
rect 7817 48976 9867 49044
rect 7817 48920 7884 48976
rect 7940 48920 8008 48976
rect 8064 48920 8132 48976
rect 8188 48920 8256 48976
rect 8312 48920 8380 48976
rect 8436 48920 8504 48976
rect 8560 48920 8628 48976
rect 8684 48920 8752 48976
rect 8808 48920 8876 48976
rect 8932 48920 9000 48976
rect 9056 48920 9124 48976
rect 9180 48920 9248 48976
rect 9304 48920 9372 48976
rect 9428 48920 9496 48976
rect 9552 48920 9620 48976
rect 9676 48920 9744 48976
rect 9800 48920 9867 48976
rect 7817 48852 9867 48920
rect 7817 48796 7884 48852
rect 7940 48796 8008 48852
rect 8064 48796 8132 48852
rect 8188 48796 8256 48852
rect 8312 48796 8380 48852
rect 8436 48796 8504 48852
rect 8560 48796 8628 48852
rect 8684 48796 8752 48852
rect 8808 48796 8876 48852
rect 8932 48796 9000 48852
rect 9056 48796 9124 48852
rect 9180 48796 9248 48852
rect 9304 48796 9372 48852
rect 9428 48796 9496 48852
rect 9552 48796 9620 48852
rect 9676 48796 9744 48852
rect 9800 48796 9867 48852
rect 7817 48728 9867 48796
rect 7817 48672 7884 48728
rect 7940 48672 8008 48728
rect 8064 48672 8132 48728
rect 8188 48672 8256 48728
rect 8312 48672 8380 48728
rect 8436 48672 8504 48728
rect 8560 48672 8628 48728
rect 8684 48672 8752 48728
rect 8808 48672 8876 48728
rect 8932 48672 9000 48728
rect 9056 48672 9124 48728
rect 9180 48672 9248 48728
rect 9304 48672 9372 48728
rect 9428 48672 9496 48728
rect 9552 48672 9620 48728
rect 9676 48672 9744 48728
rect 9800 48672 9867 48728
rect 7817 48604 9867 48672
rect 7817 48548 7884 48604
rect 7940 48548 8008 48604
rect 8064 48548 8132 48604
rect 8188 48548 8256 48604
rect 8312 48548 8380 48604
rect 8436 48548 8504 48604
rect 8560 48548 8628 48604
rect 8684 48548 8752 48604
rect 8808 48548 8876 48604
rect 8932 48548 9000 48604
rect 9056 48548 9124 48604
rect 9180 48548 9248 48604
rect 9304 48548 9372 48604
rect 9428 48548 9496 48604
rect 9552 48548 9620 48604
rect 9676 48548 9744 48604
rect 9800 48548 9867 48604
rect 7817 48480 9867 48548
rect 7817 48427 7884 48480
rect 7940 48427 8008 48480
rect 8064 48427 8132 48480
rect 8188 48427 8256 48480
rect 8312 48427 8380 48480
rect 8436 48427 8504 48480
rect 8560 48427 8628 48480
rect 8684 48427 8752 48480
rect 8808 48427 8876 48480
rect 8932 48427 9000 48480
rect 9056 48427 9124 48480
rect 9180 48427 9248 48480
rect 9304 48427 9372 48480
rect 9428 48427 9496 48480
rect 9552 48427 9620 48480
rect 9676 48427 9744 48480
rect 9800 48427 9867 48480
rect 7817 48375 7844 48427
rect 7940 48424 7952 48427
rect 7896 48375 7952 48424
rect 8004 48424 8008 48427
rect 8112 48424 8132 48427
rect 8220 48424 8256 48427
rect 8328 48424 8380 48427
rect 8004 48375 8060 48424
rect 8112 48375 8168 48424
rect 8220 48375 8276 48424
rect 8328 48375 8384 48424
rect 8436 48375 8492 48427
rect 8560 48424 8600 48427
rect 8684 48424 8708 48427
rect 8808 48424 8816 48427
rect 8544 48375 8600 48424
rect 8652 48375 8708 48424
rect 8760 48375 8816 48424
rect 8868 48424 8876 48427
rect 8976 48424 9000 48427
rect 9084 48424 9124 48427
rect 8868 48375 8924 48424
rect 8976 48375 9032 48424
rect 9084 48375 9140 48424
rect 9192 48375 9248 48427
rect 9304 48424 9356 48427
rect 9428 48424 9464 48427
rect 9552 48424 9572 48427
rect 9676 48424 9680 48427
rect 9300 48375 9356 48424
rect 9408 48375 9464 48424
rect 9516 48375 9572 48424
rect 9624 48375 9680 48424
rect 9732 48424 9744 48427
rect 9732 48375 9788 48424
rect 9840 48375 9867 48427
rect 7817 48356 9867 48375
rect 7817 48319 7884 48356
rect 7940 48319 8008 48356
rect 8064 48319 8132 48356
rect 8188 48319 8256 48356
rect 8312 48319 8380 48356
rect 8436 48319 8504 48356
rect 8560 48319 8628 48356
rect 8684 48319 8752 48356
rect 8808 48319 8876 48356
rect 8932 48319 9000 48356
rect 9056 48319 9124 48356
rect 9180 48319 9248 48356
rect 9304 48319 9372 48356
rect 9428 48319 9496 48356
rect 9552 48319 9620 48356
rect 9676 48319 9744 48356
rect 9800 48319 9867 48356
rect 7817 48267 7844 48319
rect 7940 48300 7952 48319
rect 7896 48267 7952 48300
rect 8004 48300 8008 48319
rect 8112 48300 8132 48319
rect 8220 48300 8256 48319
rect 8328 48300 8380 48319
rect 8004 48267 8060 48300
rect 8112 48267 8168 48300
rect 8220 48267 8276 48300
rect 8328 48267 8384 48300
rect 8436 48267 8492 48319
rect 8560 48300 8600 48319
rect 8684 48300 8708 48319
rect 8808 48300 8816 48319
rect 8544 48267 8600 48300
rect 8652 48267 8708 48300
rect 8760 48267 8816 48300
rect 8868 48300 8876 48319
rect 8976 48300 9000 48319
rect 9084 48300 9124 48319
rect 8868 48267 8924 48300
rect 8976 48267 9032 48300
rect 9084 48267 9140 48300
rect 9192 48267 9248 48319
rect 9304 48300 9356 48319
rect 9428 48300 9464 48319
rect 9552 48300 9572 48319
rect 9676 48300 9680 48319
rect 9300 48267 9356 48300
rect 9408 48267 9464 48300
rect 9516 48267 9572 48300
rect 9624 48267 9680 48300
rect 9732 48300 9744 48319
rect 9732 48267 9788 48300
rect 9840 48267 9867 48319
rect 7817 48232 9867 48267
rect 7817 48176 7884 48232
rect 7940 48176 8008 48232
rect 8064 48176 8132 48232
rect 8188 48176 8256 48232
rect 8312 48176 8380 48232
rect 8436 48176 8504 48232
rect 8560 48176 8628 48232
rect 8684 48176 8752 48232
rect 8808 48176 8876 48232
rect 8932 48176 9000 48232
rect 9056 48176 9124 48232
rect 9180 48176 9248 48232
rect 9304 48176 9372 48232
rect 9428 48176 9496 48232
rect 9552 48176 9620 48232
rect 9676 48176 9744 48232
rect 9800 48176 9867 48232
rect 7817 48108 9867 48176
rect 7817 48052 7884 48108
rect 7940 48052 8008 48108
rect 8064 48052 8132 48108
rect 8188 48052 8256 48108
rect 8312 48052 8380 48108
rect 8436 48052 8504 48108
rect 8560 48052 8628 48108
rect 8684 48052 8752 48108
rect 8808 48052 8876 48108
rect 8932 48052 9000 48108
rect 9056 48052 9124 48108
rect 9180 48052 9248 48108
rect 9304 48052 9372 48108
rect 9428 48052 9496 48108
rect 9552 48052 9620 48108
rect 9676 48052 9744 48108
rect 9800 48052 9867 48108
rect 7817 47163 9867 48052
rect 9927 56693 10127 57278
rect 9927 56641 9947 56693
rect 9999 56641 10055 56693
rect 10107 56641 10127 56693
rect 9927 56585 10127 56641
rect 9927 56533 9947 56585
rect 9999 56533 10055 56585
rect 10107 56533 10127 56585
rect 9927 56477 10127 56533
rect 9927 56425 9947 56477
rect 9999 56425 10055 56477
rect 10107 56425 10127 56477
rect 9927 56369 10127 56425
rect 9927 56317 9947 56369
rect 9999 56317 10055 56369
rect 10107 56317 10127 56369
rect 9927 56261 10127 56317
rect 9927 56209 9947 56261
rect 9999 56209 10055 56261
rect 10107 56209 10127 56261
rect 9927 56153 10127 56209
rect 9927 56101 9947 56153
rect 9999 56101 10055 56153
rect 10107 56101 10127 56153
rect 9927 56045 10127 56101
rect 9927 55993 9947 56045
rect 9999 55993 10055 56045
rect 10107 55993 10127 56045
rect 9927 55937 10127 55993
rect 9927 55885 9947 55937
rect 9999 55885 10055 55937
rect 10107 55885 10127 55937
rect 9927 55829 10127 55885
rect 9927 55777 9947 55829
rect 9999 55777 10055 55829
rect 10107 55777 10127 55829
rect 9927 55748 10127 55777
rect 9927 55692 9937 55748
rect 9993 55721 10061 55748
rect 9927 55669 9947 55692
rect 9999 55669 10055 55721
rect 10117 55692 10127 55748
rect 10107 55669 10127 55692
rect 9927 55624 10127 55669
rect 9927 55568 9937 55624
rect 9993 55613 10061 55624
rect 9927 55561 9947 55568
rect 9999 55561 10055 55613
rect 10117 55568 10127 55624
rect 10107 55561 10127 55568
rect 9927 55505 10127 55561
rect 9927 55500 9947 55505
rect 9927 55444 9937 55500
rect 9999 55453 10055 55505
rect 10107 55500 10127 55505
rect 9993 55444 10061 55453
rect 10117 55444 10127 55500
rect 9927 55397 10127 55444
rect 9927 55376 9947 55397
rect 9927 55320 9937 55376
rect 9999 55345 10055 55397
rect 10107 55376 10127 55397
rect 9993 55320 10061 55345
rect 10117 55320 10127 55376
rect 9927 55289 10127 55320
rect 9927 55252 9947 55289
rect 9927 55196 9937 55252
rect 9999 55237 10055 55289
rect 10107 55252 10127 55289
rect 9993 55196 10061 55237
rect 10117 55196 10127 55252
rect 9927 55181 10127 55196
rect 9927 55129 9947 55181
rect 9999 55129 10055 55181
rect 10107 55129 10127 55181
rect 9927 55128 10127 55129
rect 9927 55072 9937 55128
rect 9993 55073 10061 55128
rect 9927 55021 9947 55072
rect 9999 55021 10055 55073
rect 10117 55072 10127 55128
rect 10107 55021 10127 55072
rect 9927 55004 10127 55021
rect 9927 54948 9937 55004
rect 9993 54965 10061 55004
rect 9927 54913 9947 54948
rect 9999 54913 10055 54965
rect 10117 54948 10127 55004
rect 10107 54913 10127 54948
rect 9927 54880 10127 54913
rect 9927 54824 9937 54880
rect 9993 54857 10061 54880
rect 9927 54805 9947 54824
rect 9999 54805 10055 54857
rect 10117 54824 10127 54880
rect 10107 54805 10127 54824
rect 9927 54756 10127 54805
rect 9927 54700 9937 54756
rect 9993 54749 10061 54756
rect 9927 54697 9947 54700
rect 9999 54697 10055 54749
rect 10117 54700 10127 54756
rect 10107 54697 10127 54700
rect 9927 54641 10127 54697
rect 9927 54632 9947 54641
rect 9927 54576 9937 54632
rect 9999 54589 10055 54641
rect 10107 54632 10127 54641
rect 9993 54576 10061 54589
rect 10117 54576 10127 54632
rect 9927 54533 10127 54576
rect 9927 54508 9947 54533
rect 9927 54452 9937 54508
rect 9999 54481 10055 54533
rect 10107 54508 10127 54533
rect 9993 54452 10061 54481
rect 10117 54452 10127 54508
rect 9927 54425 10127 54452
rect 9927 54373 9947 54425
rect 9999 54373 10055 54425
rect 10107 54373 10127 54425
rect 9927 54317 10127 54373
rect 9927 54265 9947 54317
rect 9999 54265 10055 54317
rect 10107 54265 10127 54317
rect 9927 54209 10127 54265
rect 9927 54157 9947 54209
rect 9999 54157 10055 54209
rect 10107 54157 10127 54209
rect 9927 54101 10127 54157
rect 9927 54049 9947 54101
rect 9999 54049 10055 54101
rect 10107 54049 10127 54101
rect 9927 53993 10127 54049
rect 9927 53941 9947 53993
rect 9999 53941 10055 53993
rect 10107 53941 10127 53993
rect 9927 53885 10127 53941
rect 9927 53833 9947 53885
rect 9999 53833 10055 53885
rect 10107 53833 10127 53885
rect 9927 53777 10127 53833
rect 9927 53725 9947 53777
rect 9999 53725 10055 53777
rect 10107 53725 10127 53777
rect 9927 53669 10127 53725
rect 9927 53617 9947 53669
rect 9999 53617 10055 53669
rect 10107 53617 10127 53669
rect 9927 52572 10127 53617
rect 9927 52520 9947 52572
rect 9999 52520 10055 52572
rect 10107 52520 10127 52572
rect 9927 52464 10127 52520
rect 9927 52412 9947 52464
rect 9999 52412 10055 52464
rect 10107 52412 10127 52464
rect 9927 52356 10127 52412
rect 9927 52304 9947 52356
rect 9999 52304 10055 52356
rect 10107 52304 10127 52356
rect 9927 51619 10127 52304
rect 9927 51567 9947 51619
rect 9999 51567 10055 51619
rect 10107 51567 10127 51619
rect 9927 51511 10127 51567
rect 9927 51459 9947 51511
rect 9999 51459 10055 51511
rect 10107 51459 10127 51511
rect 9927 50685 10127 51459
rect 9927 50633 9947 50685
rect 9999 50633 10055 50685
rect 10107 50633 10127 50685
rect 9927 50577 10127 50633
rect 9927 50525 9947 50577
rect 9999 50525 10055 50577
rect 10107 50525 10127 50577
rect 9927 49751 10127 50525
rect 9927 49699 9947 49751
rect 9999 49699 10055 49751
rect 10107 49699 10127 49751
rect 9927 49643 10127 49699
rect 9927 49591 9947 49643
rect 9999 49591 10055 49643
rect 10107 49591 10127 49643
rect 9927 48817 10127 49591
rect 9927 48765 9947 48817
rect 9999 48765 10055 48817
rect 10107 48765 10127 48817
rect 9927 48709 10127 48765
rect 9927 48657 9947 48709
rect 9999 48657 10055 48709
rect 10107 48657 10127 48709
rect 9927 47972 10127 48657
rect 9927 47920 9947 47972
rect 9999 47920 10055 47972
rect 10107 47920 10127 47972
rect 9927 47864 10127 47920
rect 9927 47812 9947 47864
rect 9999 47812 10055 47864
rect 10107 47812 10127 47864
rect 9927 47756 10127 47812
rect 9927 47748 9947 47756
rect 9927 47692 9937 47748
rect 9999 47704 10055 47756
rect 10107 47748 10127 47756
rect 9993 47692 10061 47704
rect 10117 47692 10127 47748
rect 9927 47624 10127 47692
rect 9927 47568 9937 47624
rect 9993 47568 10061 47624
rect 10117 47568 10127 47624
rect 9927 47500 10127 47568
rect 9927 47444 9937 47500
rect 9993 47444 10061 47500
rect 10117 47444 10127 47500
rect 9927 47376 10127 47444
rect 9927 47320 9937 47376
rect 9993 47320 10061 47376
rect 10117 47320 10127 47376
rect 9927 47252 10127 47320
rect 9927 47196 9937 47252
rect 9993 47196 10061 47252
rect 10117 47196 10127 47252
rect 4851 47072 4861 47128
rect 4917 47072 4985 47128
rect 5041 47072 5051 47128
rect 4851 47004 5051 47072
rect 4851 46948 4861 47004
rect 4917 46948 4985 47004
rect 5041 46948 5051 47004
rect 4851 46880 5051 46948
rect 4851 46824 4861 46880
rect 4917 46824 4985 46880
rect 5041 46824 5051 46880
rect 4851 46756 5051 46824
rect 4851 46700 4861 46756
rect 4917 46700 4985 46756
rect 5041 46700 5051 46756
rect 4851 46632 5051 46700
rect 4851 46576 4861 46632
rect 4917 46576 4985 46632
rect 5041 46576 5051 46632
rect 4851 46508 5051 46576
rect 4851 46452 4861 46508
rect 4917 46452 4985 46508
rect 5041 46452 5051 46508
rect 4851 46442 5051 46452
rect 7265 47128 7713 47163
rect 7265 47072 7275 47128
rect 7331 47072 7399 47128
rect 7455 47072 7523 47128
rect 7579 47072 7647 47128
rect 7703 47072 7713 47128
rect 7265 47004 7713 47072
rect 7265 46948 7275 47004
rect 7331 46948 7399 47004
rect 7455 46948 7523 47004
rect 7579 46948 7647 47004
rect 7703 46948 7713 47004
rect 7265 46880 7713 46948
rect 7265 46824 7275 46880
rect 7331 46824 7399 46880
rect 7455 46824 7523 46880
rect 7579 46824 7647 46880
rect 7703 46824 7713 46880
rect 7265 46756 7713 46824
rect 7265 46700 7275 46756
rect 7331 46700 7399 46756
rect 7455 46700 7523 46756
rect 7579 46700 7647 46756
rect 7703 46700 7713 46756
rect 7265 46632 7713 46700
rect 7265 46576 7275 46632
rect 7331 46576 7399 46632
rect 7455 46576 7523 46632
rect 7579 46576 7647 46632
rect 7703 46576 7713 46632
rect 7265 46508 7713 46576
rect 7265 46452 7275 46508
rect 7331 46452 7399 46508
rect 7455 46452 7523 46508
rect 7579 46452 7647 46508
rect 7703 46452 7713 46508
rect 7265 46442 7713 46452
rect 9927 47128 10127 47196
rect 10187 57225 12237 57447
rect 12817 57499 14717 57600
rect 12817 57447 12877 57499
rect 12929 57447 12985 57499
rect 13037 57447 13093 57499
rect 13145 57447 13201 57499
rect 13253 57447 13309 57499
rect 13361 57447 13417 57499
rect 13469 57447 13525 57499
rect 13577 57447 13633 57499
rect 13685 57447 13741 57499
rect 13793 57447 13849 57499
rect 13901 57447 13957 57499
rect 14009 57447 14065 57499
rect 14117 57447 14173 57499
rect 14225 57447 14281 57499
rect 14333 57447 14389 57499
rect 14441 57447 14497 57499
rect 14549 57447 14605 57499
rect 14657 57447 14717 57499
rect 10187 57169 10254 57225
rect 10310 57169 10378 57225
rect 10434 57169 10502 57225
rect 10558 57169 10626 57225
rect 10682 57169 10750 57225
rect 10806 57169 10874 57225
rect 10930 57169 10998 57225
rect 11054 57169 11122 57225
rect 11178 57169 11246 57225
rect 11302 57169 11370 57225
rect 11426 57169 11494 57225
rect 11550 57169 11618 57225
rect 11674 57169 11742 57225
rect 11798 57169 11866 57225
rect 11922 57169 11990 57225
rect 12046 57169 12114 57225
rect 12170 57169 12237 57225
rect 10187 57104 12237 57169
rect 10187 57052 10214 57104
rect 10266 57101 10322 57104
rect 10310 57052 10322 57101
rect 10374 57101 10430 57104
rect 10482 57101 10538 57104
rect 10590 57101 10646 57104
rect 10698 57101 10754 57104
rect 10374 57052 10378 57101
rect 10482 57052 10502 57101
rect 10590 57052 10626 57101
rect 10698 57052 10750 57101
rect 10806 57052 10862 57104
rect 10914 57101 10970 57104
rect 11022 57101 11078 57104
rect 11130 57101 11186 57104
rect 10930 57052 10970 57101
rect 11054 57052 11078 57101
rect 11178 57052 11186 57101
rect 11238 57101 11294 57104
rect 11346 57101 11402 57104
rect 11454 57101 11510 57104
rect 11238 57052 11246 57101
rect 11346 57052 11370 57101
rect 11454 57052 11494 57101
rect 11562 57052 11618 57104
rect 11670 57101 11726 57104
rect 11778 57101 11834 57104
rect 11886 57101 11942 57104
rect 11994 57101 12050 57104
rect 11674 57052 11726 57101
rect 11798 57052 11834 57101
rect 11922 57052 11942 57101
rect 12046 57052 12050 57101
rect 12102 57101 12158 57104
rect 12102 57052 12114 57101
rect 12210 57052 12237 57104
rect 10187 57045 10254 57052
rect 10310 57045 10378 57052
rect 10434 57045 10502 57052
rect 10558 57045 10626 57052
rect 10682 57045 10750 57052
rect 10806 57045 10874 57052
rect 10930 57045 10998 57052
rect 11054 57045 11122 57052
rect 11178 57045 11246 57052
rect 11302 57045 11370 57052
rect 11426 57045 11494 57052
rect 11550 57045 11618 57052
rect 11674 57045 11742 57052
rect 11798 57045 11866 57052
rect 11922 57045 11990 57052
rect 12046 57045 12114 57052
rect 12170 57045 12237 57052
rect 10187 56977 12237 57045
rect 10187 56921 10254 56977
rect 10310 56921 10378 56977
rect 10434 56921 10502 56977
rect 10558 56921 10626 56977
rect 10682 56921 10750 56977
rect 10806 56921 10874 56977
rect 10930 56921 10998 56977
rect 11054 56921 11122 56977
rect 11178 56921 11246 56977
rect 11302 56921 11370 56977
rect 11426 56921 11494 56977
rect 11550 56921 11618 56977
rect 11674 56921 11742 56977
rect 11798 56921 11866 56977
rect 11922 56921 11990 56977
rect 12046 56921 12114 56977
rect 12170 56921 12237 56977
rect 10187 56853 12237 56921
rect 10187 56797 10254 56853
rect 10310 56797 10378 56853
rect 10434 56797 10502 56853
rect 10558 56797 10626 56853
rect 10682 56797 10750 56853
rect 10806 56797 10874 56853
rect 10930 56797 10998 56853
rect 11054 56797 11122 56853
rect 11178 56797 11246 56853
rect 11302 56797 11370 56853
rect 11426 56797 11494 56853
rect 11550 56797 11618 56853
rect 11674 56797 11742 56853
rect 11798 56797 11866 56853
rect 11922 56797 11990 56853
rect 12046 56797 12114 56853
rect 12170 56797 12237 56853
rect 10187 56729 12237 56797
rect 10187 56673 10254 56729
rect 10310 56673 10378 56729
rect 10434 56673 10502 56729
rect 10558 56673 10626 56729
rect 10682 56673 10750 56729
rect 10806 56673 10874 56729
rect 10930 56673 10998 56729
rect 11054 56673 11122 56729
rect 11178 56673 11246 56729
rect 11302 56673 11370 56729
rect 11426 56673 11494 56729
rect 11550 56673 11618 56729
rect 11674 56673 11742 56729
rect 11798 56673 11866 56729
rect 11922 56673 11990 56729
rect 12046 56673 12114 56729
rect 12170 56673 12237 56729
rect 10187 56643 12237 56673
rect 10187 56605 10775 56643
rect 10827 56605 10899 56643
rect 10951 56605 11023 56643
rect 11075 56605 12237 56643
rect 10187 56549 10254 56605
rect 10310 56549 10378 56605
rect 10434 56549 10502 56605
rect 10558 56549 10626 56605
rect 10682 56549 10750 56605
rect 10827 56591 10874 56605
rect 10951 56591 10998 56605
rect 11075 56591 11122 56605
rect 10806 56549 10874 56591
rect 10930 56549 10998 56591
rect 11054 56549 11122 56591
rect 11178 56549 11246 56605
rect 11302 56549 11370 56605
rect 11426 56549 11494 56605
rect 11550 56549 11618 56605
rect 11674 56549 11742 56605
rect 11798 56549 11866 56605
rect 11922 56549 11990 56605
rect 12046 56549 12114 56605
rect 12170 56549 12237 56605
rect 10187 56519 12237 56549
rect 10187 56481 10775 56519
rect 10827 56481 10899 56519
rect 10951 56481 11023 56519
rect 11075 56481 12237 56519
rect 10187 56425 10254 56481
rect 10310 56425 10378 56481
rect 10434 56425 10502 56481
rect 10558 56425 10626 56481
rect 10682 56425 10750 56481
rect 10827 56467 10874 56481
rect 10951 56467 10998 56481
rect 11075 56467 11122 56481
rect 10806 56425 10874 56467
rect 10930 56425 10998 56467
rect 11054 56425 11122 56467
rect 11178 56425 11246 56481
rect 11302 56425 11370 56481
rect 11426 56425 11494 56481
rect 11550 56425 11618 56481
rect 11674 56425 11742 56481
rect 11798 56425 11866 56481
rect 11922 56425 11990 56481
rect 12046 56425 12114 56481
rect 12170 56425 12237 56481
rect 10187 56395 12237 56425
rect 10187 56357 10775 56395
rect 10827 56357 10899 56395
rect 10951 56357 11023 56395
rect 11075 56357 12237 56395
rect 10187 56301 10254 56357
rect 10310 56301 10378 56357
rect 10434 56301 10502 56357
rect 10558 56301 10626 56357
rect 10682 56301 10750 56357
rect 10827 56343 10874 56357
rect 10951 56343 10998 56357
rect 11075 56343 11122 56357
rect 10806 56301 10874 56343
rect 10930 56301 10998 56343
rect 11054 56301 11122 56343
rect 11178 56301 11246 56357
rect 11302 56301 11370 56357
rect 11426 56301 11494 56357
rect 11550 56301 11618 56357
rect 11674 56301 11742 56357
rect 11798 56301 11866 56357
rect 11922 56301 11990 56357
rect 12046 56301 12114 56357
rect 12170 56301 12237 56357
rect 10187 56271 12237 56301
rect 10187 56233 10775 56271
rect 10827 56233 10899 56271
rect 10951 56233 11023 56271
rect 11075 56233 12237 56271
rect 10187 56177 10254 56233
rect 10310 56177 10378 56233
rect 10434 56177 10502 56233
rect 10558 56177 10626 56233
rect 10682 56177 10750 56233
rect 10827 56219 10874 56233
rect 10951 56219 10998 56233
rect 11075 56219 11122 56233
rect 10806 56177 10874 56219
rect 10930 56177 10998 56219
rect 11054 56177 11122 56219
rect 11178 56177 11246 56233
rect 11302 56177 11370 56233
rect 11426 56177 11494 56233
rect 11550 56177 11618 56233
rect 11674 56177 11742 56233
rect 11798 56177 11866 56233
rect 11922 56177 11990 56233
rect 12046 56177 12114 56233
rect 12170 56177 12237 56233
rect 10187 56147 12237 56177
rect 10187 56109 10775 56147
rect 10827 56109 10899 56147
rect 10951 56109 11023 56147
rect 11075 56109 12237 56147
rect 10187 56053 10254 56109
rect 10310 56053 10378 56109
rect 10434 56053 10502 56109
rect 10558 56053 10626 56109
rect 10682 56053 10750 56109
rect 10827 56095 10874 56109
rect 10951 56095 10998 56109
rect 11075 56095 11122 56109
rect 10806 56053 10874 56095
rect 10930 56053 10998 56095
rect 11054 56053 11122 56095
rect 11178 56053 11246 56109
rect 11302 56053 11370 56109
rect 11426 56053 11494 56109
rect 11550 56053 11618 56109
rect 11674 56053 11742 56109
rect 11798 56053 11866 56109
rect 11922 56053 11990 56109
rect 12046 56053 12114 56109
rect 12170 56053 12237 56109
rect 10187 56023 12237 56053
rect 10187 55971 10775 56023
rect 10827 55971 10899 56023
rect 10951 55971 11023 56023
rect 11075 55971 12237 56023
rect 10187 55899 12237 55971
rect 10187 55847 10775 55899
rect 10827 55847 10899 55899
rect 10951 55847 11023 55899
rect 11075 55847 12237 55899
rect 10187 55775 12237 55847
rect 10187 55723 10775 55775
rect 10827 55723 10899 55775
rect 10951 55723 11023 55775
rect 11075 55723 12237 55775
rect 10187 55651 12237 55723
rect 10187 55599 10775 55651
rect 10827 55599 10899 55651
rect 10951 55599 11023 55651
rect 11075 55599 12237 55651
rect 10187 55527 12237 55599
rect 10187 55475 10775 55527
rect 10827 55475 10899 55527
rect 10951 55475 11023 55527
rect 11075 55475 12237 55527
rect 10187 55403 12237 55475
rect 10187 55351 10775 55403
rect 10827 55351 10899 55403
rect 10951 55351 11023 55403
rect 11075 55351 12237 55403
rect 10187 55279 12237 55351
rect 10187 55227 10775 55279
rect 10827 55227 10899 55279
rect 10951 55227 11023 55279
rect 11075 55227 12237 55279
rect 10187 55155 12237 55227
rect 10187 55103 10775 55155
rect 10827 55103 10899 55155
rect 10951 55103 11023 55155
rect 11075 55103 12237 55155
rect 10187 55031 12237 55103
rect 10187 54979 10775 55031
rect 10827 54979 10899 55031
rect 10951 54979 11023 55031
rect 11075 54979 12237 55031
rect 10187 54907 12237 54979
rect 10187 54855 10775 54907
rect 10827 54855 10899 54907
rect 10951 54855 11023 54907
rect 11075 54855 12237 54907
rect 10187 54783 12237 54855
rect 10187 54731 10775 54783
rect 10827 54731 10899 54783
rect 10951 54731 11023 54783
rect 11075 54731 12237 54783
rect 10187 54659 12237 54731
rect 10187 54607 10775 54659
rect 10827 54607 10899 54659
rect 10951 54607 11023 54659
rect 11075 54607 12237 54659
rect 10187 54535 12237 54607
rect 10187 54483 10775 54535
rect 10827 54483 10899 54535
rect 10951 54483 11023 54535
rect 11075 54483 12237 54535
rect 10187 54411 12237 54483
rect 10187 54359 10775 54411
rect 10827 54359 10899 54411
rect 10951 54359 11023 54411
rect 11075 54359 12237 54411
rect 10187 54287 12237 54359
rect 10187 54235 10775 54287
rect 10827 54235 10899 54287
rect 10951 54235 11023 54287
rect 11075 54235 12237 54287
rect 10187 54163 12237 54235
rect 10187 54148 10775 54163
rect 10827 54148 10899 54163
rect 10951 54148 11023 54163
rect 11075 54148 12237 54163
rect 10187 54092 10254 54148
rect 10310 54092 10378 54148
rect 10434 54092 10502 54148
rect 10558 54092 10626 54148
rect 10682 54092 10750 54148
rect 10827 54111 10874 54148
rect 10951 54111 10998 54148
rect 11075 54111 11122 54148
rect 10806 54092 10874 54111
rect 10930 54092 10998 54111
rect 11054 54092 11122 54111
rect 11178 54092 11246 54148
rect 11302 54092 11370 54148
rect 11426 54092 11494 54148
rect 11550 54092 11618 54148
rect 11674 54092 11742 54148
rect 11798 54092 11866 54148
rect 11922 54092 11990 54148
rect 12046 54092 12114 54148
rect 12170 54092 12237 54148
rect 10187 54039 12237 54092
rect 10187 54024 10775 54039
rect 10827 54024 10899 54039
rect 10951 54024 11023 54039
rect 11075 54024 12237 54039
rect 10187 53968 10254 54024
rect 10310 53968 10378 54024
rect 10434 53968 10502 54024
rect 10558 53968 10626 54024
rect 10682 53968 10750 54024
rect 10827 53987 10874 54024
rect 10951 53987 10998 54024
rect 11075 53987 11122 54024
rect 10806 53968 10874 53987
rect 10930 53968 10998 53987
rect 11054 53968 11122 53987
rect 11178 53968 11246 54024
rect 11302 53968 11370 54024
rect 11426 53968 11494 54024
rect 11550 53968 11618 54024
rect 11674 53968 11742 54024
rect 11798 53968 11866 54024
rect 11922 53968 11990 54024
rect 12046 53968 12114 54024
rect 12170 53968 12237 54024
rect 10187 53915 12237 53968
rect 10187 53900 10775 53915
rect 10827 53900 10899 53915
rect 10951 53900 11023 53915
rect 11075 53900 12237 53915
rect 10187 53844 10254 53900
rect 10310 53844 10378 53900
rect 10434 53844 10502 53900
rect 10558 53844 10626 53900
rect 10682 53844 10750 53900
rect 10827 53863 10874 53900
rect 10951 53863 10998 53900
rect 11075 53863 11122 53900
rect 10806 53844 10874 53863
rect 10930 53844 10998 53863
rect 11054 53844 11122 53863
rect 11178 53844 11246 53900
rect 11302 53844 11370 53900
rect 11426 53844 11494 53900
rect 11550 53844 11618 53900
rect 11674 53844 11742 53900
rect 11798 53844 11866 53900
rect 11922 53844 11990 53900
rect 12046 53844 12114 53900
rect 12170 53844 12237 53900
rect 10187 53791 12237 53844
rect 10187 53776 10775 53791
rect 10827 53776 10899 53791
rect 10951 53776 11023 53791
rect 11075 53776 12237 53791
rect 10187 53720 10254 53776
rect 10310 53720 10378 53776
rect 10434 53720 10502 53776
rect 10558 53720 10626 53776
rect 10682 53720 10750 53776
rect 10827 53739 10874 53776
rect 10951 53739 10998 53776
rect 11075 53739 11122 53776
rect 10806 53720 10874 53739
rect 10930 53720 10998 53739
rect 11054 53720 11122 53739
rect 11178 53720 11246 53776
rect 11302 53720 11370 53776
rect 11426 53720 11494 53776
rect 11550 53720 11618 53776
rect 11674 53720 11742 53776
rect 11798 53720 11866 53776
rect 11922 53720 11990 53776
rect 12046 53720 12114 53776
rect 12170 53720 12237 53776
rect 10187 53667 12237 53720
rect 10187 53652 10775 53667
rect 10827 53652 10899 53667
rect 10951 53652 11023 53667
rect 11075 53652 12237 53667
rect 10187 53596 10254 53652
rect 10310 53596 10378 53652
rect 10434 53596 10502 53652
rect 10558 53596 10626 53652
rect 10682 53596 10750 53652
rect 10827 53615 10874 53652
rect 10951 53615 10998 53652
rect 11075 53615 11122 53652
rect 10806 53596 10874 53615
rect 10930 53596 10998 53615
rect 11054 53596 11122 53615
rect 11178 53596 11246 53652
rect 11302 53596 11370 53652
rect 11426 53596 11494 53652
rect 11550 53596 11618 53652
rect 11674 53596 11742 53652
rect 11798 53596 11866 53652
rect 11922 53596 11990 53652
rect 12046 53596 12114 53652
rect 12170 53596 12237 53652
rect 10187 53543 12237 53596
rect 10187 53528 10775 53543
rect 10827 53528 10899 53543
rect 10951 53528 11023 53543
rect 11075 53528 12237 53543
rect 10187 53472 10254 53528
rect 10310 53472 10378 53528
rect 10434 53472 10502 53528
rect 10558 53472 10626 53528
rect 10682 53472 10750 53528
rect 10827 53491 10874 53528
rect 10951 53491 10998 53528
rect 11075 53491 11122 53528
rect 10806 53472 10874 53491
rect 10930 53472 10998 53491
rect 11054 53472 11122 53491
rect 11178 53483 11246 53528
rect 11302 53483 11370 53528
rect 11426 53483 11494 53528
rect 11550 53483 11618 53528
rect 11674 53483 11742 53528
rect 11798 53483 11866 53528
rect 11922 53483 11990 53528
rect 12046 53483 12114 53528
rect 12170 53483 12237 53528
rect 11178 53472 11191 53483
rect 10187 53431 11191 53472
rect 11243 53472 11246 53483
rect 11351 53472 11370 53483
rect 11459 53472 11494 53483
rect 11567 53472 11618 53483
rect 11243 53431 11299 53472
rect 11351 53431 11407 53472
rect 11459 53431 11515 53472
rect 11567 53431 11623 53472
rect 11675 53431 11731 53483
rect 11798 53472 11839 53483
rect 11922 53472 11947 53483
rect 12046 53472 12055 53483
rect 11783 53431 11839 53472
rect 11891 53431 11947 53472
rect 11999 53431 12055 53472
rect 12107 53472 12114 53483
rect 12107 53431 12163 53472
rect 12215 53431 12237 53483
rect 10187 53419 12237 53431
rect 10187 53404 10775 53419
rect 10827 53404 10899 53419
rect 10951 53404 11023 53419
rect 11075 53404 12237 53419
rect 10187 53348 10254 53404
rect 10310 53348 10378 53404
rect 10434 53348 10502 53404
rect 10558 53348 10626 53404
rect 10682 53348 10750 53404
rect 10827 53367 10874 53404
rect 10951 53367 10998 53404
rect 11075 53367 11122 53404
rect 10806 53348 10874 53367
rect 10930 53348 10998 53367
rect 11054 53348 11122 53367
rect 11178 53375 11246 53404
rect 11302 53375 11370 53404
rect 11426 53375 11494 53404
rect 11550 53375 11618 53404
rect 11674 53375 11742 53404
rect 11798 53375 11866 53404
rect 11922 53375 11990 53404
rect 12046 53375 12114 53404
rect 12170 53375 12237 53404
rect 11178 53348 11191 53375
rect 10187 53323 11191 53348
rect 11243 53348 11246 53375
rect 11351 53348 11370 53375
rect 11459 53348 11494 53375
rect 11567 53348 11618 53375
rect 11243 53323 11299 53348
rect 11351 53323 11407 53348
rect 11459 53323 11515 53348
rect 11567 53323 11623 53348
rect 11675 53323 11731 53375
rect 11798 53348 11839 53375
rect 11922 53348 11947 53375
rect 12046 53348 12055 53375
rect 11783 53323 11839 53348
rect 11891 53323 11947 53348
rect 11999 53323 12055 53348
rect 12107 53348 12114 53375
rect 12107 53323 12163 53348
rect 12215 53323 12237 53375
rect 10187 53295 12237 53323
rect 10187 53280 10775 53295
rect 10827 53280 10899 53295
rect 10951 53280 11023 53295
rect 11075 53280 12237 53295
rect 10187 53224 10254 53280
rect 10310 53224 10378 53280
rect 10434 53224 10502 53280
rect 10558 53224 10626 53280
rect 10682 53224 10750 53280
rect 10827 53243 10874 53280
rect 10951 53243 10998 53280
rect 11075 53243 11122 53280
rect 10806 53224 10874 53243
rect 10930 53224 10998 53243
rect 11054 53224 11122 53243
rect 11178 53267 11246 53280
rect 11302 53267 11370 53280
rect 11426 53267 11494 53280
rect 11550 53267 11618 53280
rect 11674 53267 11742 53280
rect 11798 53267 11866 53280
rect 11922 53267 11990 53280
rect 12046 53267 12114 53280
rect 12170 53267 12237 53280
rect 11178 53224 11191 53267
rect 10187 53215 11191 53224
rect 11243 53224 11246 53267
rect 11351 53224 11370 53267
rect 11459 53224 11494 53267
rect 11567 53224 11618 53267
rect 11243 53215 11299 53224
rect 11351 53215 11407 53224
rect 11459 53215 11515 53224
rect 11567 53215 11623 53224
rect 11675 53215 11731 53267
rect 11798 53224 11839 53267
rect 11922 53224 11947 53267
rect 12046 53224 12055 53267
rect 11783 53215 11839 53224
rect 11891 53215 11947 53224
rect 11999 53215 12055 53224
rect 12107 53224 12114 53267
rect 12107 53215 12163 53224
rect 12215 53215 12237 53267
rect 10187 53156 12237 53215
rect 10187 53100 10254 53156
rect 10310 53100 10378 53156
rect 10434 53100 10502 53156
rect 10558 53100 10626 53156
rect 10682 53100 10750 53156
rect 10806 53100 10874 53156
rect 10930 53100 10998 53156
rect 11054 53100 11122 53156
rect 11178 53100 11246 53156
rect 11302 53100 11370 53156
rect 11426 53100 11494 53156
rect 11550 53100 11618 53156
rect 11674 53100 11742 53156
rect 11798 53100 11866 53156
rect 11922 53100 11990 53156
rect 12046 53100 12114 53156
rect 12170 53100 12237 53156
rect 10187 53032 12237 53100
rect 10187 52976 10254 53032
rect 10310 52976 10378 53032
rect 10434 52976 10502 53032
rect 10558 52976 10626 53032
rect 10682 52976 10750 53032
rect 10806 52976 10874 53032
rect 10930 52976 10998 53032
rect 11054 52976 11122 53032
rect 11178 52976 11246 53032
rect 11302 52976 11370 53032
rect 11426 52976 11494 53032
rect 11550 52976 11618 53032
rect 11674 52976 11742 53032
rect 11798 52976 11866 53032
rect 11922 52976 11990 53032
rect 12046 52976 12114 53032
rect 12170 52976 12237 53032
rect 10187 52908 12237 52976
rect 10187 52852 10254 52908
rect 10310 52852 10378 52908
rect 10434 52852 10502 52908
rect 10558 52852 10626 52908
rect 10682 52852 10750 52908
rect 10806 52852 10874 52908
rect 10930 52852 10998 52908
rect 11054 52852 11122 52908
rect 11178 52852 11246 52908
rect 11302 52852 11370 52908
rect 11426 52852 11494 52908
rect 11550 52852 11618 52908
rect 11674 52852 11742 52908
rect 11798 52852 11866 52908
rect 11922 52852 11990 52908
rect 12046 52852 12114 52908
rect 12170 52852 12237 52908
rect 10187 52548 12237 52852
rect 10187 52492 10254 52548
rect 10310 52492 10378 52548
rect 10434 52492 10502 52548
rect 10558 52492 10626 52548
rect 10682 52492 10750 52548
rect 10806 52492 10874 52548
rect 10930 52492 10998 52548
rect 11054 52492 11122 52548
rect 11178 52492 11246 52548
rect 11302 52492 11370 52548
rect 11426 52492 11494 52548
rect 11550 52492 11618 52548
rect 11674 52492 11742 52548
rect 11798 52492 11866 52548
rect 11922 52492 11990 52548
rect 12046 52492 12114 52548
rect 12170 52492 12237 52548
rect 10187 52424 12237 52492
rect 10187 52368 10254 52424
rect 10310 52368 10378 52424
rect 10434 52368 10502 52424
rect 10558 52368 10626 52424
rect 10682 52368 10750 52424
rect 10806 52368 10874 52424
rect 10930 52368 10998 52424
rect 11054 52368 11122 52424
rect 11178 52368 11246 52424
rect 11302 52368 11370 52424
rect 11426 52368 11494 52424
rect 11550 52368 11618 52424
rect 11674 52368 11742 52424
rect 11798 52368 11866 52424
rect 11922 52368 11990 52424
rect 12046 52368 12114 52424
rect 12170 52368 12237 52424
rect 10187 52300 12237 52368
rect 10187 52244 10254 52300
rect 10310 52244 10378 52300
rect 10434 52244 10502 52300
rect 10558 52244 10626 52300
rect 10682 52244 10750 52300
rect 10806 52244 10874 52300
rect 10930 52244 10998 52300
rect 11054 52244 11122 52300
rect 11178 52244 11246 52300
rect 11302 52244 11370 52300
rect 11426 52244 11494 52300
rect 11550 52244 11618 52300
rect 11674 52244 11742 52300
rect 11798 52244 11866 52300
rect 11922 52244 11990 52300
rect 12046 52244 12114 52300
rect 12170 52244 12237 52300
rect 10187 52176 12237 52244
rect 10187 52120 10254 52176
rect 10310 52120 10378 52176
rect 10434 52120 10502 52176
rect 10558 52120 10626 52176
rect 10682 52120 10750 52176
rect 10806 52120 10874 52176
rect 10930 52120 10998 52176
rect 11054 52120 11122 52176
rect 11178 52120 11246 52176
rect 11302 52120 11370 52176
rect 11426 52120 11494 52176
rect 11550 52120 11618 52176
rect 11674 52120 11742 52176
rect 11798 52120 11866 52176
rect 11922 52120 11990 52176
rect 12046 52120 12114 52176
rect 12170 52120 12237 52176
rect 10187 52052 12237 52120
rect 10187 52009 10254 52052
rect 10310 52009 10378 52052
rect 10434 52009 10502 52052
rect 10558 52009 10626 52052
rect 10682 52009 10750 52052
rect 10806 52009 10874 52052
rect 10930 52009 10998 52052
rect 11054 52009 11122 52052
rect 11178 52009 11246 52052
rect 11302 52009 11370 52052
rect 11426 52009 11494 52052
rect 11550 52009 11618 52052
rect 11674 52009 11742 52052
rect 11798 52009 11866 52052
rect 10187 51957 10253 52009
rect 10310 51996 10361 52009
rect 10434 51996 10469 52009
rect 10558 51996 10577 52009
rect 10682 51996 10685 52009
rect 10305 51957 10361 51996
rect 10413 51957 10469 51996
rect 10521 51957 10577 51996
rect 10629 51957 10685 51996
rect 10737 51996 10750 52009
rect 10845 51996 10874 52009
rect 10953 51996 10998 52009
rect 10737 51957 10793 51996
rect 10845 51957 10901 51996
rect 10953 51957 11009 51996
rect 11061 51957 11117 52009
rect 11178 51996 11225 52009
rect 11302 51996 11333 52009
rect 11426 51996 11441 52009
rect 11169 51957 11225 51996
rect 11277 51957 11333 51996
rect 11385 51957 11441 51996
rect 11493 51996 11494 52009
rect 11601 51996 11618 52009
rect 11709 51996 11742 52009
rect 11817 51996 11866 52009
rect 11922 51996 11990 52052
rect 12046 51996 12114 52052
rect 12170 51996 12237 52052
rect 11493 51957 11549 51996
rect 11601 51957 11657 51996
rect 11709 51957 11765 51996
rect 11817 51957 12237 51996
rect 10187 51928 12237 51957
rect 10187 51901 10254 51928
rect 10310 51901 10378 51928
rect 10434 51901 10502 51928
rect 10558 51901 10626 51928
rect 10682 51901 10750 51928
rect 10806 51901 10874 51928
rect 10930 51901 10998 51928
rect 11054 51901 11122 51928
rect 11178 51901 11246 51928
rect 11302 51901 11370 51928
rect 11426 51901 11494 51928
rect 11550 51901 11618 51928
rect 11674 51901 11742 51928
rect 11798 51901 11866 51928
rect 10187 51849 10253 51901
rect 10310 51872 10361 51901
rect 10434 51872 10469 51901
rect 10558 51872 10577 51901
rect 10682 51872 10685 51901
rect 10305 51849 10361 51872
rect 10413 51849 10469 51872
rect 10521 51849 10577 51872
rect 10629 51849 10685 51872
rect 10737 51872 10750 51901
rect 10845 51872 10874 51901
rect 10953 51872 10998 51901
rect 10737 51849 10793 51872
rect 10845 51849 10901 51872
rect 10953 51849 11009 51872
rect 11061 51849 11117 51901
rect 11178 51872 11225 51901
rect 11302 51872 11333 51901
rect 11426 51872 11441 51901
rect 11169 51849 11225 51872
rect 11277 51849 11333 51872
rect 11385 51849 11441 51872
rect 11493 51872 11494 51901
rect 11601 51872 11618 51901
rect 11709 51872 11742 51901
rect 11817 51872 11866 51901
rect 11922 51872 11990 51928
rect 12046 51872 12114 51928
rect 12170 51872 12237 51928
rect 11493 51849 11549 51872
rect 11601 51849 11657 51872
rect 11709 51849 11765 51872
rect 11817 51849 12237 51872
rect 10187 51804 12237 51849
rect 10187 51748 10254 51804
rect 10310 51748 10378 51804
rect 10434 51748 10502 51804
rect 10558 51748 10626 51804
rect 10682 51748 10750 51804
rect 10806 51748 10874 51804
rect 10930 51748 10998 51804
rect 11054 51748 11122 51804
rect 11178 51748 11246 51804
rect 11302 51748 11370 51804
rect 11426 51748 11494 51804
rect 11550 51748 11618 51804
rect 11674 51748 11742 51804
rect 11798 51748 11866 51804
rect 11922 51748 11990 51804
rect 12046 51748 12114 51804
rect 12170 51748 12237 51804
rect 10187 51680 12237 51748
rect 10187 51624 10254 51680
rect 10310 51624 10378 51680
rect 10434 51624 10502 51680
rect 10558 51624 10626 51680
rect 10682 51624 10750 51680
rect 10806 51624 10874 51680
rect 10930 51624 10998 51680
rect 11054 51624 11122 51680
rect 11178 51624 11246 51680
rect 11302 51624 11370 51680
rect 11426 51624 11494 51680
rect 11550 51624 11618 51680
rect 11674 51624 11742 51680
rect 11798 51624 11866 51680
rect 11922 51624 11990 51680
rect 12046 51624 12114 51680
rect 12170 51624 12237 51680
rect 10187 51556 12237 51624
rect 10187 51500 10254 51556
rect 10310 51500 10378 51556
rect 10434 51500 10502 51556
rect 10558 51500 10626 51556
rect 10682 51500 10750 51556
rect 10806 51500 10874 51556
rect 10930 51500 10998 51556
rect 11054 51500 11122 51556
rect 11178 51500 11246 51556
rect 11302 51500 11370 51556
rect 11426 51500 11494 51556
rect 11550 51500 11618 51556
rect 11674 51500 11742 51556
rect 11798 51500 11866 51556
rect 11922 51500 11990 51556
rect 12046 51500 12114 51556
rect 12170 51500 12237 51556
rect 10187 51432 12237 51500
rect 10187 51376 10254 51432
rect 10310 51376 10378 51432
rect 10434 51376 10502 51432
rect 10558 51376 10626 51432
rect 10682 51376 10750 51432
rect 10806 51376 10874 51432
rect 10930 51376 10998 51432
rect 11054 51376 11122 51432
rect 11178 51376 11246 51432
rect 11302 51376 11370 51432
rect 11426 51376 11494 51432
rect 11550 51376 11618 51432
rect 11674 51376 11742 51432
rect 11798 51376 11866 51432
rect 11922 51376 11990 51432
rect 12046 51376 12114 51432
rect 12170 51376 12237 51432
rect 10187 51308 12237 51376
rect 10187 51252 10254 51308
rect 10310 51252 10378 51308
rect 10434 51252 10502 51308
rect 10558 51252 10626 51308
rect 10682 51252 10750 51308
rect 10806 51252 10874 51308
rect 10930 51252 10998 51308
rect 11054 51252 11122 51308
rect 11178 51252 11246 51308
rect 11302 51252 11370 51308
rect 11426 51252 11494 51308
rect 11550 51252 11618 51308
rect 11674 51252 11742 51308
rect 11798 51252 11866 51308
rect 11922 51252 11990 51308
rect 12046 51252 12114 51308
rect 12170 51252 12237 51308
rect 10187 51206 12237 51252
rect 10187 51154 10253 51206
rect 10305 51154 10361 51206
rect 10413 51154 10469 51206
rect 10521 51154 10577 51206
rect 10629 51154 10685 51206
rect 10737 51154 10793 51206
rect 10845 51154 10901 51206
rect 10953 51154 11009 51206
rect 11061 51154 11117 51206
rect 11169 51154 11225 51206
rect 11277 51154 11333 51206
rect 11385 51154 11441 51206
rect 11493 51154 11549 51206
rect 11601 51154 11657 51206
rect 11709 51154 11765 51206
rect 11817 51154 12237 51206
rect 10187 51098 12237 51154
rect 10187 51046 10253 51098
rect 10305 51046 10361 51098
rect 10413 51046 10469 51098
rect 10521 51046 10577 51098
rect 10629 51046 10685 51098
rect 10737 51046 10793 51098
rect 10845 51046 10901 51098
rect 10953 51046 11009 51098
rect 11061 51046 11117 51098
rect 11169 51046 11225 51098
rect 11277 51046 11333 51098
rect 11385 51046 11441 51098
rect 11493 51046 11549 51098
rect 11601 51046 11657 51098
rect 11709 51046 11765 51098
rect 11817 51046 12237 51098
rect 10187 50990 12237 51046
rect 10187 50938 10253 50990
rect 10305 50938 10361 50990
rect 10413 50938 10469 50990
rect 10521 50938 10577 50990
rect 10629 50938 10685 50990
rect 10737 50938 10793 50990
rect 10845 50938 10901 50990
rect 10953 50938 11009 50990
rect 11061 50938 11117 50990
rect 11169 50938 11225 50990
rect 11277 50938 11333 50990
rect 11385 50938 11441 50990
rect 11493 50938 11549 50990
rect 11601 50938 11657 50990
rect 11709 50938 11765 50990
rect 11817 50938 12237 50990
rect 10187 50272 12237 50938
rect 10187 50220 10253 50272
rect 10305 50220 10361 50272
rect 10413 50220 10469 50272
rect 10521 50220 10577 50272
rect 10629 50220 10685 50272
rect 10737 50220 10793 50272
rect 10845 50220 10901 50272
rect 10953 50220 11009 50272
rect 11061 50220 11117 50272
rect 11169 50220 11225 50272
rect 11277 50220 11333 50272
rect 11385 50220 11441 50272
rect 11493 50220 11549 50272
rect 11601 50220 11657 50272
rect 11709 50220 11765 50272
rect 11817 50220 12237 50272
rect 10187 50164 12237 50220
rect 10187 50112 10253 50164
rect 10305 50112 10361 50164
rect 10413 50112 10469 50164
rect 10521 50112 10577 50164
rect 10629 50112 10685 50164
rect 10737 50112 10793 50164
rect 10845 50112 10901 50164
rect 10953 50112 11009 50164
rect 11061 50112 11117 50164
rect 11169 50112 11225 50164
rect 11277 50112 11333 50164
rect 11385 50112 11441 50164
rect 11493 50112 11549 50164
rect 11601 50112 11657 50164
rect 11709 50112 11765 50164
rect 11817 50112 12237 50164
rect 10187 50056 12237 50112
rect 10187 50004 10253 50056
rect 10305 50004 10361 50056
rect 10413 50004 10469 50056
rect 10521 50004 10577 50056
rect 10629 50004 10685 50056
rect 10737 50004 10793 50056
rect 10845 50004 10901 50056
rect 10953 50004 11009 50056
rect 11061 50004 11117 50056
rect 11169 50004 11225 50056
rect 11277 50004 11333 50056
rect 11385 50004 11441 50056
rect 11493 50004 11549 50056
rect 11601 50004 11657 50056
rect 11709 50004 11765 50056
rect 11817 50004 12237 50056
rect 10187 49348 12237 50004
rect 10187 49338 10254 49348
rect 10310 49338 10378 49348
rect 10434 49338 10502 49348
rect 10558 49338 10626 49348
rect 10682 49338 10750 49348
rect 10806 49338 10874 49348
rect 10930 49338 10998 49348
rect 11054 49338 11122 49348
rect 11178 49338 11246 49348
rect 11302 49338 11370 49348
rect 11426 49338 11494 49348
rect 11550 49338 11618 49348
rect 11674 49338 11742 49348
rect 11798 49338 11866 49348
rect 10187 49286 10253 49338
rect 10310 49292 10361 49338
rect 10434 49292 10469 49338
rect 10558 49292 10577 49338
rect 10682 49292 10685 49338
rect 10305 49286 10361 49292
rect 10413 49286 10469 49292
rect 10521 49286 10577 49292
rect 10629 49286 10685 49292
rect 10737 49292 10750 49338
rect 10845 49292 10874 49338
rect 10953 49292 10998 49338
rect 10737 49286 10793 49292
rect 10845 49286 10901 49292
rect 10953 49286 11009 49292
rect 11061 49286 11117 49338
rect 11178 49292 11225 49338
rect 11302 49292 11333 49338
rect 11426 49292 11441 49338
rect 11169 49286 11225 49292
rect 11277 49286 11333 49292
rect 11385 49286 11441 49292
rect 11493 49292 11494 49338
rect 11601 49292 11618 49338
rect 11709 49292 11742 49338
rect 11817 49292 11866 49338
rect 11922 49292 11990 49348
rect 12046 49292 12114 49348
rect 12170 49292 12237 49348
rect 11493 49286 11549 49292
rect 11601 49286 11657 49292
rect 11709 49286 11765 49292
rect 11817 49286 12237 49292
rect 10187 49230 12237 49286
rect 10187 49178 10253 49230
rect 10305 49224 10361 49230
rect 10413 49224 10469 49230
rect 10521 49224 10577 49230
rect 10629 49224 10685 49230
rect 10310 49178 10361 49224
rect 10434 49178 10469 49224
rect 10558 49178 10577 49224
rect 10682 49178 10685 49224
rect 10737 49224 10793 49230
rect 10845 49224 10901 49230
rect 10953 49224 11009 49230
rect 10737 49178 10750 49224
rect 10845 49178 10874 49224
rect 10953 49178 10998 49224
rect 11061 49178 11117 49230
rect 11169 49224 11225 49230
rect 11277 49224 11333 49230
rect 11385 49224 11441 49230
rect 11178 49178 11225 49224
rect 11302 49178 11333 49224
rect 11426 49178 11441 49224
rect 11493 49224 11549 49230
rect 11601 49224 11657 49230
rect 11709 49224 11765 49230
rect 11817 49224 12237 49230
rect 11493 49178 11494 49224
rect 11601 49178 11618 49224
rect 11709 49178 11742 49224
rect 11817 49178 11866 49224
rect 10187 49168 10254 49178
rect 10310 49168 10378 49178
rect 10434 49168 10502 49178
rect 10558 49168 10626 49178
rect 10682 49168 10750 49178
rect 10806 49168 10874 49178
rect 10930 49168 10998 49178
rect 11054 49168 11122 49178
rect 11178 49168 11246 49178
rect 11302 49168 11370 49178
rect 11426 49168 11494 49178
rect 11550 49168 11618 49178
rect 11674 49168 11742 49178
rect 11798 49168 11866 49178
rect 11922 49168 11990 49224
rect 12046 49168 12114 49224
rect 12170 49168 12237 49224
rect 10187 49122 12237 49168
rect 10187 49070 10253 49122
rect 10305 49100 10361 49122
rect 10413 49100 10469 49122
rect 10521 49100 10577 49122
rect 10629 49100 10685 49122
rect 10310 49070 10361 49100
rect 10434 49070 10469 49100
rect 10558 49070 10577 49100
rect 10682 49070 10685 49100
rect 10737 49100 10793 49122
rect 10845 49100 10901 49122
rect 10953 49100 11009 49122
rect 10737 49070 10750 49100
rect 10845 49070 10874 49100
rect 10953 49070 10998 49100
rect 11061 49070 11117 49122
rect 11169 49100 11225 49122
rect 11277 49100 11333 49122
rect 11385 49100 11441 49122
rect 11178 49070 11225 49100
rect 11302 49070 11333 49100
rect 11426 49070 11441 49100
rect 11493 49100 11549 49122
rect 11601 49100 11657 49122
rect 11709 49100 11765 49122
rect 11817 49100 12237 49122
rect 11493 49070 11494 49100
rect 11601 49070 11618 49100
rect 11709 49070 11742 49100
rect 11817 49070 11866 49100
rect 10187 49044 10254 49070
rect 10310 49044 10378 49070
rect 10434 49044 10502 49070
rect 10558 49044 10626 49070
rect 10682 49044 10750 49070
rect 10806 49044 10874 49070
rect 10930 49044 10998 49070
rect 11054 49044 11122 49070
rect 11178 49044 11246 49070
rect 11302 49044 11370 49070
rect 11426 49044 11494 49070
rect 11550 49044 11618 49070
rect 11674 49044 11742 49070
rect 11798 49044 11866 49070
rect 11922 49044 11990 49100
rect 12046 49044 12114 49100
rect 12170 49044 12237 49100
rect 10187 48976 12237 49044
rect 10187 48920 10254 48976
rect 10310 48920 10378 48976
rect 10434 48920 10502 48976
rect 10558 48920 10626 48976
rect 10682 48920 10750 48976
rect 10806 48920 10874 48976
rect 10930 48920 10998 48976
rect 11054 48920 11122 48976
rect 11178 48920 11246 48976
rect 11302 48920 11370 48976
rect 11426 48920 11494 48976
rect 11550 48920 11618 48976
rect 11674 48920 11742 48976
rect 11798 48920 11866 48976
rect 11922 48920 11990 48976
rect 12046 48920 12114 48976
rect 12170 48920 12237 48976
rect 10187 48852 12237 48920
rect 10187 48796 10254 48852
rect 10310 48796 10378 48852
rect 10434 48796 10502 48852
rect 10558 48796 10626 48852
rect 10682 48796 10750 48852
rect 10806 48796 10874 48852
rect 10930 48796 10998 48852
rect 11054 48796 11122 48852
rect 11178 48796 11246 48852
rect 11302 48796 11370 48852
rect 11426 48796 11494 48852
rect 11550 48796 11618 48852
rect 11674 48796 11742 48852
rect 11798 48796 11866 48852
rect 11922 48796 11990 48852
rect 12046 48796 12114 48852
rect 12170 48796 12237 48852
rect 10187 48728 12237 48796
rect 10187 48672 10254 48728
rect 10310 48672 10378 48728
rect 10434 48672 10502 48728
rect 10558 48672 10626 48728
rect 10682 48672 10750 48728
rect 10806 48672 10874 48728
rect 10930 48672 10998 48728
rect 11054 48672 11122 48728
rect 11178 48672 11246 48728
rect 11302 48672 11370 48728
rect 11426 48672 11494 48728
rect 11550 48672 11618 48728
rect 11674 48672 11742 48728
rect 11798 48672 11866 48728
rect 11922 48672 11990 48728
rect 12046 48672 12114 48728
rect 12170 48672 12237 48728
rect 10187 48604 12237 48672
rect 10187 48548 10254 48604
rect 10310 48548 10378 48604
rect 10434 48548 10502 48604
rect 10558 48548 10626 48604
rect 10682 48548 10750 48604
rect 10806 48548 10874 48604
rect 10930 48548 10998 48604
rect 11054 48548 11122 48604
rect 11178 48548 11246 48604
rect 11302 48548 11370 48604
rect 11426 48548 11494 48604
rect 11550 48548 11618 48604
rect 11674 48548 11742 48604
rect 11798 48548 11866 48604
rect 11922 48548 11990 48604
rect 12046 48548 12114 48604
rect 12170 48548 12237 48604
rect 10187 48480 12237 48548
rect 10187 48427 10254 48480
rect 10310 48427 10378 48480
rect 10434 48427 10502 48480
rect 10558 48427 10626 48480
rect 10682 48427 10750 48480
rect 10806 48427 10874 48480
rect 10930 48427 10998 48480
rect 11054 48427 11122 48480
rect 11178 48427 11246 48480
rect 11302 48427 11370 48480
rect 11426 48427 11494 48480
rect 11550 48427 11618 48480
rect 11674 48427 11742 48480
rect 11798 48427 11866 48480
rect 10187 48375 10253 48427
rect 10310 48424 10361 48427
rect 10434 48424 10469 48427
rect 10558 48424 10577 48427
rect 10682 48424 10685 48427
rect 10305 48375 10361 48424
rect 10413 48375 10469 48424
rect 10521 48375 10577 48424
rect 10629 48375 10685 48424
rect 10737 48424 10750 48427
rect 10845 48424 10874 48427
rect 10953 48424 10998 48427
rect 10737 48375 10793 48424
rect 10845 48375 10901 48424
rect 10953 48375 11009 48424
rect 11061 48375 11117 48427
rect 11178 48424 11225 48427
rect 11302 48424 11333 48427
rect 11426 48424 11441 48427
rect 11169 48375 11225 48424
rect 11277 48375 11333 48424
rect 11385 48375 11441 48424
rect 11493 48424 11494 48427
rect 11601 48424 11618 48427
rect 11709 48424 11742 48427
rect 11817 48424 11866 48427
rect 11922 48424 11990 48480
rect 12046 48424 12114 48480
rect 12170 48424 12237 48480
rect 11493 48375 11549 48424
rect 11601 48375 11657 48424
rect 11709 48375 11765 48424
rect 11817 48375 12237 48424
rect 10187 48356 12237 48375
rect 10187 48319 10254 48356
rect 10310 48319 10378 48356
rect 10434 48319 10502 48356
rect 10558 48319 10626 48356
rect 10682 48319 10750 48356
rect 10806 48319 10874 48356
rect 10930 48319 10998 48356
rect 11054 48319 11122 48356
rect 11178 48319 11246 48356
rect 11302 48319 11370 48356
rect 11426 48319 11494 48356
rect 11550 48319 11618 48356
rect 11674 48319 11742 48356
rect 11798 48319 11866 48356
rect 10187 48267 10253 48319
rect 10310 48300 10361 48319
rect 10434 48300 10469 48319
rect 10558 48300 10577 48319
rect 10682 48300 10685 48319
rect 10305 48267 10361 48300
rect 10413 48267 10469 48300
rect 10521 48267 10577 48300
rect 10629 48267 10685 48300
rect 10737 48300 10750 48319
rect 10845 48300 10874 48319
rect 10953 48300 10998 48319
rect 10737 48267 10793 48300
rect 10845 48267 10901 48300
rect 10953 48267 11009 48300
rect 11061 48267 11117 48319
rect 11178 48300 11225 48319
rect 11302 48300 11333 48319
rect 11426 48300 11441 48319
rect 11169 48267 11225 48300
rect 11277 48267 11333 48300
rect 11385 48267 11441 48300
rect 11493 48300 11494 48319
rect 11601 48300 11618 48319
rect 11709 48300 11742 48319
rect 11817 48300 11866 48319
rect 11922 48300 11990 48356
rect 12046 48300 12114 48356
rect 12170 48300 12237 48356
rect 11493 48267 11549 48300
rect 11601 48267 11657 48300
rect 11709 48267 11765 48300
rect 11817 48267 12237 48300
rect 10187 48232 12237 48267
rect 10187 48176 10254 48232
rect 10310 48176 10378 48232
rect 10434 48176 10502 48232
rect 10558 48176 10626 48232
rect 10682 48176 10750 48232
rect 10806 48176 10874 48232
rect 10930 48176 10998 48232
rect 11054 48176 11122 48232
rect 11178 48176 11246 48232
rect 11302 48176 11370 48232
rect 11426 48176 11494 48232
rect 11550 48176 11618 48232
rect 11674 48176 11742 48232
rect 11798 48176 11866 48232
rect 11922 48176 11990 48232
rect 12046 48176 12114 48232
rect 12170 48176 12237 48232
rect 10187 48108 12237 48176
rect 10187 48052 10254 48108
rect 10310 48052 10378 48108
rect 10434 48052 10502 48108
rect 10558 48052 10626 48108
rect 10682 48052 10750 48108
rect 10806 48052 10874 48108
rect 10930 48052 10998 48108
rect 11054 48052 11122 48108
rect 11178 48052 11246 48108
rect 11302 48052 11370 48108
rect 11426 48052 11494 48108
rect 11550 48052 11618 48108
rect 11674 48052 11742 48108
rect 11798 48052 11866 48108
rect 11922 48052 11990 48108
rect 12046 48052 12114 48108
rect 12170 48052 12237 48108
rect 10187 47163 12237 48052
rect 12297 56741 12497 57278
rect 12297 56689 12317 56741
rect 12369 56689 12425 56741
rect 12477 56689 12497 56741
rect 12297 55748 12497 56689
rect 12297 55692 12307 55748
rect 12363 55692 12431 55748
rect 12487 55692 12497 55748
rect 12297 55624 12497 55692
rect 12297 55568 12307 55624
rect 12363 55568 12431 55624
rect 12487 55568 12497 55624
rect 12297 55500 12497 55568
rect 12297 55444 12307 55500
rect 12363 55444 12431 55500
rect 12487 55444 12497 55500
rect 12297 55376 12497 55444
rect 12297 55320 12307 55376
rect 12363 55320 12431 55376
rect 12487 55320 12497 55376
rect 12297 55252 12497 55320
rect 12297 55196 12307 55252
rect 12363 55196 12431 55252
rect 12487 55196 12497 55252
rect 12297 55128 12497 55196
rect 12297 55072 12307 55128
rect 12363 55072 12431 55128
rect 12487 55072 12497 55128
rect 12297 55004 12497 55072
rect 12297 54948 12307 55004
rect 12363 54948 12431 55004
rect 12487 54948 12497 55004
rect 12297 54880 12497 54948
rect 12297 54824 12307 54880
rect 12363 54824 12431 54880
rect 12487 54824 12497 54880
rect 12297 54756 12497 54824
rect 12297 54700 12307 54756
rect 12363 54700 12431 54756
rect 12487 54700 12497 54756
rect 12297 54632 12497 54700
rect 12297 54576 12307 54632
rect 12363 54576 12431 54632
rect 12487 54576 12497 54632
rect 12297 54508 12497 54576
rect 12297 54452 12307 54508
rect 12363 54452 12431 54508
rect 12487 54452 12497 54508
rect 12297 53621 12497 54452
rect 12297 53569 12317 53621
rect 12369 53569 12425 53621
rect 12477 53569 12497 53621
rect 12297 52594 12497 53569
rect 12297 52542 12336 52594
rect 12388 52542 12497 52594
rect 12297 52486 12497 52542
rect 12297 52434 12336 52486
rect 12388 52434 12497 52486
rect 12297 52378 12497 52434
rect 12297 52326 12336 52378
rect 12388 52326 12497 52378
rect 12297 52270 12497 52326
rect 12297 52218 12336 52270
rect 12388 52218 12497 52270
rect 12297 52162 12497 52218
rect 12297 52110 12336 52162
rect 12388 52110 12497 52162
rect 12297 52054 12497 52110
rect 12297 52002 12336 52054
rect 12388 52002 12497 52054
rect 12297 51946 12497 52002
rect 12297 51894 12336 51946
rect 12388 51894 12497 51946
rect 12297 51838 12497 51894
rect 12297 51786 12336 51838
rect 12388 51786 12497 51838
rect 12297 51730 12497 51786
rect 12297 51678 12336 51730
rect 12388 51678 12497 51730
rect 12297 51622 12497 51678
rect 12297 51570 12336 51622
rect 12388 51570 12497 51622
rect 12297 51514 12497 51570
rect 12297 51462 12336 51514
rect 12388 51462 12497 51514
rect 12297 51406 12497 51462
rect 12297 51354 12336 51406
rect 12388 51354 12497 51406
rect 12297 51298 12497 51354
rect 12297 51246 12336 51298
rect 12388 51246 12497 51298
rect 12297 51190 12497 51246
rect 12297 51138 12336 51190
rect 12388 51138 12497 51190
rect 12297 51082 12497 51138
rect 12297 51030 12336 51082
rect 12388 51030 12497 51082
rect 12297 50974 12497 51030
rect 12297 50922 12336 50974
rect 12388 50922 12497 50974
rect 12297 50866 12497 50922
rect 12297 50814 12336 50866
rect 12388 50814 12497 50866
rect 12297 50758 12497 50814
rect 12297 50706 12336 50758
rect 12388 50706 12497 50758
rect 12297 50650 12497 50706
rect 12297 50598 12336 50650
rect 12388 50598 12497 50650
rect 12297 50542 12497 50598
rect 12297 50490 12336 50542
rect 12388 50490 12497 50542
rect 12297 50434 12497 50490
rect 12297 50382 12336 50434
rect 12388 50382 12497 50434
rect 12297 50326 12497 50382
rect 12297 50274 12336 50326
rect 12388 50274 12497 50326
rect 12297 50218 12497 50274
rect 12297 50166 12336 50218
rect 12388 50166 12497 50218
rect 12297 50110 12497 50166
rect 12297 50058 12336 50110
rect 12388 50058 12497 50110
rect 12297 50002 12497 50058
rect 12297 49950 12336 50002
rect 12388 49950 12497 50002
rect 12297 49894 12497 49950
rect 12297 49842 12336 49894
rect 12388 49842 12497 49894
rect 12297 49786 12497 49842
rect 12297 49734 12336 49786
rect 12388 49734 12497 49786
rect 12297 49678 12497 49734
rect 12297 49626 12336 49678
rect 12388 49626 12497 49678
rect 12297 49570 12497 49626
rect 12297 49518 12336 49570
rect 12388 49518 12497 49570
rect 12297 49462 12497 49518
rect 12297 49410 12336 49462
rect 12388 49410 12497 49462
rect 12297 49354 12497 49410
rect 12297 49302 12336 49354
rect 12388 49302 12497 49354
rect 12297 49246 12497 49302
rect 12297 49194 12336 49246
rect 12388 49194 12497 49246
rect 12297 49138 12497 49194
rect 12297 49086 12336 49138
rect 12388 49086 12497 49138
rect 12297 49030 12497 49086
rect 12297 48978 12336 49030
rect 12388 48978 12497 49030
rect 12297 48922 12497 48978
rect 12297 48870 12336 48922
rect 12388 48870 12497 48922
rect 12297 48814 12497 48870
rect 12297 48762 12336 48814
rect 12388 48762 12497 48814
rect 12297 48706 12497 48762
rect 12297 48654 12336 48706
rect 12388 48654 12497 48706
rect 12297 48598 12497 48654
rect 12297 48546 12336 48598
rect 12388 48546 12497 48598
rect 12297 48490 12497 48546
rect 12297 48438 12336 48490
rect 12388 48438 12497 48490
rect 12297 48382 12497 48438
rect 12297 48330 12336 48382
rect 12388 48330 12497 48382
rect 12297 48274 12497 48330
rect 12297 48222 12336 48274
rect 12388 48222 12497 48274
rect 12297 48166 12497 48222
rect 12297 48114 12336 48166
rect 12388 48114 12497 48166
rect 12297 48058 12497 48114
rect 12297 48006 12336 48058
rect 12388 48006 12497 48058
rect 12297 47950 12497 48006
rect 12297 47898 12336 47950
rect 12388 47898 12497 47950
rect 12297 47842 12497 47898
rect 12297 47790 12336 47842
rect 12388 47790 12497 47842
rect 12297 47748 12497 47790
rect 12297 47692 12307 47748
rect 12363 47734 12431 47748
rect 12388 47692 12431 47734
rect 12487 47692 12497 47748
rect 12297 47682 12336 47692
rect 12388 47682 12497 47692
rect 12297 47624 12497 47682
rect 12297 47568 12307 47624
rect 12363 47568 12431 47624
rect 12487 47568 12497 47624
rect 12297 47500 12497 47568
rect 12297 47444 12307 47500
rect 12363 47444 12431 47500
rect 12487 47444 12497 47500
rect 12297 47376 12497 47444
rect 12297 47320 12307 47376
rect 12363 47320 12431 47376
rect 12487 47320 12497 47376
rect 12297 47252 12497 47320
rect 12297 47196 12307 47252
rect 12363 47196 12431 47252
rect 12487 47196 12497 47252
rect 9927 47072 9937 47128
rect 9993 47072 10061 47128
rect 10117 47072 10127 47128
rect 9927 47004 10127 47072
rect 9927 46948 9937 47004
rect 9993 46948 10061 47004
rect 10117 46948 10127 47004
rect 9927 46880 10127 46948
rect 9927 46824 9937 46880
rect 9993 46824 10061 46880
rect 10117 46824 10127 46880
rect 9927 46756 10127 46824
rect 9927 46700 9937 46756
rect 9993 46700 10061 46756
rect 10117 46700 10127 46756
rect 9927 46632 10127 46700
rect 9927 46576 9937 46632
rect 9993 46576 10061 46632
rect 10117 46576 10127 46632
rect 9927 46508 10127 46576
rect 9927 46452 9937 46508
rect 9993 46452 10061 46508
rect 10117 46452 10127 46508
rect 9927 46442 10127 46452
rect 12297 47128 12497 47196
rect 12817 57225 14717 57447
rect 12817 57169 12871 57225
rect 12927 57169 12995 57225
rect 13051 57169 13119 57225
rect 13175 57169 13243 57225
rect 13299 57169 13367 57225
rect 13423 57169 13491 57225
rect 13547 57169 13615 57225
rect 13671 57169 13739 57225
rect 13795 57169 13863 57225
rect 13919 57169 13987 57225
rect 14043 57169 14111 57225
rect 14167 57169 14235 57225
rect 14291 57169 14359 57225
rect 14415 57169 14483 57225
rect 14539 57169 14607 57225
rect 14663 57169 14717 57225
rect 12817 57104 14717 57169
rect 12817 57101 12931 57104
rect 12817 57045 12871 57101
rect 12927 57052 12931 57101
rect 12983 57101 13039 57104
rect 13091 57101 13147 57104
rect 13199 57101 13255 57104
rect 12983 57052 12995 57101
rect 13091 57052 13119 57101
rect 13199 57052 13243 57101
rect 13307 57052 13363 57104
rect 13415 57101 13471 57104
rect 13523 57101 13579 57104
rect 13631 57101 13687 57104
rect 13423 57052 13471 57101
rect 13547 57052 13579 57101
rect 13671 57052 13687 57101
rect 13739 57101 13795 57104
rect 12927 57045 12995 57052
rect 13051 57045 13119 57052
rect 13175 57045 13243 57052
rect 13299 57045 13367 57052
rect 13423 57045 13491 57052
rect 13547 57045 13615 57052
rect 13671 57045 13739 57052
rect 13847 57101 13903 57104
rect 13955 57101 14011 57104
rect 14063 57101 14119 57104
rect 13847 57052 13863 57101
rect 13955 57052 13987 57101
rect 14063 57052 14111 57101
rect 14171 57052 14227 57104
rect 14279 57101 14335 57104
rect 14387 57101 14443 57104
rect 14495 57101 14551 57104
rect 14291 57052 14335 57101
rect 14415 57052 14443 57101
rect 14539 57052 14551 57101
rect 14603 57101 14717 57104
rect 14603 57052 14607 57101
rect 13795 57045 13863 57052
rect 13919 57045 13987 57052
rect 14043 57045 14111 57052
rect 14167 57045 14235 57052
rect 14291 57045 14359 57052
rect 14415 57045 14483 57052
rect 14539 57045 14607 57052
rect 14663 57045 14717 57101
rect 12817 56977 14717 57045
rect 12817 56921 12871 56977
rect 12927 56921 12995 56977
rect 13051 56921 13119 56977
rect 13175 56921 13243 56977
rect 13299 56921 13367 56977
rect 13423 56921 13491 56977
rect 13547 56921 13615 56977
rect 13671 56921 13739 56977
rect 13795 56921 13863 56977
rect 13919 56921 13987 56977
rect 14043 56921 14111 56977
rect 14167 56921 14235 56977
rect 14291 56921 14359 56977
rect 14415 56921 14483 56977
rect 14539 56921 14607 56977
rect 14663 56921 14717 56977
rect 12817 56853 14717 56921
rect 12817 56797 12871 56853
rect 12927 56797 12995 56853
rect 13051 56797 13119 56853
rect 13175 56797 13243 56853
rect 13299 56797 13367 56853
rect 13423 56797 13491 56853
rect 13547 56797 13615 56853
rect 13671 56797 13739 56853
rect 13795 56797 13863 56853
rect 13919 56797 13987 56853
rect 14043 56797 14111 56853
rect 14167 56797 14235 56853
rect 14291 56797 14359 56853
rect 14415 56797 14483 56853
rect 14539 56797 14607 56853
rect 14663 56797 14717 56853
rect 12817 56729 14717 56797
rect 12817 56673 12871 56729
rect 12927 56673 12995 56729
rect 13051 56673 13119 56729
rect 13175 56673 13243 56729
rect 13299 56673 13367 56729
rect 13423 56673 13491 56729
rect 13547 56673 13615 56729
rect 13671 56673 13739 56729
rect 13795 56673 13863 56729
rect 13919 56673 13987 56729
rect 14043 56673 14111 56729
rect 14167 56673 14235 56729
rect 14291 56673 14359 56729
rect 14415 56673 14483 56729
rect 14539 56673 14607 56729
rect 14663 56673 14717 56729
rect 12817 56643 14717 56673
rect 12817 56605 14185 56643
rect 14237 56605 14309 56643
rect 14361 56605 14433 56643
rect 14485 56605 14557 56643
rect 14609 56605 14717 56643
rect 12817 56549 12871 56605
rect 12927 56549 12995 56605
rect 13051 56549 13119 56605
rect 13175 56549 13243 56605
rect 13299 56549 13367 56605
rect 13423 56549 13491 56605
rect 13547 56549 13615 56605
rect 13671 56549 13739 56605
rect 13795 56549 13863 56605
rect 13919 56549 13987 56605
rect 14043 56549 14111 56605
rect 14167 56591 14185 56605
rect 14291 56591 14309 56605
rect 14415 56591 14433 56605
rect 14539 56591 14557 56605
rect 14167 56549 14235 56591
rect 14291 56549 14359 56591
rect 14415 56549 14483 56591
rect 14539 56549 14607 56591
rect 14663 56549 14717 56605
rect 12817 56519 14717 56549
rect 12817 56481 14185 56519
rect 14237 56481 14309 56519
rect 14361 56481 14433 56519
rect 14485 56481 14557 56519
rect 14609 56481 14717 56519
rect 12817 56425 12871 56481
rect 12927 56425 12995 56481
rect 13051 56425 13119 56481
rect 13175 56425 13243 56481
rect 13299 56425 13367 56481
rect 13423 56425 13491 56481
rect 13547 56425 13615 56481
rect 13671 56425 13739 56481
rect 13795 56425 13863 56481
rect 13919 56425 13987 56481
rect 14043 56425 14111 56481
rect 14167 56467 14185 56481
rect 14291 56467 14309 56481
rect 14415 56467 14433 56481
rect 14539 56467 14557 56481
rect 14167 56425 14235 56467
rect 14291 56425 14359 56467
rect 14415 56425 14483 56467
rect 14539 56425 14607 56467
rect 14663 56425 14717 56481
rect 12817 56395 14717 56425
rect 12817 56357 14185 56395
rect 14237 56357 14309 56395
rect 14361 56357 14433 56395
rect 14485 56357 14557 56395
rect 14609 56357 14717 56395
rect 12817 56301 12871 56357
rect 12927 56301 12995 56357
rect 13051 56301 13119 56357
rect 13175 56301 13243 56357
rect 13299 56301 13367 56357
rect 13423 56301 13491 56357
rect 13547 56301 13615 56357
rect 13671 56301 13739 56357
rect 13795 56301 13863 56357
rect 13919 56301 13987 56357
rect 14043 56301 14111 56357
rect 14167 56343 14185 56357
rect 14291 56343 14309 56357
rect 14415 56343 14433 56357
rect 14539 56343 14557 56357
rect 14167 56301 14235 56343
rect 14291 56301 14359 56343
rect 14415 56301 14483 56343
rect 14539 56301 14607 56343
rect 14663 56301 14717 56357
rect 12817 56271 14717 56301
rect 12817 56233 14185 56271
rect 14237 56233 14309 56271
rect 14361 56233 14433 56271
rect 14485 56233 14557 56271
rect 14609 56233 14717 56271
rect 12817 56177 12871 56233
rect 12927 56177 12995 56233
rect 13051 56177 13119 56233
rect 13175 56177 13243 56233
rect 13299 56177 13367 56233
rect 13423 56177 13491 56233
rect 13547 56177 13615 56233
rect 13671 56177 13739 56233
rect 13795 56177 13863 56233
rect 13919 56177 13987 56233
rect 14043 56177 14111 56233
rect 14167 56219 14185 56233
rect 14291 56219 14309 56233
rect 14415 56219 14433 56233
rect 14539 56219 14557 56233
rect 14167 56177 14235 56219
rect 14291 56177 14359 56219
rect 14415 56177 14483 56219
rect 14539 56177 14607 56219
rect 14663 56177 14717 56233
rect 12817 56147 14717 56177
rect 12817 56109 14185 56147
rect 14237 56109 14309 56147
rect 14361 56109 14433 56147
rect 14485 56109 14557 56147
rect 14609 56109 14717 56147
rect 12817 56053 12871 56109
rect 12927 56053 12995 56109
rect 13051 56053 13119 56109
rect 13175 56053 13243 56109
rect 13299 56053 13367 56109
rect 13423 56053 13491 56109
rect 13547 56053 13615 56109
rect 13671 56053 13739 56109
rect 13795 56053 13863 56109
rect 13919 56053 13987 56109
rect 14043 56053 14111 56109
rect 14167 56095 14185 56109
rect 14291 56095 14309 56109
rect 14415 56095 14433 56109
rect 14539 56095 14557 56109
rect 14167 56053 14235 56095
rect 14291 56053 14359 56095
rect 14415 56053 14483 56095
rect 14539 56053 14607 56095
rect 14663 56053 14717 56109
rect 12817 56023 14717 56053
rect 12817 55971 14185 56023
rect 14237 55971 14309 56023
rect 14361 55971 14433 56023
rect 14485 55971 14557 56023
rect 14609 55971 14717 56023
rect 14892 57261 14989 57271
rect 14892 56017 14902 57261
rect 14958 56017 14989 57261
rect 14892 56007 14989 56017
rect 12817 55899 14717 55971
rect 12817 55847 14185 55899
rect 14237 55847 14309 55899
rect 14361 55847 14433 55899
rect 14485 55847 14557 55899
rect 14609 55847 14717 55899
rect 12817 55775 14717 55847
rect 12817 55723 14185 55775
rect 14237 55723 14309 55775
rect 14361 55723 14433 55775
rect 14485 55723 14557 55775
rect 14609 55723 14717 55775
rect 12817 55651 14717 55723
rect 12817 55599 14185 55651
rect 14237 55599 14309 55651
rect 14361 55599 14433 55651
rect 14485 55599 14557 55651
rect 14609 55599 14717 55651
rect 12817 55527 14717 55599
rect 12817 55475 14185 55527
rect 14237 55475 14309 55527
rect 14361 55475 14433 55527
rect 14485 55475 14557 55527
rect 14609 55475 14717 55527
rect 12817 55403 14717 55475
rect 12817 55351 14185 55403
rect 14237 55351 14309 55403
rect 14361 55351 14433 55403
rect 14485 55351 14557 55403
rect 14609 55351 14717 55403
rect 12817 55279 14717 55351
rect 12817 55227 14185 55279
rect 14237 55227 14309 55279
rect 14361 55227 14433 55279
rect 14485 55227 14557 55279
rect 14609 55227 14717 55279
rect 12817 55155 14717 55227
rect 12817 55103 14185 55155
rect 14237 55103 14309 55155
rect 14361 55103 14433 55155
rect 14485 55103 14557 55155
rect 14609 55103 14717 55155
rect 12817 55031 14717 55103
rect 12817 54979 14185 55031
rect 14237 54979 14309 55031
rect 14361 54979 14433 55031
rect 14485 54979 14557 55031
rect 14609 54979 14717 55031
rect 12817 54907 14717 54979
rect 12817 54855 14185 54907
rect 14237 54855 14309 54907
rect 14361 54855 14433 54907
rect 14485 54855 14557 54907
rect 14609 54855 14717 54907
rect 12817 54783 14717 54855
rect 12817 54731 14185 54783
rect 14237 54731 14309 54783
rect 14361 54731 14433 54783
rect 14485 54731 14557 54783
rect 14609 54731 14717 54783
rect 12817 54659 14717 54731
rect 12817 54607 14185 54659
rect 14237 54607 14309 54659
rect 14361 54607 14433 54659
rect 14485 54607 14557 54659
rect 14609 54607 14717 54659
rect 12817 54535 14717 54607
rect 12817 54483 14185 54535
rect 14237 54483 14309 54535
rect 14361 54483 14433 54535
rect 14485 54483 14557 54535
rect 14609 54483 14717 54535
rect 12817 54411 14717 54483
rect 12817 54359 14185 54411
rect 14237 54359 14309 54411
rect 14361 54359 14433 54411
rect 14485 54359 14557 54411
rect 14609 54359 14717 54411
rect 12817 54287 14717 54359
rect 12817 54235 14185 54287
rect 14237 54235 14309 54287
rect 14361 54235 14433 54287
rect 14485 54235 14557 54287
rect 14609 54235 14717 54287
rect 12817 54163 14717 54235
rect 12817 54148 14185 54163
rect 14237 54148 14309 54163
rect 14361 54148 14433 54163
rect 14485 54148 14557 54163
rect 14609 54148 14717 54163
rect 12817 54092 12871 54148
rect 12927 54092 12995 54148
rect 13051 54092 13119 54148
rect 13175 54092 13243 54148
rect 13299 54092 13367 54148
rect 13423 54092 13491 54148
rect 13547 54092 13615 54148
rect 13671 54092 13739 54148
rect 13795 54092 13863 54148
rect 13919 54092 13987 54148
rect 14043 54092 14111 54148
rect 14167 54111 14185 54148
rect 14291 54111 14309 54148
rect 14415 54111 14433 54148
rect 14539 54111 14557 54148
rect 14167 54092 14235 54111
rect 14291 54092 14359 54111
rect 14415 54092 14483 54111
rect 14539 54092 14607 54111
rect 14663 54092 14717 54148
rect 12817 54039 14717 54092
rect 12817 54024 14185 54039
rect 14237 54024 14309 54039
rect 14361 54024 14433 54039
rect 14485 54024 14557 54039
rect 14609 54024 14717 54039
rect 12817 53968 12871 54024
rect 12927 53968 12995 54024
rect 13051 53968 13119 54024
rect 13175 53968 13243 54024
rect 13299 53968 13367 54024
rect 13423 53968 13491 54024
rect 13547 53968 13615 54024
rect 13671 53968 13739 54024
rect 13795 53968 13863 54024
rect 13919 53968 13987 54024
rect 14043 53968 14111 54024
rect 14167 53987 14185 54024
rect 14291 53987 14309 54024
rect 14415 53987 14433 54024
rect 14539 53987 14557 54024
rect 14167 53968 14235 53987
rect 14291 53968 14359 53987
rect 14415 53968 14483 53987
rect 14539 53968 14607 53987
rect 14663 53968 14717 54024
rect 12817 53915 14717 53968
rect 12817 53900 14185 53915
rect 14237 53900 14309 53915
rect 14361 53900 14433 53915
rect 14485 53900 14557 53915
rect 14609 53900 14717 53915
rect 12817 53844 12871 53900
rect 12927 53844 12995 53900
rect 13051 53844 13119 53900
rect 13175 53844 13243 53900
rect 13299 53844 13367 53900
rect 13423 53844 13491 53900
rect 13547 53844 13615 53900
rect 13671 53844 13739 53900
rect 13795 53844 13863 53900
rect 13919 53844 13987 53900
rect 14043 53844 14111 53900
rect 14167 53863 14185 53900
rect 14291 53863 14309 53900
rect 14415 53863 14433 53900
rect 14539 53863 14557 53900
rect 14167 53844 14235 53863
rect 14291 53844 14359 53863
rect 14415 53844 14483 53863
rect 14539 53844 14607 53863
rect 14663 53844 14717 53900
rect 12817 53791 14717 53844
rect 12817 53776 14185 53791
rect 14237 53776 14309 53791
rect 14361 53776 14433 53791
rect 14485 53776 14557 53791
rect 14609 53776 14717 53791
rect 12817 53720 12871 53776
rect 12927 53720 12995 53776
rect 13051 53720 13119 53776
rect 13175 53720 13243 53776
rect 13299 53720 13367 53776
rect 13423 53720 13491 53776
rect 13547 53720 13615 53776
rect 13671 53720 13739 53776
rect 13795 53720 13863 53776
rect 13919 53720 13987 53776
rect 14043 53720 14111 53776
rect 14167 53739 14185 53776
rect 14291 53739 14309 53776
rect 14415 53739 14433 53776
rect 14539 53739 14557 53776
rect 14167 53720 14235 53739
rect 14291 53720 14359 53739
rect 14415 53720 14483 53739
rect 14539 53720 14607 53739
rect 14663 53720 14717 53776
rect 12817 53667 14717 53720
rect 12817 53652 14185 53667
rect 14237 53652 14309 53667
rect 14361 53652 14433 53667
rect 14485 53652 14557 53667
rect 14609 53652 14717 53667
rect 12817 53596 12871 53652
rect 12927 53596 12995 53652
rect 13051 53596 13119 53652
rect 13175 53596 13243 53652
rect 13299 53596 13367 53652
rect 13423 53596 13491 53652
rect 13547 53596 13615 53652
rect 13671 53596 13739 53652
rect 13795 53596 13863 53652
rect 13919 53596 13987 53652
rect 14043 53596 14111 53652
rect 14167 53615 14185 53652
rect 14291 53615 14309 53652
rect 14415 53615 14433 53652
rect 14539 53615 14557 53652
rect 14167 53596 14235 53615
rect 14291 53596 14359 53615
rect 14415 53596 14483 53615
rect 14539 53596 14607 53615
rect 14663 53596 14717 53652
rect 12817 53543 14717 53596
rect 12817 53528 14185 53543
rect 14237 53528 14309 53543
rect 14361 53528 14433 53543
rect 14485 53528 14557 53543
rect 14609 53528 14717 53543
rect 12817 53483 12871 53528
rect 12927 53483 12995 53528
rect 13051 53483 13119 53528
rect 13175 53483 13243 53528
rect 13299 53483 13367 53528
rect 13423 53483 13491 53528
rect 13547 53483 13615 53528
rect 13671 53483 13739 53528
rect 13795 53483 13863 53528
rect 13919 53483 13987 53528
rect 14043 53483 14111 53528
rect 12817 53431 12869 53483
rect 12927 53472 12977 53483
rect 13051 53472 13085 53483
rect 13175 53472 13193 53483
rect 13299 53472 13301 53483
rect 12921 53431 12977 53472
rect 13029 53431 13085 53472
rect 13137 53431 13193 53472
rect 13245 53431 13301 53472
rect 13353 53472 13367 53483
rect 13461 53472 13491 53483
rect 13569 53472 13615 53483
rect 13353 53431 13409 53472
rect 13461 53431 13517 53472
rect 13569 53431 13625 53472
rect 13677 53431 13733 53483
rect 13795 53472 13841 53483
rect 13919 53472 13949 53483
rect 14043 53472 14057 53483
rect 13785 53431 13841 53472
rect 13893 53431 13949 53472
rect 14001 53431 14057 53472
rect 14109 53472 14111 53483
rect 14167 53491 14185 53528
rect 14291 53491 14309 53528
rect 14415 53491 14433 53528
rect 14539 53491 14557 53528
rect 14167 53472 14235 53491
rect 14291 53472 14359 53491
rect 14415 53472 14483 53491
rect 14539 53472 14607 53491
rect 14663 53472 14717 53528
rect 14109 53431 14717 53472
rect 12817 53419 14717 53431
rect 12817 53404 14185 53419
rect 14237 53404 14309 53419
rect 14361 53404 14433 53419
rect 14485 53404 14557 53419
rect 14609 53404 14717 53419
rect 12817 53375 12871 53404
rect 12927 53375 12995 53404
rect 13051 53375 13119 53404
rect 13175 53375 13243 53404
rect 13299 53375 13367 53404
rect 13423 53375 13491 53404
rect 13547 53375 13615 53404
rect 13671 53375 13739 53404
rect 13795 53375 13863 53404
rect 13919 53375 13987 53404
rect 14043 53375 14111 53404
rect 12817 53323 12869 53375
rect 12927 53348 12977 53375
rect 13051 53348 13085 53375
rect 13175 53348 13193 53375
rect 13299 53348 13301 53375
rect 12921 53323 12977 53348
rect 13029 53323 13085 53348
rect 13137 53323 13193 53348
rect 13245 53323 13301 53348
rect 13353 53348 13367 53375
rect 13461 53348 13491 53375
rect 13569 53348 13615 53375
rect 13353 53323 13409 53348
rect 13461 53323 13517 53348
rect 13569 53323 13625 53348
rect 13677 53323 13733 53375
rect 13795 53348 13841 53375
rect 13919 53348 13949 53375
rect 14043 53348 14057 53375
rect 13785 53323 13841 53348
rect 13893 53323 13949 53348
rect 14001 53323 14057 53348
rect 14109 53348 14111 53375
rect 14167 53367 14185 53404
rect 14291 53367 14309 53404
rect 14415 53367 14433 53404
rect 14539 53367 14557 53404
rect 14167 53348 14235 53367
rect 14291 53348 14359 53367
rect 14415 53348 14483 53367
rect 14539 53348 14607 53367
rect 14663 53348 14717 53404
rect 14109 53323 14717 53348
rect 12817 53295 14717 53323
rect 12817 53280 14185 53295
rect 14237 53280 14309 53295
rect 14361 53280 14433 53295
rect 14485 53280 14557 53295
rect 14609 53280 14717 53295
rect 12817 53267 12871 53280
rect 12927 53267 12995 53280
rect 13051 53267 13119 53280
rect 13175 53267 13243 53280
rect 13299 53267 13367 53280
rect 13423 53267 13491 53280
rect 13547 53267 13615 53280
rect 13671 53267 13739 53280
rect 13795 53267 13863 53280
rect 13919 53267 13987 53280
rect 14043 53267 14111 53280
rect 12817 53215 12869 53267
rect 12927 53224 12977 53267
rect 13051 53224 13085 53267
rect 13175 53224 13193 53267
rect 13299 53224 13301 53267
rect 12921 53215 12977 53224
rect 13029 53215 13085 53224
rect 13137 53215 13193 53224
rect 13245 53215 13301 53224
rect 13353 53224 13367 53267
rect 13461 53224 13491 53267
rect 13569 53224 13615 53267
rect 13353 53215 13409 53224
rect 13461 53215 13517 53224
rect 13569 53215 13625 53224
rect 13677 53215 13733 53267
rect 13795 53224 13841 53267
rect 13919 53224 13949 53267
rect 14043 53224 14057 53267
rect 13785 53215 13841 53224
rect 13893 53215 13949 53224
rect 14001 53215 14057 53224
rect 14109 53224 14111 53267
rect 14167 53243 14185 53280
rect 14291 53243 14309 53280
rect 14415 53243 14433 53280
rect 14539 53243 14557 53280
rect 14167 53224 14235 53243
rect 14291 53224 14359 53243
rect 14415 53224 14483 53243
rect 14539 53224 14607 53243
rect 14663 53224 14717 53280
rect 14109 53215 14717 53224
rect 12817 53156 14717 53215
rect 12817 53100 12871 53156
rect 12927 53100 12995 53156
rect 13051 53100 13119 53156
rect 13175 53100 13243 53156
rect 13299 53100 13367 53156
rect 13423 53100 13491 53156
rect 13547 53100 13615 53156
rect 13671 53100 13739 53156
rect 13795 53100 13863 53156
rect 13919 53100 13987 53156
rect 14043 53100 14111 53156
rect 14167 53100 14235 53156
rect 14291 53100 14359 53156
rect 14415 53100 14483 53156
rect 14539 53100 14607 53156
rect 14663 53100 14717 53156
rect 12817 53032 14717 53100
rect 12817 52976 12871 53032
rect 12927 52976 12995 53032
rect 13051 52976 13119 53032
rect 13175 52976 13243 53032
rect 13299 52976 13367 53032
rect 13423 52976 13491 53032
rect 13547 52976 13615 53032
rect 13671 52976 13739 53032
rect 13795 52976 13863 53032
rect 13919 52976 13987 53032
rect 14043 52976 14111 53032
rect 14167 52976 14235 53032
rect 14291 52976 14359 53032
rect 14415 52976 14483 53032
rect 14539 52976 14607 53032
rect 14663 52976 14717 53032
rect 12817 52908 14717 52976
rect 12817 52852 12871 52908
rect 12927 52852 12995 52908
rect 13051 52852 13119 52908
rect 13175 52852 13243 52908
rect 13299 52852 13367 52908
rect 13423 52852 13491 52908
rect 13547 52852 13615 52908
rect 13671 52852 13739 52908
rect 13795 52852 13863 52908
rect 13919 52852 13987 52908
rect 14043 52852 14111 52908
rect 14167 52852 14235 52908
rect 14291 52852 14359 52908
rect 14415 52852 14483 52908
rect 14539 52852 14607 52908
rect 14663 52852 14717 52908
rect 12817 52548 14717 52852
rect 14892 54176 14989 54186
rect 14892 52824 14902 54176
rect 14958 52824 14989 54176
rect 14892 52814 14989 52824
rect 12817 52492 12871 52548
rect 12927 52492 12995 52548
rect 13051 52492 13119 52548
rect 13175 52492 13243 52548
rect 13299 52492 13367 52548
rect 13423 52492 13491 52548
rect 13547 52492 13615 52548
rect 13671 52492 13739 52548
rect 13795 52492 13863 52548
rect 13919 52492 13987 52548
rect 14043 52492 14111 52548
rect 14167 52492 14235 52548
rect 14291 52492 14359 52548
rect 14415 52492 14483 52548
rect 14539 52492 14607 52548
rect 14663 52492 14717 52548
rect 12817 52424 14717 52492
rect 12817 52368 12871 52424
rect 12927 52368 12995 52424
rect 13051 52368 13119 52424
rect 13175 52368 13243 52424
rect 13299 52368 13367 52424
rect 13423 52368 13491 52424
rect 13547 52368 13615 52424
rect 13671 52368 13739 52424
rect 13795 52368 13863 52424
rect 13919 52368 13987 52424
rect 14043 52368 14111 52424
rect 14167 52368 14235 52424
rect 14291 52368 14359 52424
rect 14415 52368 14483 52424
rect 14539 52368 14607 52424
rect 14663 52368 14717 52424
rect 12817 52300 14717 52368
rect 12817 52244 12871 52300
rect 12927 52244 12995 52300
rect 13051 52244 13119 52300
rect 13175 52244 13243 52300
rect 13299 52244 13367 52300
rect 13423 52244 13491 52300
rect 13547 52244 13615 52300
rect 13671 52244 13739 52300
rect 13795 52244 13863 52300
rect 13919 52244 13987 52300
rect 14043 52244 14111 52300
rect 14167 52244 14235 52300
rect 14291 52244 14359 52300
rect 14415 52244 14483 52300
rect 14539 52244 14607 52300
rect 14663 52244 14717 52300
rect 12817 52176 14717 52244
rect 12817 52120 12871 52176
rect 12927 52120 12995 52176
rect 13051 52120 13119 52176
rect 13175 52120 13243 52176
rect 13299 52120 13367 52176
rect 13423 52120 13491 52176
rect 13547 52120 13615 52176
rect 13671 52120 13739 52176
rect 13795 52120 13863 52176
rect 13919 52120 13987 52176
rect 14043 52120 14111 52176
rect 14167 52120 14235 52176
rect 14291 52120 14359 52176
rect 14415 52120 14483 52176
rect 14539 52120 14607 52176
rect 14663 52120 14717 52176
rect 12817 52052 14717 52120
rect 12817 51996 12871 52052
rect 12927 51996 12995 52052
rect 13051 51996 13119 52052
rect 13175 51996 13243 52052
rect 13299 51996 13367 52052
rect 13423 51996 13491 52052
rect 13547 51996 13615 52052
rect 13671 51996 13739 52052
rect 13795 51996 13863 52052
rect 13919 51996 13987 52052
rect 14043 51996 14111 52052
rect 14167 51996 14235 52052
rect 14291 51996 14359 52052
rect 14415 51996 14483 52052
rect 14539 51996 14607 52052
rect 14663 51996 14717 52052
rect 12817 51928 14717 51996
rect 12817 51872 12871 51928
rect 12927 51872 12995 51928
rect 13051 51872 13119 51928
rect 13175 51872 13243 51928
rect 13299 51872 13367 51928
rect 13423 51872 13491 51928
rect 13547 51872 13615 51928
rect 13671 51872 13739 51928
rect 13795 51872 13863 51928
rect 13919 51872 13987 51928
rect 14043 51872 14111 51928
rect 14167 51872 14235 51928
rect 14291 51872 14359 51928
rect 14415 51872 14483 51928
rect 14539 51872 14607 51928
rect 14663 51872 14717 51928
rect 12817 51804 14717 51872
rect 12817 51748 12871 51804
rect 12927 51748 12995 51804
rect 13051 51748 13119 51804
rect 13175 51748 13243 51804
rect 13299 51748 13367 51804
rect 13423 51748 13491 51804
rect 13547 51748 13615 51804
rect 13671 51748 13739 51804
rect 13795 51748 13863 51804
rect 13919 51748 13987 51804
rect 14043 51748 14111 51804
rect 14167 51748 14235 51804
rect 14291 51748 14359 51804
rect 14415 51748 14483 51804
rect 14539 51748 14607 51804
rect 14663 51748 14717 51804
rect 12817 51680 14717 51748
rect 12817 51624 12871 51680
rect 12927 51624 12995 51680
rect 13051 51624 13119 51680
rect 13175 51624 13243 51680
rect 13299 51624 13367 51680
rect 13423 51624 13491 51680
rect 13547 51624 13615 51680
rect 13671 51624 13739 51680
rect 13795 51624 13863 51680
rect 13919 51624 13987 51680
rect 14043 51624 14111 51680
rect 14167 51624 14235 51680
rect 14291 51624 14359 51680
rect 14415 51624 14483 51680
rect 14539 51624 14607 51680
rect 14663 51624 14717 51680
rect 12817 51556 14717 51624
rect 12817 51500 12871 51556
rect 12927 51500 12995 51556
rect 13051 51500 13119 51556
rect 13175 51500 13243 51556
rect 13299 51500 13367 51556
rect 13423 51500 13491 51556
rect 13547 51500 13615 51556
rect 13671 51500 13739 51556
rect 13795 51500 13863 51556
rect 13919 51500 13987 51556
rect 14043 51500 14111 51556
rect 14167 51500 14235 51556
rect 14291 51500 14359 51556
rect 14415 51500 14483 51556
rect 14539 51500 14607 51556
rect 14663 51500 14717 51556
rect 12817 51432 14717 51500
rect 12817 51376 12871 51432
rect 12927 51376 12995 51432
rect 13051 51376 13119 51432
rect 13175 51376 13243 51432
rect 13299 51376 13367 51432
rect 13423 51376 13491 51432
rect 13547 51376 13615 51432
rect 13671 51376 13739 51432
rect 13795 51376 13863 51432
rect 13919 51376 13987 51432
rect 14043 51376 14111 51432
rect 14167 51376 14235 51432
rect 14291 51376 14359 51432
rect 14415 51376 14483 51432
rect 14539 51376 14607 51432
rect 14663 51376 14717 51432
rect 12817 51308 14717 51376
rect 12817 51252 12871 51308
rect 12927 51252 12995 51308
rect 13051 51252 13119 51308
rect 13175 51252 13243 51308
rect 13299 51252 13367 51308
rect 13423 51252 13491 51308
rect 13547 51252 13615 51308
rect 13671 51252 13739 51308
rect 13795 51252 13863 51308
rect 13919 51252 13987 51308
rect 14043 51252 14111 51308
rect 14167 51252 14235 51308
rect 14291 51252 14359 51308
rect 14415 51252 14483 51308
rect 14539 51252 14607 51308
rect 14663 51252 14717 51308
rect 12817 49348 14717 51252
rect 14892 52576 14989 52600
rect 14892 51224 14902 52576
rect 14958 51224 14989 52576
rect 14892 51200 14989 51224
rect 12817 49292 12871 49348
rect 12927 49292 12995 49348
rect 13051 49292 13119 49348
rect 13175 49292 13243 49348
rect 13299 49292 13367 49348
rect 13423 49292 13491 49348
rect 13547 49292 13615 49348
rect 13671 49292 13739 49348
rect 13795 49292 13863 49348
rect 13919 49292 13987 49348
rect 14043 49292 14111 49348
rect 14167 49292 14235 49348
rect 14291 49292 14359 49348
rect 14415 49292 14483 49348
rect 14539 49292 14607 49348
rect 14663 49292 14717 49348
rect 12817 49224 14717 49292
rect 12817 49168 12871 49224
rect 12927 49168 12995 49224
rect 13051 49168 13119 49224
rect 13175 49168 13243 49224
rect 13299 49168 13367 49224
rect 13423 49168 13491 49224
rect 13547 49168 13615 49224
rect 13671 49168 13739 49224
rect 13795 49168 13863 49224
rect 13919 49168 13987 49224
rect 14043 49168 14111 49224
rect 14167 49168 14235 49224
rect 14291 49168 14359 49224
rect 14415 49168 14483 49224
rect 14539 49168 14607 49224
rect 14663 49168 14717 49224
rect 12817 49100 14717 49168
rect 12817 49044 12871 49100
rect 12927 49044 12995 49100
rect 13051 49044 13119 49100
rect 13175 49044 13243 49100
rect 13299 49044 13367 49100
rect 13423 49044 13491 49100
rect 13547 49044 13615 49100
rect 13671 49044 13739 49100
rect 13795 49044 13863 49100
rect 13919 49044 13987 49100
rect 14043 49044 14111 49100
rect 14167 49044 14235 49100
rect 14291 49044 14359 49100
rect 14415 49044 14483 49100
rect 14539 49044 14607 49100
rect 14663 49044 14717 49100
rect 12817 48976 14717 49044
rect 12817 48920 12871 48976
rect 12927 48920 12995 48976
rect 13051 48920 13119 48976
rect 13175 48920 13243 48976
rect 13299 48920 13367 48976
rect 13423 48920 13491 48976
rect 13547 48920 13615 48976
rect 13671 48920 13739 48976
rect 13795 48920 13863 48976
rect 13919 48920 13987 48976
rect 14043 48920 14111 48976
rect 14167 48920 14235 48976
rect 14291 48920 14359 48976
rect 14415 48920 14483 48976
rect 14539 48920 14607 48976
rect 14663 48920 14717 48976
rect 12817 48852 14717 48920
rect 12817 48796 12871 48852
rect 12927 48796 12995 48852
rect 13051 48796 13119 48852
rect 13175 48796 13243 48852
rect 13299 48796 13367 48852
rect 13423 48796 13491 48852
rect 13547 48796 13615 48852
rect 13671 48796 13739 48852
rect 13795 48796 13863 48852
rect 13919 48796 13987 48852
rect 14043 48796 14111 48852
rect 14167 48796 14235 48852
rect 14291 48796 14359 48852
rect 14415 48796 14483 48852
rect 14539 48796 14607 48852
rect 14663 48796 14717 48852
rect 12817 48728 14717 48796
rect 12817 48672 12871 48728
rect 12927 48672 12995 48728
rect 13051 48672 13119 48728
rect 13175 48672 13243 48728
rect 13299 48672 13367 48728
rect 13423 48672 13491 48728
rect 13547 48672 13615 48728
rect 13671 48672 13739 48728
rect 13795 48672 13863 48728
rect 13919 48672 13987 48728
rect 14043 48672 14111 48728
rect 14167 48672 14235 48728
rect 14291 48672 14359 48728
rect 14415 48672 14483 48728
rect 14539 48672 14607 48728
rect 14663 48672 14717 48728
rect 12817 48604 14717 48672
rect 12817 48548 12871 48604
rect 12927 48548 12995 48604
rect 13051 48548 13119 48604
rect 13175 48548 13243 48604
rect 13299 48548 13367 48604
rect 13423 48548 13491 48604
rect 13547 48548 13615 48604
rect 13671 48548 13739 48604
rect 13795 48548 13863 48604
rect 13919 48548 13987 48604
rect 14043 48548 14111 48604
rect 14167 48548 14235 48604
rect 14291 48548 14359 48604
rect 14415 48548 14483 48604
rect 14539 48548 14607 48604
rect 14663 48548 14717 48604
rect 12817 48480 14717 48548
rect 12817 48424 12871 48480
rect 12927 48424 12995 48480
rect 13051 48424 13119 48480
rect 13175 48424 13243 48480
rect 13299 48424 13367 48480
rect 13423 48424 13491 48480
rect 13547 48424 13615 48480
rect 13671 48424 13739 48480
rect 13795 48424 13863 48480
rect 13919 48424 13987 48480
rect 14043 48424 14111 48480
rect 14167 48424 14235 48480
rect 14291 48424 14359 48480
rect 14415 48424 14483 48480
rect 14539 48424 14607 48480
rect 14663 48424 14717 48480
rect 12817 48356 14717 48424
rect 12817 48300 12871 48356
rect 12927 48300 12995 48356
rect 13051 48300 13119 48356
rect 13175 48300 13243 48356
rect 13299 48300 13367 48356
rect 13423 48300 13491 48356
rect 13547 48300 13615 48356
rect 13671 48300 13739 48356
rect 13795 48300 13863 48356
rect 13919 48300 13987 48356
rect 14043 48300 14111 48356
rect 14167 48300 14235 48356
rect 14291 48300 14359 48356
rect 14415 48300 14483 48356
rect 14539 48300 14607 48356
rect 14663 48300 14717 48356
rect 12817 48232 14717 48300
rect 12817 48176 12871 48232
rect 12927 48176 12995 48232
rect 13051 48176 13119 48232
rect 13175 48176 13243 48232
rect 13299 48176 13367 48232
rect 13423 48176 13491 48232
rect 13547 48176 13615 48232
rect 13671 48176 13739 48232
rect 13795 48176 13863 48232
rect 13919 48176 13987 48232
rect 14043 48176 14111 48232
rect 14167 48176 14235 48232
rect 14291 48176 14359 48232
rect 14415 48176 14483 48232
rect 14539 48176 14607 48232
rect 14663 48176 14717 48232
rect 12817 48108 14717 48176
rect 12817 48052 12871 48108
rect 12927 48052 12995 48108
rect 13051 48052 13119 48108
rect 13175 48052 13243 48108
rect 13299 48052 13367 48108
rect 13423 48052 13491 48108
rect 13547 48052 13615 48108
rect 13671 48052 13739 48108
rect 13795 48052 13863 48108
rect 13919 48052 13987 48108
rect 14043 48052 14111 48108
rect 14167 48052 14235 48108
rect 14291 48052 14359 48108
rect 14415 48052 14483 48108
rect 14539 48052 14607 48108
rect 14663 48052 14717 48108
rect 12817 47163 14717 48052
rect 14892 49376 14989 49386
rect 14892 48024 14902 49376
rect 14958 48024 14989 49376
rect 14892 48014 14989 48024
rect 12297 47072 12307 47128
rect 12363 47072 12431 47128
rect 12487 47072 12497 47128
rect 12297 47004 12497 47072
rect 12297 46948 12307 47004
rect 12363 46948 12431 47004
rect 12487 46948 12497 47004
rect 12297 46880 12497 46948
rect 12297 46824 12307 46880
rect 12363 46824 12431 46880
rect 12487 46824 12497 46880
rect 12297 46756 12497 46824
rect 12297 46700 12307 46756
rect 12363 46700 12431 46756
rect 12487 46700 12497 46756
rect 12297 46632 12497 46700
rect 12297 46576 12307 46632
rect 12363 46576 12431 46632
rect 12487 46576 12497 46632
rect 12297 46508 12497 46576
rect 12297 46452 12307 46508
rect 12363 46452 12431 46508
rect 12487 46452 12497 46508
rect 12297 46442 12497 46452
rect 14892 46176 14989 46186
rect 2798 46148 4734 46158
rect 2798 46092 2808 46148
rect 2864 46092 2932 46148
rect 2988 46092 3056 46148
rect 3112 46092 3180 46148
rect 3236 46092 3304 46148
rect 3360 46092 3428 46148
rect 3484 46092 3552 46148
rect 3608 46092 3676 46148
rect 3732 46092 3800 46148
rect 3856 46092 3924 46148
rect 3980 46092 4048 46148
rect 4104 46092 4172 46148
rect 4228 46092 4296 46148
rect 4352 46092 4420 46148
rect 4476 46092 4544 46148
rect 4600 46092 4668 46148
rect 4724 46092 4734 46148
rect 2798 46024 4734 46092
rect 2798 45968 2808 46024
rect 2864 45968 2932 46024
rect 2988 45968 3056 46024
rect 3112 45968 3180 46024
rect 3236 45968 3304 46024
rect 3360 45968 3428 46024
rect 3484 45968 3552 46024
rect 3608 45968 3676 46024
rect 3732 45968 3800 46024
rect 3856 45968 3924 46024
rect 3980 45968 4048 46024
rect 4104 45968 4172 46024
rect 4228 45968 4296 46024
rect 4352 45968 4420 46024
rect 4476 45968 4544 46024
rect 4600 45968 4668 46024
rect 4724 45968 4734 46024
rect 2798 45900 4734 45968
rect 2798 45844 2808 45900
rect 2864 45844 2932 45900
rect 2988 45844 3056 45900
rect 3112 45844 3180 45900
rect 3236 45844 3304 45900
rect 3360 45844 3428 45900
rect 3484 45844 3552 45900
rect 3608 45844 3676 45900
rect 3732 45844 3800 45900
rect 3856 45844 3924 45900
rect 3980 45844 4048 45900
rect 4104 45844 4172 45900
rect 4228 45844 4296 45900
rect 4352 45844 4420 45900
rect 4476 45844 4544 45900
rect 4600 45844 4668 45900
rect 4724 45844 4734 45900
rect 2798 45776 4734 45844
rect 2798 45720 2808 45776
rect 2864 45720 2932 45776
rect 2988 45720 3056 45776
rect 3112 45720 3180 45776
rect 3236 45720 3304 45776
rect 3360 45720 3428 45776
rect 3484 45720 3552 45776
rect 3608 45720 3676 45776
rect 3732 45720 3800 45776
rect 3856 45720 3924 45776
rect 3980 45720 4048 45776
rect 4104 45720 4172 45776
rect 4228 45720 4296 45776
rect 4352 45720 4420 45776
rect 4476 45720 4544 45776
rect 4600 45720 4668 45776
rect 4724 45720 4734 45776
rect 2798 45652 4734 45720
rect 2798 45596 2808 45652
rect 2864 45596 2932 45652
rect 2988 45596 3056 45652
rect 3112 45596 3180 45652
rect 3236 45596 3304 45652
rect 3360 45596 3428 45652
rect 3484 45596 3552 45652
rect 3608 45596 3676 45652
rect 3732 45596 3800 45652
rect 3856 45596 3924 45652
rect 3980 45596 4048 45652
rect 4104 45596 4172 45652
rect 4228 45596 4296 45652
rect 4352 45596 4420 45652
rect 4476 45596 4544 45652
rect 4600 45596 4668 45652
rect 4724 45596 4734 45652
rect 2798 45528 4734 45596
rect 2798 45472 2808 45528
rect 2864 45472 2932 45528
rect 2988 45472 3056 45528
rect 3112 45472 3180 45528
rect 3236 45472 3304 45528
rect 3360 45472 3428 45528
rect 3484 45472 3552 45528
rect 3608 45472 3676 45528
rect 3732 45472 3800 45528
rect 3856 45472 3924 45528
rect 3980 45472 4048 45528
rect 4104 45472 4172 45528
rect 4228 45472 4296 45528
rect 4352 45472 4420 45528
rect 4476 45472 4544 45528
rect 4600 45472 4668 45528
rect 4724 45472 4734 45528
rect 2798 45404 4734 45472
rect 2798 45348 2808 45404
rect 2864 45348 2932 45404
rect 2988 45348 3056 45404
rect 3112 45348 3180 45404
rect 3236 45348 3304 45404
rect 3360 45348 3428 45404
rect 3484 45348 3552 45404
rect 3608 45348 3676 45404
rect 3732 45348 3800 45404
rect 3856 45348 3924 45404
rect 3980 45348 4048 45404
rect 4104 45348 4172 45404
rect 4228 45348 4296 45404
rect 4352 45348 4420 45404
rect 4476 45348 4544 45404
rect 4600 45348 4668 45404
rect 4724 45348 4734 45404
rect 2798 45280 4734 45348
rect 2798 45224 2808 45280
rect 2864 45224 2932 45280
rect 2988 45224 3056 45280
rect 3112 45224 3180 45280
rect 3236 45224 3304 45280
rect 3360 45224 3428 45280
rect 3484 45224 3552 45280
rect 3608 45224 3676 45280
rect 3732 45224 3800 45280
rect 3856 45224 3924 45280
rect 3980 45224 4048 45280
rect 4104 45224 4172 45280
rect 4228 45224 4296 45280
rect 4352 45224 4420 45280
rect 4476 45224 4544 45280
rect 4600 45224 4668 45280
rect 4724 45224 4734 45280
rect 2798 45156 4734 45224
rect 2798 45100 2808 45156
rect 2864 45100 2932 45156
rect 2988 45100 3056 45156
rect 3112 45100 3180 45156
rect 3236 45100 3304 45156
rect 3360 45100 3428 45156
rect 3484 45100 3552 45156
rect 3608 45100 3676 45156
rect 3732 45100 3800 45156
rect 3856 45100 3924 45156
rect 3980 45100 4048 45156
rect 4104 45100 4172 45156
rect 4228 45100 4296 45156
rect 4352 45100 4420 45156
rect 4476 45100 4544 45156
rect 4600 45100 4668 45156
rect 4724 45100 4734 45156
rect 2798 45032 4734 45100
rect 2798 44976 2808 45032
rect 2864 44976 2932 45032
rect 2988 44976 3056 45032
rect 3112 44976 3180 45032
rect 3236 44976 3304 45032
rect 3360 44976 3428 45032
rect 3484 44976 3552 45032
rect 3608 44976 3676 45032
rect 3732 44976 3800 45032
rect 3856 44976 3924 45032
rect 3980 44976 4048 45032
rect 4104 44976 4172 45032
rect 4228 44976 4296 45032
rect 4352 44976 4420 45032
rect 4476 44976 4544 45032
rect 4600 44976 4668 45032
rect 4724 44976 4734 45032
rect 2798 44908 4734 44976
rect 2798 44852 2808 44908
rect 2864 44852 2932 44908
rect 2988 44852 3056 44908
rect 3112 44852 3180 44908
rect 3236 44852 3304 44908
rect 3360 44852 3428 44908
rect 3484 44852 3552 44908
rect 3608 44852 3676 44908
rect 3732 44852 3800 44908
rect 3856 44852 3924 44908
rect 3980 44852 4048 44908
rect 4104 44852 4172 44908
rect 4228 44852 4296 44908
rect 4352 44852 4420 44908
rect 4476 44852 4544 44908
rect 4600 44852 4668 44908
rect 4724 44852 4734 44908
rect 2798 44842 4734 44852
rect 5168 46148 7104 46158
rect 5168 46092 5178 46148
rect 5234 46092 5302 46148
rect 5358 46092 5426 46148
rect 5482 46092 5550 46148
rect 5606 46092 5674 46148
rect 5730 46092 5798 46148
rect 5854 46092 5922 46148
rect 5978 46092 6046 46148
rect 6102 46092 6170 46148
rect 6226 46092 6294 46148
rect 6350 46092 6418 46148
rect 6474 46092 6542 46148
rect 6598 46092 6666 46148
rect 6722 46092 6790 46148
rect 6846 46092 6914 46148
rect 6970 46092 7038 46148
rect 7094 46092 7104 46148
rect 5168 46024 7104 46092
rect 5168 45968 5178 46024
rect 5234 45968 5302 46024
rect 5358 45968 5426 46024
rect 5482 45968 5550 46024
rect 5606 45968 5674 46024
rect 5730 45968 5798 46024
rect 5854 45968 5922 46024
rect 5978 45968 6046 46024
rect 6102 45968 6170 46024
rect 6226 45968 6294 46024
rect 6350 45968 6418 46024
rect 6474 45968 6542 46024
rect 6598 45968 6666 46024
rect 6722 45968 6790 46024
rect 6846 45968 6914 46024
rect 6970 45968 7038 46024
rect 7094 45968 7104 46024
rect 5168 45900 7104 45968
rect 5168 45844 5178 45900
rect 5234 45844 5302 45900
rect 5358 45844 5426 45900
rect 5482 45844 5550 45900
rect 5606 45844 5674 45900
rect 5730 45844 5798 45900
rect 5854 45844 5922 45900
rect 5978 45844 6046 45900
rect 6102 45844 6170 45900
rect 6226 45844 6294 45900
rect 6350 45844 6418 45900
rect 6474 45844 6542 45900
rect 6598 45844 6666 45900
rect 6722 45844 6790 45900
rect 6846 45844 6914 45900
rect 6970 45844 7038 45900
rect 7094 45844 7104 45900
rect 5168 45776 7104 45844
rect 5168 45720 5178 45776
rect 5234 45720 5302 45776
rect 5358 45720 5426 45776
rect 5482 45720 5550 45776
rect 5606 45720 5674 45776
rect 5730 45720 5798 45776
rect 5854 45720 5922 45776
rect 5978 45720 6046 45776
rect 6102 45720 6170 45776
rect 6226 45720 6294 45776
rect 6350 45720 6418 45776
rect 6474 45720 6542 45776
rect 6598 45720 6666 45776
rect 6722 45720 6790 45776
rect 6846 45720 6914 45776
rect 6970 45720 7038 45776
rect 7094 45720 7104 45776
rect 5168 45652 7104 45720
rect 5168 45596 5178 45652
rect 5234 45596 5302 45652
rect 5358 45596 5426 45652
rect 5482 45596 5550 45652
rect 5606 45596 5674 45652
rect 5730 45596 5798 45652
rect 5854 45596 5922 45652
rect 5978 45596 6046 45652
rect 6102 45596 6170 45652
rect 6226 45596 6294 45652
rect 6350 45596 6418 45652
rect 6474 45596 6542 45652
rect 6598 45596 6666 45652
rect 6722 45596 6790 45652
rect 6846 45596 6914 45652
rect 6970 45596 7038 45652
rect 7094 45596 7104 45652
rect 5168 45528 7104 45596
rect 5168 45472 5178 45528
rect 5234 45472 5302 45528
rect 5358 45472 5426 45528
rect 5482 45472 5550 45528
rect 5606 45472 5674 45528
rect 5730 45472 5798 45528
rect 5854 45472 5922 45528
rect 5978 45472 6046 45528
rect 6102 45472 6170 45528
rect 6226 45472 6294 45528
rect 6350 45472 6418 45528
rect 6474 45472 6542 45528
rect 6598 45472 6666 45528
rect 6722 45472 6790 45528
rect 6846 45472 6914 45528
rect 6970 45472 7038 45528
rect 7094 45472 7104 45528
rect 5168 45404 7104 45472
rect 5168 45348 5178 45404
rect 5234 45348 5302 45404
rect 5358 45348 5426 45404
rect 5482 45348 5550 45404
rect 5606 45348 5674 45404
rect 5730 45348 5798 45404
rect 5854 45348 5922 45404
rect 5978 45348 6046 45404
rect 6102 45348 6170 45404
rect 6226 45348 6294 45404
rect 6350 45348 6418 45404
rect 6474 45348 6542 45404
rect 6598 45348 6666 45404
rect 6722 45348 6790 45404
rect 6846 45348 6914 45404
rect 6970 45348 7038 45404
rect 7094 45348 7104 45404
rect 5168 45280 7104 45348
rect 5168 45224 5178 45280
rect 5234 45224 5302 45280
rect 5358 45224 5426 45280
rect 5482 45224 5550 45280
rect 5606 45224 5674 45280
rect 5730 45224 5798 45280
rect 5854 45224 5922 45280
rect 5978 45224 6046 45280
rect 6102 45224 6170 45280
rect 6226 45224 6294 45280
rect 6350 45224 6418 45280
rect 6474 45224 6542 45280
rect 6598 45224 6666 45280
rect 6722 45224 6790 45280
rect 6846 45224 6914 45280
rect 6970 45224 7038 45280
rect 7094 45224 7104 45280
rect 5168 45156 7104 45224
rect 5168 45100 5178 45156
rect 5234 45100 5302 45156
rect 5358 45100 5426 45156
rect 5482 45100 5550 45156
rect 5606 45100 5674 45156
rect 5730 45100 5798 45156
rect 5854 45100 5922 45156
rect 5978 45100 6046 45156
rect 6102 45100 6170 45156
rect 6226 45100 6294 45156
rect 6350 45100 6418 45156
rect 6474 45100 6542 45156
rect 6598 45100 6666 45156
rect 6722 45100 6790 45156
rect 6846 45100 6914 45156
rect 6970 45100 7038 45156
rect 7094 45100 7104 45156
rect 5168 45032 7104 45100
rect 5168 44976 5178 45032
rect 5234 44976 5302 45032
rect 5358 44976 5426 45032
rect 5482 44976 5550 45032
rect 5606 44976 5674 45032
rect 5730 44976 5798 45032
rect 5854 44976 5922 45032
rect 5978 44976 6046 45032
rect 6102 44976 6170 45032
rect 6226 44976 6294 45032
rect 6350 44976 6418 45032
rect 6474 44976 6542 45032
rect 6598 44976 6666 45032
rect 6722 44976 6790 45032
rect 6846 44976 6914 45032
rect 6970 44976 7038 45032
rect 7094 44976 7104 45032
rect 5168 44908 7104 44976
rect 5168 44852 5178 44908
rect 5234 44852 5302 44908
rect 5358 44852 5426 44908
rect 5482 44852 5550 44908
rect 5606 44852 5674 44908
rect 5730 44852 5798 44908
rect 5854 44852 5922 44908
rect 5978 44852 6046 44908
rect 6102 44852 6170 44908
rect 6226 44852 6294 44908
rect 6350 44852 6418 44908
rect 6474 44852 6542 44908
rect 6598 44852 6666 44908
rect 6722 44852 6790 44908
rect 6846 44852 6914 44908
rect 6970 44852 7038 44908
rect 7094 44852 7104 44908
rect 5168 44842 7104 44852
rect 7874 46148 9810 46158
rect 7874 46092 7884 46148
rect 7940 46092 8008 46148
rect 8064 46092 8132 46148
rect 8188 46092 8256 46148
rect 8312 46092 8380 46148
rect 8436 46092 8504 46148
rect 8560 46092 8628 46148
rect 8684 46092 8752 46148
rect 8808 46092 8876 46148
rect 8932 46092 9000 46148
rect 9056 46092 9124 46148
rect 9180 46092 9248 46148
rect 9304 46092 9372 46148
rect 9428 46092 9496 46148
rect 9552 46092 9620 46148
rect 9676 46092 9744 46148
rect 9800 46092 9810 46148
rect 7874 46024 9810 46092
rect 7874 45968 7884 46024
rect 7940 45968 8008 46024
rect 8064 45968 8132 46024
rect 8188 45968 8256 46024
rect 8312 45968 8380 46024
rect 8436 45968 8504 46024
rect 8560 45968 8628 46024
rect 8684 45968 8752 46024
rect 8808 45968 8876 46024
rect 8932 45968 9000 46024
rect 9056 45968 9124 46024
rect 9180 45968 9248 46024
rect 9304 45968 9372 46024
rect 9428 45968 9496 46024
rect 9552 45968 9620 46024
rect 9676 45968 9744 46024
rect 9800 45968 9810 46024
rect 7874 45900 9810 45968
rect 7874 45844 7884 45900
rect 7940 45844 8008 45900
rect 8064 45844 8132 45900
rect 8188 45844 8256 45900
rect 8312 45844 8380 45900
rect 8436 45844 8504 45900
rect 8560 45844 8628 45900
rect 8684 45844 8752 45900
rect 8808 45844 8876 45900
rect 8932 45844 9000 45900
rect 9056 45844 9124 45900
rect 9180 45844 9248 45900
rect 9304 45844 9372 45900
rect 9428 45844 9496 45900
rect 9552 45844 9620 45900
rect 9676 45844 9744 45900
rect 9800 45844 9810 45900
rect 7874 45776 9810 45844
rect 7874 45720 7884 45776
rect 7940 45720 8008 45776
rect 8064 45720 8132 45776
rect 8188 45720 8256 45776
rect 8312 45720 8380 45776
rect 8436 45720 8504 45776
rect 8560 45720 8628 45776
rect 8684 45720 8752 45776
rect 8808 45720 8876 45776
rect 8932 45720 9000 45776
rect 9056 45720 9124 45776
rect 9180 45720 9248 45776
rect 9304 45720 9372 45776
rect 9428 45720 9496 45776
rect 9552 45720 9620 45776
rect 9676 45720 9744 45776
rect 9800 45720 9810 45776
rect 7874 45652 9810 45720
rect 7874 45596 7884 45652
rect 7940 45596 8008 45652
rect 8064 45596 8132 45652
rect 8188 45596 8256 45652
rect 8312 45596 8380 45652
rect 8436 45596 8504 45652
rect 8560 45596 8628 45652
rect 8684 45596 8752 45652
rect 8808 45596 8876 45652
rect 8932 45596 9000 45652
rect 9056 45596 9124 45652
rect 9180 45596 9248 45652
rect 9304 45596 9372 45652
rect 9428 45596 9496 45652
rect 9552 45596 9620 45652
rect 9676 45596 9744 45652
rect 9800 45596 9810 45652
rect 7874 45528 9810 45596
rect 7874 45472 7884 45528
rect 7940 45472 8008 45528
rect 8064 45472 8132 45528
rect 8188 45472 8256 45528
rect 8312 45472 8380 45528
rect 8436 45472 8504 45528
rect 8560 45472 8628 45528
rect 8684 45472 8752 45528
rect 8808 45472 8876 45528
rect 8932 45472 9000 45528
rect 9056 45472 9124 45528
rect 9180 45472 9248 45528
rect 9304 45472 9372 45528
rect 9428 45472 9496 45528
rect 9552 45472 9620 45528
rect 9676 45472 9744 45528
rect 9800 45472 9810 45528
rect 7874 45404 9810 45472
rect 7874 45348 7884 45404
rect 7940 45348 8008 45404
rect 8064 45348 8132 45404
rect 8188 45348 8256 45404
rect 8312 45348 8380 45404
rect 8436 45348 8504 45404
rect 8560 45348 8628 45404
rect 8684 45348 8752 45404
rect 8808 45348 8876 45404
rect 8932 45348 9000 45404
rect 9056 45348 9124 45404
rect 9180 45348 9248 45404
rect 9304 45348 9372 45404
rect 9428 45348 9496 45404
rect 9552 45348 9620 45404
rect 9676 45348 9744 45404
rect 9800 45348 9810 45404
rect 7874 45280 9810 45348
rect 7874 45224 7884 45280
rect 7940 45224 8008 45280
rect 8064 45224 8132 45280
rect 8188 45224 8256 45280
rect 8312 45224 8380 45280
rect 8436 45224 8504 45280
rect 8560 45224 8628 45280
rect 8684 45224 8752 45280
rect 8808 45224 8876 45280
rect 8932 45224 9000 45280
rect 9056 45224 9124 45280
rect 9180 45224 9248 45280
rect 9304 45224 9372 45280
rect 9428 45224 9496 45280
rect 9552 45224 9620 45280
rect 9676 45224 9744 45280
rect 9800 45224 9810 45280
rect 7874 45156 9810 45224
rect 7874 45100 7884 45156
rect 7940 45100 8008 45156
rect 8064 45100 8132 45156
rect 8188 45100 8256 45156
rect 8312 45100 8380 45156
rect 8436 45100 8504 45156
rect 8560 45100 8628 45156
rect 8684 45100 8752 45156
rect 8808 45100 8876 45156
rect 8932 45100 9000 45156
rect 9056 45100 9124 45156
rect 9180 45100 9248 45156
rect 9304 45100 9372 45156
rect 9428 45100 9496 45156
rect 9552 45100 9620 45156
rect 9676 45100 9744 45156
rect 9800 45100 9810 45156
rect 7874 45032 9810 45100
rect 7874 44976 7884 45032
rect 7940 44976 8008 45032
rect 8064 44976 8132 45032
rect 8188 44976 8256 45032
rect 8312 44976 8380 45032
rect 8436 44976 8504 45032
rect 8560 44976 8628 45032
rect 8684 44976 8752 45032
rect 8808 44976 8876 45032
rect 8932 44976 9000 45032
rect 9056 44976 9124 45032
rect 9180 44976 9248 45032
rect 9304 44976 9372 45032
rect 9428 44976 9496 45032
rect 9552 44976 9620 45032
rect 9676 44976 9744 45032
rect 9800 44976 9810 45032
rect 7874 44908 9810 44976
rect 7874 44852 7884 44908
rect 7940 44852 8008 44908
rect 8064 44852 8132 44908
rect 8188 44852 8256 44908
rect 8312 44852 8380 44908
rect 8436 44852 8504 44908
rect 8560 44852 8628 44908
rect 8684 44852 8752 44908
rect 8808 44852 8876 44908
rect 8932 44852 9000 44908
rect 9056 44852 9124 44908
rect 9180 44852 9248 44908
rect 9304 44852 9372 44908
rect 9428 44852 9496 44908
rect 9552 44852 9620 44908
rect 9676 44852 9744 44908
rect 9800 44852 9810 44908
rect 7874 44842 9810 44852
rect 10244 46148 12180 46158
rect 10244 46092 10254 46148
rect 10310 46092 10378 46148
rect 10434 46092 10502 46148
rect 10558 46092 10626 46148
rect 10682 46092 10750 46148
rect 10806 46092 10874 46148
rect 10930 46092 10998 46148
rect 11054 46092 11122 46148
rect 11178 46092 11246 46148
rect 11302 46092 11370 46148
rect 11426 46092 11494 46148
rect 11550 46092 11618 46148
rect 11674 46092 11742 46148
rect 11798 46092 11866 46148
rect 11922 46092 11990 46148
rect 12046 46092 12114 46148
rect 12170 46092 12180 46148
rect 10244 46024 12180 46092
rect 10244 45968 10254 46024
rect 10310 45968 10378 46024
rect 10434 45968 10502 46024
rect 10558 45968 10626 46024
rect 10682 45968 10750 46024
rect 10806 45968 10874 46024
rect 10930 45968 10998 46024
rect 11054 45968 11122 46024
rect 11178 45968 11246 46024
rect 11302 45968 11370 46024
rect 11426 45968 11494 46024
rect 11550 45968 11618 46024
rect 11674 45968 11742 46024
rect 11798 45968 11866 46024
rect 11922 45968 11990 46024
rect 12046 45968 12114 46024
rect 12170 45968 12180 46024
rect 10244 45900 12180 45968
rect 10244 45844 10254 45900
rect 10310 45844 10378 45900
rect 10434 45844 10502 45900
rect 10558 45844 10626 45900
rect 10682 45844 10750 45900
rect 10806 45844 10874 45900
rect 10930 45844 10998 45900
rect 11054 45844 11122 45900
rect 11178 45844 11246 45900
rect 11302 45844 11370 45900
rect 11426 45844 11494 45900
rect 11550 45844 11618 45900
rect 11674 45844 11742 45900
rect 11798 45844 11866 45900
rect 11922 45844 11990 45900
rect 12046 45844 12114 45900
rect 12170 45844 12180 45900
rect 10244 45776 12180 45844
rect 10244 45720 10254 45776
rect 10310 45720 10378 45776
rect 10434 45720 10502 45776
rect 10558 45720 10626 45776
rect 10682 45720 10750 45776
rect 10806 45720 10874 45776
rect 10930 45720 10998 45776
rect 11054 45720 11122 45776
rect 11178 45720 11246 45776
rect 11302 45720 11370 45776
rect 11426 45720 11494 45776
rect 11550 45720 11618 45776
rect 11674 45720 11742 45776
rect 11798 45720 11866 45776
rect 11922 45720 11990 45776
rect 12046 45720 12114 45776
rect 12170 45720 12180 45776
rect 10244 45652 12180 45720
rect 10244 45596 10254 45652
rect 10310 45596 10378 45652
rect 10434 45596 10502 45652
rect 10558 45596 10626 45652
rect 10682 45596 10750 45652
rect 10806 45596 10874 45652
rect 10930 45596 10998 45652
rect 11054 45596 11122 45652
rect 11178 45596 11246 45652
rect 11302 45596 11370 45652
rect 11426 45596 11494 45652
rect 11550 45596 11618 45652
rect 11674 45596 11742 45652
rect 11798 45596 11866 45652
rect 11922 45596 11990 45652
rect 12046 45596 12114 45652
rect 12170 45596 12180 45652
rect 10244 45528 12180 45596
rect 10244 45472 10254 45528
rect 10310 45472 10378 45528
rect 10434 45472 10502 45528
rect 10558 45472 10626 45528
rect 10682 45472 10750 45528
rect 10806 45472 10874 45528
rect 10930 45472 10998 45528
rect 11054 45472 11122 45528
rect 11178 45472 11246 45528
rect 11302 45472 11370 45528
rect 11426 45472 11494 45528
rect 11550 45472 11618 45528
rect 11674 45472 11742 45528
rect 11798 45472 11866 45528
rect 11922 45472 11990 45528
rect 12046 45472 12114 45528
rect 12170 45472 12180 45528
rect 10244 45404 12180 45472
rect 10244 45348 10254 45404
rect 10310 45348 10378 45404
rect 10434 45348 10502 45404
rect 10558 45348 10626 45404
rect 10682 45348 10750 45404
rect 10806 45348 10874 45404
rect 10930 45348 10998 45404
rect 11054 45348 11122 45404
rect 11178 45348 11246 45404
rect 11302 45348 11370 45404
rect 11426 45348 11494 45404
rect 11550 45348 11618 45404
rect 11674 45348 11742 45404
rect 11798 45348 11866 45404
rect 11922 45348 11990 45404
rect 12046 45348 12114 45404
rect 12170 45348 12180 45404
rect 10244 45280 12180 45348
rect 10244 45224 10254 45280
rect 10310 45224 10378 45280
rect 10434 45224 10502 45280
rect 10558 45224 10626 45280
rect 10682 45224 10750 45280
rect 10806 45224 10874 45280
rect 10930 45224 10998 45280
rect 11054 45224 11122 45280
rect 11178 45224 11246 45280
rect 11302 45224 11370 45280
rect 11426 45224 11494 45280
rect 11550 45224 11618 45280
rect 11674 45224 11742 45280
rect 11798 45224 11866 45280
rect 11922 45224 11990 45280
rect 12046 45224 12114 45280
rect 12170 45224 12180 45280
rect 10244 45156 12180 45224
rect 10244 45100 10254 45156
rect 10310 45100 10378 45156
rect 10434 45100 10502 45156
rect 10558 45100 10626 45156
rect 10682 45100 10750 45156
rect 10806 45100 10874 45156
rect 10930 45100 10998 45156
rect 11054 45100 11122 45156
rect 11178 45100 11246 45156
rect 11302 45100 11370 45156
rect 11426 45100 11494 45156
rect 11550 45100 11618 45156
rect 11674 45100 11742 45156
rect 11798 45100 11866 45156
rect 11922 45100 11990 45156
rect 12046 45100 12114 45156
rect 12170 45100 12180 45156
rect 10244 45032 12180 45100
rect 10244 44976 10254 45032
rect 10310 44976 10378 45032
rect 10434 44976 10502 45032
rect 10558 44976 10626 45032
rect 10682 44976 10750 45032
rect 10806 44976 10874 45032
rect 10930 44976 10998 45032
rect 11054 44976 11122 45032
rect 11178 44976 11246 45032
rect 11302 44976 11370 45032
rect 11426 44976 11494 45032
rect 11550 44976 11618 45032
rect 11674 44976 11742 45032
rect 11798 44976 11866 45032
rect 11922 44976 11990 45032
rect 12046 44976 12114 45032
rect 12170 44976 12180 45032
rect 10244 44908 12180 44976
rect 10244 44852 10254 44908
rect 10310 44852 10378 44908
rect 10434 44852 10502 44908
rect 10558 44852 10626 44908
rect 10682 44852 10750 44908
rect 10806 44852 10874 44908
rect 10930 44852 10998 44908
rect 11054 44852 11122 44908
rect 11178 44852 11246 44908
rect 11302 44852 11370 44908
rect 11426 44852 11494 44908
rect 11550 44852 11618 44908
rect 11674 44852 11742 44908
rect 11798 44852 11866 44908
rect 11922 44852 11990 44908
rect 12046 44852 12114 44908
rect 12170 44852 12180 44908
rect 10244 44842 12180 44852
rect 12861 46148 14673 46158
rect 12861 46092 12871 46148
rect 12927 46092 12995 46148
rect 13051 46092 13119 46148
rect 13175 46092 13243 46148
rect 13299 46092 13367 46148
rect 13423 46092 13491 46148
rect 13547 46092 13615 46148
rect 13671 46092 13739 46148
rect 13795 46092 13863 46148
rect 13919 46092 13987 46148
rect 14043 46092 14111 46148
rect 14167 46092 14235 46148
rect 14291 46092 14359 46148
rect 14415 46092 14483 46148
rect 14539 46092 14607 46148
rect 14663 46092 14673 46148
rect 12861 46024 14673 46092
rect 12861 45968 12871 46024
rect 12927 45968 12995 46024
rect 13051 45968 13119 46024
rect 13175 45968 13243 46024
rect 13299 45968 13367 46024
rect 13423 45968 13491 46024
rect 13547 45968 13615 46024
rect 13671 45968 13739 46024
rect 13795 45968 13863 46024
rect 13919 45968 13987 46024
rect 14043 45968 14111 46024
rect 14167 45968 14235 46024
rect 14291 45968 14359 46024
rect 14415 45968 14483 46024
rect 14539 45968 14607 46024
rect 14663 45968 14673 46024
rect 12861 45900 14673 45968
rect 12861 45844 12871 45900
rect 12927 45844 12995 45900
rect 13051 45844 13119 45900
rect 13175 45844 13243 45900
rect 13299 45844 13367 45900
rect 13423 45844 13491 45900
rect 13547 45844 13615 45900
rect 13671 45844 13739 45900
rect 13795 45844 13863 45900
rect 13919 45844 13987 45900
rect 14043 45844 14111 45900
rect 14167 45844 14235 45900
rect 14291 45844 14359 45900
rect 14415 45844 14483 45900
rect 14539 45844 14607 45900
rect 14663 45844 14673 45900
rect 12861 45776 14673 45844
rect 12861 45720 12871 45776
rect 12927 45720 12995 45776
rect 13051 45720 13119 45776
rect 13175 45720 13243 45776
rect 13299 45720 13367 45776
rect 13423 45720 13491 45776
rect 13547 45720 13615 45776
rect 13671 45720 13739 45776
rect 13795 45720 13863 45776
rect 13919 45720 13987 45776
rect 14043 45720 14111 45776
rect 14167 45720 14235 45776
rect 14291 45720 14359 45776
rect 14415 45720 14483 45776
rect 14539 45720 14607 45776
rect 14663 45720 14673 45776
rect 12861 45652 14673 45720
rect 12861 45596 12871 45652
rect 12927 45596 12995 45652
rect 13051 45596 13119 45652
rect 13175 45596 13243 45652
rect 13299 45596 13367 45652
rect 13423 45596 13491 45652
rect 13547 45596 13615 45652
rect 13671 45596 13739 45652
rect 13795 45596 13863 45652
rect 13919 45596 13987 45652
rect 14043 45596 14111 45652
rect 14167 45596 14235 45652
rect 14291 45596 14359 45652
rect 14415 45596 14483 45652
rect 14539 45596 14607 45652
rect 14663 45596 14673 45652
rect 12861 45528 14673 45596
rect 12861 45472 12871 45528
rect 12927 45472 12995 45528
rect 13051 45472 13119 45528
rect 13175 45472 13243 45528
rect 13299 45472 13367 45528
rect 13423 45472 13491 45528
rect 13547 45472 13615 45528
rect 13671 45472 13739 45528
rect 13795 45472 13863 45528
rect 13919 45472 13987 45528
rect 14043 45472 14111 45528
rect 14167 45472 14235 45528
rect 14291 45472 14359 45528
rect 14415 45472 14483 45528
rect 14539 45472 14607 45528
rect 14663 45472 14673 45528
rect 12861 45404 14673 45472
rect 12861 45348 12871 45404
rect 12927 45348 12995 45404
rect 13051 45348 13119 45404
rect 13175 45348 13243 45404
rect 13299 45348 13367 45404
rect 13423 45348 13491 45404
rect 13547 45348 13615 45404
rect 13671 45348 13739 45404
rect 13795 45348 13863 45404
rect 13919 45348 13987 45404
rect 14043 45348 14111 45404
rect 14167 45348 14235 45404
rect 14291 45348 14359 45404
rect 14415 45348 14483 45404
rect 14539 45348 14607 45404
rect 14663 45348 14673 45404
rect 12861 45280 14673 45348
rect 12861 45224 12871 45280
rect 12927 45224 12995 45280
rect 13051 45224 13119 45280
rect 13175 45224 13243 45280
rect 13299 45224 13367 45280
rect 13423 45224 13491 45280
rect 13547 45224 13615 45280
rect 13671 45224 13739 45280
rect 13795 45224 13863 45280
rect 13919 45224 13987 45280
rect 14043 45224 14111 45280
rect 14167 45224 14235 45280
rect 14291 45224 14359 45280
rect 14415 45224 14483 45280
rect 14539 45224 14607 45280
rect 14663 45224 14673 45280
rect 12861 45156 14673 45224
rect 12861 45100 12871 45156
rect 12927 45100 12995 45156
rect 13051 45100 13119 45156
rect 13175 45100 13243 45156
rect 13299 45100 13367 45156
rect 13423 45100 13491 45156
rect 13547 45100 13615 45156
rect 13671 45100 13739 45156
rect 13795 45100 13863 45156
rect 13919 45100 13987 45156
rect 14043 45100 14111 45156
rect 14167 45100 14235 45156
rect 14291 45100 14359 45156
rect 14415 45100 14483 45156
rect 14539 45100 14607 45156
rect 14663 45100 14673 45156
rect 12861 45032 14673 45100
rect 12861 44976 12871 45032
rect 12927 44976 12995 45032
rect 13051 44976 13119 45032
rect 13175 44976 13243 45032
rect 13299 44976 13367 45032
rect 13423 44976 13491 45032
rect 13547 44976 13615 45032
rect 13671 44976 13739 45032
rect 13795 44976 13863 45032
rect 13919 44976 13987 45032
rect 14043 44976 14111 45032
rect 14167 44976 14235 45032
rect 14291 44976 14359 45032
rect 14415 44976 14483 45032
rect 14539 44976 14607 45032
rect 14663 44976 14673 45032
rect 12861 44908 14673 44976
rect 12861 44852 12871 44908
rect 12927 44852 12995 44908
rect 13051 44852 13119 44908
rect 13175 44852 13243 44908
rect 13299 44852 13367 44908
rect 13423 44852 13491 44908
rect 13547 44852 13615 44908
rect 13671 44852 13739 44908
rect 13795 44852 13863 44908
rect 13919 44852 13987 44908
rect 14043 44852 14111 44908
rect 14167 44852 14235 44908
rect 14291 44852 14359 44908
rect 14415 44852 14483 44908
rect 14539 44852 14607 44908
rect 14663 44852 14673 44908
rect 12861 44842 14673 44852
rect 14892 44824 14902 46176
rect 14958 44824 14989 46176
rect 14892 44814 14989 44824
rect 2481 44548 2681 44558
rect 2481 44492 2491 44548
rect 2547 44492 2615 44548
rect 2671 44492 2681 44548
rect 2481 44424 2681 44492
rect 2481 44368 2491 44424
rect 2547 44368 2615 44424
rect 2671 44368 2681 44424
rect 2481 44300 2681 44368
rect 2481 44244 2491 44300
rect 2547 44244 2615 44300
rect 2671 44244 2681 44300
rect 2481 44176 2681 44244
rect 2481 44120 2491 44176
rect 2547 44120 2615 44176
rect 2671 44120 2681 44176
rect 2481 44052 2681 44120
rect 2481 43996 2491 44052
rect 2547 43996 2615 44052
rect 2671 43996 2681 44052
rect 2481 43928 2681 43996
rect 2481 43872 2491 43928
rect 2547 43872 2615 43928
rect 2671 43872 2681 43928
rect 2481 43804 2681 43872
rect 2481 43748 2491 43804
rect 2547 43748 2615 43804
rect 2671 43748 2681 43804
rect 2481 43680 2681 43748
rect 2481 43624 2491 43680
rect 2547 43624 2615 43680
rect 2671 43624 2681 43680
rect 2481 43556 2681 43624
rect 2481 43500 2491 43556
rect 2547 43500 2615 43556
rect 2671 43500 2681 43556
rect 2481 43432 2681 43500
rect 2481 43376 2491 43432
rect 2547 43376 2615 43432
rect 2671 43376 2681 43432
rect 2481 43308 2681 43376
rect 2481 43252 2491 43308
rect 2547 43252 2615 43308
rect 2671 43252 2681 43308
rect 2481 43242 2681 43252
rect 4851 44548 5051 44558
rect 4851 44492 4861 44548
rect 4917 44492 4985 44548
rect 5041 44492 5051 44548
rect 4851 44424 5051 44492
rect 4851 44368 4861 44424
rect 4917 44368 4985 44424
rect 5041 44368 5051 44424
rect 4851 44300 5051 44368
rect 4851 44244 4861 44300
rect 4917 44244 4985 44300
rect 5041 44244 5051 44300
rect 4851 44176 5051 44244
rect 4851 44120 4861 44176
rect 4917 44120 4985 44176
rect 5041 44120 5051 44176
rect 4851 44052 5051 44120
rect 4851 43996 4861 44052
rect 4917 43996 4985 44052
rect 5041 43996 5051 44052
rect 4851 43928 5051 43996
rect 4851 43872 4861 43928
rect 4917 43872 4985 43928
rect 5041 43872 5051 43928
rect 4851 43804 5051 43872
rect 4851 43748 4861 43804
rect 4917 43748 4985 43804
rect 5041 43748 5051 43804
rect 4851 43680 5051 43748
rect 4851 43624 4861 43680
rect 4917 43624 4985 43680
rect 5041 43624 5051 43680
rect 4851 43556 5051 43624
rect 4851 43500 4861 43556
rect 4917 43500 4985 43556
rect 5041 43500 5051 43556
rect 4851 43432 5051 43500
rect 4851 43376 4861 43432
rect 4917 43376 4985 43432
rect 5041 43376 5051 43432
rect 4851 43308 5051 43376
rect 4851 43252 4861 43308
rect 4917 43252 4985 43308
rect 5041 43252 5051 43308
rect 4851 43242 5051 43252
rect 7265 44548 7713 44558
rect 7265 44492 7275 44548
rect 7331 44492 7399 44548
rect 7455 44492 7523 44548
rect 7579 44492 7647 44548
rect 7703 44492 7713 44548
rect 7265 44424 7713 44492
rect 7265 44368 7275 44424
rect 7331 44368 7399 44424
rect 7455 44368 7523 44424
rect 7579 44368 7647 44424
rect 7703 44368 7713 44424
rect 7265 44300 7713 44368
rect 7265 44244 7275 44300
rect 7331 44244 7399 44300
rect 7455 44244 7523 44300
rect 7579 44244 7647 44300
rect 7703 44244 7713 44300
rect 7265 44176 7713 44244
rect 7265 44120 7275 44176
rect 7331 44120 7399 44176
rect 7455 44120 7523 44176
rect 7579 44120 7647 44176
rect 7703 44120 7713 44176
rect 7265 44052 7713 44120
rect 7265 43996 7275 44052
rect 7331 43996 7399 44052
rect 7455 43996 7523 44052
rect 7579 43996 7647 44052
rect 7703 43996 7713 44052
rect 7265 43928 7713 43996
rect 7265 43872 7275 43928
rect 7331 43872 7399 43928
rect 7455 43872 7523 43928
rect 7579 43872 7647 43928
rect 7703 43872 7713 43928
rect 7265 43804 7713 43872
rect 7265 43748 7275 43804
rect 7331 43748 7399 43804
rect 7455 43748 7523 43804
rect 7579 43748 7647 43804
rect 7703 43748 7713 43804
rect 7265 43680 7713 43748
rect 7265 43624 7275 43680
rect 7331 43624 7399 43680
rect 7455 43624 7523 43680
rect 7579 43624 7647 43680
rect 7703 43624 7713 43680
rect 7265 43556 7713 43624
rect 7265 43500 7275 43556
rect 7331 43500 7399 43556
rect 7455 43500 7523 43556
rect 7579 43500 7647 43556
rect 7703 43500 7713 43556
rect 7265 43432 7713 43500
rect 7265 43376 7275 43432
rect 7331 43376 7399 43432
rect 7455 43376 7523 43432
rect 7579 43376 7647 43432
rect 7703 43376 7713 43432
rect 7265 43308 7713 43376
rect 7265 43252 7275 43308
rect 7331 43252 7399 43308
rect 7455 43252 7523 43308
rect 7579 43252 7647 43308
rect 7703 43252 7713 43308
rect 7265 43242 7713 43252
rect 9927 44548 10127 44558
rect 9927 44492 9937 44548
rect 9993 44492 10061 44548
rect 10117 44492 10127 44548
rect 9927 44424 10127 44492
rect 9927 44368 9937 44424
rect 9993 44368 10061 44424
rect 10117 44368 10127 44424
rect 9927 44300 10127 44368
rect 9927 44244 9937 44300
rect 9993 44244 10061 44300
rect 10117 44244 10127 44300
rect 9927 44176 10127 44244
rect 9927 44120 9937 44176
rect 9993 44120 10061 44176
rect 10117 44120 10127 44176
rect 9927 44052 10127 44120
rect 9927 43996 9937 44052
rect 9993 43996 10061 44052
rect 10117 43996 10127 44052
rect 9927 43928 10127 43996
rect 9927 43872 9937 43928
rect 9993 43872 10061 43928
rect 10117 43872 10127 43928
rect 9927 43804 10127 43872
rect 9927 43748 9937 43804
rect 9993 43748 10061 43804
rect 10117 43748 10127 43804
rect 9927 43680 10127 43748
rect 9927 43624 9937 43680
rect 9993 43624 10061 43680
rect 10117 43624 10127 43680
rect 9927 43556 10127 43624
rect 9927 43500 9937 43556
rect 9993 43500 10061 43556
rect 10117 43500 10127 43556
rect 9927 43432 10127 43500
rect 9927 43376 9937 43432
rect 9993 43376 10061 43432
rect 10117 43376 10127 43432
rect 9927 43308 10127 43376
rect 9927 43252 9937 43308
rect 9993 43252 10061 43308
rect 10117 43252 10127 43308
rect 9927 43242 10127 43252
rect 12297 44548 12497 44558
rect 12297 44492 12307 44548
rect 12363 44492 12431 44548
rect 12487 44492 12497 44548
rect 12297 44424 12497 44492
rect 12297 44368 12307 44424
rect 12363 44368 12431 44424
rect 12487 44368 12497 44424
rect 12297 44300 12497 44368
rect 12297 44244 12307 44300
rect 12363 44244 12431 44300
rect 12487 44244 12497 44300
rect 12297 44176 12497 44244
rect 12297 44120 12307 44176
rect 12363 44120 12431 44176
rect 12487 44120 12497 44176
rect 12297 44052 12497 44120
rect 12297 43996 12307 44052
rect 12363 43996 12431 44052
rect 12487 43996 12497 44052
rect 12297 43928 12497 43996
rect 12297 43872 12307 43928
rect 12363 43872 12431 43928
rect 12487 43872 12497 43928
rect 12297 43804 12497 43872
rect 12297 43748 12307 43804
rect 12363 43748 12431 43804
rect 12487 43748 12497 43804
rect 12297 43680 12497 43748
rect 12297 43624 12307 43680
rect 12363 43624 12431 43680
rect 12487 43624 12497 43680
rect 12297 43556 12497 43624
rect 12297 43500 12307 43556
rect 12363 43500 12431 43556
rect 12487 43500 12497 43556
rect 12297 43432 12497 43500
rect 12297 43376 12307 43432
rect 12363 43376 12431 43432
rect 12487 43376 12497 43432
rect 12297 43308 12497 43376
rect 12297 43252 12307 43308
rect 12363 43252 12431 43308
rect 12487 43252 12497 43308
rect 12297 43242 12497 43252
rect 2481 42948 2681 42958
rect 2481 42892 2491 42948
rect 2547 42892 2615 42948
rect 2671 42892 2681 42948
rect 2481 42824 2681 42892
rect 2481 42768 2491 42824
rect 2547 42768 2615 42824
rect 2671 42768 2681 42824
rect 2481 42700 2681 42768
rect 2481 42644 2491 42700
rect 2547 42644 2615 42700
rect 2671 42644 2681 42700
rect 2481 42576 2681 42644
rect 2481 42520 2491 42576
rect 2547 42520 2615 42576
rect 2671 42520 2681 42576
rect 2481 42452 2681 42520
rect 2481 42396 2491 42452
rect 2547 42396 2615 42452
rect 2671 42396 2681 42452
rect 2481 42328 2681 42396
rect 2481 42272 2491 42328
rect 2547 42272 2615 42328
rect 2671 42272 2681 42328
rect 2481 42204 2681 42272
rect 2481 42148 2491 42204
rect 2547 42148 2615 42204
rect 2671 42148 2681 42204
rect 2481 42080 2681 42148
rect 2481 42024 2491 42080
rect 2547 42024 2615 42080
rect 2671 42024 2681 42080
rect 2481 41956 2681 42024
rect 2481 41900 2491 41956
rect 2547 41900 2615 41956
rect 2671 41900 2681 41956
rect 2481 41832 2681 41900
rect 2481 41776 2491 41832
rect 2547 41776 2615 41832
rect 2671 41776 2681 41832
rect 2481 41708 2681 41776
rect 2481 41652 2491 41708
rect 2547 41652 2615 41708
rect 2671 41652 2681 41708
rect 2481 41642 2681 41652
rect 4851 42948 5051 42958
rect 4851 42892 4861 42948
rect 4917 42892 4985 42948
rect 5041 42892 5051 42948
rect 4851 42824 5051 42892
rect 4851 42768 4861 42824
rect 4917 42768 4985 42824
rect 5041 42768 5051 42824
rect 4851 42700 5051 42768
rect 4851 42644 4861 42700
rect 4917 42644 4985 42700
rect 5041 42644 5051 42700
rect 4851 42576 5051 42644
rect 4851 42520 4861 42576
rect 4917 42520 4985 42576
rect 5041 42520 5051 42576
rect 4851 42452 5051 42520
rect 4851 42396 4861 42452
rect 4917 42396 4985 42452
rect 5041 42396 5051 42452
rect 4851 42328 5051 42396
rect 4851 42272 4861 42328
rect 4917 42272 4985 42328
rect 5041 42272 5051 42328
rect 4851 42204 5051 42272
rect 4851 42148 4861 42204
rect 4917 42148 4985 42204
rect 5041 42148 5051 42204
rect 4851 42080 5051 42148
rect 4851 42024 4861 42080
rect 4917 42024 4985 42080
rect 5041 42024 5051 42080
rect 4851 41956 5051 42024
rect 4851 41900 4861 41956
rect 4917 41900 4985 41956
rect 5041 41900 5051 41956
rect 4851 41832 5051 41900
rect 4851 41776 4861 41832
rect 4917 41776 4985 41832
rect 5041 41776 5051 41832
rect 4851 41708 5051 41776
rect 4851 41652 4861 41708
rect 4917 41652 4985 41708
rect 5041 41652 5051 41708
rect 4851 41642 5051 41652
rect 7265 42948 7713 42958
rect 7265 42892 7275 42948
rect 7331 42892 7399 42948
rect 7455 42892 7523 42948
rect 7579 42892 7647 42948
rect 7703 42892 7713 42948
rect 7265 42824 7713 42892
rect 7265 42768 7275 42824
rect 7331 42768 7399 42824
rect 7455 42768 7523 42824
rect 7579 42768 7647 42824
rect 7703 42768 7713 42824
rect 7265 42700 7713 42768
rect 7265 42644 7275 42700
rect 7331 42644 7399 42700
rect 7455 42644 7523 42700
rect 7579 42644 7647 42700
rect 7703 42644 7713 42700
rect 7265 42576 7713 42644
rect 7265 42520 7275 42576
rect 7331 42520 7399 42576
rect 7455 42520 7523 42576
rect 7579 42520 7647 42576
rect 7703 42520 7713 42576
rect 7265 42452 7713 42520
rect 7265 42396 7275 42452
rect 7331 42396 7399 42452
rect 7455 42396 7523 42452
rect 7579 42396 7647 42452
rect 7703 42396 7713 42452
rect 7265 42328 7713 42396
rect 7265 42272 7275 42328
rect 7331 42272 7399 42328
rect 7455 42272 7523 42328
rect 7579 42272 7647 42328
rect 7703 42272 7713 42328
rect 7265 42204 7713 42272
rect 7265 42148 7275 42204
rect 7331 42148 7399 42204
rect 7455 42148 7523 42204
rect 7579 42148 7647 42204
rect 7703 42148 7713 42204
rect 7265 42080 7713 42148
rect 7265 42024 7275 42080
rect 7331 42024 7399 42080
rect 7455 42024 7523 42080
rect 7579 42024 7647 42080
rect 7703 42024 7713 42080
rect 7265 41956 7713 42024
rect 7265 41900 7275 41956
rect 7331 41900 7399 41956
rect 7455 41900 7523 41956
rect 7579 41900 7647 41956
rect 7703 41900 7713 41956
rect 7265 41832 7713 41900
rect 7265 41776 7275 41832
rect 7331 41776 7399 41832
rect 7455 41776 7523 41832
rect 7579 41776 7647 41832
rect 7703 41776 7713 41832
rect 7265 41708 7713 41776
rect 7265 41652 7275 41708
rect 7331 41652 7399 41708
rect 7455 41652 7523 41708
rect 7579 41652 7647 41708
rect 7703 41652 7713 41708
rect 7265 41642 7713 41652
rect 9927 42948 10127 42958
rect 9927 42892 9937 42948
rect 9993 42892 10061 42948
rect 10117 42892 10127 42948
rect 9927 42824 10127 42892
rect 9927 42768 9937 42824
rect 9993 42768 10061 42824
rect 10117 42768 10127 42824
rect 9927 42700 10127 42768
rect 9927 42644 9937 42700
rect 9993 42644 10061 42700
rect 10117 42644 10127 42700
rect 9927 42576 10127 42644
rect 9927 42520 9937 42576
rect 9993 42520 10061 42576
rect 10117 42520 10127 42576
rect 9927 42452 10127 42520
rect 9927 42396 9937 42452
rect 9993 42396 10061 42452
rect 10117 42396 10127 42452
rect 9927 42328 10127 42396
rect 9927 42272 9937 42328
rect 9993 42272 10061 42328
rect 10117 42272 10127 42328
rect 9927 42204 10127 42272
rect 9927 42148 9937 42204
rect 9993 42148 10061 42204
rect 10117 42148 10127 42204
rect 9927 42080 10127 42148
rect 9927 42024 9937 42080
rect 9993 42024 10061 42080
rect 10117 42024 10127 42080
rect 9927 41956 10127 42024
rect 9927 41900 9937 41956
rect 9993 41900 10061 41956
rect 10117 41900 10127 41956
rect 9927 41832 10127 41900
rect 9927 41776 9937 41832
rect 9993 41776 10061 41832
rect 10117 41776 10127 41832
rect 9927 41708 10127 41776
rect 9927 41652 9937 41708
rect 9993 41652 10061 41708
rect 10117 41652 10127 41708
rect 9927 41642 10127 41652
rect 12297 42948 12497 42958
rect 12297 42892 12307 42948
rect 12363 42892 12431 42948
rect 12487 42892 12497 42948
rect 12297 42824 12497 42892
rect 12297 42768 12307 42824
rect 12363 42768 12431 42824
rect 12487 42768 12497 42824
rect 12297 42700 12497 42768
rect 12297 42644 12307 42700
rect 12363 42644 12431 42700
rect 12487 42644 12497 42700
rect 12297 42576 12497 42644
rect 12297 42520 12307 42576
rect 12363 42520 12431 42576
rect 12487 42520 12497 42576
rect 12297 42452 12497 42520
rect 12297 42396 12307 42452
rect 12363 42396 12431 42452
rect 12487 42396 12497 42452
rect 12297 42328 12497 42396
rect 12297 42272 12307 42328
rect 12363 42272 12431 42328
rect 12487 42272 12497 42328
rect 12297 42204 12497 42272
rect 12297 42148 12307 42204
rect 12363 42148 12431 42204
rect 12487 42148 12497 42204
rect 12297 42080 12497 42148
rect 12297 42024 12307 42080
rect 12363 42024 12431 42080
rect 12487 42024 12497 42080
rect 12297 41956 12497 42024
rect 12297 41900 12307 41956
rect 12363 41900 12431 41956
rect 12487 41900 12497 41956
rect 12297 41832 12497 41900
rect 12297 41776 12307 41832
rect 12363 41776 12431 41832
rect 12487 41776 12497 41832
rect 12297 41708 12497 41776
rect 12297 41652 12307 41708
rect 12363 41652 12431 41708
rect 12487 41652 12497 41708
rect 12297 41642 12497 41652
rect 2481 41348 2681 41358
rect 2481 41292 2491 41348
rect 2547 41292 2615 41348
rect 2671 41292 2681 41348
rect 2481 41224 2681 41292
rect 2481 41168 2491 41224
rect 2547 41168 2615 41224
rect 2671 41168 2681 41224
rect 2481 41100 2681 41168
rect 2481 41044 2491 41100
rect 2547 41044 2615 41100
rect 2671 41044 2681 41100
rect 2481 40976 2681 41044
rect 2481 40920 2491 40976
rect 2547 40920 2615 40976
rect 2671 40920 2681 40976
rect 2481 40852 2681 40920
rect 2481 40796 2491 40852
rect 2547 40796 2615 40852
rect 2671 40796 2681 40852
rect 2481 40728 2681 40796
rect 2481 40672 2491 40728
rect 2547 40672 2615 40728
rect 2671 40672 2681 40728
rect 2481 40604 2681 40672
rect 2481 40548 2491 40604
rect 2547 40548 2615 40604
rect 2671 40548 2681 40604
rect 2481 40480 2681 40548
rect 2481 40424 2491 40480
rect 2547 40424 2615 40480
rect 2671 40424 2681 40480
rect 2481 40356 2681 40424
rect 2481 40300 2491 40356
rect 2547 40300 2615 40356
rect 2671 40300 2681 40356
rect 2481 40232 2681 40300
rect 2481 40176 2491 40232
rect 2547 40176 2615 40232
rect 2671 40176 2681 40232
rect 2481 40108 2681 40176
rect 2481 40052 2491 40108
rect 2547 40052 2615 40108
rect 2671 40052 2681 40108
rect 2481 40042 2681 40052
rect 4851 41348 5051 41358
rect 4851 41292 4861 41348
rect 4917 41292 4985 41348
rect 5041 41292 5051 41348
rect 4851 41224 5051 41292
rect 4851 41168 4861 41224
rect 4917 41168 4985 41224
rect 5041 41168 5051 41224
rect 4851 41100 5051 41168
rect 4851 41044 4861 41100
rect 4917 41044 4985 41100
rect 5041 41044 5051 41100
rect 4851 40976 5051 41044
rect 4851 40920 4861 40976
rect 4917 40920 4985 40976
rect 5041 40920 5051 40976
rect 4851 40852 5051 40920
rect 4851 40796 4861 40852
rect 4917 40796 4985 40852
rect 5041 40796 5051 40852
rect 4851 40728 5051 40796
rect 4851 40672 4861 40728
rect 4917 40672 4985 40728
rect 5041 40672 5051 40728
rect 4851 40604 5051 40672
rect 4851 40548 4861 40604
rect 4917 40548 4985 40604
rect 5041 40548 5051 40604
rect 4851 40480 5051 40548
rect 4851 40424 4861 40480
rect 4917 40424 4985 40480
rect 5041 40424 5051 40480
rect 4851 40356 5051 40424
rect 4851 40300 4861 40356
rect 4917 40300 4985 40356
rect 5041 40300 5051 40356
rect 4851 40232 5051 40300
rect 4851 40176 4861 40232
rect 4917 40176 4985 40232
rect 5041 40176 5051 40232
rect 4851 40108 5051 40176
rect 4851 40052 4861 40108
rect 4917 40052 4985 40108
rect 5041 40052 5051 40108
rect 4851 40042 5051 40052
rect 7265 41348 7713 41358
rect 7265 41292 7275 41348
rect 7331 41292 7399 41348
rect 7455 41292 7523 41348
rect 7579 41292 7647 41348
rect 7703 41292 7713 41348
rect 7265 41224 7713 41292
rect 7265 41168 7275 41224
rect 7331 41168 7399 41224
rect 7455 41168 7523 41224
rect 7579 41168 7647 41224
rect 7703 41168 7713 41224
rect 7265 41100 7713 41168
rect 7265 41044 7275 41100
rect 7331 41044 7399 41100
rect 7455 41044 7523 41100
rect 7579 41044 7647 41100
rect 7703 41044 7713 41100
rect 7265 40976 7713 41044
rect 7265 40920 7275 40976
rect 7331 40920 7399 40976
rect 7455 40920 7523 40976
rect 7579 40920 7647 40976
rect 7703 40920 7713 40976
rect 7265 40852 7713 40920
rect 7265 40796 7275 40852
rect 7331 40796 7399 40852
rect 7455 40796 7523 40852
rect 7579 40796 7647 40852
rect 7703 40796 7713 40852
rect 7265 40728 7713 40796
rect 7265 40672 7275 40728
rect 7331 40672 7399 40728
rect 7455 40672 7523 40728
rect 7579 40672 7647 40728
rect 7703 40672 7713 40728
rect 7265 40604 7713 40672
rect 7265 40548 7275 40604
rect 7331 40548 7399 40604
rect 7455 40548 7523 40604
rect 7579 40548 7647 40604
rect 7703 40548 7713 40604
rect 7265 40480 7713 40548
rect 7265 40424 7275 40480
rect 7331 40424 7399 40480
rect 7455 40424 7523 40480
rect 7579 40424 7647 40480
rect 7703 40424 7713 40480
rect 7265 40356 7713 40424
rect 7265 40300 7275 40356
rect 7331 40300 7399 40356
rect 7455 40300 7523 40356
rect 7579 40300 7647 40356
rect 7703 40300 7713 40356
rect 7265 40232 7713 40300
rect 7265 40176 7275 40232
rect 7331 40176 7399 40232
rect 7455 40176 7523 40232
rect 7579 40176 7647 40232
rect 7703 40176 7713 40232
rect 7265 40108 7713 40176
rect 7265 40052 7275 40108
rect 7331 40052 7399 40108
rect 7455 40052 7523 40108
rect 7579 40052 7647 40108
rect 7703 40052 7713 40108
rect 7265 40042 7713 40052
rect 9927 41348 10127 41358
rect 9927 41292 9937 41348
rect 9993 41292 10061 41348
rect 10117 41292 10127 41348
rect 9927 41224 10127 41292
rect 9927 41168 9937 41224
rect 9993 41168 10061 41224
rect 10117 41168 10127 41224
rect 9927 41100 10127 41168
rect 9927 41044 9937 41100
rect 9993 41044 10061 41100
rect 10117 41044 10127 41100
rect 9927 40976 10127 41044
rect 9927 40920 9937 40976
rect 9993 40920 10061 40976
rect 10117 40920 10127 40976
rect 9927 40852 10127 40920
rect 9927 40796 9937 40852
rect 9993 40796 10061 40852
rect 10117 40796 10127 40852
rect 9927 40728 10127 40796
rect 9927 40672 9937 40728
rect 9993 40672 10061 40728
rect 10117 40672 10127 40728
rect 9927 40604 10127 40672
rect 9927 40548 9937 40604
rect 9993 40548 10061 40604
rect 10117 40548 10127 40604
rect 9927 40480 10127 40548
rect 9927 40424 9937 40480
rect 9993 40424 10061 40480
rect 10117 40424 10127 40480
rect 9927 40356 10127 40424
rect 9927 40300 9937 40356
rect 9993 40300 10061 40356
rect 10117 40300 10127 40356
rect 9927 40232 10127 40300
rect 9927 40176 9937 40232
rect 9993 40176 10061 40232
rect 10117 40176 10127 40232
rect 9927 40108 10127 40176
rect 9927 40052 9937 40108
rect 9993 40052 10061 40108
rect 10117 40052 10127 40108
rect 9927 40042 10127 40052
rect 12297 41348 12497 41358
rect 12297 41292 12307 41348
rect 12363 41292 12431 41348
rect 12487 41292 12497 41348
rect 12297 41224 12497 41292
rect 12297 41168 12307 41224
rect 12363 41168 12431 41224
rect 12487 41168 12497 41224
rect 12297 41100 12497 41168
rect 12297 41044 12307 41100
rect 12363 41044 12431 41100
rect 12487 41044 12497 41100
rect 12297 40976 12497 41044
rect 12297 40920 12307 40976
rect 12363 40920 12431 40976
rect 12487 40920 12497 40976
rect 12297 40852 12497 40920
rect 12297 40796 12307 40852
rect 12363 40796 12431 40852
rect 12487 40796 12497 40852
rect 12297 40728 12497 40796
rect 12297 40672 12307 40728
rect 12363 40672 12431 40728
rect 12487 40672 12497 40728
rect 12297 40604 12497 40672
rect 12297 40548 12307 40604
rect 12363 40548 12431 40604
rect 12487 40548 12497 40604
rect 12297 40480 12497 40548
rect 12297 40424 12307 40480
rect 12363 40424 12431 40480
rect 12487 40424 12497 40480
rect 12297 40356 12497 40424
rect 12297 40300 12307 40356
rect 12363 40300 12431 40356
rect 12487 40300 12497 40356
rect 12297 40232 12497 40300
rect 12297 40176 12307 40232
rect 12363 40176 12431 40232
rect 12487 40176 12497 40232
rect 12297 40108 12497 40176
rect 12297 40052 12307 40108
rect 12363 40052 12431 40108
rect 12487 40052 12497 40108
rect 12297 40042 12497 40052
rect 2292 39671 2302 39727
rect 2358 39671 2368 39727
rect 2292 39595 2368 39671
rect 2292 39539 2302 39595
rect 2358 39539 2368 39595
rect 2292 39463 2368 39539
rect 2292 39407 2302 39463
rect 2358 39407 2368 39463
rect 2292 39331 2368 39407
rect 2292 39275 2302 39331
rect 2358 39275 2368 39331
rect 2292 39199 2368 39275
rect 2292 39143 2302 39199
rect 2358 39143 2368 39199
rect 2292 39067 2368 39143
rect 2292 39011 2302 39067
rect 2358 39011 2368 39067
rect 2292 38935 2368 39011
rect 2292 38879 2302 38935
rect 2358 38879 2368 38935
rect 2292 38803 2368 38879
rect 2292 38747 2302 38803
rect 2358 38747 2368 38803
rect 2292 38671 2368 38747
rect 2292 38615 2302 38671
rect 2358 38615 2368 38671
rect 2292 38539 2368 38615
rect 2292 38483 2302 38539
rect 2358 38483 2368 38539
rect 2292 38400 2368 38483
rect -11 38176 86 38200
rect -11 36824 20 38176
rect 76 36824 86 38176
rect 14892 38176 14989 38200
rect 305 38148 2117 38158
rect 305 38092 315 38148
rect 371 38092 439 38148
rect 495 38092 563 38148
rect 619 38092 687 38148
rect 743 38092 811 38148
rect 867 38092 935 38148
rect 991 38092 1059 38148
rect 1115 38092 1183 38148
rect 1239 38092 1307 38148
rect 1363 38092 1431 38148
rect 1487 38092 1555 38148
rect 1611 38092 1679 38148
rect 1735 38092 1803 38148
rect 1859 38092 1927 38148
rect 1983 38092 2051 38148
rect 2107 38092 2117 38148
rect 305 38024 2117 38092
rect 305 37968 315 38024
rect 371 37968 439 38024
rect 495 37968 563 38024
rect 619 37968 687 38024
rect 743 37968 811 38024
rect 867 37968 935 38024
rect 991 37968 1059 38024
rect 1115 37968 1183 38024
rect 1239 37968 1307 38024
rect 1363 37968 1431 38024
rect 1487 37968 1555 38024
rect 1611 37968 1679 38024
rect 1735 37968 1803 38024
rect 1859 37968 1927 38024
rect 1983 37968 2051 38024
rect 2107 37968 2117 38024
rect 305 37900 2117 37968
rect 305 37844 315 37900
rect 371 37844 439 37900
rect 495 37844 563 37900
rect 619 37844 687 37900
rect 743 37844 811 37900
rect 867 37844 935 37900
rect 991 37844 1059 37900
rect 1115 37844 1183 37900
rect 1239 37844 1307 37900
rect 1363 37844 1431 37900
rect 1487 37844 1555 37900
rect 1611 37844 1679 37900
rect 1735 37844 1803 37900
rect 1859 37844 1927 37900
rect 1983 37844 2051 37900
rect 2107 37844 2117 37900
rect 305 37776 2117 37844
rect 305 37720 315 37776
rect 371 37720 439 37776
rect 495 37720 563 37776
rect 619 37720 687 37776
rect 743 37720 811 37776
rect 867 37720 935 37776
rect 991 37720 1059 37776
rect 1115 37720 1183 37776
rect 1239 37720 1307 37776
rect 1363 37720 1431 37776
rect 1487 37720 1555 37776
rect 1611 37720 1679 37776
rect 1735 37720 1803 37776
rect 1859 37720 1927 37776
rect 1983 37720 2051 37776
rect 2107 37720 2117 37776
rect 305 37652 2117 37720
rect 305 37596 315 37652
rect 371 37596 439 37652
rect 495 37596 563 37652
rect 619 37596 687 37652
rect 743 37596 811 37652
rect 867 37596 935 37652
rect 991 37596 1059 37652
rect 1115 37596 1183 37652
rect 1239 37596 1307 37652
rect 1363 37596 1431 37652
rect 1487 37596 1555 37652
rect 1611 37596 1679 37652
rect 1735 37596 1803 37652
rect 1859 37596 1927 37652
rect 1983 37596 2051 37652
rect 2107 37596 2117 37652
rect 305 37528 2117 37596
rect 305 37472 315 37528
rect 371 37472 439 37528
rect 495 37472 563 37528
rect 619 37472 687 37528
rect 743 37472 811 37528
rect 867 37472 935 37528
rect 991 37472 1059 37528
rect 1115 37472 1183 37528
rect 1239 37472 1307 37528
rect 1363 37472 1431 37528
rect 1487 37472 1555 37528
rect 1611 37472 1679 37528
rect 1735 37472 1803 37528
rect 1859 37472 1927 37528
rect 1983 37472 2051 37528
rect 2107 37472 2117 37528
rect 305 37404 2117 37472
rect 305 37348 315 37404
rect 371 37348 439 37404
rect 495 37348 563 37404
rect 619 37348 687 37404
rect 743 37348 811 37404
rect 867 37348 935 37404
rect 991 37348 1059 37404
rect 1115 37348 1183 37404
rect 1239 37348 1307 37404
rect 1363 37348 1431 37404
rect 1487 37348 1555 37404
rect 1611 37348 1679 37404
rect 1735 37348 1803 37404
rect 1859 37348 1927 37404
rect 1983 37348 2051 37404
rect 2107 37348 2117 37404
rect 305 37280 2117 37348
rect 305 37224 315 37280
rect 371 37224 439 37280
rect 495 37224 563 37280
rect 619 37224 687 37280
rect 743 37224 811 37280
rect 867 37224 935 37280
rect 991 37224 1059 37280
rect 1115 37224 1183 37280
rect 1239 37224 1307 37280
rect 1363 37224 1431 37280
rect 1487 37224 1555 37280
rect 1611 37224 1679 37280
rect 1735 37224 1803 37280
rect 1859 37224 1927 37280
rect 1983 37224 2051 37280
rect 2107 37224 2117 37280
rect 305 37156 2117 37224
rect 305 37100 315 37156
rect 371 37100 439 37156
rect 495 37100 563 37156
rect 619 37100 687 37156
rect 743 37100 811 37156
rect 867 37100 935 37156
rect 991 37100 1059 37156
rect 1115 37100 1183 37156
rect 1239 37100 1307 37156
rect 1363 37100 1431 37156
rect 1487 37100 1555 37156
rect 1611 37100 1679 37156
rect 1735 37100 1803 37156
rect 1859 37100 1927 37156
rect 1983 37100 2051 37156
rect 2107 37100 2117 37156
rect 305 37032 2117 37100
rect 305 36976 315 37032
rect 371 36976 439 37032
rect 495 36976 563 37032
rect 619 36976 687 37032
rect 743 36976 811 37032
rect 867 36976 935 37032
rect 991 36976 1059 37032
rect 1115 36976 1183 37032
rect 1239 36976 1307 37032
rect 1363 36976 1431 37032
rect 1487 36976 1555 37032
rect 1611 36976 1679 37032
rect 1735 36976 1803 37032
rect 1859 36976 1927 37032
rect 1983 36976 2051 37032
rect 2107 36976 2117 37032
rect 305 36908 2117 36976
rect 305 36852 315 36908
rect 371 36852 439 36908
rect 495 36852 563 36908
rect 619 36852 687 36908
rect 743 36852 811 36908
rect 867 36852 935 36908
rect 991 36852 1059 36908
rect 1115 36852 1183 36908
rect 1239 36852 1307 36908
rect 1363 36852 1431 36908
rect 1487 36852 1555 36908
rect 1611 36852 1679 36908
rect 1735 36852 1803 36908
rect 1859 36852 1927 36908
rect 1983 36852 2051 36908
rect 2107 36852 2117 36908
rect 305 36842 2117 36852
rect 2798 38148 4734 38158
rect 2798 38092 2808 38148
rect 2864 38092 2932 38148
rect 2988 38092 3056 38148
rect 3112 38092 3180 38148
rect 3236 38092 3304 38148
rect 3360 38092 3428 38148
rect 3484 38092 3552 38148
rect 3608 38092 3676 38148
rect 3732 38092 3800 38148
rect 3856 38092 3924 38148
rect 3980 38092 4048 38148
rect 4104 38092 4172 38148
rect 4228 38092 4296 38148
rect 4352 38092 4420 38148
rect 4476 38092 4544 38148
rect 4600 38092 4668 38148
rect 4724 38092 4734 38148
rect 2798 38024 4734 38092
rect 2798 37968 2808 38024
rect 2864 37968 2932 38024
rect 2988 37968 3056 38024
rect 3112 37968 3180 38024
rect 3236 37968 3304 38024
rect 3360 37968 3428 38024
rect 3484 37968 3552 38024
rect 3608 37968 3676 38024
rect 3732 37968 3800 38024
rect 3856 37968 3924 38024
rect 3980 37968 4048 38024
rect 4104 37968 4172 38024
rect 4228 37968 4296 38024
rect 4352 37968 4420 38024
rect 4476 37968 4544 38024
rect 4600 37968 4668 38024
rect 4724 37968 4734 38024
rect 2798 37900 4734 37968
rect 2798 37844 2808 37900
rect 2864 37844 2932 37900
rect 2988 37844 3056 37900
rect 3112 37844 3180 37900
rect 3236 37844 3304 37900
rect 3360 37844 3428 37900
rect 3484 37844 3552 37900
rect 3608 37844 3676 37900
rect 3732 37844 3800 37900
rect 3856 37844 3924 37900
rect 3980 37844 4048 37900
rect 4104 37844 4172 37900
rect 4228 37844 4296 37900
rect 4352 37844 4420 37900
rect 4476 37844 4544 37900
rect 4600 37844 4668 37900
rect 4724 37844 4734 37900
rect 2798 37776 4734 37844
rect 2798 37720 2808 37776
rect 2864 37720 2932 37776
rect 2988 37720 3056 37776
rect 3112 37720 3180 37776
rect 3236 37720 3304 37776
rect 3360 37720 3428 37776
rect 3484 37720 3552 37776
rect 3608 37720 3676 37776
rect 3732 37720 3800 37776
rect 3856 37720 3924 37776
rect 3980 37720 4048 37776
rect 4104 37720 4172 37776
rect 4228 37720 4296 37776
rect 4352 37720 4420 37776
rect 4476 37720 4544 37776
rect 4600 37720 4668 37776
rect 4724 37720 4734 37776
rect 2798 37652 4734 37720
rect 2798 37596 2808 37652
rect 2864 37596 2932 37652
rect 2988 37596 3056 37652
rect 3112 37596 3180 37652
rect 3236 37596 3304 37652
rect 3360 37596 3428 37652
rect 3484 37596 3552 37652
rect 3608 37596 3676 37652
rect 3732 37596 3800 37652
rect 3856 37596 3924 37652
rect 3980 37596 4048 37652
rect 4104 37596 4172 37652
rect 4228 37596 4296 37652
rect 4352 37596 4420 37652
rect 4476 37596 4544 37652
rect 4600 37596 4668 37652
rect 4724 37596 4734 37652
rect 2798 37528 4734 37596
rect 2798 37472 2808 37528
rect 2864 37472 2932 37528
rect 2988 37472 3056 37528
rect 3112 37472 3180 37528
rect 3236 37472 3304 37528
rect 3360 37472 3428 37528
rect 3484 37472 3552 37528
rect 3608 37472 3676 37528
rect 3732 37472 3800 37528
rect 3856 37472 3924 37528
rect 3980 37472 4048 37528
rect 4104 37472 4172 37528
rect 4228 37472 4296 37528
rect 4352 37472 4420 37528
rect 4476 37472 4544 37528
rect 4600 37472 4668 37528
rect 4724 37472 4734 37528
rect 2798 37404 4734 37472
rect 2798 37348 2808 37404
rect 2864 37348 2932 37404
rect 2988 37348 3056 37404
rect 3112 37348 3180 37404
rect 3236 37348 3304 37404
rect 3360 37348 3428 37404
rect 3484 37348 3552 37404
rect 3608 37348 3676 37404
rect 3732 37348 3800 37404
rect 3856 37348 3924 37404
rect 3980 37348 4048 37404
rect 4104 37348 4172 37404
rect 4228 37348 4296 37404
rect 4352 37348 4420 37404
rect 4476 37348 4544 37404
rect 4600 37348 4668 37404
rect 4724 37348 4734 37404
rect 2798 37280 4734 37348
rect 2798 37224 2808 37280
rect 2864 37224 2932 37280
rect 2988 37224 3056 37280
rect 3112 37224 3180 37280
rect 3236 37224 3304 37280
rect 3360 37224 3428 37280
rect 3484 37224 3552 37280
rect 3608 37224 3676 37280
rect 3732 37224 3800 37280
rect 3856 37224 3924 37280
rect 3980 37224 4048 37280
rect 4104 37224 4172 37280
rect 4228 37224 4296 37280
rect 4352 37224 4420 37280
rect 4476 37224 4544 37280
rect 4600 37224 4668 37280
rect 4724 37224 4734 37280
rect 2798 37156 4734 37224
rect 2798 37100 2808 37156
rect 2864 37100 2932 37156
rect 2988 37100 3056 37156
rect 3112 37100 3180 37156
rect 3236 37100 3304 37156
rect 3360 37100 3428 37156
rect 3484 37100 3552 37156
rect 3608 37100 3676 37156
rect 3732 37100 3800 37156
rect 3856 37100 3924 37156
rect 3980 37100 4048 37156
rect 4104 37100 4172 37156
rect 4228 37100 4296 37156
rect 4352 37100 4420 37156
rect 4476 37100 4544 37156
rect 4600 37100 4668 37156
rect 4724 37100 4734 37156
rect 2798 37032 4734 37100
rect 2798 36976 2808 37032
rect 2864 36976 2932 37032
rect 2988 36976 3056 37032
rect 3112 36976 3180 37032
rect 3236 36976 3304 37032
rect 3360 36976 3428 37032
rect 3484 36976 3552 37032
rect 3608 36976 3676 37032
rect 3732 36976 3800 37032
rect 3856 36976 3924 37032
rect 3980 36976 4048 37032
rect 4104 36976 4172 37032
rect 4228 36976 4296 37032
rect 4352 36976 4420 37032
rect 4476 36976 4544 37032
rect 4600 36976 4668 37032
rect 4724 36976 4734 37032
rect 2798 36908 4734 36976
rect 2798 36852 2808 36908
rect 2864 36852 2932 36908
rect 2988 36852 3056 36908
rect 3112 36852 3180 36908
rect 3236 36852 3304 36908
rect 3360 36852 3428 36908
rect 3484 36852 3552 36908
rect 3608 36852 3676 36908
rect 3732 36852 3800 36908
rect 3856 36852 3924 36908
rect 3980 36852 4048 36908
rect 4104 36852 4172 36908
rect 4228 36852 4296 36908
rect 4352 36852 4420 36908
rect 4476 36852 4544 36908
rect 4600 36852 4668 36908
rect 4724 36852 4734 36908
rect 2798 36842 4734 36852
rect 5168 38148 7104 38158
rect 5168 38092 5178 38148
rect 5234 38092 5302 38148
rect 5358 38092 5426 38148
rect 5482 38092 5550 38148
rect 5606 38092 5674 38148
rect 5730 38092 5798 38148
rect 5854 38092 5922 38148
rect 5978 38092 6046 38148
rect 6102 38092 6170 38148
rect 6226 38092 6294 38148
rect 6350 38092 6418 38148
rect 6474 38092 6542 38148
rect 6598 38092 6666 38148
rect 6722 38092 6790 38148
rect 6846 38092 6914 38148
rect 6970 38092 7038 38148
rect 7094 38092 7104 38148
rect 5168 38024 7104 38092
rect 5168 37968 5178 38024
rect 5234 37968 5302 38024
rect 5358 37968 5426 38024
rect 5482 37968 5550 38024
rect 5606 37968 5674 38024
rect 5730 37968 5798 38024
rect 5854 37968 5922 38024
rect 5978 37968 6046 38024
rect 6102 37968 6170 38024
rect 6226 37968 6294 38024
rect 6350 37968 6418 38024
rect 6474 37968 6542 38024
rect 6598 37968 6666 38024
rect 6722 37968 6790 38024
rect 6846 37968 6914 38024
rect 6970 37968 7038 38024
rect 7094 37968 7104 38024
rect 5168 37900 7104 37968
rect 5168 37844 5178 37900
rect 5234 37844 5302 37900
rect 5358 37844 5426 37900
rect 5482 37844 5550 37900
rect 5606 37844 5674 37900
rect 5730 37844 5798 37900
rect 5854 37844 5922 37900
rect 5978 37844 6046 37900
rect 6102 37844 6170 37900
rect 6226 37844 6294 37900
rect 6350 37844 6418 37900
rect 6474 37844 6542 37900
rect 6598 37844 6666 37900
rect 6722 37844 6790 37900
rect 6846 37844 6914 37900
rect 6970 37844 7038 37900
rect 7094 37844 7104 37900
rect 5168 37776 7104 37844
rect 5168 37720 5178 37776
rect 5234 37720 5302 37776
rect 5358 37720 5426 37776
rect 5482 37720 5550 37776
rect 5606 37720 5674 37776
rect 5730 37720 5798 37776
rect 5854 37720 5922 37776
rect 5978 37720 6046 37776
rect 6102 37720 6170 37776
rect 6226 37720 6294 37776
rect 6350 37720 6418 37776
rect 6474 37720 6542 37776
rect 6598 37720 6666 37776
rect 6722 37720 6790 37776
rect 6846 37720 6914 37776
rect 6970 37720 7038 37776
rect 7094 37720 7104 37776
rect 5168 37652 7104 37720
rect 5168 37596 5178 37652
rect 5234 37596 5302 37652
rect 5358 37596 5426 37652
rect 5482 37596 5550 37652
rect 5606 37596 5674 37652
rect 5730 37596 5798 37652
rect 5854 37596 5922 37652
rect 5978 37596 6046 37652
rect 6102 37596 6170 37652
rect 6226 37596 6294 37652
rect 6350 37596 6418 37652
rect 6474 37596 6542 37652
rect 6598 37596 6666 37652
rect 6722 37596 6790 37652
rect 6846 37596 6914 37652
rect 6970 37596 7038 37652
rect 7094 37596 7104 37652
rect 5168 37528 7104 37596
rect 5168 37472 5178 37528
rect 5234 37472 5302 37528
rect 5358 37472 5426 37528
rect 5482 37472 5550 37528
rect 5606 37472 5674 37528
rect 5730 37472 5798 37528
rect 5854 37472 5922 37528
rect 5978 37472 6046 37528
rect 6102 37472 6170 37528
rect 6226 37472 6294 37528
rect 6350 37472 6418 37528
rect 6474 37472 6542 37528
rect 6598 37472 6666 37528
rect 6722 37472 6790 37528
rect 6846 37472 6914 37528
rect 6970 37472 7038 37528
rect 7094 37472 7104 37528
rect 5168 37404 7104 37472
rect 5168 37348 5178 37404
rect 5234 37348 5302 37404
rect 5358 37348 5426 37404
rect 5482 37348 5550 37404
rect 5606 37348 5674 37404
rect 5730 37348 5798 37404
rect 5854 37348 5922 37404
rect 5978 37348 6046 37404
rect 6102 37348 6170 37404
rect 6226 37348 6294 37404
rect 6350 37348 6418 37404
rect 6474 37348 6542 37404
rect 6598 37348 6666 37404
rect 6722 37348 6790 37404
rect 6846 37348 6914 37404
rect 6970 37348 7038 37404
rect 7094 37348 7104 37404
rect 5168 37280 7104 37348
rect 5168 37224 5178 37280
rect 5234 37224 5302 37280
rect 5358 37224 5426 37280
rect 5482 37224 5550 37280
rect 5606 37224 5674 37280
rect 5730 37224 5798 37280
rect 5854 37224 5922 37280
rect 5978 37224 6046 37280
rect 6102 37224 6170 37280
rect 6226 37224 6294 37280
rect 6350 37224 6418 37280
rect 6474 37224 6542 37280
rect 6598 37224 6666 37280
rect 6722 37224 6790 37280
rect 6846 37224 6914 37280
rect 6970 37224 7038 37280
rect 7094 37224 7104 37280
rect 5168 37156 7104 37224
rect 5168 37100 5178 37156
rect 5234 37100 5302 37156
rect 5358 37100 5426 37156
rect 5482 37100 5550 37156
rect 5606 37100 5674 37156
rect 5730 37100 5798 37156
rect 5854 37100 5922 37156
rect 5978 37100 6046 37156
rect 6102 37100 6170 37156
rect 6226 37100 6294 37156
rect 6350 37100 6418 37156
rect 6474 37100 6542 37156
rect 6598 37100 6666 37156
rect 6722 37100 6790 37156
rect 6846 37100 6914 37156
rect 6970 37100 7038 37156
rect 7094 37100 7104 37156
rect 5168 37032 7104 37100
rect 5168 36976 5178 37032
rect 5234 36976 5302 37032
rect 5358 36976 5426 37032
rect 5482 36976 5550 37032
rect 5606 36976 5674 37032
rect 5730 36976 5798 37032
rect 5854 36976 5922 37032
rect 5978 36976 6046 37032
rect 6102 36976 6170 37032
rect 6226 36976 6294 37032
rect 6350 36976 6418 37032
rect 6474 36976 6542 37032
rect 6598 36976 6666 37032
rect 6722 36976 6790 37032
rect 6846 36976 6914 37032
rect 6970 36976 7038 37032
rect 7094 36976 7104 37032
rect 5168 36908 7104 36976
rect 5168 36852 5178 36908
rect 5234 36852 5302 36908
rect 5358 36852 5426 36908
rect 5482 36852 5550 36908
rect 5606 36852 5674 36908
rect 5730 36852 5798 36908
rect 5854 36852 5922 36908
rect 5978 36852 6046 36908
rect 6102 36852 6170 36908
rect 6226 36852 6294 36908
rect 6350 36852 6418 36908
rect 6474 36852 6542 36908
rect 6598 36852 6666 36908
rect 6722 36852 6790 36908
rect 6846 36852 6914 36908
rect 6970 36852 7038 36908
rect 7094 36852 7104 36908
rect 5168 36842 7104 36852
rect 7874 38148 9810 38158
rect 7874 38092 7884 38148
rect 7940 38092 8008 38148
rect 8064 38092 8132 38148
rect 8188 38092 8256 38148
rect 8312 38092 8380 38148
rect 8436 38092 8504 38148
rect 8560 38092 8628 38148
rect 8684 38092 8752 38148
rect 8808 38092 8876 38148
rect 8932 38092 9000 38148
rect 9056 38092 9124 38148
rect 9180 38092 9248 38148
rect 9304 38092 9372 38148
rect 9428 38092 9496 38148
rect 9552 38092 9620 38148
rect 9676 38092 9744 38148
rect 9800 38092 9810 38148
rect 7874 38024 9810 38092
rect 7874 37968 7884 38024
rect 7940 37968 8008 38024
rect 8064 37968 8132 38024
rect 8188 37968 8256 38024
rect 8312 37968 8380 38024
rect 8436 37968 8504 38024
rect 8560 37968 8628 38024
rect 8684 37968 8752 38024
rect 8808 37968 8876 38024
rect 8932 37968 9000 38024
rect 9056 37968 9124 38024
rect 9180 37968 9248 38024
rect 9304 37968 9372 38024
rect 9428 37968 9496 38024
rect 9552 37968 9620 38024
rect 9676 37968 9744 38024
rect 9800 37968 9810 38024
rect 7874 37900 9810 37968
rect 7874 37844 7884 37900
rect 7940 37844 8008 37900
rect 8064 37844 8132 37900
rect 8188 37844 8256 37900
rect 8312 37844 8380 37900
rect 8436 37844 8504 37900
rect 8560 37844 8628 37900
rect 8684 37844 8752 37900
rect 8808 37844 8876 37900
rect 8932 37844 9000 37900
rect 9056 37844 9124 37900
rect 9180 37844 9248 37900
rect 9304 37844 9372 37900
rect 9428 37844 9496 37900
rect 9552 37844 9620 37900
rect 9676 37844 9744 37900
rect 9800 37844 9810 37900
rect 7874 37776 9810 37844
rect 7874 37720 7884 37776
rect 7940 37720 8008 37776
rect 8064 37720 8132 37776
rect 8188 37720 8256 37776
rect 8312 37720 8380 37776
rect 8436 37720 8504 37776
rect 8560 37720 8628 37776
rect 8684 37720 8752 37776
rect 8808 37720 8876 37776
rect 8932 37720 9000 37776
rect 9056 37720 9124 37776
rect 9180 37720 9248 37776
rect 9304 37720 9372 37776
rect 9428 37720 9496 37776
rect 9552 37720 9620 37776
rect 9676 37720 9744 37776
rect 9800 37720 9810 37776
rect 7874 37652 9810 37720
rect 7874 37596 7884 37652
rect 7940 37596 8008 37652
rect 8064 37596 8132 37652
rect 8188 37596 8256 37652
rect 8312 37596 8380 37652
rect 8436 37596 8504 37652
rect 8560 37596 8628 37652
rect 8684 37596 8752 37652
rect 8808 37596 8876 37652
rect 8932 37596 9000 37652
rect 9056 37596 9124 37652
rect 9180 37596 9248 37652
rect 9304 37596 9372 37652
rect 9428 37596 9496 37652
rect 9552 37596 9620 37652
rect 9676 37596 9744 37652
rect 9800 37596 9810 37652
rect 7874 37528 9810 37596
rect 7874 37472 7884 37528
rect 7940 37472 8008 37528
rect 8064 37472 8132 37528
rect 8188 37472 8256 37528
rect 8312 37472 8380 37528
rect 8436 37472 8504 37528
rect 8560 37472 8628 37528
rect 8684 37472 8752 37528
rect 8808 37472 8876 37528
rect 8932 37472 9000 37528
rect 9056 37472 9124 37528
rect 9180 37472 9248 37528
rect 9304 37472 9372 37528
rect 9428 37472 9496 37528
rect 9552 37472 9620 37528
rect 9676 37472 9744 37528
rect 9800 37472 9810 37528
rect 7874 37404 9810 37472
rect 7874 37348 7884 37404
rect 7940 37348 8008 37404
rect 8064 37348 8132 37404
rect 8188 37348 8256 37404
rect 8312 37348 8380 37404
rect 8436 37348 8504 37404
rect 8560 37348 8628 37404
rect 8684 37348 8752 37404
rect 8808 37348 8876 37404
rect 8932 37348 9000 37404
rect 9056 37348 9124 37404
rect 9180 37348 9248 37404
rect 9304 37348 9372 37404
rect 9428 37348 9496 37404
rect 9552 37348 9620 37404
rect 9676 37348 9744 37404
rect 9800 37348 9810 37404
rect 7874 37280 9810 37348
rect 7874 37224 7884 37280
rect 7940 37224 8008 37280
rect 8064 37224 8132 37280
rect 8188 37224 8256 37280
rect 8312 37224 8380 37280
rect 8436 37224 8504 37280
rect 8560 37224 8628 37280
rect 8684 37224 8752 37280
rect 8808 37224 8876 37280
rect 8932 37224 9000 37280
rect 9056 37224 9124 37280
rect 9180 37224 9248 37280
rect 9304 37224 9372 37280
rect 9428 37224 9496 37280
rect 9552 37224 9620 37280
rect 9676 37224 9744 37280
rect 9800 37224 9810 37280
rect 7874 37156 9810 37224
rect 7874 37100 7884 37156
rect 7940 37100 8008 37156
rect 8064 37100 8132 37156
rect 8188 37100 8256 37156
rect 8312 37100 8380 37156
rect 8436 37100 8504 37156
rect 8560 37100 8628 37156
rect 8684 37100 8752 37156
rect 8808 37100 8876 37156
rect 8932 37100 9000 37156
rect 9056 37100 9124 37156
rect 9180 37100 9248 37156
rect 9304 37100 9372 37156
rect 9428 37100 9496 37156
rect 9552 37100 9620 37156
rect 9676 37100 9744 37156
rect 9800 37100 9810 37156
rect 7874 37032 9810 37100
rect 7874 36976 7884 37032
rect 7940 36976 8008 37032
rect 8064 36976 8132 37032
rect 8188 36976 8256 37032
rect 8312 36976 8380 37032
rect 8436 36976 8504 37032
rect 8560 36976 8628 37032
rect 8684 36976 8752 37032
rect 8808 36976 8876 37032
rect 8932 36976 9000 37032
rect 9056 36976 9124 37032
rect 9180 36976 9248 37032
rect 9304 36976 9372 37032
rect 9428 36976 9496 37032
rect 9552 36976 9620 37032
rect 9676 36976 9744 37032
rect 9800 36976 9810 37032
rect 7874 36908 9810 36976
rect 7874 36852 7884 36908
rect 7940 36852 8008 36908
rect 8064 36852 8132 36908
rect 8188 36852 8256 36908
rect 8312 36852 8380 36908
rect 8436 36852 8504 36908
rect 8560 36852 8628 36908
rect 8684 36852 8752 36908
rect 8808 36852 8876 36908
rect 8932 36852 9000 36908
rect 9056 36852 9124 36908
rect 9180 36852 9248 36908
rect 9304 36852 9372 36908
rect 9428 36852 9496 36908
rect 9552 36852 9620 36908
rect 9676 36852 9744 36908
rect 9800 36852 9810 36908
rect 7874 36842 9810 36852
rect 10244 38148 12180 38158
rect 10244 38092 10254 38148
rect 10310 38092 10378 38148
rect 10434 38092 10502 38148
rect 10558 38092 10626 38148
rect 10682 38092 10750 38148
rect 10806 38092 10874 38148
rect 10930 38092 10998 38148
rect 11054 38092 11122 38148
rect 11178 38092 11246 38148
rect 11302 38092 11370 38148
rect 11426 38092 11494 38148
rect 11550 38092 11618 38148
rect 11674 38092 11742 38148
rect 11798 38092 11866 38148
rect 11922 38092 11990 38148
rect 12046 38092 12114 38148
rect 12170 38092 12180 38148
rect 10244 38024 12180 38092
rect 10244 37968 10254 38024
rect 10310 37968 10378 38024
rect 10434 37968 10502 38024
rect 10558 37968 10626 38024
rect 10682 37968 10750 38024
rect 10806 37968 10874 38024
rect 10930 37968 10998 38024
rect 11054 37968 11122 38024
rect 11178 37968 11246 38024
rect 11302 37968 11370 38024
rect 11426 37968 11494 38024
rect 11550 37968 11618 38024
rect 11674 37968 11742 38024
rect 11798 37968 11866 38024
rect 11922 37968 11990 38024
rect 12046 37968 12114 38024
rect 12170 37968 12180 38024
rect 10244 37900 12180 37968
rect 10244 37844 10254 37900
rect 10310 37844 10378 37900
rect 10434 37844 10502 37900
rect 10558 37844 10626 37900
rect 10682 37844 10750 37900
rect 10806 37844 10874 37900
rect 10930 37844 10998 37900
rect 11054 37844 11122 37900
rect 11178 37844 11246 37900
rect 11302 37844 11370 37900
rect 11426 37844 11494 37900
rect 11550 37844 11618 37900
rect 11674 37844 11742 37900
rect 11798 37844 11866 37900
rect 11922 37844 11990 37900
rect 12046 37844 12114 37900
rect 12170 37844 12180 37900
rect 10244 37776 12180 37844
rect 10244 37720 10254 37776
rect 10310 37720 10378 37776
rect 10434 37720 10502 37776
rect 10558 37720 10626 37776
rect 10682 37720 10750 37776
rect 10806 37720 10874 37776
rect 10930 37720 10998 37776
rect 11054 37720 11122 37776
rect 11178 37720 11246 37776
rect 11302 37720 11370 37776
rect 11426 37720 11494 37776
rect 11550 37720 11618 37776
rect 11674 37720 11742 37776
rect 11798 37720 11866 37776
rect 11922 37720 11990 37776
rect 12046 37720 12114 37776
rect 12170 37720 12180 37776
rect 10244 37652 12180 37720
rect 10244 37596 10254 37652
rect 10310 37596 10378 37652
rect 10434 37596 10502 37652
rect 10558 37596 10626 37652
rect 10682 37596 10750 37652
rect 10806 37596 10874 37652
rect 10930 37596 10998 37652
rect 11054 37596 11122 37652
rect 11178 37596 11246 37652
rect 11302 37596 11370 37652
rect 11426 37596 11494 37652
rect 11550 37596 11618 37652
rect 11674 37596 11742 37652
rect 11798 37596 11866 37652
rect 11922 37596 11990 37652
rect 12046 37596 12114 37652
rect 12170 37596 12180 37652
rect 10244 37528 12180 37596
rect 10244 37472 10254 37528
rect 10310 37472 10378 37528
rect 10434 37472 10502 37528
rect 10558 37472 10626 37528
rect 10682 37472 10750 37528
rect 10806 37472 10874 37528
rect 10930 37472 10998 37528
rect 11054 37472 11122 37528
rect 11178 37472 11246 37528
rect 11302 37472 11370 37528
rect 11426 37472 11494 37528
rect 11550 37472 11618 37528
rect 11674 37472 11742 37528
rect 11798 37472 11866 37528
rect 11922 37472 11990 37528
rect 12046 37472 12114 37528
rect 12170 37472 12180 37528
rect 10244 37404 12180 37472
rect 10244 37348 10254 37404
rect 10310 37348 10378 37404
rect 10434 37348 10502 37404
rect 10558 37348 10626 37404
rect 10682 37348 10750 37404
rect 10806 37348 10874 37404
rect 10930 37348 10998 37404
rect 11054 37348 11122 37404
rect 11178 37348 11246 37404
rect 11302 37348 11370 37404
rect 11426 37348 11494 37404
rect 11550 37348 11618 37404
rect 11674 37348 11742 37404
rect 11798 37348 11866 37404
rect 11922 37348 11990 37404
rect 12046 37348 12114 37404
rect 12170 37348 12180 37404
rect 10244 37280 12180 37348
rect 10244 37224 10254 37280
rect 10310 37224 10378 37280
rect 10434 37224 10502 37280
rect 10558 37224 10626 37280
rect 10682 37224 10750 37280
rect 10806 37224 10874 37280
rect 10930 37224 10998 37280
rect 11054 37224 11122 37280
rect 11178 37224 11246 37280
rect 11302 37224 11370 37280
rect 11426 37224 11494 37280
rect 11550 37224 11618 37280
rect 11674 37224 11742 37280
rect 11798 37224 11866 37280
rect 11922 37224 11990 37280
rect 12046 37224 12114 37280
rect 12170 37224 12180 37280
rect 10244 37156 12180 37224
rect 10244 37100 10254 37156
rect 10310 37100 10378 37156
rect 10434 37100 10502 37156
rect 10558 37100 10626 37156
rect 10682 37100 10750 37156
rect 10806 37100 10874 37156
rect 10930 37100 10998 37156
rect 11054 37100 11122 37156
rect 11178 37100 11246 37156
rect 11302 37100 11370 37156
rect 11426 37100 11494 37156
rect 11550 37100 11618 37156
rect 11674 37100 11742 37156
rect 11798 37100 11866 37156
rect 11922 37100 11990 37156
rect 12046 37100 12114 37156
rect 12170 37100 12180 37156
rect 10244 37032 12180 37100
rect 10244 36976 10254 37032
rect 10310 36976 10378 37032
rect 10434 36976 10502 37032
rect 10558 36976 10626 37032
rect 10682 36976 10750 37032
rect 10806 36976 10874 37032
rect 10930 36976 10998 37032
rect 11054 36976 11122 37032
rect 11178 36976 11246 37032
rect 11302 36976 11370 37032
rect 11426 36976 11494 37032
rect 11550 36976 11618 37032
rect 11674 36976 11742 37032
rect 11798 36976 11866 37032
rect 11922 36976 11990 37032
rect 12046 36976 12114 37032
rect 12170 36976 12180 37032
rect 10244 36908 12180 36976
rect 10244 36852 10254 36908
rect 10310 36852 10378 36908
rect 10434 36852 10502 36908
rect 10558 36852 10626 36908
rect 10682 36852 10750 36908
rect 10806 36852 10874 36908
rect 10930 36852 10998 36908
rect 11054 36852 11122 36908
rect 11178 36852 11246 36908
rect 11302 36852 11370 36908
rect 11426 36852 11494 36908
rect 11550 36852 11618 36908
rect 11674 36852 11742 36908
rect 11798 36852 11866 36908
rect 11922 36852 11990 36908
rect 12046 36852 12114 36908
rect 12170 36852 12180 36908
rect 10244 36842 12180 36852
rect 12861 38148 14673 38158
rect 12861 38092 12871 38148
rect 12927 38092 12995 38148
rect 13051 38092 13119 38148
rect 13175 38092 13243 38148
rect 13299 38092 13367 38148
rect 13423 38092 13491 38148
rect 13547 38092 13615 38148
rect 13671 38092 13739 38148
rect 13795 38092 13863 38148
rect 13919 38092 13987 38148
rect 14043 38092 14111 38148
rect 14167 38092 14235 38148
rect 14291 38092 14359 38148
rect 14415 38092 14483 38148
rect 14539 38092 14607 38148
rect 14663 38092 14673 38148
rect 12861 38024 14673 38092
rect 12861 37968 12871 38024
rect 12927 37968 12995 38024
rect 13051 37968 13119 38024
rect 13175 37968 13243 38024
rect 13299 37968 13367 38024
rect 13423 37968 13491 38024
rect 13547 37968 13615 38024
rect 13671 37968 13739 38024
rect 13795 37968 13863 38024
rect 13919 37968 13987 38024
rect 14043 37968 14111 38024
rect 14167 37968 14235 38024
rect 14291 37968 14359 38024
rect 14415 37968 14483 38024
rect 14539 37968 14607 38024
rect 14663 37968 14673 38024
rect 12861 37900 14673 37968
rect 12861 37844 12871 37900
rect 12927 37844 12995 37900
rect 13051 37844 13119 37900
rect 13175 37844 13243 37900
rect 13299 37844 13367 37900
rect 13423 37844 13491 37900
rect 13547 37844 13615 37900
rect 13671 37844 13739 37900
rect 13795 37844 13863 37900
rect 13919 37844 13987 37900
rect 14043 37844 14111 37900
rect 14167 37844 14235 37900
rect 14291 37844 14359 37900
rect 14415 37844 14483 37900
rect 14539 37844 14607 37900
rect 14663 37844 14673 37900
rect 12861 37776 14673 37844
rect 12861 37720 12871 37776
rect 12927 37720 12995 37776
rect 13051 37720 13119 37776
rect 13175 37720 13243 37776
rect 13299 37720 13367 37776
rect 13423 37720 13491 37776
rect 13547 37720 13615 37776
rect 13671 37720 13739 37776
rect 13795 37720 13863 37776
rect 13919 37720 13987 37776
rect 14043 37720 14111 37776
rect 14167 37720 14235 37776
rect 14291 37720 14359 37776
rect 14415 37720 14483 37776
rect 14539 37720 14607 37776
rect 14663 37720 14673 37776
rect 12861 37652 14673 37720
rect 12861 37596 12871 37652
rect 12927 37596 12995 37652
rect 13051 37596 13119 37652
rect 13175 37596 13243 37652
rect 13299 37596 13367 37652
rect 13423 37596 13491 37652
rect 13547 37596 13615 37652
rect 13671 37596 13739 37652
rect 13795 37596 13863 37652
rect 13919 37596 13987 37652
rect 14043 37596 14111 37652
rect 14167 37596 14235 37652
rect 14291 37596 14359 37652
rect 14415 37596 14483 37652
rect 14539 37596 14607 37652
rect 14663 37596 14673 37652
rect 12861 37528 14673 37596
rect 12861 37472 12871 37528
rect 12927 37472 12995 37528
rect 13051 37472 13119 37528
rect 13175 37472 13243 37528
rect 13299 37472 13367 37528
rect 13423 37472 13491 37528
rect 13547 37472 13615 37528
rect 13671 37472 13739 37528
rect 13795 37472 13863 37528
rect 13919 37472 13987 37528
rect 14043 37472 14111 37528
rect 14167 37472 14235 37528
rect 14291 37472 14359 37528
rect 14415 37472 14483 37528
rect 14539 37472 14607 37528
rect 14663 37472 14673 37528
rect 12861 37404 14673 37472
rect 12861 37348 12871 37404
rect 12927 37348 12995 37404
rect 13051 37348 13119 37404
rect 13175 37348 13243 37404
rect 13299 37348 13367 37404
rect 13423 37348 13491 37404
rect 13547 37348 13615 37404
rect 13671 37348 13739 37404
rect 13795 37348 13863 37404
rect 13919 37348 13987 37404
rect 14043 37348 14111 37404
rect 14167 37348 14235 37404
rect 14291 37348 14359 37404
rect 14415 37348 14483 37404
rect 14539 37348 14607 37404
rect 14663 37348 14673 37404
rect 12861 37280 14673 37348
rect 12861 37224 12871 37280
rect 12927 37224 12995 37280
rect 13051 37224 13119 37280
rect 13175 37224 13243 37280
rect 13299 37224 13367 37280
rect 13423 37224 13491 37280
rect 13547 37224 13615 37280
rect 13671 37224 13739 37280
rect 13795 37224 13863 37280
rect 13919 37224 13987 37280
rect 14043 37224 14111 37280
rect 14167 37224 14235 37280
rect 14291 37224 14359 37280
rect 14415 37224 14483 37280
rect 14539 37224 14607 37280
rect 14663 37224 14673 37280
rect 12861 37156 14673 37224
rect 12861 37100 12871 37156
rect 12927 37100 12995 37156
rect 13051 37100 13119 37156
rect 13175 37100 13243 37156
rect 13299 37100 13367 37156
rect 13423 37100 13491 37156
rect 13547 37100 13615 37156
rect 13671 37100 13739 37156
rect 13795 37100 13863 37156
rect 13919 37100 13987 37156
rect 14043 37100 14111 37156
rect 14167 37100 14235 37156
rect 14291 37100 14359 37156
rect 14415 37100 14483 37156
rect 14539 37100 14607 37156
rect 14663 37100 14673 37156
rect 12861 37032 14673 37100
rect 12861 36976 12871 37032
rect 12927 36976 12995 37032
rect 13051 36976 13119 37032
rect 13175 36976 13243 37032
rect 13299 36976 13367 37032
rect 13423 36976 13491 37032
rect 13547 36976 13615 37032
rect 13671 36976 13739 37032
rect 13795 36976 13863 37032
rect 13919 36976 13987 37032
rect 14043 36976 14111 37032
rect 14167 36976 14235 37032
rect 14291 36976 14359 37032
rect 14415 36976 14483 37032
rect 14539 36976 14607 37032
rect 14663 36976 14673 37032
rect 12861 36908 14673 36976
rect 12861 36852 12871 36908
rect 12927 36852 12995 36908
rect 13051 36852 13119 36908
rect 13175 36852 13243 36908
rect 13299 36852 13367 36908
rect 13423 36852 13491 36908
rect 13547 36852 13615 36908
rect 13671 36852 13739 36908
rect 13795 36852 13863 36908
rect 13919 36852 13987 36908
rect 14043 36852 14111 36908
rect 14167 36852 14235 36908
rect 14291 36852 14359 36908
rect 14415 36852 14483 36908
rect 14539 36852 14607 36908
rect 14663 36852 14673 36908
rect 12861 36842 14673 36852
rect -11 36800 86 36824
rect 14892 36824 14902 38176
rect 14958 36824 14989 38176
rect 14892 36800 14989 36824
rect -11 36586 86 36596
rect -11 33614 20 36586
rect 76 33614 86 36586
rect 14892 36586 14989 36596
rect 305 36554 2117 36564
rect 305 36498 315 36554
rect 371 36498 439 36554
rect 495 36498 563 36554
rect 619 36498 687 36554
rect 743 36498 811 36554
rect 867 36498 935 36554
rect 991 36498 1059 36554
rect 1115 36498 1183 36554
rect 1239 36498 1307 36554
rect 1363 36498 1431 36554
rect 1487 36498 1555 36554
rect 1611 36498 1679 36554
rect 1735 36498 1803 36554
rect 1859 36498 1927 36554
rect 1983 36498 2051 36554
rect 2107 36498 2117 36554
rect 305 36430 2117 36498
rect 305 36374 315 36430
rect 371 36374 439 36430
rect 495 36374 563 36430
rect 619 36374 687 36430
rect 743 36374 811 36430
rect 867 36374 935 36430
rect 991 36374 1059 36430
rect 1115 36374 1183 36430
rect 1239 36374 1307 36430
rect 1363 36374 1431 36430
rect 1487 36374 1555 36430
rect 1611 36374 1679 36430
rect 1735 36374 1803 36430
rect 1859 36374 1927 36430
rect 1983 36374 2051 36430
rect 2107 36374 2117 36430
rect 305 36306 2117 36374
rect 305 36250 315 36306
rect 371 36250 439 36306
rect 495 36250 563 36306
rect 619 36250 687 36306
rect 743 36250 811 36306
rect 867 36250 935 36306
rect 991 36250 1059 36306
rect 1115 36250 1183 36306
rect 1239 36250 1307 36306
rect 1363 36250 1431 36306
rect 1487 36250 1555 36306
rect 1611 36250 1679 36306
rect 1735 36250 1803 36306
rect 1859 36250 1927 36306
rect 1983 36250 2051 36306
rect 2107 36250 2117 36306
rect 305 36182 2117 36250
rect 305 36126 315 36182
rect 371 36126 439 36182
rect 495 36126 563 36182
rect 619 36126 687 36182
rect 743 36126 811 36182
rect 867 36126 935 36182
rect 991 36126 1059 36182
rect 1115 36126 1183 36182
rect 1239 36126 1307 36182
rect 1363 36126 1431 36182
rect 1487 36126 1555 36182
rect 1611 36126 1679 36182
rect 1735 36126 1803 36182
rect 1859 36126 1927 36182
rect 1983 36126 2051 36182
rect 2107 36126 2117 36182
rect 305 36058 2117 36126
rect 305 36002 315 36058
rect 371 36002 439 36058
rect 495 36002 563 36058
rect 619 36002 687 36058
rect 743 36002 811 36058
rect 867 36002 935 36058
rect 991 36002 1059 36058
rect 1115 36002 1183 36058
rect 1239 36002 1307 36058
rect 1363 36002 1431 36058
rect 1487 36002 1555 36058
rect 1611 36002 1679 36058
rect 1735 36002 1803 36058
rect 1859 36002 1927 36058
rect 1983 36002 2051 36058
rect 2107 36002 2117 36058
rect 305 35934 2117 36002
rect 305 35878 315 35934
rect 371 35878 439 35934
rect 495 35878 563 35934
rect 619 35878 687 35934
rect 743 35878 811 35934
rect 867 35878 935 35934
rect 991 35878 1059 35934
rect 1115 35878 1183 35934
rect 1239 35878 1307 35934
rect 1363 35878 1431 35934
rect 1487 35878 1555 35934
rect 1611 35878 1679 35934
rect 1735 35878 1803 35934
rect 1859 35878 1927 35934
rect 1983 35878 2051 35934
rect 2107 35878 2117 35934
rect 305 35810 2117 35878
rect 305 35754 315 35810
rect 371 35754 439 35810
rect 495 35754 563 35810
rect 619 35754 687 35810
rect 743 35754 811 35810
rect 867 35754 935 35810
rect 991 35754 1059 35810
rect 1115 35754 1183 35810
rect 1239 35754 1307 35810
rect 1363 35754 1431 35810
rect 1487 35754 1555 35810
rect 1611 35754 1679 35810
rect 1735 35754 1803 35810
rect 1859 35754 1927 35810
rect 1983 35754 2051 35810
rect 2107 35754 2117 35810
rect 305 35686 2117 35754
rect 305 35630 315 35686
rect 371 35630 439 35686
rect 495 35630 563 35686
rect 619 35630 687 35686
rect 743 35630 811 35686
rect 867 35630 935 35686
rect 991 35630 1059 35686
rect 1115 35630 1183 35686
rect 1239 35630 1307 35686
rect 1363 35630 1431 35686
rect 1487 35630 1555 35686
rect 1611 35630 1679 35686
rect 1735 35630 1803 35686
rect 1859 35630 1927 35686
rect 1983 35630 2051 35686
rect 2107 35630 2117 35686
rect 305 35562 2117 35630
rect 305 35506 315 35562
rect 371 35506 439 35562
rect 495 35506 563 35562
rect 619 35506 687 35562
rect 743 35506 811 35562
rect 867 35506 935 35562
rect 991 35506 1059 35562
rect 1115 35506 1183 35562
rect 1239 35506 1307 35562
rect 1363 35506 1431 35562
rect 1487 35506 1555 35562
rect 1611 35506 1679 35562
rect 1735 35506 1803 35562
rect 1859 35506 1927 35562
rect 1983 35506 2051 35562
rect 2107 35506 2117 35562
rect 305 35438 2117 35506
rect 305 35382 315 35438
rect 371 35382 439 35438
rect 495 35382 563 35438
rect 619 35382 687 35438
rect 743 35382 811 35438
rect 867 35382 935 35438
rect 991 35382 1059 35438
rect 1115 35382 1183 35438
rect 1239 35382 1307 35438
rect 1363 35382 1431 35438
rect 1487 35382 1555 35438
rect 1611 35382 1679 35438
rect 1735 35382 1803 35438
rect 1859 35382 1927 35438
rect 1983 35382 2051 35438
rect 2107 35382 2117 35438
rect 305 35314 2117 35382
rect 305 35258 315 35314
rect 371 35258 439 35314
rect 495 35258 563 35314
rect 619 35258 687 35314
rect 743 35258 811 35314
rect 867 35258 935 35314
rect 991 35258 1059 35314
rect 1115 35258 1183 35314
rect 1239 35258 1307 35314
rect 1363 35258 1431 35314
rect 1487 35258 1555 35314
rect 1611 35258 1679 35314
rect 1735 35258 1803 35314
rect 1859 35258 1927 35314
rect 1983 35258 2051 35314
rect 2107 35258 2117 35314
rect 305 35190 2117 35258
rect 305 35134 315 35190
rect 371 35134 439 35190
rect 495 35134 563 35190
rect 619 35134 687 35190
rect 743 35134 811 35190
rect 867 35134 935 35190
rect 991 35134 1059 35190
rect 1115 35134 1183 35190
rect 1239 35134 1307 35190
rect 1363 35134 1431 35190
rect 1487 35134 1555 35190
rect 1611 35134 1679 35190
rect 1735 35134 1803 35190
rect 1859 35134 1927 35190
rect 1983 35134 2051 35190
rect 2107 35134 2117 35190
rect 305 35066 2117 35134
rect 305 35010 315 35066
rect 371 35010 439 35066
rect 495 35010 563 35066
rect 619 35010 687 35066
rect 743 35010 811 35066
rect 867 35010 935 35066
rect 991 35010 1059 35066
rect 1115 35010 1183 35066
rect 1239 35010 1307 35066
rect 1363 35010 1431 35066
rect 1487 35010 1555 35066
rect 1611 35010 1679 35066
rect 1735 35010 1803 35066
rect 1859 35010 1927 35066
rect 1983 35010 2051 35066
rect 2107 35010 2117 35066
rect 305 34942 2117 35010
rect 305 34886 315 34942
rect 371 34886 439 34942
rect 495 34886 563 34942
rect 619 34886 687 34942
rect 743 34886 811 34942
rect 867 34886 935 34942
rect 991 34886 1059 34942
rect 1115 34886 1183 34942
rect 1239 34886 1307 34942
rect 1363 34886 1431 34942
rect 1487 34886 1555 34942
rect 1611 34886 1679 34942
rect 1735 34886 1803 34942
rect 1859 34886 1927 34942
rect 1983 34886 2051 34942
rect 2107 34886 2117 34942
rect 305 34818 2117 34886
rect 305 34762 315 34818
rect 371 34762 439 34818
rect 495 34762 563 34818
rect 619 34762 687 34818
rect 743 34762 811 34818
rect 867 34762 935 34818
rect 991 34762 1059 34818
rect 1115 34762 1183 34818
rect 1239 34762 1307 34818
rect 1363 34762 1431 34818
rect 1487 34762 1555 34818
rect 1611 34762 1679 34818
rect 1735 34762 1803 34818
rect 1859 34762 1927 34818
rect 1983 34762 2051 34818
rect 2107 34762 2117 34818
rect 305 34694 2117 34762
rect 305 34638 315 34694
rect 371 34638 439 34694
rect 495 34638 563 34694
rect 619 34638 687 34694
rect 743 34638 811 34694
rect 867 34638 935 34694
rect 991 34638 1059 34694
rect 1115 34638 1183 34694
rect 1239 34638 1307 34694
rect 1363 34638 1431 34694
rect 1487 34638 1555 34694
rect 1611 34638 1679 34694
rect 1735 34638 1803 34694
rect 1859 34638 1927 34694
rect 1983 34638 2051 34694
rect 2107 34638 2117 34694
rect 305 34570 2117 34638
rect 305 34514 315 34570
rect 371 34514 439 34570
rect 495 34514 563 34570
rect 619 34514 687 34570
rect 743 34514 811 34570
rect 867 34514 935 34570
rect 991 34514 1059 34570
rect 1115 34514 1183 34570
rect 1239 34514 1307 34570
rect 1363 34514 1431 34570
rect 1487 34514 1555 34570
rect 1611 34514 1679 34570
rect 1735 34514 1803 34570
rect 1859 34514 1927 34570
rect 1983 34514 2051 34570
rect 2107 34514 2117 34570
rect 305 34446 2117 34514
rect 305 34390 315 34446
rect 371 34390 439 34446
rect 495 34390 563 34446
rect 619 34390 687 34446
rect 743 34390 811 34446
rect 867 34390 935 34446
rect 991 34390 1059 34446
rect 1115 34390 1183 34446
rect 1239 34390 1307 34446
rect 1363 34390 1431 34446
rect 1487 34390 1555 34446
rect 1611 34390 1679 34446
rect 1735 34390 1803 34446
rect 1859 34390 1927 34446
rect 1983 34390 2051 34446
rect 2107 34390 2117 34446
rect 305 34322 2117 34390
rect 305 34266 315 34322
rect 371 34266 439 34322
rect 495 34266 563 34322
rect 619 34266 687 34322
rect 743 34266 811 34322
rect 867 34266 935 34322
rect 991 34266 1059 34322
rect 1115 34266 1183 34322
rect 1239 34266 1307 34322
rect 1363 34266 1431 34322
rect 1487 34266 1555 34322
rect 1611 34266 1679 34322
rect 1735 34266 1803 34322
rect 1859 34266 1927 34322
rect 1983 34266 2051 34322
rect 2107 34266 2117 34322
rect 305 34198 2117 34266
rect 305 34142 315 34198
rect 371 34142 439 34198
rect 495 34142 563 34198
rect 619 34142 687 34198
rect 743 34142 811 34198
rect 867 34142 935 34198
rect 991 34142 1059 34198
rect 1115 34142 1183 34198
rect 1239 34142 1307 34198
rect 1363 34142 1431 34198
rect 1487 34142 1555 34198
rect 1611 34142 1679 34198
rect 1735 34142 1803 34198
rect 1859 34142 1927 34198
rect 1983 34142 2051 34198
rect 2107 34142 2117 34198
rect 305 34074 2117 34142
rect 305 34018 315 34074
rect 371 34018 439 34074
rect 495 34018 563 34074
rect 619 34018 687 34074
rect 743 34018 811 34074
rect 867 34018 935 34074
rect 991 34018 1059 34074
rect 1115 34018 1183 34074
rect 1239 34018 1307 34074
rect 1363 34018 1431 34074
rect 1487 34018 1555 34074
rect 1611 34018 1679 34074
rect 1735 34018 1803 34074
rect 1859 34018 1927 34074
rect 1983 34018 2051 34074
rect 2107 34018 2117 34074
rect 305 33950 2117 34018
rect 305 33894 315 33950
rect 371 33894 439 33950
rect 495 33894 563 33950
rect 619 33894 687 33950
rect 743 33894 811 33950
rect 867 33894 935 33950
rect 991 33894 1059 33950
rect 1115 33894 1183 33950
rect 1239 33894 1307 33950
rect 1363 33894 1431 33950
rect 1487 33894 1555 33950
rect 1611 33894 1679 33950
rect 1735 33894 1803 33950
rect 1859 33894 1927 33950
rect 1983 33894 2051 33950
rect 2107 33894 2117 33950
rect 305 33826 2117 33894
rect 305 33770 315 33826
rect 371 33770 439 33826
rect 495 33770 563 33826
rect 619 33770 687 33826
rect 743 33770 811 33826
rect 867 33770 935 33826
rect 991 33770 1059 33826
rect 1115 33770 1183 33826
rect 1239 33770 1307 33826
rect 1363 33770 1431 33826
rect 1487 33770 1555 33826
rect 1611 33770 1679 33826
rect 1735 33770 1803 33826
rect 1859 33770 1927 33826
rect 1983 33770 2051 33826
rect 2107 33770 2117 33826
rect 305 33702 2117 33770
rect 305 33646 315 33702
rect 371 33646 439 33702
rect 495 33646 563 33702
rect 619 33646 687 33702
rect 743 33646 811 33702
rect 867 33646 935 33702
rect 991 33646 1059 33702
rect 1115 33646 1183 33702
rect 1239 33646 1307 33702
rect 1363 33646 1431 33702
rect 1487 33646 1555 33702
rect 1611 33646 1679 33702
rect 1735 33646 1803 33702
rect 1859 33646 1927 33702
rect 1983 33646 2051 33702
rect 2107 33646 2117 33702
rect 305 33636 2117 33646
rect 2798 36554 4734 36564
rect 2798 36498 2808 36554
rect 2864 36498 2932 36554
rect 2988 36498 3056 36554
rect 3112 36498 3180 36554
rect 3236 36498 3304 36554
rect 3360 36498 3428 36554
rect 3484 36498 3552 36554
rect 3608 36498 3676 36554
rect 3732 36498 3800 36554
rect 3856 36498 3924 36554
rect 3980 36498 4048 36554
rect 4104 36498 4172 36554
rect 4228 36498 4296 36554
rect 4352 36498 4420 36554
rect 4476 36498 4544 36554
rect 4600 36498 4668 36554
rect 4724 36498 4734 36554
rect 2798 36430 4734 36498
rect 2798 36374 2808 36430
rect 2864 36374 2932 36430
rect 2988 36374 3056 36430
rect 3112 36374 3180 36430
rect 3236 36374 3304 36430
rect 3360 36374 3428 36430
rect 3484 36374 3552 36430
rect 3608 36374 3676 36430
rect 3732 36374 3800 36430
rect 3856 36374 3924 36430
rect 3980 36374 4048 36430
rect 4104 36374 4172 36430
rect 4228 36374 4296 36430
rect 4352 36374 4420 36430
rect 4476 36374 4544 36430
rect 4600 36374 4668 36430
rect 4724 36374 4734 36430
rect 2798 36306 4734 36374
rect 2798 36250 2808 36306
rect 2864 36250 2932 36306
rect 2988 36250 3056 36306
rect 3112 36250 3180 36306
rect 3236 36250 3304 36306
rect 3360 36250 3428 36306
rect 3484 36250 3552 36306
rect 3608 36250 3676 36306
rect 3732 36250 3800 36306
rect 3856 36250 3924 36306
rect 3980 36250 4048 36306
rect 4104 36250 4172 36306
rect 4228 36250 4296 36306
rect 4352 36250 4420 36306
rect 4476 36250 4544 36306
rect 4600 36250 4668 36306
rect 4724 36250 4734 36306
rect 2798 36182 4734 36250
rect 2798 36126 2808 36182
rect 2864 36126 2932 36182
rect 2988 36126 3056 36182
rect 3112 36126 3180 36182
rect 3236 36126 3304 36182
rect 3360 36126 3428 36182
rect 3484 36126 3552 36182
rect 3608 36126 3676 36182
rect 3732 36126 3800 36182
rect 3856 36126 3924 36182
rect 3980 36126 4048 36182
rect 4104 36126 4172 36182
rect 4228 36126 4296 36182
rect 4352 36126 4420 36182
rect 4476 36126 4544 36182
rect 4600 36126 4668 36182
rect 4724 36126 4734 36182
rect 2798 36058 4734 36126
rect 2798 36002 2808 36058
rect 2864 36002 2932 36058
rect 2988 36002 3056 36058
rect 3112 36002 3180 36058
rect 3236 36002 3304 36058
rect 3360 36002 3428 36058
rect 3484 36002 3552 36058
rect 3608 36002 3676 36058
rect 3732 36002 3800 36058
rect 3856 36002 3924 36058
rect 3980 36002 4048 36058
rect 4104 36002 4172 36058
rect 4228 36002 4296 36058
rect 4352 36002 4420 36058
rect 4476 36002 4544 36058
rect 4600 36002 4668 36058
rect 4724 36002 4734 36058
rect 2798 35934 4734 36002
rect 2798 35878 2808 35934
rect 2864 35878 2932 35934
rect 2988 35878 3056 35934
rect 3112 35878 3180 35934
rect 3236 35878 3304 35934
rect 3360 35878 3428 35934
rect 3484 35878 3552 35934
rect 3608 35878 3676 35934
rect 3732 35878 3800 35934
rect 3856 35878 3924 35934
rect 3980 35878 4048 35934
rect 4104 35878 4172 35934
rect 4228 35878 4296 35934
rect 4352 35878 4420 35934
rect 4476 35878 4544 35934
rect 4600 35878 4668 35934
rect 4724 35878 4734 35934
rect 2798 35810 4734 35878
rect 2798 35754 2808 35810
rect 2864 35754 2932 35810
rect 2988 35754 3056 35810
rect 3112 35754 3180 35810
rect 3236 35754 3304 35810
rect 3360 35754 3428 35810
rect 3484 35754 3552 35810
rect 3608 35754 3676 35810
rect 3732 35754 3800 35810
rect 3856 35754 3924 35810
rect 3980 35754 4048 35810
rect 4104 35754 4172 35810
rect 4228 35754 4296 35810
rect 4352 35754 4420 35810
rect 4476 35754 4544 35810
rect 4600 35754 4668 35810
rect 4724 35754 4734 35810
rect 2798 35686 4734 35754
rect 2798 35630 2808 35686
rect 2864 35630 2932 35686
rect 2988 35630 3056 35686
rect 3112 35630 3180 35686
rect 3236 35630 3304 35686
rect 3360 35630 3428 35686
rect 3484 35630 3552 35686
rect 3608 35630 3676 35686
rect 3732 35630 3800 35686
rect 3856 35630 3924 35686
rect 3980 35630 4048 35686
rect 4104 35630 4172 35686
rect 4228 35630 4296 35686
rect 4352 35630 4420 35686
rect 4476 35630 4544 35686
rect 4600 35630 4668 35686
rect 4724 35630 4734 35686
rect 2798 35562 4734 35630
rect 2798 35506 2808 35562
rect 2864 35506 2932 35562
rect 2988 35506 3056 35562
rect 3112 35506 3180 35562
rect 3236 35506 3304 35562
rect 3360 35506 3428 35562
rect 3484 35506 3552 35562
rect 3608 35506 3676 35562
rect 3732 35506 3800 35562
rect 3856 35506 3924 35562
rect 3980 35506 4048 35562
rect 4104 35506 4172 35562
rect 4228 35506 4296 35562
rect 4352 35506 4420 35562
rect 4476 35506 4544 35562
rect 4600 35506 4668 35562
rect 4724 35506 4734 35562
rect 2798 35438 4734 35506
rect 2798 35382 2808 35438
rect 2864 35382 2932 35438
rect 2988 35382 3056 35438
rect 3112 35382 3180 35438
rect 3236 35382 3304 35438
rect 3360 35382 3428 35438
rect 3484 35382 3552 35438
rect 3608 35382 3676 35438
rect 3732 35382 3800 35438
rect 3856 35382 3924 35438
rect 3980 35382 4048 35438
rect 4104 35382 4172 35438
rect 4228 35382 4296 35438
rect 4352 35382 4420 35438
rect 4476 35382 4544 35438
rect 4600 35382 4668 35438
rect 4724 35382 4734 35438
rect 2798 35314 4734 35382
rect 2798 35258 2808 35314
rect 2864 35258 2932 35314
rect 2988 35258 3056 35314
rect 3112 35258 3180 35314
rect 3236 35258 3304 35314
rect 3360 35258 3428 35314
rect 3484 35258 3552 35314
rect 3608 35258 3676 35314
rect 3732 35258 3800 35314
rect 3856 35258 3924 35314
rect 3980 35258 4048 35314
rect 4104 35258 4172 35314
rect 4228 35258 4296 35314
rect 4352 35258 4420 35314
rect 4476 35258 4544 35314
rect 4600 35258 4668 35314
rect 4724 35258 4734 35314
rect 2798 35190 4734 35258
rect 2798 35134 2808 35190
rect 2864 35134 2932 35190
rect 2988 35134 3056 35190
rect 3112 35134 3180 35190
rect 3236 35134 3304 35190
rect 3360 35134 3428 35190
rect 3484 35134 3552 35190
rect 3608 35134 3676 35190
rect 3732 35134 3800 35190
rect 3856 35134 3924 35190
rect 3980 35134 4048 35190
rect 4104 35134 4172 35190
rect 4228 35134 4296 35190
rect 4352 35134 4420 35190
rect 4476 35134 4544 35190
rect 4600 35134 4668 35190
rect 4724 35134 4734 35190
rect 2798 35066 4734 35134
rect 2798 35010 2808 35066
rect 2864 35010 2932 35066
rect 2988 35010 3056 35066
rect 3112 35010 3180 35066
rect 3236 35010 3304 35066
rect 3360 35010 3428 35066
rect 3484 35010 3552 35066
rect 3608 35010 3676 35066
rect 3732 35010 3800 35066
rect 3856 35010 3924 35066
rect 3980 35010 4048 35066
rect 4104 35010 4172 35066
rect 4228 35010 4296 35066
rect 4352 35010 4420 35066
rect 4476 35010 4544 35066
rect 4600 35010 4668 35066
rect 4724 35010 4734 35066
rect 2798 34942 4734 35010
rect 2798 34886 2808 34942
rect 2864 34886 2932 34942
rect 2988 34886 3056 34942
rect 3112 34886 3180 34942
rect 3236 34886 3304 34942
rect 3360 34886 3428 34942
rect 3484 34886 3552 34942
rect 3608 34886 3676 34942
rect 3732 34886 3800 34942
rect 3856 34886 3924 34942
rect 3980 34886 4048 34942
rect 4104 34886 4172 34942
rect 4228 34886 4296 34942
rect 4352 34886 4420 34942
rect 4476 34886 4544 34942
rect 4600 34886 4668 34942
rect 4724 34886 4734 34942
rect 2798 34818 4734 34886
rect 2798 34762 2808 34818
rect 2864 34762 2932 34818
rect 2988 34762 3056 34818
rect 3112 34762 3180 34818
rect 3236 34762 3304 34818
rect 3360 34762 3428 34818
rect 3484 34762 3552 34818
rect 3608 34762 3676 34818
rect 3732 34762 3800 34818
rect 3856 34762 3924 34818
rect 3980 34762 4048 34818
rect 4104 34762 4172 34818
rect 4228 34762 4296 34818
rect 4352 34762 4420 34818
rect 4476 34762 4544 34818
rect 4600 34762 4668 34818
rect 4724 34762 4734 34818
rect 2798 34694 4734 34762
rect 2798 34638 2808 34694
rect 2864 34638 2932 34694
rect 2988 34638 3056 34694
rect 3112 34638 3180 34694
rect 3236 34638 3304 34694
rect 3360 34638 3428 34694
rect 3484 34638 3552 34694
rect 3608 34638 3676 34694
rect 3732 34638 3800 34694
rect 3856 34638 3924 34694
rect 3980 34638 4048 34694
rect 4104 34638 4172 34694
rect 4228 34638 4296 34694
rect 4352 34638 4420 34694
rect 4476 34638 4544 34694
rect 4600 34638 4668 34694
rect 4724 34638 4734 34694
rect 2798 34570 4734 34638
rect 2798 34514 2808 34570
rect 2864 34514 2932 34570
rect 2988 34514 3056 34570
rect 3112 34514 3180 34570
rect 3236 34514 3304 34570
rect 3360 34514 3428 34570
rect 3484 34514 3552 34570
rect 3608 34514 3676 34570
rect 3732 34514 3800 34570
rect 3856 34514 3924 34570
rect 3980 34514 4048 34570
rect 4104 34514 4172 34570
rect 4228 34514 4296 34570
rect 4352 34514 4420 34570
rect 4476 34514 4544 34570
rect 4600 34514 4668 34570
rect 4724 34514 4734 34570
rect 2798 34446 4734 34514
rect 2798 34390 2808 34446
rect 2864 34390 2932 34446
rect 2988 34390 3056 34446
rect 3112 34390 3180 34446
rect 3236 34390 3304 34446
rect 3360 34390 3428 34446
rect 3484 34390 3552 34446
rect 3608 34390 3676 34446
rect 3732 34390 3800 34446
rect 3856 34390 3924 34446
rect 3980 34390 4048 34446
rect 4104 34390 4172 34446
rect 4228 34390 4296 34446
rect 4352 34390 4420 34446
rect 4476 34390 4544 34446
rect 4600 34390 4668 34446
rect 4724 34390 4734 34446
rect 2798 34322 4734 34390
rect 2798 34266 2808 34322
rect 2864 34266 2932 34322
rect 2988 34266 3056 34322
rect 3112 34266 3180 34322
rect 3236 34266 3304 34322
rect 3360 34266 3428 34322
rect 3484 34266 3552 34322
rect 3608 34266 3676 34322
rect 3732 34266 3800 34322
rect 3856 34266 3924 34322
rect 3980 34266 4048 34322
rect 4104 34266 4172 34322
rect 4228 34266 4296 34322
rect 4352 34266 4420 34322
rect 4476 34266 4544 34322
rect 4600 34266 4668 34322
rect 4724 34266 4734 34322
rect 2798 34198 4734 34266
rect 2798 34142 2808 34198
rect 2864 34142 2932 34198
rect 2988 34142 3056 34198
rect 3112 34142 3180 34198
rect 3236 34142 3304 34198
rect 3360 34142 3428 34198
rect 3484 34142 3552 34198
rect 3608 34142 3676 34198
rect 3732 34142 3800 34198
rect 3856 34142 3924 34198
rect 3980 34142 4048 34198
rect 4104 34142 4172 34198
rect 4228 34142 4296 34198
rect 4352 34142 4420 34198
rect 4476 34142 4544 34198
rect 4600 34142 4668 34198
rect 4724 34142 4734 34198
rect 2798 34074 4734 34142
rect 2798 34018 2808 34074
rect 2864 34018 2932 34074
rect 2988 34018 3056 34074
rect 3112 34018 3180 34074
rect 3236 34018 3304 34074
rect 3360 34018 3428 34074
rect 3484 34018 3552 34074
rect 3608 34018 3676 34074
rect 3732 34018 3800 34074
rect 3856 34018 3924 34074
rect 3980 34018 4048 34074
rect 4104 34018 4172 34074
rect 4228 34018 4296 34074
rect 4352 34018 4420 34074
rect 4476 34018 4544 34074
rect 4600 34018 4668 34074
rect 4724 34018 4734 34074
rect 2798 33950 4734 34018
rect 2798 33894 2808 33950
rect 2864 33894 2932 33950
rect 2988 33894 3056 33950
rect 3112 33894 3180 33950
rect 3236 33894 3304 33950
rect 3360 33894 3428 33950
rect 3484 33894 3552 33950
rect 3608 33894 3676 33950
rect 3732 33894 3800 33950
rect 3856 33894 3924 33950
rect 3980 33894 4048 33950
rect 4104 33894 4172 33950
rect 4228 33894 4296 33950
rect 4352 33894 4420 33950
rect 4476 33894 4544 33950
rect 4600 33894 4668 33950
rect 4724 33894 4734 33950
rect 2798 33826 4734 33894
rect 2798 33770 2808 33826
rect 2864 33770 2932 33826
rect 2988 33770 3056 33826
rect 3112 33770 3180 33826
rect 3236 33770 3304 33826
rect 3360 33770 3428 33826
rect 3484 33770 3552 33826
rect 3608 33770 3676 33826
rect 3732 33770 3800 33826
rect 3856 33770 3924 33826
rect 3980 33770 4048 33826
rect 4104 33770 4172 33826
rect 4228 33770 4296 33826
rect 4352 33770 4420 33826
rect 4476 33770 4544 33826
rect 4600 33770 4668 33826
rect 4724 33770 4734 33826
rect 2798 33702 4734 33770
rect 2798 33646 2808 33702
rect 2864 33646 2932 33702
rect 2988 33646 3056 33702
rect 3112 33646 3180 33702
rect 3236 33646 3304 33702
rect 3360 33646 3428 33702
rect 3484 33646 3552 33702
rect 3608 33646 3676 33702
rect 3732 33646 3800 33702
rect 3856 33646 3924 33702
rect 3980 33646 4048 33702
rect 4104 33646 4172 33702
rect 4228 33646 4296 33702
rect 4352 33646 4420 33702
rect 4476 33646 4544 33702
rect 4600 33646 4668 33702
rect 4724 33646 4734 33702
rect 2798 33636 4734 33646
rect 5168 36554 7104 36564
rect 5168 36498 5178 36554
rect 5234 36498 5302 36554
rect 5358 36498 5426 36554
rect 5482 36498 5550 36554
rect 5606 36498 5674 36554
rect 5730 36498 5798 36554
rect 5854 36498 5922 36554
rect 5978 36498 6046 36554
rect 6102 36498 6170 36554
rect 6226 36498 6294 36554
rect 6350 36498 6418 36554
rect 6474 36498 6542 36554
rect 6598 36498 6666 36554
rect 6722 36498 6790 36554
rect 6846 36498 6914 36554
rect 6970 36498 7038 36554
rect 7094 36498 7104 36554
rect 5168 36430 7104 36498
rect 5168 36374 5178 36430
rect 5234 36374 5302 36430
rect 5358 36374 5426 36430
rect 5482 36374 5550 36430
rect 5606 36374 5674 36430
rect 5730 36374 5798 36430
rect 5854 36374 5922 36430
rect 5978 36374 6046 36430
rect 6102 36374 6170 36430
rect 6226 36374 6294 36430
rect 6350 36374 6418 36430
rect 6474 36374 6542 36430
rect 6598 36374 6666 36430
rect 6722 36374 6790 36430
rect 6846 36374 6914 36430
rect 6970 36374 7038 36430
rect 7094 36374 7104 36430
rect 5168 36306 7104 36374
rect 5168 36250 5178 36306
rect 5234 36250 5302 36306
rect 5358 36250 5426 36306
rect 5482 36250 5550 36306
rect 5606 36250 5674 36306
rect 5730 36250 5798 36306
rect 5854 36250 5922 36306
rect 5978 36250 6046 36306
rect 6102 36250 6170 36306
rect 6226 36250 6294 36306
rect 6350 36250 6418 36306
rect 6474 36250 6542 36306
rect 6598 36250 6666 36306
rect 6722 36250 6790 36306
rect 6846 36250 6914 36306
rect 6970 36250 7038 36306
rect 7094 36250 7104 36306
rect 5168 36182 7104 36250
rect 5168 36126 5178 36182
rect 5234 36126 5302 36182
rect 5358 36126 5426 36182
rect 5482 36126 5550 36182
rect 5606 36126 5674 36182
rect 5730 36126 5798 36182
rect 5854 36126 5922 36182
rect 5978 36126 6046 36182
rect 6102 36126 6170 36182
rect 6226 36126 6294 36182
rect 6350 36126 6418 36182
rect 6474 36126 6542 36182
rect 6598 36126 6666 36182
rect 6722 36126 6790 36182
rect 6846 36126 6914 36182
rect 6970 36126 7038 36182
rect 7094 36126 7104 36182
rect 5168 36058 7104 36126
rect 5168 36002 5178 36058
rect 5234 36002 5302 36058
rect 5358 36002 5426 36058
rect 5482 36002 5550 36058
rect 5606 36002 5674 36058
rect 5730 36002 5798 36058
rect 5854 36002 5922 36058
rect 5978 36002 6046 36058
rect 6102 36002 6170 36058
rect 6226 36002 6294 36058
rect 6350 36002 6418 36058
rect 6474 36002 6542 36058
rect 6598 36002 6666 36058
rect 6722 36002 6790 36058
rect 6846 36002 6914 36058
rect 6970 36002 7038 36058
rect 7094 36002 7104 36058
rect 5168 35934 7104 36002
rect 5168 35878 5178 35934
rect 5234 35878 5302 35934
rect 5358 35878 5426 35934
rect 5482 35878 5550 35934
rect 5606 35878 5674 35934
rect 5730 35878 5798 35934
rect 5854 35878 5922 35934
rect 5978 35878 6046 35934
rect 6102 35878 6170 35934
rect 6226 35878 6294 35934
rect 6350 35878 6418 35934
rect 6474 35878 6542 35934
rect 6598 35878 6666 35934
rect 6722 35878 6790 35934
rect 6846 35878 6914 35934
rect 6970 35878 7038 35934
rect 7094 35878 7104 35934
rect 5168 35810 7104 35878
rect 5168 35754 5178 35810
rect 5234 35754 5302 35810
rect 5358 35754 5426 35810
rect 5482 35754 5550 35810
rect 5606 35754 5674 35810
rect 5730 35754 5798 35810
rect 5854 35754 5922 35810
rect 5978 35754 6046 35810
rect 6102 35754 6170 35810
rect 6226 35754 6294 35810
rect 6350 35754 6418 35810
rect 6474 35754 6542 35810
rect 6598 35754 6666 35810
rect 6722 35754 6790 35810
rect 6846 35754 6914 35810
rect 6970 35754 7038 35810
rect 7094 35754 7104 35810
rect 5168 35686 7104 35754
rect 5168 35630 5178 35686
rect 5234 35630 5302 35686
rect 5358 35630 5426 35686
rect 5482 35630 5550 35686
rect 5606 35630 5674 35686
rect 5730 35630 5798 35686
rect 5854 35630 5922 35686
rect 5978 35630 6046 35686
rect 6102 35630 6170 35686
rect 6226 35630 6294 35686
rect 6350 35630 6418 35686
rect 6474 35630 6542 35686
rect 6598 35630 6666 35686
rect 6722 35630 6790 35686
rect 6846 35630 6914 35686
rect 6970 35630 7038 35686
rect 7094 35630 7104 35686
rect 5168 35562 7104 35630
rect 5168 35506 5178 35562
rect 5234 35506 5302 35562
rect 5358 35506 5426 35562
rect 5482 35506 5550 35562
rect 5606 35506 5674 35562
rect 5730 35506 5798 35562
rect 5854 35506 5922 35562
rect 5978 35506 6046 35562
rect 6102 35506 6170 35562
rect 6226 35506 6294 35562
rect 6350 35506 6418 35562
rect 6474 35506 6542 35562
rect 6598 35506 6666 35562
rect 6722 35506 6790 35562
rect 6846 35506 6914 35562
rect 6970 35506 7038 35562
rect 7094 35506 7104 35562
rect 5168 35438 7104 35506
rect 5168 35382 5178 35438
rect 5234 35382 5302 35438
rect 5358 35382 5426 35438
rect 5482 35382 5550 35438
rect 5606 35382 5674 35438
rect 5730 35382 5798 35438
rect 5854 35382 5922 35438
rect 5978 35382 6046 35438
rect 6102 35382 6170 35438
rect 6226 35382 6294 35438
rect 6350 35382 6418 35438
rect 6474 35382 6542 35438
rect 6598 35382 6666 35438
rect 6722 35382 6790 35438
rect 6846 35382 6914 35438
rect 6970 35382 7038 35438
rect 7094 35382 7104 35438
rect 5168 35314 7104 35382
rect 5168 35258 5178 35314
rect 5234 35258 5302 35314
rect 5358 35258 5426 35314
rect 5482 35258 5550 35314
rect 5606 35258 5674 35314
rect 5730 35258 5798 35314
rect 5854 35258 5922 35314
rect 5978 35258 6046 35314
rect 6102 35258 6170 35314
rect 6226 35258 6294 35314
rect 6350 35258 6418 35314
rect 6474 35258 6542 35314
rect 6598 35258 6666 35314
rect 6722 35258 6790 35314
rect 6846 35258 6914 35314
rect 6970 35258 7038 35314
rect 7094 35258 7104 35314
rect 5168 35190 7104 35258
rect 5168 35134 5178 35190
rect 5234 35134 5302 35190
rect 5358 35134 5426 35190
rect 5482 35134 5550 35190
rect 5606 35134 5674 35190
rect 5730 35134 5798 35190
rect 5854 35134 5922 35190
rect 5978 35134 6046 35190
rect 6102 35134 6170 35190
rect 6226 35134 6294 35190
rect 6350 35134 6418 35190
rect 6474 35134 6542 35190
rect 6598 35134 6666 35190
rect 6722 35134 6790 35190
rect 6846 35134 6914 35190
rect 6970 35134 7038 35190
rect 7094 35134 7104 35190
rect 5168 35066 7104 35134
rect 5168 35010 5178 35066
rect 5234 35010 5302 35066
rect 5358 35010 5426 35066
rect 5482 35010 5550 35066
rect 5606 35010 5674 35066
rect 5730 35010 5798 35066
rect 5854 35010 5922 35066
rect 5978 35010 6046 35066
rect 6102 35010 6170 35066
rect 6226 35010 6294 35066
rect 6350 35010 6418 35066
rect 6474 35010 6542 35066
rect 6598 35010 6666 35066
rect 6722 35010 6790 35066
rect 6846 35010 6914 35066
rect 6970 35010 7038 35066
rect 7094 35010 7104 35066
rect 5168 34942 7104 35010
rect 5168 34886 5178 34942
rect 5234 34886 5302 34942
rect 5358 34886 5426 34942
rect 5482 34886 5550 34942
rect 5606 34886 5674 34942
rect 5730 34886 5798 34942
rect 5854 34886 5922 34942
rect 5978 34886 6046 34942
rect 6102 34886 6170 34942
rect 6226 34886 6294 34942
rect 6350 34886 6418 34942
rect 6474 34886 6542 34942
rect 6598 34886 6666 34942
rect 6722 34886 6790 34942
rect 6846 34886 6914 34942
rect 6970 34886 7038 34942
rect 7094 34886 7104 34942
rect 5168 34818 7104 34886
rect 5168 34762 5178 34818
rect 5234 34762 5302 34818
rect 5358 34762 5426 34818
rect 5482 34762 5550 34818
rect 5606 34762 5674 34818
rect 5730 34762 5798 34818
rect 5854 34762 5922 34818
rect 5978 34762 6046 34818
rect 6102 34762 6170 34818
rect 6226 34762 6294 34818
rect 6350 34762 6418 34818
rect 6474 34762 6542 34818
rect 6598 34762 6666 34818
rect 6722 34762 6790 34818
rect 6846 34762 6914 34818
rect 6970 34762 7038 34818
rect 7094 34762 7104 34818
rect 5168 34694 7104 34762
rect 5168 34638 5178 34694
rect 5234 34638 5302 34694
rect 5358 34638 5426 34694
rect 5482 34638 5550 34694
rect 5606 34638 5674 34694
rect 5730 34638 5798 34694
rect 5854 34638 5922 34694
rect 5978 34638 6046 34694
rect 6102 34638 6170 34694
rect 6226 34638 6294 34694
rect 6350 34638 6418 34694
rect 6474 34638 6542 34694
rect 6598 34638 6666 34694
rect 6722 34638 6790 34694
rect 6846 34638 6914 34694
rect 6970 34638 7038 34694
rect 7094 34638 7104 34694
rect 5168 34570 7104 34638
rect 5168 34514 5178 34570
rect 5234 34514 5302 34570
rect 5358 34514 5426 34570
rect 5482 34514 5550 34570
rect 5606 34514 5674 34570
rect 5730 34514 5798 34570
rect 5854 34514 5922 34570
rect 5978 34514 6046 34570
rect 6102 34514 6170 34570
rect 6226 34514 6294 34570
rect 6350 34514 6418 34570
rect 6474 34514 6542 34570
rect 6598 34514 6666 34570
rect 6722 34514 6790 34570
rect 6846 34514 6914 34570
rect 6970 34514 7038 34570
rect 7094 34514 7104 34570
rect 5168 34446 7104 34514
rect 5168 34390 5178 34446
rect 5234 34390 5302 34446
rect 5358 34390 5426 34446
rect 5482 34390 5550 34446
rect 5606 34390 5674 34446
rect 5730 34390 5798 34446
rect 5854 34390 5922 34446
rect 5978 34390 6046 34446
rect 6102 34390 6170 34446
rect 6226 34390 6294 34446
rect 6350 34390 6418 34446
rect 6474 34390 6542 34446
rect 6598 34390 6666 34446
rect 6722 34390 6790 34446
rect 6846 34390 6914 34446
rect 6970 34390 7038 34446
rect 7094 34390 7104 34446
rect 5168 34322 7104 34390
rect 5168 34266 5178 34322
rect 5234 34266 5302 34322
rect 5358 34266 5426 34322
rect 5482 34266 5550 34322
rect 5606 34266 5674 34322
rect 5730 34266 5798 34322
rect 5854 34266 5922 34322
rect 5978 34266 6046 34322
rect 6102 34266 6170 34322
rect 6226 34266 6294 34322
rect 6350 34266 6418 34322
rect 6474 34266 6542 34322
rect 6598 34266 6666 34322
rect 6722 34266 6790 34322
rect 6846 34266 6914 34322
rect 6970 34266 7038 34322
rect 7094 34266 7104 34322
rect 5168 34198 7104 34266
rect 5168 34142 5178 34198
rect 5234 34142 5302 34198
rect 5358 34142 5426 34198
rect 5482 34142 5550 34198
rect 5606 34142 5674 34198
rect 5730 34142 5798 34198
rect 5854 34142 5922 34198
rect 5978 34142 6046 34198
rect 6102 34142 6170 34198
rect 6226 34142 6294 34198
rect 6350 34142 6418 34198
rect 6474 34142 6542 34198
rect 6598 34142 6666 34198
rect 6722 34142 6790 34198
rect 6846 34142 6914 34198
rect 6970 34142 7038 34198
rect 7094 34142 7104 34198
rect 5168 34074 7104 34142
rect 5168 34018 5178 34074
rect 5234 34018 5302 34074
rect 5358 34018 5426 34074
rect 5482 34018 5550 34074
rect 5606 34018 5674 34074
rect 5730 34018 5798 34074
rect 5854 34018 5922 34074
rect 5978 34018 6046 34074
rect 6102 34018 6170 34074
rect 6226 34018 6294 34074
rect 6350 34018 6418 34074
rect 6474 34018 6542 34074
rect 6598 34018 6666 34074
rect 6722 34018 6790 34074
rect 6846 34018 6914 34074
rect 6970 34018 7038 34074
rect 7094 34018 7104 34074
rect 5168 33950 7104 34018
rect 5168 33894 5178 33950
rect 5234 33894 5302 33950
rect 5358 33894 5426 33950
rect 5482 33894 5550 33950
rect 5606 33894 5674 33950
rect 5730 33894 5798 33950
rect 5854 33894 5922 33950
rect 5978 33894 6046 33950
rect 6102 33894 6170 33950
rect 6226 33894 6294 33950
rect 6350 33894 6418 33950
rect 6474 33894 6542 33950
rect 6598 33894 6666 33950
rect 6722 33894 6790 33950
rect 6846 33894 6914 33950
rect 6970 33894 7038 33950
rect 7094 33894 7104 33950
rect 5168 33826 7104 33894
rect 5168 33770 5178 33826
rect 5234 33770 5302 33826
rect 5358 33770 5426 33826
rect 5482 33770 5550 33826
rect 5606 33770 5674 33826
rect 5730 33770 5798 33826
rect 5854 33770 5922 33826
rect 5978 33770 6046 33826
rect 6102 33770 6170 33826
rect 6226 33770 6294 33826
rect 6350 33770 6418 33826
rect 6474 33770 6542 33826
rect 6598 33770 6666 33826
rect 6722 33770 6790 33826
rect 6846 33770 6914 33826
rect 6970 33770 7038 33826
rect 7094 33770 7104 33826
rect 5168 33702 7104 33770
rect 5168 33646 5178 33702
rect 5234 33646 5302 33702
rect 5358 33646 5426 33702
rect 5482 33646 5550 33702
rect 5606 33646 5674 33702
rect 5730 33646 5798 33702
rect 5854 33646 5922 33702
rect 5978 33646 6046 33702
rect 6102 33646 6170 33702
rect 6226 33646 6294 33702
rect 6350 33646 6418 33702
rect 6474 33646 6542 33702
rect 6598 33646 6666 33702
rect 6722 33646 6790 33702
rect 6846 33646 6914 33702
rect 6970 33646 7038 33702
rect 7094 33646 7104 33702
rect 5168 33636 7104 33646
rect 7874 36554 9810 36564
rect 7874 36498 7884 36554
rect 7940 36498 8008 36554
rect 8064 36498 8132 36554
rect 8188 36498 8256 36554
rect 8312 36498 8380 36554
rect 8436 36498 8504 36554
rect 8560 36498 8628 36554
rect 8684 36498 8752 36554
rect 8808 36498 8876 36554
rect 8932 36498 9000 36554
rect 9056 36498 9124 36554
rect 9180 36498 9248 36554
rect 9304 36498 9372 36554
rect 9428 36498 9496 36554
rect 9552 36498 9620 36554
rect 9676 36498 9744 36554
rect 9800 36498 9810 36554
rect 7874 36430 9810 36498
rect 7874 36374 7884 36430
rect 7940 36374 8008 36430
rect 8064 36374 8132 36430
rect 8188 36374 8256 36430
rect 8312 36374 8380 36430
rect 8436 36374 8504 36430
rect 8560 36374 8628 36430
rect 8684 36374 8752 36430
rect 8808 36374 8876 36430
rect 8932 36374 9000 36430
rect 9056 36374 9124 36430
rect 9180 36374 9248 36430
rect 9304 36374 9372 36430
rect 9428 36374 9496 36430
rect 9552 36374 9620 36430
rect 9676 36374 9744 36430
rect 9800 36374 9810 36430
rect 7874 36306 9810 36374
rect 7874 36250 7884 36306
rect 7940 36250 8008 36306
rect 8064 36250 8132 36306
rect 8188 36250 8256 36306
rect 8312 36250 8380 36306
rect 8436 36250 8504 36306
rect 8560 36250 8628 36306
rect 8684 36250 8752 36306
rect 8808 36250 8876 36306
rect 8932 36250 9000 36306
rect 9056 36250 9124 36306
rect 9180 36250 9248 36306
rect 9304 36250 9372 36306
rect 9428 36250 9496 36306
rect 9552 36250 9620 36306
rect 9676 36250 9744 36306
rect 9800 36250 9810 36306
rect 7874 36182 9810 36250
rect 7874 36126 7884 36182
rect 7940 36126 8008 36182
rect 8064 36126 8132 36182
rect 8188 36126 8256 36182
rect 8312 36126 8380 36182
rect 8436 36126 8504 36182
rect 8560 36126 8628 36182
rect 8684 36126 8752 36182
rect 8808 36126 8876 36182
rect 8932 36126 9000 36182
rect 9056 36126 9124 36182
rect 9180 36126 9248 36182
rect 9304 36126 9372 36182
rect 9428 36126 9496 36182
rect 9552 36126 9620 36182
rect 9676 36126 9744 36182
rect 9800 36126 9810 36182
rect 7874 36058 9810 36126
rect 7874 36002 7884 36058
rect 7940 36002 8008 36058
rect 8064 36002 8132 36058
rect 8188 36002 8256 36058
rect 8312 36002 8380 36058
rect 8436 36002 8504 36058
rect 8560 36002 8628 36058
rect 8684 36002 8752 36058
rect 8808 36002 8876 36058
rect 8932 36002 9000 36058
rect 9056 36002 9124 36058
rect 9180 36002 9248 36058
rect 9304 36002 9372 36058
rect 9428 36002 9496 36058
rect 9552 36002 9620 36058
rect 9676 36002 9744 36058
rect 9800 36002 9810 36058
rect 7874 35934 9810 36002
rect 7874 35878 7884 35934
rect 7940 35878 8008 35934
rect 8064 35878 8132 35934
rect 8188 35878 8256 35934
rect 8312 35878 8380 35934
rect 8436 35878 8504 35934
rect 8560 35878 8628 35934
rect 8684 35878 8752 35934
rect 8808 35878 8876 35934
rect 8932 35878 9000 35934
rect 9056 35878 9124 35934
rect 9180 35878 9248 35934
rect 9304 35878 9372 35934
rect 9428 35878 9496 35934
rect 9552 35878 9620 35934
rect 9676 35878 9744 35934
rect 9800 35878 9810 35934
rect 7874 35810 9810 35878
rect 7874 35754 7884 35810
rect 7940 35754 8008 35810
rect 8064 35754 8132 35810
rect 8188 35754 8256 35810
rect 8312 35754 8380 35810
rect 8436 35754 8504 35810
rect 8560 35754 8628 35810
rect 8684 35754 8752 35810
rect 8808 35754 8876 35810
rect 8932 35754 9000 35810
rect 9056 35754 9124 35810
rect 9180 35754 9248 35810
rect 9304 35754 9372 35810
rect 9428 35754 9496 35810
rect 9552 35754 9620 35810
rect 9676 35754 9744 35810
rect 9800 35754 9810 35810
rect 7874 35686 9810 35754
rect 7874 35630 7884 35686
rect 7940 35630 8008 35686
rect 8064 35630 8132 35686
rect 8188 35630 8256 35686
rect 8312 35630 8380 35686
rect 8436 35630 8504 35686
rect 8560 35630 8628 35686
rect 8684 35630 8752 35686
rect 8808 35630 8876 35686
rect 8932 35630 9000 35686
rect 9056 35630 9124 35686
rect 9180 35630 9248 35686
rect 9304 35630 9372 35686
rect 9428 35630 9496 35686
rect 9552 35630 9620 35686
rect 9676 35630 9744 35686
rect 9800 35630 9810 35686
rect 7874 35562 9810 35630
rect 7874 35506 7884 35562
rect 7940 35506 8008 35562
rect 8064 35506 8132 35562
rect 8188 35506 8256 35562
rect 8312 35506 8380 35562
rect 8436 35506 8504 35562
rect 8560 35506 8628 35562
rect 8684 35506 8752 35562
rect 8808 35506 8876 35562
rect 8932 35506 9000 35562
rect 9056 35506 9124 35562
rect 9180 35506 9248 35562
rect 9304 35506 9372 35562
rect 9428 35506 9496 35562
rect 9552 35506 9620 35562
rect 9676 35506 9744 35562
rect 9800 35506 9810 35562
rect 7874 35438 9810 35506
rect 7874 35382 7884 35438
rect 7940 35382 8008 35438
rect 8064 35382 8132 35438
rect 8188 35382 8256 35438
rect 8312 35382 8380 35438
rect 8436 35382 8504 35438
rect 8560 35382 8628 35438
rect 8684 35382 8752 35438
rect 8808 35382 8876 35438
rect 8932 35382 9000 35438
rect 9056 35382 9124 35438
rect 9180 35382 9248 35438
rect 9304 35382 9372 35438
rect 9428 35382 9496 35438
rect 9552 35382 9620 35438
rect 9676 35382 9744 35438
rect 9800 35382 9810 35438
rect 7874 35314 9810 35382
rect 7874 35258 7884 35314
rect 7940 35258 8008 35314
rect 8064 35258 8132 35314
rect 8188 35258 8256 35314
rect 8312 35258 8380 35314
rect 8436 35258 8504 35314
rect 8560 35258 8628 35314
rect 8684 35258 8752 35314
rect 8808 35258 8876 35314
rect 8932 35258 9000 35314
rect 9056 35258 9124 35314
rect 9180 35258 9248 35314
rect 9304 35258 9372 35314
rect 9428 35258 9496 35314
rect 9552 35258 9620 35314
rect 9676 35258 9744 35314
rect 9800 35258 9810 35314
rect 7874 35190 9810 35258
rect 7874 35134 7884 35190
rect 7940 35134 8008 35190
rect 8064 35134 8132 35190
rect 8188 35134 8256 35190
rect 8312 35134 8380 35190
rect 8436 35134 8504 35190
rect 8560 35134 8628 35190
rect 8684 35134 8752 35190
rect 8808 35134 8876 35190
rect 8932 35134 9000 35190
rect 9056 35134 9124 35190
rect 9180 35134 9248 35190
rect 9304 35134 9372 35190
rect 9428 35134 9496 35190
rect 9552 35134 9620 35190
rect 9676 35134 9744 35190
rect 9800 35134 9810 35190
rect 7874 35066 9810 35134
rect 7874 35010 7884 35066
rect 7940 35010 8008 35066
rect 8064 35010 8132 35066
rect 8188 35010 8256 35066
rect 8312 35010 8380 35066
rect 8436 35010 8504 35066
rect 8560 35010 8628 35066
rect 8684 35010 8752 35066
rect 8808 35010 8876 35066
rect 8932 35010 9000 35066
rect 9056 35010 9124 35066
rect 9180 35010 9248 35066
rect 9304 35010 9372 35066
rect 9428 35010 9496 35066
rect 9552 35010 9620 35066
rect 9676 35010 9744 35066
rect 9800 35010 9810 35066
rect 7874 34942 9810 35010
rect 7874 34886 7884 34942
rect 7940 34886 8008 34942
rect 8064 34886 8132 34942
rect 8188 34886 8256 34942
rect 8312 34886 8380 34942
rect 8436 34886 8504 34942
rect 8560 34886 8628 34942
rect 8684 34886 8752 34942
rect 8808 34886 8876 34942
rect 8932 34886 9000 34942
rect 9056 34886 9124 34942
rect 9180 34886 9248 34942
rect 9304 34886 9372 34942
rect 9428 34886 9496 34942
rect 9552 34886 9620 34942
rect 9676 34886 9744 34942
rect 9800 34886 9810 34942
rect 7874 34818 9810 34886
rect 7874 34762 7884 34818
rect 7940 34762 8008 34818
rect 8064 34762 8132 34818
rect 8188 34762 8256 34818
rect 8312 34762 8380 34818
rect 8436 34762 8504 34818
rect 8560 34762 8628 34818
rect 8684 34762 8752 34818
rect 8808 34762 8876 34818
rect 8932 34762 9000 34818
rect 9056 34762 9124 34818
rect 9180 34762 9248 34818
rect 9304 34762 9372 34818
rect 9428 34762 9496 34818
rect 9552 34762 9620 34818
rect 9676 34762 9744 34818
rect 9800 34762 9810 34818
rect 7874 34694 9810 34762
rect 7874 34638 7884 34694
rect 7940 34638 8008 34694
rect 8064 34638 8132 34694
rect 8188 34638 8256 34694
rect 8312 34638 8380 34694
rect 8436 34638 8504 34694
rect 8560 34638 8628 34694
rect 8684 34638 8752 34694
rect 8808 34638 8876 34694
rect 8932 34638 9000 34694
rect 9056 34638 9124 34694
rect 9180 34638 9248 34694
rect 9304 34638 9372 34694
rect 9428 34638 9496 34694
rect 9552 34638 9620 34694
rect 9676 34638 9744 34694
rect 9800 34638 9810 34694
rect 7874 34570 9810 34638
rect 7874 34514 7884 34570
rect 7940 34514 8008 34570
rect 8064 34514 8132 34570
rect 8188 34514 8256 34570
rect 8312 34514 8380 34570
rect 8436 34514 8504 34570
rect 8560 34514 8628 34570
rect 8684 34514 8752 34570
rect 8808 34514 8876 34570
rect 8932 34514 9000 34570
rect 9056 34514 9124 34570
rect 9180 34514 9248 34570
rect 9304 34514 9372 34570
rect 9428 34514 9496 34570
rect 9552 34514 9620 34570
rect 9676 34514 9744 34570
rect 9800 34514 9810 34570
rect 7874 34446 9810 34514
rect 7874 34390 7884 34446
rect 7940 34390 8008 34446
rect 8064 34390 8132 34446
rect 8188 34390 8256 34446
rect 8312 34390 8380 34446
rect 8436 34390 8504 34446
rect 8560 34390 8628 34446
rect 8684 34390 8752 34446
rect 8808 34390 8876 34446
rect 8932 34390 9000 34446
rect 9056 34390 9124 34446
rect 9180 34390 9248 34446
rect 9304 34390 9372 34446
rect 9428 34390 9496 34446
rect 9552 34390 9620 34446
rect 9676 34390 9744 34446
rect 9800 34390 9810 34446
rect 7874 34322 9810 34390
rect 7874 34266 7884 34322
rect 7940 34266 8008 34322
rect 8064 34266 8132 34322
rect 8188 34266 8256 34322
rect 8312 34266 8380 34322
rect 8436 34266 8504 34322
rect 8560 34266 8628 34322
rect 8684 34266 8752 34322
rect 8808 34266 8876 34322
rect 8932 34266 9000 34322
rect 9056 34266 9124 34322
rect 9180 34266 9248 34322
rect 9304 34266 9372 34322
rect 9428 34266 9496 34322
rect 9552 34266 9620 34322
rect 9676 34266 9744 34322
rect 9800 34266 9810 34322
rect 7874 34198 9810 34266
rect 7874 34142 7884 34198
rect 7940 34142 8008 34198
rect 8064 34142 8132 34198
rect 8188 34142 8256 34198
rect 8312 34142 8380 34198
rect 8436 34142 8504 34198
rect 8560 34142 8628 34198
rect 8684 34142 8752 34198
rect 8808 34142 8876 34198
rect 8932 34142 9000 34198
rect 9056 34142 9124 34198
rect 9180 34142 9248 34198
rect 9304 34142 9372 34198
rect 9428 34142 9496 34198
rect 9552 34142 9620 34198
rect 9676 34142 9744 34198
rect 9800 34142 9810 34198
rect 7874 34074 9810 34142
rect 7874 34018 7884 34074
rect 7940 34018 8008 34074
rect 8064 34018 8132 34074
rect 8188 34018 8256 34074
rect 8312 34018 8380 34074
rect 8436 34018 8504 34074
rect 8560 34018 8628 34074
rect 8684 34018 8752 34074
rect 8808 34018 8876 34074
rect 8932 34018 9000 34074
rect 9056 34018 9124 34074
rect 9180 34018 9248 34074
rect 9304 34018 9372 34074
rect 9428 34018 9496 34074
rect 9552 34018 9620 34074
rect 9676 34018 9744 34074
rect 9800 34018 9810 34074
rect 7874 33950 9810 34018
rect 7874 33894 7884 33950
rect 7940 33894 8008 33950
rect 8064 33894 8132 33950
rect 8188 33894 8256 33950
rect 8312 33894 8380 33950
rect 8436 33894 8504 33950
rect 8560 33894 8628 33950
rect 8684 33894 8752 33950
rect 8808 33894 8876 33950
rect 8932 33894 9000 33950
rect 9056 33894 9124 33950
rect 9180 33894 9248 33950
rect 9304 33894 9372 33950
rect 9428 33894 9496 33950
rect 9552 33894 9620 33950
rect 9676 33894 9744 33950
rect 9800 33894 9810 33950
rect 7874 33826 9810 33894
rect 7874 33770 7884 33826
rect 7940 33770 8008 33826
rect 8064 33770 8132 33826
rect 8188 33770 8256 33826
rect 8312 33770 8380 33826
rect 8436 33770 8504 33826
rect 8560 33770 8628 33826
rect 8684 33770 8752 33826
rect 8808 33770 8876 33826
rect 8932 33770 9000 33826
rect 9056 33770 9124 33826
rect 9180 33770 9248 33826
rect 9304 33770 9372 33826
rect 9428 33770 9496 33826
rect 9552 33770 9620 33826
rect 9676 33770 9744 33826
rect 9800 33770 9810 33826
rect 7874 33702 9810 33770
rect 7874 33646 7884 33702
rect 7940 33646 8008 33702
rect 8064 33646 8132 33702
rect 8188 33646 8256 33702
rect 8312 33646 8380 33702
rect 8436 33646 8504 33702
rect 8560 33646 8628 33702
rect 8684 33646 8752 33702
rect 8808 33646 8876 33702
rect 8932 33646 9000 33702
rect 9056 33646 9124 33702
rect 9180 33646 9248 33702
rect 9304 33646 9372 33702
rect 9428 33646 9496 33702
rect 9552 33646 9620 33702
rect 9676 33646 9744 33702
rect 9800 33646 9810 33702
rect 7874 33636 9810 33646
rect 10244 36554 12180 36564
rect 10244 36498 10254 36554
rect 10310 36498 10378 36554
rect 10434 36498 10502 36554
rect 10558 36498 10626 36554
rect 10682 36498 10750 36554
rect 10806 36498 10874 36554
rect 10930 36498 10998 36554
rect 11054 36498 11122 36554
rect 11178 36498 11246 36554
rect 11302 36498 11370 36554
rect 11426 36498 11494 36554
rect 11550 36498 11618 36554
rect 11674 36498 11742 36554
rect 11798 36498 11866 36554
rect 11922 36498 11990 36554
rect 12046 36498 12114 36554
rect 12170 36498 12180 36554
rect 10244 36430 12180 36498
rect 10244 36374 10254 36430
rect 10310 36374 10378 36430
rect 10434 36374 10502 36430
rect 10558 36374 10626 36430
rect 10682 36374 10750 36430
rect 10806 36374 10874 36430
rect 10930 36374 10998 36430
rect 11054 36374 11122 36430
rect 11178 36374 11246 36430
rect 11302 36374 11370 36430
rect 11426 36374 11494 36430
rect 11550 36374 11618 36430
rect 11674 36374 11742 36430
rect 11798 36374 11866 36430
rect 11922 36374 11990 36430
rect 12046 36374 12114 36430
rect 12170 36374 12180 36430
rect 10244 36306 12180 36374
rect 10244 36250 10254 36306
rect 10310 36250 10378 36306
rect 10434 36250 10502 36306
rect 10558 36250 10626 36306
rect 10682 36250 10750 36306
rect 10806 36250 10874 36306
rect 10930 36250 10998 36306
rect 11054 36250 11122 36306
rect 11178 36250 11246 36306
rect 11302 36250 11370 36306
rect 11426 36250 11494 36306
rect 11550 36250 11618 36306
rect 11674 36250 11742 36306
rect 11798 36250 11866 36306
rect 11922 36250 11990 36306
rect 12046 36250 12114 36306
rect 12170 36250 12180 36306
rect 10244 36182 12180 36250
rect 10244 36126 10254 36182
rect 10310 36126 10378 36182
rect 10434 36126 10502 36182
rect 10558 36126 10626 36182
rect 10682 36126 10750 36182
rect 10806 36126 10874 36182
rect 10930 36126 10998 36182
rect 11054 36126 11122 36182
rect 11178 36126 11246 36182
rect 11302 36126 11370 36182
rect 11426 36126 11494 36182
rect 11550 36126 11618 36182
rect 11674 36126 11742 36182
rect 11798 36126 11866 36182
rect 11922 36126 11990 36182
rect 12046 36126 12114 36182
rect 12170 36126 12180 36182
rect 10244 36058 12180 36126
rect 10244 36002 10254 36058
rect 10310 36002 10378 36058
rect 10434 36002 10502 36058
rect 10558 36002 10626 36058
rect 10682 36002 10750 36058
rect 10806 36002 10874 36058
rect 10930 36002 10998 36058
rect 11054 36002 11122 36058
rect 11178 36002 11246 36058
rect 11302 36002 11370 36058
rect 11426 36002 11494 36058
rect 11550 36002 11618 36058
rect 11674 36002 11742 36058
rect 11798 36002 11866 36058
rect 11922 36002 11990 36058
rect 12046 36002 12114 36058
rect 12170 36002 12180 36058
rect 10244 35934 12180 36002
rect 10244 35878 10254 35934
rect 10310 35878 10378 35934
rect 10434 35878 10502 35934
rect 10558 35878 10626 35934
rect 10682 35878 10750 35934
rect 10806 35878 10874 35934
rect 10930 35878 10998 35934
rect 11054 35878 11122 35934
rect 11178 35878 11246 35934
rect 11302 35878 11370 35934
rect 11426 35878 11494 35934
rect 11550 35878 11618 35934
rect 11674 35878 11742 35934
rect 11798 35878 11866 35934
rect 11922 35878 11990 35934
rect 12046 35878 12114 35934
rect 12170 35878 12180 35934
rect 10244 35810 12180 35878
rect 10244 35754 10254 35810
rect 10310 35754 10378 35810
rect 10434 35754 10502 35810
rect 10558 35754 10626 35810
rect 10682 35754 10750 35810
rect 10806 35754 10874 35810
rect 10930 35754 10998 35810
rect 11054 35754 11122 35810
rect 11178 35754 11246 35810
rect 11302 35754 11370 35810
rect 11426 35754 11494 35810
rect 11550 35754 11618 35810
rect 11674 35754 11742 35810
rect 11798 35754 11866 35810
rect 11922 35754 11990 35810
rect 12046 35754 12114 35810
rect 12170 35754 12180 35810
rect 10244 35686 12180 35754
rect 10244 35630 10254 35686
rect 10310 35630 10378 35686
rect 10434 35630 10502 35686
rect 10558 35630 10626 35686
rect 10682 35630 10750 35686
rect 10806 35630 10874 35686
rect 10930 35630 10998 35686
rect 11054 35630 11122 35686
rect 11178 35630 11246 35686
rect 11302 35630 11370 35686
rect 11426 35630 11494 35686
rect 11550 35630 11618 35686
rect 11674 35630 11742 35686
rect 11798 35630 11866 35686
rect 11922 35630 11990 35686
rect 12046 35630 12114 35686
rect 12170 35630 12180 35686
rect 10244 35562 12180 35630
rect 10244 35506 10254 35562
rect 10310 35506 10378 35562
rect 10434 35506 10502 35562
rect 10558 35506 10626 35562
rect 10682 35506 10750 35562
rect 10806 35506 10874 35562
rect 10930 35506 10998 35562
rect 11054 35506 11122 35562
rect 11178 35506 11246 35562
rect 11302 35506 11370 35562
rect 11426 35506 11494 35562
rect 11550 35506 11618 35562
rect 11674 35506 11742 35562
rect 11798 35506 11866 35562
rect 11922 35506 11990 35562
rect 12046 35506 12114 35562
rect 12170 35506 12180 35562
rect 10244 35438 12180 35506
rect 10244 35382 10254 35438
rect 10310 35382 10378 35438
rect 10434 35382 10502 35438
rect 10558 35382 10626 35438
rect 10682 35382 10750 35438
rect 10806 35382 10874 35438
rect 10930 35382 10998 35438
rect 11054 35382 11122 35438
rect 11178 35382 11246 35438
rect 11302 35382 11370 35438
rect 11426 35382 11494 35438
rect 11550 35382 11618 35438
rect 11674 35382 11742 35438
rect 11798 35382 11866 35438
rect 11922 35382 11990 35438
rect 12046 35382 12114 35438
rect 12170 35382 12180 35438
rect 10244 35314 12180 35382
rect 10244 35258 10254 35314
rect 10310 35258 10378 35314
rect 10434 35258 10502 35314
rect 10558 35258 10626 35314
rect 10682 35258 10750 35314
rect 10806 35258 10874 35314
rect 10930 35258 10998 35314
rect 11054 35258 11122 35314
rect 11178 35258 11246 35314
rect 11302 35258 11370 35314
rect 11426 35258 11494 35314
rect 11550 35258 11618 35314
rect 11674 35258 11742 35314
rect 11798 35258 11866 35314
rect 11922 35258 11990 35314
rect 12046 35258 12114 35314
rect 12170 35258 12180 35314
rect 10244 35190 12180 35258
rect 10244 35134 10254 35190
rect 10310 35134 10378 35190
rect 10434 35134 10502 35190
rect 10558 35134 10626 35190
rect 10682 35134 10750 35190
rect 10806 35134 10874 35190
rect 10930 35134 10998 35190
rect 11054 35134 11122 35190
rect 11178 35134 11246 35190
rect 11302 35134 11370 35190
rect 11426 35134 11494 35190
rect 11550 35134 11618 35190
rect 11674 35134 11742 35190
rect 11798 35134 11866 35190
rect 11922 35134 11990 35190
rect 12046 35134 12114 35190
rect 12170 35134 12180 35190
rect 10244 35066 12180 35134
rect 10244 35010 10254 35066
rect 10310 35010 10378 35066
rect 10434 35010 10502 35066
rect 10558 35010 10626 35066
rect 10682 35010 10750 35066
rect 10806 35010 10874 35066
rect 10930 35010 10998 35066
rect 11054 35010 11122 35066
rect 11178 35010 11246 35066
rect 11302 35010 11370 35066
rect 11426 35010 11494 35066
rect 11550 35010 11618 35066
rect 11674 35010 11742 35066
rect 11798 35010 11866 35066
rect 11922 35010 11990 35066
rect 12046 35010 12114 35066
rect 12170 35010 12180 35066
rect 10244 34942 12180 35010
rect 10244 34886 10254 34942
rect 10310 34886 10378 34942
rect 10434 34886 10502 34942
rect 10558 34886 10626 34942
rect 10682 34886 10750 34942
rect 10806 34886 10874 34942
rect 10930 34886 10998 34942
rect 11054 34886 11122 34942
rect 11178 34886 11246 34942
rect 11302 34886 11370 34942
rect 11426 34886 11494 34942
rect 11550 34886 11618 34942
rect 11674 34886 11742 34942
rect 11798 34886 11866 34942
rect 11922 34886 11990 34942
rect 12046 34886 12114 34942
rect 12170 34886 12180 34942
rect 10244 34818 12180 34886
rect 10244 34762 10254 34818
rect 10310 34762 10378 34818
rect 10434 34762 10502 34818
rect 10558 34762 10626 34818
rect 10682 34762 10750 34818
rect 10806 34762 10874 34818
rect 10930 34762 10998 34818
rect 11054 34762 11122 34818
rect 11178 34762 11246 34818
rect 11302 34762 11370 34818
rect 11426 34762 11494 34818
rect 11550 34762 11618 34818
rect 11674 34762 11742 34818
rect 11798 34762 11866 34818
rect 11922 34762 11990 34818
rect 12046 34762 12114 34818
rect 12170 34762 12180 34818
rect 10244 34694 12180 34762
rect 10244 34638 10254 34694
rect 10310 34638 10378 34694
rect 10434 34638 10502 34694
rect 10558 34638 10626 34694
rect 10682 34638 10750 34694
rect 10806 34638 10874 34694
rect 10930 34638 10998 34694
rect 11054 34638 11122 34694
rect 11178 34638 11246 34694
rect 11302 34638 11370 34694
rect 11426 34638 11494 34694
rect 11550 34638 11618 34694
rect 11674 34638 11742 34694
rect 11798 34638 11866 34694
rect 11922 34638 11990 34694
rect 12046 34638 12114 34694
rect 12170 34638 12180 34694
rect 10244 34570 12180 34638
rect 10244 34514 10254 34570
rect 10310 34514 10378 34570
rect 10434 34514 10502 34570
rect 10558 34514 10626 34570
rect 10682 34514 10750 34570
rect 10806 34514 10874 34570
rect 10930 34514 10998 34570
rect 11054 34514 11122 34570
rect 11178 34514 11246 34570
rect 11302 34514 11370 34570
rect 11426 34514 11494 34570
rect 11550 34514 11618 34570
rect 11674 34514 11742 34570
rect 11798 34514 11866 34570
rect 11922 34514 11990 34570
rect 12046 34514 12114 34570
rect 12170 34514 12180 34570
rect 10244 34446 12180 34514
rect 10244 34390 10254 34446
rect 10310 34390 10378 34446
rect 10434 34390 10502 34446
rect 10558 34390 10626 34446
rect 10682 34390 10750 34446
rect 10806 34390 10874 34446
rect 10930 34390 10998 34446
rect 11054 34390 11122 34446
rect 11178 34390 11246 34446
rect 11302 34390 11370 34446
rect 11426 34390 11494 34446
rect 11550 34390 11618 34446
rect 11674 34390 11742 34446
rect 11798 34390 11866 34446
rect 11922 34390 11990 34446
rect 12046 34390 12114 34446
rect 12170 34390 12180 34446
rect 10244 34322 12180 34390
rect 10244 34266 10254 34322
rect 10310 34266 10378 34322
rect 10434 34266 10502 34322
rect 10558 34266 10626 34322
rect 10682 34266 10750 34322
rect 10806 34266 10874 34322
rect 10930 34266 10998 34322
rect 11054 34266 11122 34322
rect 11178 34266 11246 34322
rect 11302 34266 11370 34322
rect 11426 34266 11494 34322
rect 11550 34266 11618 34322
rect 11674 34266 11742 34322
rect 11798 34266 11866 34322
rect 11922 34266 11990 34322
rect 12046 34266 12114 34322
rect 12170 34266 12180 34322
rect 10244 34198 12180 34266
rect 10244 34142 10254 34198
rect 10310 34142 10378 34198
rect 10434 34142 10502 34198
rect 10558 34142 10626 34198
rect 10682 34142 10750 34198
rect 10806 34142 10874 34198
rect 10930 34142 10998 34198
rect 11054 34142 11122 34198
rect 11178 34142 11246 34198
rect 11302 34142 11370 34198
rect 11426 34142 11494 34198
rect 11550 34142 11618 34198
rect 11674 34142 11742 34198
rect 11798 34142 11866 34198
rect 11922 34142 11990 34198
rect 12046 34142 12114 34198
rect 12170 34142 12180 34198
rect 10244 34074 12180 34142
rect 10244 34018 10254 34074
rect 10310 34018 10378 34074
rect 10434 34018 10502 34074
rect 10558 34018 10626 34074
rect 10682 34018 10750 34074
rect 10806 34018 10874 34074
rect 10930 34018 10998 34074
rect 11054 34018 11122 34074
rect 11178 34018 11246 34074
rect 11302 34018 11370 34074
rect 11426 34018 11494 34074
rect 11550 34018 11618 34074
rect 11674 34018 11742 34074
rect 11798 34018 11866 34074
rect 11922 34018 11990 34074
rect 12046 34018 12114 34074
rect 12170 34018 12180 34074
rect 10244 33950 12180 34018
rect 10244 33894 10254 33950
rect 10310 33894 10378 33950
rect 10434 33894 10502 33950
rect 10558 33894 10626 33950
rect 10682 33894 10750 33950
rect 10806 33894 10874 33950
rect 10930 33894 10998 33950
rect 11054 33894 11122 33950
rect 11178 33894 11246 33950
rect 11302 33894 11370 33950
rect 11426 33894 11494 33950
rect 11550 33894 11618 33950
rect 11674 33894 11742 33950
rect 11798 33894 11866 33950
rect 11922 33894 11990 33950
rect 12046 33894 12114 33950
rect 12170 33894 12180 33950
rect 10244 33826 12180 33894
rect 10244 33770 10254 33826
rect 10310 33770 10378 33826
rect 10434 33770 10502 33826
rect 10558 33770 10626 33826
rect 10682 33770 10750 33826
rect 10806 33770 10874 33826
rect 10930 33770 10998 33826
rect 11054 33770 11122 33826
rect 11178 33770 11246 33826
rect 11302 33770 11370 33826
rect 11426 33770 11494 33826
rect 11550 33770 11618 33826
rect 11674 33770 11742 33826
rect 11798 33770 11866 33826
rect 11922 33770 11990 33826
rect 12046 33770 12114 33826
rect 12170 33770 12180 33826
rect 10244 33702 12180 33770
rect 10244 33646 10254 33702
rect 10310 33646 10378 33702
rect 10434 33646 10502 33702
rect 10558 33646 10626 33702
rect 10682 33646 10750 33702
rect 10806 33646 10874 33702
rect 10930 33646 10998 33702
rect 11054 33646 11122 33702
rect 11178 33646 11246 33702
rect 11302 33646 11370 33702
rect 11426 33646 11494 33702
rect 11550 33646 11618 33702
rect 11674 33646 11742 33702
rect 11798 33646 11866 33702
rect 11922 33646 11990 33702
rect 12046 33646 12114 33702
rect 12170 33646 12180 33702
rect 10244 33636 12180 33646
rect 12861 36554 14673 36564
rect 12861 36498 12871 36554
rect 12927 36498 12995 36554
rect 13051 36498 13119 36554
rect 13175 36498 13243 36554
rect 13299 36498 13367 36554
rect 13423 36498 13491 36554
rect 13547 36498 13615 36554
rect 13671 36498 13739 36554
rect 13795 36498 13863 36554
rect 13919 36498 13987 36554
rect 14043 36498 14111 36554
rect 14167 36498 14235 36554
rect 14291 36498 14359 36554
rect 14415 36498 14483 36554
rect 14539 36498 14607 36554
rect 14663 36498 14673 36554
rect 12861 36430 14673 36498
rect 12861 36374 12871 36430
rect 12927 36374 12995 36430
rect 13051 36374 13119 36430
rect 13175 36374 13243 36430
rect 13299 36374 13367 36430
rect 13423 36374 13491 36430
rect 13547 36374 13615 36430
rect 13671 36374 13739 36430
rect 13795 36374 13863 36430
rect 13919 36374 13987 36430
rect 14043 36374 14111 36430
rect 14167 36374 14235 36430
rect 14291 36374 14359 36430
rect 14415 36374 14483 36430
rect 14539 36374 14607 36430
rect 14663 36374 14673 36430
rect 12861 36306 14673 36374
rect 12861 36250 12871 36306
rect 12927 36250 12995 36306
rect 13051 36250 13119 36306
rect 13175 36250 13243 36306
rect 13299 36250 13367 36306
rect 13423 36250 13491 36306
rect 13547 36250 13615 36306
rect 13671 36250 13739 36306
rect 13795 36250 13863 36306
rect 13919 36250 13987 36306
rect 14043 36250 14111 36306
rect 14167 36250 14235 36306
rect 14291 36250 14359 36306
rect 14415 36250 14483 36306
rect 14539 36250 14607 36306
rect 14663 36250 14673 36306
rect 12861 36182 14673 36250
rect 12861 36126 12871 36182
rect 12927 36126 12995 36182
rect 13051 36126 13119 36182
rect 13175 36126 13243 36182
rect 13299 36126 13367 36182
rect 13423 36126 13491 36182
rect 13547 36126 13615 36182
rect 13671 36126 13739 36182
rect 13795 36126 13863 36182
rect 13919 36126 13987 36182
rect 14043 36126 14111 36182
rect 14167 36126 14235 36182
rect 14291 36126 14359 36182
rect 14415 36126 14483 36182
rect 14539 36126 14607 36182
rect 14663 36126 14673 36182
rect 12861 36058 14673 36126
rect 12861 36002 12871 36058
rect 12927 36002 12995 36058
rect 13051 36002 13119 36058
rect 13175 36002 13243 36058
rect 13299 36002 13367 36058
rect 13423 36002 13491 36058
rect 13547 36002 13615 36058
rect 13671 36002 13739 36058
rect 13795 36002 13863 36058
rect 13919 36002 13987 36058
rect 14043 36002 14111 36058
rect 14167 36002 14235 36058
rect 14291 36002 14359 36058
rect 14415 36002 14483 36058
rect 14539 36002 14607 36058
rect 14663 36002 14673 36058
rect 12861 35934 14673 36002
rect 12861 35878 12871 35934
rect 12927 35878 12995 35934
rect 13051 35878 13119 35934
rect 13175 35878 13243 35934
rect 13299 35878 13367 35934
rect 13423 35878 13491 35934
rect 13547 35878 13615 35934
rect 13671 35878 13739 35934
rect 13795 35878 13863 35934
rect 13919 35878 13987 35934
rect 14043 35878 14111 35934
rect 14167 35878 14235 35934
rect 14291 35878 14359 35934
rect 14415 35878 14483 35934
rect 14539 35878 14607 35934
rect 14663 35878 14673 35934
rect 12861 35810 14673 35878
rect 12861 35754 12871 35810
rect 12927 35754 12995 35810
rect 13051 35754 13119 35810
rect 13175 35754 13243 35810
rect 13299 35754 13367 35810
rect 13423 35754 13491 35810
rect 13547 35754 13615 35810
rect 13671 35754 13739 35810
rect 13795 35754 13863 35810
rect 13919 35754 13987 35810
rect 14043 35754 14111 35810
rect 14167 35754 14235 35810
rect 14291 35754 14359 35810
rect 14415 35754 14483 35810
rect 14539 35754 14607 35810
rect 14663 35754 14673 35810
rect 12861 35686 14673 35754
rect 12861 35630 12871 35686
rect 12927 35630 12995 35686
rect 13051 35630 13119 35686
rect 13175 35630 13243 35686
rect 13299 35630 13367 35686
rect 13423 35630 13491 35686
rect 13547 35630 13615 35686
rect 13671 35630 13739 35686
rect 13795 35630 13863 35686
rect 13919 35630 13987 35686
rect 14043 35630 14111 35686
rect 14167 35630 14235 35686
rect 14291 35630 14359 35686
rect 14415 35630 14483 35686
rect 14539 35630 14607 35686
rect 14663 35630 14673 35686
rect 12861 35562 14673 35630
rect 12861 35506 12871 35562
rect 12927 35506 12995 35562
rect 13051 35506 13119 35562
rect 13175 35506 13243 35562
rect 13299 35506 13367 35562
rect 13423 35506 13491 35562
rect 13547 35506 13615 35562
rect 13671 35506 13739 35562
rect 13795 35506 13863 35562
rect 13919 35506 13987 35562
rect 14043 35506 14111 35562
rect 14167 35506 14235 35562
rect 14291 35506 14359 35562
rect 14415 35506 14483 35562
rect 14539 35506 14607 35562
rect 14663 35506 14673 35562
rect 12861 35438 14673 35506
rect 12861 35382 12871 35438
rect 12927 35382 12995 35438
rect 13051 35382 13119 35438
rect 13175 35382 13243 35438
rect 13299 35382 13367 35438
rect 13423 35382 13491 35438
rect 13547 35382 13615 35438
rect 13671 35382 13739 35438
rect 13795 35382 13863 35438
rect 13919 35382 13987 35438
rect 14043 35382 14111 35438
rect 14167 35382 14235 35438
rect 14291 35382 14359 35438
rect 14415 35382 14483 35438
rect 14539 35382 14607 35438
rect 14663 35382 14673 35438
rect 12861 35314 14673 35382
rect 12861 35258 12871 35314
rect 12927 35258 12995 35314
rect 13051 35258 13119 35314
rect 13175 35258 13243 35314
rect 13299 35258 13367 35314
rect 13423 35258 13491 35314
rect 13547 35258 13615 35314
rect 13671 35258 13739 35314
rect 13795 35258 13863 35314
rect 13919 35258 13987 35314
rect 14043 35258 14111 35314
rect 14167 35258 14235 35314
rect 14291 35258 14359 35314
rect 14415 35258 14483 35314
rect 14539 35258 14607 35314
rect 14663 35258 14673 35314
rect 12861 35190 14673 35258
rect 12861 35134 12871 35190
rect 12927 35134 12995 35190
rect 13051 35134 13119 35190
rect 13175 35134 13243 35190
rect 13299 35134 13367 35190
rect 13423 35134 13491 35190
rect 13547 35134 13615 35190
rect 13671 35134 13739 35190
rect 13795 35134 13863 35190
rect 13919 35134 13987 35190
rect 14043 35134 14111 35190
rect 14167 35134 14235 35190
rect 14291 35134 14359 35190
rect 14415 35134 14483 35190
rect 14539 35134 14607 35190
rect 14663 35134 14673 35190
rect 12861 35066 14673 35134
rect 12861 35010 12871 35066
rect 12927 35010 12995 35066
rect 13051 35010 13119 35066
rect 13175 35010 13243 35066
rect 13299 35010 13367 35066
rect 13423 35010 13491 35066
rect 13547 35010 13615 35066
rect 13671 35010 13739 35066
rect 13795 35010 13863 35066
rect 13919 35010 13987 35066
rect 14043 35010 14111 35066
rect 14167 35010 14235 35066
rect 14291 35010 14359 35066
rect 14415 35010 14483 35066
rect 14539 35010 14607 35066
rect 14663 35010 14673 35066
rect 12861 34942 14673 35010
rect 12861 34886 12871 34942
rect 12927 34886 12995 34942
rect 13051 34886 13119 34942
rect 13175 34886 13243 34942
rect 13299 34886 13367 34942
rect 13423 34886 13491 34942
rect 13547 34886 13615 34942
rect 13671 34886 13739 34942
rect 13795 34886 13863 34942
rect 13919 34886 13987 34942
rect 14043 34886 14111 34942
rect 14167 34886 14235 34942
rect 14291 34886 14359 34942
rect 14415 34886 14483 34942
rect 14539 34886 14607 34942
rect 14663 34886 14673 34942
rect 12861 34818 14673 34886
rect 12861 34762 12871 34818
rect 12927 34762 12995 34818
rect 13051 34762 13119 34818
rect 13175 34762 13243 34818
rect 13299 34762 13367 34818
rect 13423 34762 13491 34818
rect 13547 34762 13615 34818
rect 13671 34762 13739 34818
rect 13795 34762 13863 34818
rect 13919 34762 13987 34818
rect 14043 34762 14111 34818
rect 14167 34762 14235 34818
rect 14291 34762 14359 34818
rect 14415 34762 14483 34818
rect 14539 34762 14607 34818
rect 14663 34762 14673 34818
rect 12861 34694 14673 34762
rect 12861 34638 12871 34694
rect 12927 34638 12995 34694
rect 13051 34638 13119 34694
rect 13175 34638 13243 34694
rect 13299 34638 13367 34694
rect 13423 34638 13491 34694
rect 13547 34638 13615 34694
rect 13671 34638 13739 34694
rect 13795 34638 13863 34694
rect 13919 34638 13987 34694
rect 14043 34638 14111 34694
rect 14167 34638 14235 34694
rect 14291 34638 14359 34694
rect 14415 34638 14483 34694
rect 14539 34638 14607 34694
rect 14663 34638 14673 34694
rect 12861 34570 14673 34638
rect 12861 34514 12871 34570
rect 12927 34514 12995 34570
rect 13051 34514 13119 34570
rect 13175 34514 13243 34570
rect 13299 34514 13367 34570
rect 13423 34514 13491 34570
rect 13547 34514 13615 34570
rect 13671 34514 13739 34570
rect 13795 34514 13863 34570
rect 13919 34514 13987 34570
rect 14043 34514 14111 34570
rect 14167 34514 14235 34570
rect 14291 34514 14359 34570
rect 14415 34514 14483 34570
rect 14539 34514 14607 34570
rect 14663 34514 14673 34570
rect 12861 34446 14673 34514
rect 12861 34390 12871 34446
rect 12927 34390 12995 34446
rect 13051 34390 13119 34446
rect 13175 34390 13243 34446
rect 13299 34390 13367 34446
rect 13423 34390 13491 34446
rect 13547 34390 13615 34446
rect 13671 34390 13739 34446
rect 13795 34390 13863 34446
rect 13919 34390 13987 34446
rect 14043 34390 14111 34446
rect 14167 34390 14235 34446
rect 14291 34390 14359 34446
rect 14415 34390 14483 34446
rect 14539 34390 14607 34446
rect 14663 34390 14673 34446
rect 12861 34322 14673 34390
rect 12861 34266 12871 34322
rect 12927 34266 12995 34322
rect 13051 34266 13119 34322
rect 13175 34266 13243 34322
rect 13299 34266 13367 34322
rect 13423 34266 13491 34322
rect 13547 34266 13615 34322
rect 13671 34266 13739 34322
rect 13795 34266 13863 34322
rect 13919 34266 13987 34322
rect 14043 34266 14111 34322
rect 14167 34266 14235 34322
rect 14291 34266 14359 34322
rect 14415 34266 14483 34322
rect 14539 34266 14607 34322
rect 14663 34266 14673 34322
rect 12861 34198 14673 34266
rect 12861 34142 12871 34198
rect 12927 34142 12995 34198
rect 13051 34142 13119 34198
rect 13175 34142 13243 34198
rect 13299 34142 13367 34198
rect 13423 34142 13491 34198
rect 13547 34142 13615 34198
rect 13671 34142 13739 34198
rect 13795 34142 13863 34198
rect 13919 34142 13987 34198
rect 14043 34142 14111 34198
rect 14167 34142 14235 34198
rect 14291 34142 14359 34198
rect 14415 34142 14483 34198
rect 14539 34142 14607 34198
rect 14663 34142 14673 34198
rect 12861 34074 14673 34142
rect 12861 34018 12871 34074
rect 12927 34018 12995 34074
rect 13051 34018 13119 34074
rect 13175 34018 13243 34074
rect 13299 34018 13367 34074
rect 13423 34018 13491 34074
rect 13547 34018 13615 34074
rect 13671 34018 13739 34074
rect 13795 34018 13863 34074
rect 13919 34018 13987 34074
rect 14043 34018 14111 34074
rect 14167 34018 14235 34074
rect 14291 34018 14359 34074
rect 14415 34018 14483 34074
rect 14539 34018 14607 34074
rect 14663 34018 14673 34074
rect 12861 33950 14673 34018
rect 12861 33894 12871 33950
rect 12927 33894 12995 33950
rect 13051 33894 13119 33950
rect 13175 33894 13243 33950
rect 13299 33894 13367 33950
rect 13423 33894 13491 33950
rect 13547 33894 13615 33950
rect 13671 33894 13739 33950
rect 13795 33894 13863 33950
rect 13919 33894 13987 33950
rect 14043 33894 14111 33950
rect 14167 33894 14235 33950
rect 14291 33894 14359 33950
rect 14415 33894 14483 33950
rect 14539 33894 14607 33950
rect 14663 33894 14673 33950
rect 12861 33826 14673 33894
rect 12861 33770 12871 33826
rect 12927 33770 12995 33826
rect 13051 33770 13119 33826
rect 13175 33770 13243 33826
rect 13299 33770 13367 33826
rect 13423 33770 13491 33826
rect 13547 33770 13615 33826
rect 13671 33770 13739 33826
rect 13795 33770 13863 33826
rect 13919 33770 13987 33826
rect 14043 33770 14111 33826
rect 14167 33770 14235 33826
rect 14291 33770 14359 33826
rect 14415 33770 14483 33826
rect 14539 33770 14607 33826
rect 14663 33770 14673 33826
rect 12861 33702 14673 33770
rect 12861 33646 12871 33702
rect 12927 33646 12995 33702
rect 13051 33646 13119 33702
rect 13175 33646 13243 33702
rect 13299 33646 13367 33702
rect 13423 33646 13491 33702
rect 13547 33646 13615 33702
rect 13671 33646 13739 33702
rect 13795 33646 13863 33702
rect 13919 33646 13987 33702
rect 14043 33646 14111 33702
rect 14167 33646 14235 33702
rect 14291 33646 14359 33702
rect 14415 33646 14483 33702
rect 14539 33646 14607 33702
rect 14663 33646 14673 33702
rect 12861 33636 14673 33646
rect -11 33604 86 33614
rect 14892 33614 14902 36586
rect 14958 33614 14989 36586
rect 14892 33604 14989 33614
rect 2481 33354 2681 33364
rect 2481 33298 2491 33354
rect 2547 33298 2615 33354
rect 2671 33298 2681 33354
rect 2481 33230 2681 33298
rect 2481 33174 2491 33230
rect 2547 33174 2615 33230
rect 2671 33174 2681 33230
rect 2481 33106 2681 33174
rect 2481 33050 2491 33106
rect 2547 33050 2615 33106
rect 2671 33050 2681 33106
rect 2481 32982 2681 33050
rect 2481 32926 2491 32982
rect 2547 32926 2615 32982
rect 2671 32926 2681 32982
rect 2481 32858 2681 32926
rect 2481 32802 2491 32858
rect 2547 32802 2615 32858
rect 2671 32802 2681 32858
rect 2481 32734 2681 32802
rect 2481 32678 2491 32734
rect 2547 32678 2615 32734
rect 2671 32678 2681 32734
rect 2481 32610 2681 32678
rect 2481 32554 2491 32610
rect 2547 32554 2615 32610
rect 2671 32554 2681 32610
rect 2481 32486 2681 32554
rect 2481 32430 2491 32486
rect 2547 32430 2615 32486
rect 2671 32430 2681 32486
rect 2481 32362 2681 32430
rect 2481 32306 2491 32362
rect 2547 32306 2615 32362
rect 2671 32306 2681 32362
rect 2481 32238 2681 32306
rect 2481 32182 2491 32238
rect 2547 32182 2615 32238
rect 2671 32182 2681 32238
rect 2481 32114 2681 32182
rect 2481 32058 2491 32114
rect 2547 32058 2615 32114
rect 2671 32058 2681 32114
rect 2481 31990 2681 32058
rect 2481 31934 2491 31990
rect 2547 31934 2615 31990
rect 2671 31934 2681 31990
rect 2481 31866 2681 31934
rect 2481 31810 2491 31866
rect 2547 31810 2615 31866
rect 2671 31810 2681 31866
rect 2481 31742 2681 31810
rect 2481 31686 2491 31742
rect 2547 31686 2615 31742
rect 2671 31686 2681 31742
rect 2481 31618 2681 31686
rect 2481 31562 2491 31618
rect 2547 31562 2615 31618
rect 2671 31562 2681 31618
rect 2481 31494 2681 31562
rect 2481 31438 2491 31494
rect 2547 31438 2615 31494
rect 2671 31438 2681 31494
rect 2481 31370 2681 31438
rect 2481 31314 2491 31370
rect 2547 31314 2615 31370
rect 2671 31314 2681 31370
rect 2481 31246 2681 31314
rect 2481 31190 2491 31246
rect 2547 31190 2615 31246
rect 2671 31190 2681 31246
rect 2481 31122 2681 31190
rect 2481 31066 2491 31122
rect 2547 31066 2615 31122
rect 2671 31066 2681 31122
rect 2481 30998 2681 31066
rect 2481 30942 2491 30998
rect 2547 30942 2615 30998
rect 2671 30942 2681 30998
rect 2481 30874 2681 30942
rect 2481 30818 2491 30874
rect 2547 30818 2615 30874
rect 2671 30818 2681 30874
rect 2481 30750 2681 30818
rect 2481 30694 2491 30750
rect 2547 30694 2615 30750
rect 2671 30694 2681 30750
rect 2481 30626 2681 30694
rect 2481 30570 2491 30626
rect 2547 30570 2615 30626
rect 2671 30570 2681 30626
rect 2481 30502 2681 30570
rect 2481 30446 2491 30502
rect 2547 30446 2615 30502
rect 2671 30446 2681 30502
rect 2481 30436 2681 30446
rect 4851 33354 5051 33364
rect 4851 33298 4861 33354
rect 4917 33298 4985 33354
rect 5041 33298 5051 33354
rect 4851 33230 5051 33298
rect 4851 33174 4861 33230
rect 4917 33174 4985 33230
rect 5041 33174 5051 33230
rect 4851 33106 5051 33174
rect 4851 33050 4861 33106
rect 4917 33050 4985 33106
rect 5041 33050 5051 33106
rect 4851 32982 5051 33050
rect 4851 32926 4861 32982
rect 4917 32926 4985 32982
rect 5041 32926 5051 32982
rect 4851 32858 5051 32926
rect 4851 32802 4861 32858
rect 4917 32802 4985 32858
rect 5041 32802 5051 32858
rect 4851 32734 5051 32802
rect 4851 32678 4861 32734
rect 4917 32678 4985 32734
rect 5041 32678 5051 32734
rect 4851 32610 5051 32678
rect 4851 32554 4861 32610
rect 4917 32554 4985 32610
rect 5041 32554 5051 32610
rect 4851 32486 5051 32554
rect 4851 32430 4861 32486
rect 4917 32430 4985 32486
rect 5041 32430 5051 32486
rect 4851 32362 5051 32430
rect 4851 32306 4861 32362
rect 4917 32306 4985 32362
rect 5041 32306 5051 32362
rect 4851 32238 5051 32306
rect 4851 32182 4861 32238
rect 4917 32182 4985 32238
rect 5041 32182 5051 32238
rect 4851 32114 5051 32182
rect 4851 32058 4861 32114
rect 4917 32058 4985 32114
rect 5041 32058 5051 32114
rect 4851 31990 5051 32058
rect 4851 31934 4861 31990
rect 4917 31934 4985 31990
rect 5041 31934 5051 31990
rect 4851 31866 5051 31934
rect 4851 31810 4861 31866
rect 4917 31810 4985 31866
rect 5041 31810 5051 31866
rect 4851 31742 5051 31810
rect 4851 31686 4861 31742
rect 4917 31686 4985 31742
rect 5041 31686 5051 31742
rect 4851 31618 5051 31686
rect 4851 31562 4861 31618
rect 4917 31562 4985 31618
rect 5041 31562 5051 31618
rect 4851 31494 5051 31562
rect 4851 31438 4861 31494
rect 4917 31438 4985 31494
rect 5041 31438 5051 31494
rect 4851 31370 5051 31438
rect 4851 31314 4861 31370
rect 4917 31314 4985 31370
rect 5041 31314 5051 31370
rect 4851 31246 5051 31314
rect 4851 31190 4861 31246
rect 4917 31190 4985 31246
rect 5041 31190 5051 31246
rect 4851 31122 5051 31190
rect 4851 31066 4861 31122
rect 4917 31066 4985 31122
rect 5041 31066 5051 31122
rect 4851 30998 5051 31066
rect 4851 30942 4861 30998
rect 4917 30942 4985 30998
rect 5041 30942 5051 30998
rect 4851 30874 5051 30942
rect 4851 30818 4861 30874
rect 4917 30818 4985 30874
rect 5041 30818 5051 30874
rect 4851 30750 5051 30818
rect 4851 30694 4861 30750
rect 4917 30694 4985 30750
rect 5041 30694 5051 30750
rect 4851 30626 5051 30694
rect 4851 30570 4861 30626
rect 4917 30570 4985 30626
rect 5041 30570 5051 30626
rect 4851 30502 5051 30570
rect 4851 30446 4861 30502
rect 4917 30446 4985 30502
rect 5041 30446 5051 30502
rect 4851 30436 5051 30446
rect 7265 33354 7713 33364
rect 7265 33298 7275 33354
rect 7331 33298 7399 33354
rect 7455 33298 7523 33354
rect 7579 33298 7647 33354
rect 7703 33298 7713 33354
rect 7265 33230 7713 33298
rect 7265 33174 7275 33230
rect 7331 33174 7399 33230
rect 7455 33174 7523 33230
rect 7579 33174 7647 33230
rect 7703 33174 7713 33230
rect 7265 33106 7713 33174
rect 7265 33050 7275 33106
rect 7331 33050 7399 33106
rect 7455 33050 7523 33106
rect 7579 33050 7647 33106
rect 7703 33050 7713 33106
rect 7265 32982 7713 33050
rect 7265 32926 7275 32982
rect 7331 32926 7399 32982
rect 7455 32926 7523 32982
rect 7579 32926 7647 32982
rect 7703 32926 7713 32982
rect 7265 32858 7713 32926
rect 7265 32802 7275 32858
rect 7331 32802 7399 32858
rect 7455 32802 7523 32858
rect 7579 32802 7647 32858
rect 7703 32802 7713 32858
rect 7265 32734 7713 32802
rect 7265 32678 7275 32734
rect 7331 32678 7399 32734
rect 7455 32678 7523 32734
rect 7579 32678 7647 32734
rect 7703 32678 7713 32734
rect 7265 32610 7713 32678
rect 7265 32554 7275 32610
rect 7331 32554 7399 32610
rect 7455 32554 7523 32610
rect 7579 32554 7647 32610
rect 7703 32554 7713 32610
rect 7265 32486 7713 32554
rect 7265 32430 7275 32486
rect 7331 32430 7399 32486
rect 7455 32430 7523 32486
rect 7579 32430 7647 32486
rect 7703 32430 7713 32486
rect 7265 32362 7713 32430
rect 7265 32306 7275 32362
rect 7331 32306 7399 32362
rect 7455 32306 7523 32362
rect 7579 32306 7647 32362
rect 7703 32306 7713 32362
rect 7265 32238 7713 32306
rect 7265 32182 7275 32238
rect 7331 32182 7399 32238
rect 7455 32182 7523 32238
rect 7579 32182 7647 32238
rect 7703 32182 7713 32238
rect 7265 32114 7713 32182
rect 7265 32058 7275 32114
rect 7331 32058 7399 32114
rect 7455 32058 7523 32114
rect 7579 32058 7647 32114
rect 7703 32058 7713 32114
rect 7265 31990 7713 32058
rect 7265 31934 7275 31990
rect 7331 31934 7399 31990
rect 7455 31934 7523 31990
rect 7579 31934 7647 31990
rect 7703 31934 7713 31990
rect 7265 31866 7713 31934
rect 7265 31810 7275 31866
rect 7331 31810 7399 31866
rect 7455 31810 7523 31866
rect 7579 31810 7647 31866
rect 7703 31810 7713 31866
rect 7265 31742 7713 31810
rect 7265 31686 7275 31742
rect 7331 31686 7399 31742
rect 7455 31686 7523 31742
rect 7579 31686 7647 31742
rect 7703 31686 7713 31742
rect 7265 31618 7713 31686
rect 7265 31562 7275 31618
rect 7331 31562 7399 31618
rect 7455 31562 7523 31618
rect 7579 31562 7647 31618
rect 7703 31562 7713 31618
rect 7265 31494 7713 31562
rect 7265 31438 7275 31494
rect 7331 31438 7399 31494
rect 7455 31438 7523 31494
rect 7579 31438 7647 31494
rect 7703 31438 7713 31494
rect 7265 31370 7713 31438
rect 7265 31314 7275 31370
rect 7331 31314 7399 31370
rect 7455 31314 7523 31370
rect 7579 31314 7647 31370
rect 7703 31314 7713 31370
rect 7265 31246 7713 31314
rect 7265 31190 7275 31246
rect 7331 31190 7399 31246
rect 7455 31190 7523 31246
rect 7579 31190 7647 31246
rect 7703 31190 7713 31246
rect 7265 31122 7713 31190
rect 7265 31066 7275 31122
rect 7331 31066 7399 31122
rect 7455 31066 7523 31122
rect 7579 31066 7647 31122
rect 7703 31066 7713 31122
rect 7265 30998 7713 31066
rect 7265 30942 7275 30998
rect 7331 30942 7399 30998
rect 7455 30942 7523 30998
rect 7579 30942 7647 30998
rect 7703 30942 7713 30998
rect 7265 30874 7713 30942
rect 7265 30818 7275 30874
rect 7331 30818 7399 30874
rect 7455 30818 7523 30874
rect 7579 30818 7647 30874
rect 7703 30818 7713 30874
rect 7265 30750 7713 30818
rect 7265 30694 7275 30750
rect 7331 30694 7399 30750
rect 7455 30694 7523 30750
rect 7579 30694 7647 30750
rect 7703 30694 7713 30750
rect 7265 30626 7713 30694
rect 7265 30570 7275 30626
rect 7331 30570 7399 30626
rect 7455 30570 7523 30626
rect 7579 30570 7647 30626
rect 7703 30570 7713 30626
rect 7265 30502 7713 30570
rect 7265 30446 7275 30502
rect 7331 30446 7399 30502
rect 7455 30446 7523 30502
rect 7579 30446 7647 30502
rect 7703 30446 7713 30502
rect 7265 30436 7713 30446
rect 9927 33354 10127 33364
rect 9927 33298 9937 33354
rect 9993 33298 10061 33354
rect 10117 33298 10127 33354
rect 9927 33230 10127 33298
rect 9927 33174 9937 33230
rect 9993 33174 10061 33230
rect 10117 33174 10127 33230
rect 9927 33106 10127 33174
rect 9927 33050 9937 33106
rect 9993 33050 10061 33106
rect 10117 33050 10127 33106
rect 9927 32982 10127 33050
rect 9927 32926 9937 32982
rect 9993 32926 10061 32982
rect 10117 32926 10127 32982
rect 9927 32858 10127 32926
rect 9927 32802 9937 32858
rect 9993 32802 10061 32858
rect 10117 32802 10127 32858
rect 9927 32734 10127 32802
rect 9927 32678 9937 32734
rect 9993 32678 10061 32734
rect 10117 32678 10127 32734
rect 9927 32610 10127 32678
rect 9927 32554 9937 32610
rect 9993 32554 10061 32610
rect 10117 32554 10127 32610
rect 9927 32486 10127 32554
rect 9927 32430 9937 32486
rect 9993 32430 10061 32486
rect 10117 32430 10127 32486
rect 9927 32362 10127 32430
rect 9927 32306 9937 32362
rect 9993 32306 10061 32362
rect 10117 32306 10127 32362
rect 9927 32238 10127 32306
rect 9927 32182 9937 32238
rect 9993 32182 10061 32238
rect 10117 32182 10127 32238
rect 9927 32114 10127 32182
rect 9927 32058 9937 32114
rect 9993 32058 10061 32114
rect 10117 32058 10127 32114
rect 9927 31990 10127 32058
rect 9927 31934 9937 31990
rect 9993 31934 10061 31990
rect 10117 31934 10127 31990
rect 9927 31866 10127 31934
rect 9927 31810 9937 31866
rect 9993 31810 10061 31866
rect 10117 31810 10127 31866
rect 9927 31742 10127 31810
rect 9927 31686 9937 31742
rect 9993 31686 10061 31742
rect 10117 31686 10127 31742
rect 9927 31618 10127 31686
rect 9927 31562 9937 31618
rect 9993 31562 10061 31618
rect 10117 31562 10127 31618
rect 9927 31494 10127 31562
rect 9927 31438 9937 31494
rect 9993 31438 10061 31494
rect 10117 31438 10127 31494
rect 9927 31370 10127 31438
rect 9927 31314 9937 31370
rect 9993 31314 10061 31370
rect 10117 31314 10127 31370
rect 9927 31246 10127 31314
rect 9927 31190 9937 31246
rect 9993 31190 10061 31246
rect 10117 31190 10127 31246
rect 9927 31122 10127 31190
rect 9927 31066 9937 31122
rect 9993 31066 10061 31122
rect 10117 31066 10127 31122
rect 9927 30998 10127 31066
rect 9927 30942 9937 30998
rect 9993 30942 10061 30998
rect 10117 30942 10127 30998
rect 9927 30874 10127 30942
rect 9927 30818 9937 30874
rect 9993 30818 10061 30874
rect 10117 30818 10127 30874
rect 9927 30750 10127 30818
rect 9927 30694 9937 30750
rect 9993 30694 10061 30750
rect 10117 30694 10127 30750
rect 9927 30626 10127 30694
rect 9927 30570 9937 30626
rect 9993 30570 10061 30626
rect 10117 30570 10127 30626
rect 9927 30502 10127 30570
rect 9927 30446 9937 30502
rect 9993 30446 10061 30502
rect 10117 30446 10127 30502
rect 9927 30436 10127 30446
rect 12297 33354 12497 33364
rect 12297 33298 12307 33354
rect 12363 33298 12431 33354
rect 12487 33298 12497 33354
rect 12297 33230 12497 33298
rect 12297 33174 12307 33230
rect 12363 33174 12431 33230
rect 12487 33174 12497 33230
rect 12297 33106 12497 33174
rect 12297 33050 12307 33106
rect 12363 33050 12431 33106
rect 12487 33050 12497 33106
rect 12297 32982 12497 33050
rect 12297 32926 12307 32982
rect 12363 32926 12431 32982
rect 12487 32926 12497 32982
rect 12297 32858 12497 32926
rect 12297 32802 12307 32858
rect 12363 32802 12431 32858
rect 12487 32802 12497 32858
rect 12297 32734 12497 32802
rect 12297 32678 12307 32734
rect 12363 32678 12431 32734
rect 12487 32678 12497 32734
rect 12297 32610 12497 32678
rect 12297 32554 12307 32610
rect 12363 32554 12431 32610
rect 12487 32554 12497 32610
rect 12297 32486 12497 32554
rect 12297 32430 12307 32486
rect 12363 32430 12431 32486
rect 12487 32430 12497 32486
rect 12297 32362 12497 32430
rect 12297 32306 12307 32362
rect 12363 32306 12431 32362
rect 12487 32306 12497 32362
rect 12297 32238 12497 32306
rect 12297 32182 12307 32238
rect 12363 32182 12431 32238
rect 12487 32182 12497 32238
rect 12297 32114 12497 32182
rect 12297 32058 12307 32114
rect 12363 32058 12431 32114
rect 12487 32058 12497 32114
rect 12297 31990 12497 32058
rect 12297 31934 12307 31990
rect 12363 31934 12431 31990
rect 12487 31934 12497 31990
rect 12297 31866 12497 31934
rect 12297 31810 12307 31866
rect 12363 31810 12431 31866
rect 12487 31810 12497 31866
rect 12297 31742 12497 31810
rect 12297 31686 12307 31742
rect 12363 31686 12431 31742
rect 12487 31686 12497 31742
rect 12297 31618 12497 31686
rect 12297 31562 12307 31618
rect 12363 31562 12431 31618
rect 12487 31562 12497 31618
rect 12297 31494 12497 31562
rect 12297 31438 12307 31494
rect 12363 31438 12431 31494
rect 12487 31438 12497 31494
rect 12297 31370 12497 31438
rect 12297 31314 12307 31370
rect 12363 31314 12431 31370
rect 12487 31314 12497 31370
rect 12297 31246 12497 31314
rect 12297 31190 12307 31246
rect 12363 31190 12431 31246
rect 12487 31190 12497 31246
rect 12297 31122 12497 31190
rect 12297 31066 12307 31122
rect 12363 31066 12431 31122
rect 12487 31066 12497 31122
rect 12297 30998 12497 31066
rect 12297 30942 12307 30998
rect 12363 30942 12431 30998
rect 12487 30942 12497 30998
rect 12297 30874 12497 30942
rect 12297 30818 12307 30874
rect 12363 30818 12431 30874
rect 12487 30818 12497 30874
rect 12297 30750 12497 30818
rect 12297 30694 12307 30750
rect 12363 30694 12431 30750
rect 12487 30694 12497 30750
rect 12297 30626 12497 30694
rect 12297 30570 12307 30626
rect 12363 30570 12431 30626
rect 12487 30570 12497 30626
rect 12297 30502 12497 30570
rect 12297 30446 12307 30502
rect 12363 30446 12431 30502
rect 12487 30446 12497 30502
rect 12297 30436 12497 30446
rect 2481 30148 2681 30158
rect 2481 30092 2491 30148
rect 2547 30092 2615 30148
rect 2671 30092 2681 30148
rect 2481 30024 2681 30092
rect 2481 29968 2491 30024
rect 2547 29968 2615 30024
rect 2671 29968 2681 30024
rect 2481 29900 2681 29968
rect 2481 29844 2491 29900
rect 2547 29844 2615 29900
rect 2671 29844 2681 29900
rect 2481 29776 2681 29844
rect 2481 29720 2491 29776
rect 2547 29720 2615 29776
rect 2671 29720 2681 29776
rect 2481 29652 2681 29720
rect 2481 29596 2491 29652
rect 2547 29596 2615 29652
rect 2671 29596 2681 29652
rect 2481 29528 2681 29596
rect 2481 29472 2491 29528
rect 2547 29472 2615 29528
rect 2671 29472 2681 29528
rect 2481 29404 2681 29472
rect 2481 29348 2491 29404
rect 2547 29348 2615 29404
rect 2671 29348 2681 29404
rect 2481 29280 2681 29348
rect 2481 29224 2491 29280
rect 2547 29224 2615 29280
rect 2671 29224 2681 29280
rect 2481 29156 2681 29224
rect 2481 29100 2491 29156
rect 2547 29100 2615 29156
rect 2671 29100 2681 29156
rect 2481 29032 2681 29100
rect 2481 28976 2491 29032
rect 2547 28976 2615 29032
rect 2671 28976 2681 29032
rect 2481 28908 2681 28976
rect 2481 28852 2491 28908
rect 2547 28852 2615 28908
rect 2671 28852 2681 28908
rect 2481 28842 2681 28852
rect 4851 30148 5051 30158
rect 4851 30092 4861 30148
rect 4917 30092 4985 30148
rect 5041 30092 5051 30148
rect 4851 30024 5051 30092
rect 4851 29968 4861 30024
rect 4917 29968 4985 30024
rect 5041 29968 5051 30024
rect 4851 29900 5051 29968
rect 4851 29844 4861 29900
rect 4917 29844 4985 29900
rect 5041 29844 5051 29900
rect 4851 29776 5051 29844
rect 4851 29720 4861 29776
rect 4917 29720 4985 29776
rect 5041 29720 5051 29776
rect 4851 29652 5051 29720
rect 4851 29596 4861 29652
rect 4917 29596 4985 29652
rect 5041 29596 5051 29652
rect 4851 29528 5051 29596
rect 4851 29472 4861 29528
rect 4917 29472 4985 29528
rect 5041 29472 5051 29528
rect 4851 29404 5051 29472
rect 4851 29348 4861 29404
rect 4917 29348 4985 29404
rect 5041 29348 5051 29404
rect 4851 29280 5051 29348
rect 4851 29224 4861 29280
rect 4917 29224 4985 29280
rect 5041 29224 5051 29280
rect 4851 29156 5051 29224
rect 4851 29100 4861 29156
rect 4917 29100 4985 29156
rect 5041 29100 5051 29156
rect 4851 29032 5051 29100
rect 4851 28976 4861 29032
rect 4917 28976 4985 29032
rect 5041 28976 5051 29032
rect 4851 28908 5051 28976
rect 4851 28852 4861 28908
rect 4917 28852 4985 28908
rect 5041 28852 5051 28908
rect 4851 28842 5051 28852
rect 7265 30148 7713 30158
rect 7265 30092 7275 30148
rect 7331 30092 7399 30148
rect 7455 30092 7523 30148
rect 7579 30092 7647 30148
rect 7703 30092 7713 30148
rect 7265 30024 7713 30092
rect 7265 29968 7275 30024
rect 7331 29968 7399 30024
rect 7455 29968 7523 30024
rect 7579 29968 7647 30024
rect 7703 29968 7713 30024
rect 7265 29900 7713 29968
rect 7265 29844 7275 29900
rect 7331 29844 7399 29900
rect 7455 29844 7523 29900
rect 7579 29844 7647 29900
rect 7703 29844 7713 29900
rect 7265 29776 7713 29844
rect 7265 29720 7275 29776
rect 7331 29720 7399 29776
rect 7455 29720 7523 29776
rect 7579 29720 7647 29776
rect 7703 29720 7713 29776
rect 7265 29652 7713 29720
rect 7265 29596 7275 29652
rect 7331 29596 7399 29652
rect 7455 29596 7523 29652
rect 7579 29596 7647 29652
rect 7703 29596 7713 29652
rect 7265 29528 7713 29596
rect 7265 29472 7275 29528
rect 7331 29472 7399 29528
rect 7455 29472 7523 29528
rect 7579 29472 7647 29528
rect 7703 29472 7713 29528
rect 7265 29404 7713 29472
rect 7265 29348 7275 29404
rect 7331 29348 7399 29404
rect 7455 29348 7523 29404
rect 7579 29348 7647 29404
rect 7703 29348 7713 29404
rect 7265 29280 7713 29348
rect 7265 29224 7275 29280
rect 7331 29224 7399 29280
rect 7455 29224 7523 29280
rect 7579 29224 7647 29280
rect 7703 29224 7713 29280
rect 7265 29156 7713 29224
rect 7265 29100 7275 29156
rect 7331 29100 7399 29156
rect 7455 29100 7523 29156
rect 7579 29100 7647 29156
rect 7703 29100 7713 29156
rect 7265 29032 7713 29100
rect 7265 28976 7275 29032
rect 7331 28976 7399 29032
rect 7455 28976 7523 29032
rect 7579 28976 7647 29032
rect 7703 28976 7713 29032
rect 7265 28908 7713 28976
rect 7265 28852 7275 28908
rect 7331 28852 7399 28908
rect 7455 28852 7523 28908
rect 7579 28852 7647 28908
rect 7703 28852 7713 28908
rect 7265 28842 7713 28852
rect 9927 30148 10127 30158
rect 9927 30092 9937 30148
rect 9993 30092 10061 30148
rect 10117 30092 10127 30148
rect 9927 30024 10127 30092
rect 9927 29968 9937 30024
rect 9993 29968 10061 30024
rect 10117 29968 10127 30024
rect 9927 29900 10127 29968
rect 9927 29844 9937 29900
rect 9993 29844 10061 29900
rect 10117 29844 10127 29900
rect 9927 29776 10127 29844
rect 9927 29720 9937 29776
rect 9993 29720 10061 29776
rect 10117 29720 10127 29776
rect 9927 29652 10127 29720
rect 9927 29596 9937 29652
rect 9993 29596 10061 29652
rect 10117 29596 10127 29652
rect 9927 29528 10127 29596
rect 9927 29472 9937 29528
rect 9993 29472 10061 29528
rect 10117 29472 10127 29528
rect 9927 29404 10127 29472
rect 9927 29348 9937 29404
rect 9993 29348 10061 29404
rect 10117 29348 10127 29404
rect 9927 29280 10127 29348
rect 9927 29224 9937 29280
rect 9993 29224 10061 29280
rect 10117 29224 10127 29280
rect 9927 29156 10127 29224
rect 9927 29100 9937 29156
rect 9993 29100 10061 29156
rect 10117 29100 10127 29156
rect 9927 29032 10127 29100
rect 9927 28976 9937 29032
rect 9993 28976 10061 29032
rect 10117 28976 10127 29032
rect 9927 28908 10127 28976
rect 9927 28852 9937 28908
rect 9993 28852 10061 28908
rect 10117 28852 10127 28908
rect 9927 28842 10127 28852
rect 12297 30148 12497 30158
rect 12297 30092 12307 30148
rect 12363 30092 12431 30148
rect 12487 30092 12497 30148
rect 12297 30024 12497 30092
rect 12297 29968 12307 30024
rect 12363 29968 12431 30024
rect 12487 29968 12497 30024
rect 12297 29900 12497 29968
rect 12297 29844 12307 29900
rect 12363 29844 12431 29900
rect 12487 29844 12497 29900
rect 12297 29776 12497 29844
rect 12297 29720 12307 29776
rect 12363 29720 12431 29776
rect 12487 29720 12497 29776
rect 12297 29652 12497 29720
rect 12297 29596 12307 29652
rect 12363 29596 12431 29652
rect 12487 29596 12497 29652
rect 12297 29528 12497 29596
rect 12297 29472 12307 29528
rect 12363 29472 12431 29528
rect 12487 29472 12497 29528
rect 12297 29404 12497 29472
rect 12297 29348 12307 29404
rect 12363 29348 12431 29404
rect 12487 29348 12497 29404
rect 12297 29280 12497 29348
rect 12297 29224 12307 29280
rect 12363 29224 12431 29280
rect 12487 29224 12497 29280
rect 12297 29156 12497 29224
rect 12297 29100 12307 29156
rect 12363 29100 12431 29156
rect 12487 29100 12497 29156
rect 12297 29032 12497 29100
rect 12297 28976 12307 29032
rect 12363 28976 12431 29032
rect 12487 28976 12497 29032
rect 12297 28908 12497 28976
rect 12297 28852 12307 28908
rect 12363 28852 12431 28908
rect 12487 28852 12497 28908
rect 12297 28842 12497 28852
rect -11 28576 86 28586
rect -11 27224 20 28576
rect 76 27224 86 28576
rect 14892 28576 14989 28586
rect 305 28548 2117 28558
rect 305 28492 315 28548
rect 371 28492 439 28548
rect 495 28492 563 28548
rect 619 28492 687 28548
rect 743 28492 811 28548
rect 867 28492 935 28548
rect 991 28492 1059 28548
rect 1115 28492 1183 28548
rect 1239 28492 1307 28548
rect 1363 28492 1431 28548
rect 1487 28492 1555 28548
rect 1611 28492 1679 28548
rect 1735 28492 1803 28548
rect 1859 28492 1927 28548
rect 1983 28492 2051 28548
rect 2107 28492 2117 28548
rect 305 28424 2117 28492
rect 305 28368 315 28424
rect 371 28368 439 28424
rect 495 28368 563 28424
rect 619 28368 687 28424
rect 743 28368 811 28424
rect 867 28368 935 28424
rect 991 28368 1059 28424
rect 1115 28368 1183 28424
rect 1239 28368 1307 28424
rect 1363 28368 1431 28424
rect 1487 28368 1555 28424
rect 1611 28368 1679 28424
rect 1735 28368 1803 28424
rect 1859 28368 1927 28424
rect 1983 28368 2051 28424
rect 2107 28368 2117 28424
rect 305 28300 2117 28368
rect 305 28244 315 28300
rect 371 28244 439 28300
rect 495 28244 563 28300
rect 619 28244 687 28300
rect 743 28244 811 28300
rect 867 28244 935 28300
rect 991 28244 1059 28300
rect 1115 28244 1183 28300
rect 1239 28244 1307 28300
rect 1363 28244 1431 28300
rect 1487 28244 1555 28300
rect 1611 28244 1679 28300
rect 1735 28244 1803 28300
rect 1859 28244 1927 28300
rect 1983 28244 2051 28300
rect 2107 28244 2117 28300
rect 305 28176 2117 28244
rect 305 28120 315 28176
rect 371 28120 439 28176
rect 495 28120 563 28176
rect 619 28120 687 28176
rect 743 28120 811 28176
rect 867 28120 935 28176
rect 991 28120 1059 28176
rect 1115 28120 1183 28176
rect 1239 28120 1307 28176
rect 1363 28120 1431 28176
rect 1487 28120 1555 28176
rect 1611 28120 1679 28176
rect 1735 28120 1803 28176
rect 1859 28120 1927 28176
rect 1983 28120 2051 28176
rect 2107 28120 2117 28176
rect 305 28052 2117 28120
rect 305 27996 315 28052
rect 371 27996 439 28052
rect 495 27996 563 28052
rect 619 27996 687 28052
rect 743 27996 811 28052
rect 867 27996 935 28052
rect 991 27996 1059 28052
rect 1115 27996 1183 28052
rect 1239 27996 1307 28052
rect 1363 27996 1431 28052
rect 1487 27996 1555 28052
rect 1611 27996 1679 28052
rect 1735 27996 1803 28052
rect 1859 27996 1927 28052
rect 1983 27996 2051 28052
rect 2107 27996 2117 28052
rect 305 27928 2117 27996
rect 305 27872 315 27928
rect 371 27872 439 27928
rect 495 27872 563 27928
rect 619 27872 687 27928
rect 743 27872 811 27928
rect 867 27872 935 27928
rect 991 27872 1059 27928
rect 1115 27872 1183 27928
rect 1239 27872 1307 27928
rect 1363 27872 1431 27928
rect 1487 27872 1555 27928
rect 1611 27872 1679 27928
rect 1735 27872 1803 27928
rect 1859 27872 1927 27928
rect 1983 27872 2051 27928
rect 2107 27872 2117 27928
rect 305 27804 2117 27872
rect 305 27748 315 27804
rect 371 27748 439 27804
rect 495 27748 563 27804
rect 619 27748 687 27804
rect 743 27748 811 27804
rect 867 27748 935 27804
rect 991 27748 1059 27804
rect 1115 27748 1183 27804
rect 1239 27748 1307 27804
rect 1363 27748 1431 27804
rect 1487 27748 1555 27804
rect 1611 27748 1679 27804
rect 1735 27748 1803 27804
rect 1859 27748 1927 27804
rect 1983 27748 2051 27804
rect 2107 27748 2117 27804
rect 305 27680 2117 27748
rect 305 27624 315 27680
rect 371 27624 439 27680
rect 495 27624 563 27680
rect 619 27624 687 27680
rect 743 27624 811 27680
rect 867 27624 935 27680
rect 991 27624 1059 27680
rect 1115 27624 1183 27680
rect 1239 27624 1307 27680
rect 1363 27624 1431 27680
rect 1487 27624 1555 27680
rect 1611 27624 1679 27680
rect 1735 27624 1803 27680
rect 1859 27624 1927 27680
rect 1983 27624 2051 27680
rect 2107 27624 2117 27680
rect 305 27556 2117 27624
rect 305 27500 315 27556
rect 371 27500 439 27556
rect 495 27500 563 27556
rect 619 27500 687 27556
rect 743 27500 811 27556
rect 867 27500 935 27556
rect 991 27500 1059 27556
rect 1115 27500 1183 27556
rect 1239 27500 1307 27556
rect 1363 27500 1431 27556
rect 1487 27500 1555 27556
rect 1611 27500 1679 27556
rect 1735 27500 1803 27556
rect 1859 27500 1927 27556
rect 1983 27500 2051 27556
rect 2107 27500 2117 27556
rect 305 27432 2117 27500
rect 305 27376 315 27432
rect 371 27376 439 27432
rect 495 27376 563 27432
rect 619 27376 687 27432
rect 743 27376 811 27432
rect 867 27376 935 27432
rect 991 27376 1059 27432
rect 1115 27376 1183 27432
rect 1239 27376 1307 27432
rect 1363 27376 1431 27432
rect 1487 27376 1555 27432
rect 1611 27376 1679 27432
rect 1735 27376 1803 27432
rect 1859 27376 1927 27432
rect 1983 27376 2051 27432
rect 2107 27376 2117 27432
rect 305 27308 2117 27376
rect 305 27252 315 27308
rect 371 27252 439 27308
rect 495 27252 563 27308
rect 619 27252 687 27308
rect 743 27252 811 27308
rect 867 27252 935 27308
rect 991 27252 1059 27308
rect 1115 27252 1183 27308
rect 1239 27252 1307 27308
rect 1363 27252 1431 27308
rect 1487 27252 1555 27308
rect 1611 27252 1679 27308
rect 1735 27252 1803 27308
rect 1859 27252 1927 27308
rect 1983 27252 2051 27308
rect 2107 27252 2117 27308
rect 305 27242 2117 27252
rect 2798 28548 4734 28558
rect 2798 28492 2808 28548
rect 2864 28492 2932 28548
rect 2988 28492 3056 28548
rect 3112 28492 3180 28548
rect 3236 28492 3304 28548
rect 3360 28492 3428 28548
rect 3484 28492 3552 28548
rect 3608 28492 3676 28548
rect 3732 28492 3800 28548
rect 3856 28492 3924 28548
rect 3980 28492 4048 28548
rect 4104 28492 4172 28548
rect 4228 28492 4296 28548
rect 4352 28492 4420 28548
rect 4476 28492 4544 28548
rect 4600 28492 4668 28548
rect 4724 28492 4734 28548
rect 2798 28424 4734 28492
rect 2798 28368 2808 28424
rect 2864 28368 2932 28424
rect 2988 28368 3056 28424
rect 3112 28368 3180 28424
rect 3236 28368 3304 28424
rect 3360 28368 3428 28424
rect 3484 28368 3552 28424
rect 3608 28368 3676 28424
rect 3732 28368 3800 28424
rect 3856 28368 3924 28424
rect 3980 28368 4048 28424
rect 4104 28368 4172 28424
rect 4228 28368 4296 28424
rect 4352 28368 4420 28424
rect 4476 28368 4544 28424
rect 4600 28368 4668 28424
rect 4724 28368 4734 28424
rect 2798 28300 4734 28368
rect 2798 28244 2808 28300
rect 2864 28244 2932 28300
rect 2988 28244 3056 28300
rect 3112 28244 3180 28300
rect 3236 28244 3304 28300
rect 3360 28244 3428 28300
rect 3484 28244 3552 28300
rect 3608 28244 3676 28300
rect 3732 28244 3800 28300
rect 3856 28244 3924 28300
rect 3980 28244 4048 28300
rect 4104 28244 4172 28300
rect 4228 28244 4296 28300
rect 4352 28244 4420 28300
rect 4476 28244 4544 28300
rect 4600 28244 4668 28300
rect 4724 28244 4734 28300
rect 2798 28176 4734 28244
rect 2798 28120 2808 28176
rect 2864 28120 2932 28176
rect 2988 28120 3056 28176
rect 3112 28120 3180 28176
rect 3236 28120 3304 28176
rect 3360 28120 3428 28176
rect 3484 28120 3552 28176
rect 3608 28120 3676 28176
rect 3732 28120 3800 28176
rect 3856 28120 3924 28176
rect 3980 28120 4048 28176
rect 4104 28120 4172 28176
rect 4228 28120 4296 28176
rect 4352 28120 4420 28176
rect 4476 28120 4544 28176
rect 4600 28120 4668 28176
rect 4724 28120 4734 28176
rect 2798 28052 4734 28120
rect 2798 27996 2808 28052
rect 2864 27996 2932 28052
rect 2988 27996 3056 28052
rect 3112 27996 3180 28052
rect 3236 27996 3304 28052
rect 3360 27996 3428 28052
rect 3484 27996 3552 28052
rect 3608 27996 3676 28052
rect 3732 27996 3800 28052
rect 3856 27996 3924 28052
rect 3980 27996 4048 28052
rect 4104 27996 4172 28052
rect 4228 27996 4296 28052
rect 4352 27996 4420 28052
rect 4476 27996 4544 28052
rect 4600 27996 4668 28052
rect 4724 27996 4734 28052
rect 2798 27928 4734 27996
rect 2798 27872 2808 27928
rect 2864 27872 2932 27928
rect 2988 27872 3056 27928
rect 3112 27872 3180 27928
rect 3236 27872 3304 27928
rect 3360 27872 3428 27928
rect 3484 27872 3552 27928
rect 3608 27872 3676 27928
rect 3732 27872 3800 27928
rect 3856 27872 3924 27928
rect 3980 27872 4048 27928
rect 4104 27872 4172 27928
rect 4228 27872 4296 27928
rect 4352 27872 4420 27928
rect 4476 27872 4544 27928
rect 4600 27872 4668 27928
rect 4724 27872 4734 27928
rect 2798 27804 4734 27872
rect 2798 27748 2808 27804
rect 2864 27748 2932 27804
rect 2988 27748 3056 27804
rect 3112 27748 3180 27804
rect 3236 27748 3304 27804
rect 3360 27748 3428 27804
rect 3484 27748 3552 27804
rect 3608 27748 3676 27804
rect 3732 27748 3800 27804
rect 3856 27748 3924 27804
rect 3980 27748 4048 27804
rect 4104 27748 4172 27804
rect 4228 27748 4296 27804
rect 4352 27748 4420 27804
rect 4476 27748 4544 27804
rect 4600 27748 4668 27804
rect 4724 27748 4734 27804
rect 2798 27680 4734 27748
rect 2798 27624 2808 27680
rect 2864 27624 2932 27680
rect 2988 27624 3056 27680
rect 3112 27624 3180 27680
rect 3236 27624 3304 27680
rect 3360 27624 3428 27680
rect 3484 27624 3552 27680
rect 3608 27624 3676 27680
rect 3732 27624 3800 27680
rect 3856 27624 3924 27680
rect 3980 27624 4048 27680
rect 4104 27624 4172 27680
rect 4228 27624 4296 27680
rect 4352 27624 4420 27680
rect 4476 27624 4544 27680
rect 4600 27624 4668 27680
rect 4724 27624 4734 27680
rect 2798 27556 4734 27624
rect 2798 27500 2808 27556
rect 2864 27500 2932 27556
rect 2988 27500 3056 27556
rect 3112 27500 3180 27556
rect 3236 27500 3304 27556
rect 3360 27500 3428 27556
rect 3484 27500 3552 27556
rect 3608 27500 3676 27556
rect 3732 27500 3800 27556
rect 3856 27500 3924 27556
rect 3980 27500 4048 27556
rect 4104 27500 4172 27556
rect 4228 27500 4296 27556
rect 4352 27500 4420 27556
rect 4476 27500 4544 27556
rect 4600 27500 4668 27556
rect 4724 27500 4734 27556
rect 2798 27432 4734 27500
rect 2798 27376 2808 27432
rect 2864 27376 2932 27432
rect 2988 27376 3056 27432
rect 3112 27376 3180 27432
rect 3236 27376 3304 27432
rect 3360 27376 3428 27432
rect 3484 27376 3552 27432
rect 3608 27376 3676 27432
rect 3732 27376 3800 27432
rect 3856 27376 3924 27432
rect 3980 27376 4048 27432
rect 4104 27376 4172 27432
rect 4228 27376 4296 27432
rect 4352 27376 4420 27432
rect 4476 27376 4544 27432
rect 4600 27376 4668 27432
rect 4724 27376 4734 27432
rect 2798 27308 4734 27376
rect 2798 27252 2808 27308
rect 2864 27252 2932 27308
rect 2988 27252 3056 27308
rect 3112 27252 3180 27308
rect 3236 27252 3304 27308
rect 3360 27252 3428 27308
rect 3484 27252 3552 27308
rect 3608 27252 3676 27308
rect 3732 27252 3800 27308
rect 3856 27252 3924 27308
rect 3980 27252 4048 27308
rect 4104 27252 4172 27308
rect 4228 27252 4296 27308
rect 4352 27252 4420 27308
rect 4476 27252 4544 27308
rect 4600 27252 4668 27308
rect 4724 27252 4734 27308
rect 2798 27242 4734 27252
rect 5168 28548 7104 28558
rect 5168 28492 5178 28548
rect 5234 28492 5302 28548
rect 5358 28492 5426 28548
rect 5482 28492 5550 28548
rect 5606 28492 5674 28548
rect 5730 28492 5798 28548
rect 5854 28492 5922 28548
rect 5978 28492 6046 28548
rect 6102 28492 6170 28548
rect 6226 28492 6294 28548
rect 6350 28492 6418 28548
rect 6474 28492 6542 28548
rect 6598 28492 6666 28548
rect 6722 28492 6790 28548
rect 6846 28492 6914 28548
rect 6970 28492 7038 28548
rect 7094 28492 7104 28548
rect 5168 28424 7104 28492
rect 5168 28368 5178 28424
rect 5234 28368 5302 28424
rect 5358 28368 5426 28424
rect 5482 28368 5550 28424
rect 5606 28368 5674 28424
rect 5730 28368 5798 28424
rect 5854 28368 5922 28424
rect 5978 28368 6046 28424
rect 6102 28368 6170 28424
rect 6226 28368 6294 28424
rect 6350 28368 6418 28424
rect 6474 28368 6542 28424
rect 6598 28368 6666 28424
rect 6722 28368 6790 28424
rect 6846 28368 6914 28424
rect 6970 28368 7038 28424
rect 7094 28368 7104 28424
rect 5168 28300 7104 28368
rect 5168 28244 5178 28300
rect 5234 28244 5302 28300
rect 5358 28244 5426 28300
rect 5482 28244 5550 28300
rect 5606 28244 5674 28300
rect 5730 28244 5798 28300
rect 5854 28244 5922 28300
rect 5978 28244 6046 28300
rect 6102 28244 6170 28300
rect 6226 28244 6294 28300
rect 6350 28244 6418 28300
rect 6474 28244 6542 28300
rect 6598 28244 6666 28300
rect 6722 28244 6790 28300
rect 6846 28244 6914 28300
rect 6970 28244 7038 28300
rect 7094 28244 7104 28300
rect 5168 28176 7104 28244
rect 5168 28120 5178 28176
rect 5234 28120 5302 28176
rect 5358 28120 5426 28176
rect 5482 28120 5550 28176
rect 5606 28120 5674 28176
rect 5730 28120 5798 28176
rect 5854 28120 5922 28176
rect 5978 28120 6046 28176
rect 6102 28120 6170 28176
rect 6226 28120 6294 28176
rect 6350 28120 6418 28176
rect 6474 28120 6542 28176
rect 6598 28120 6666 28176
rect 6722 28120 6790 28176
rect 6846 28120 6914 28176
rect 6970 28120 7038 28176
rect 7094 28120 7104 28176
rect 5168 28052 7104 28120
rect 5168 27996 5178 28052
rect 5234 27996 5302 28052
rect 5358 27996 5426 28052
rect 5482 27996 5550 28052
rect 5606 27996 5674 28052
rect 5730 27996 5798 28052
rect 5854 27996 5922 28052
rect 5978 27996 6046 28052
rect 6102 27996 6170 28052
rect 6226 27996 6294 28052
rect 6350 27996 6418 28052
rect 6474 27996 6542 28052
rect 6598 27996 6666 28052
rect 6722 27996 6790 28052
rect 6846 27996 6914 28052
rect 6970 27996 7038 28052
rect 7094 27996 7104 28052
rect 5168 27928 7104 27996
rect 5168 27872 5178 27928
rect 5234 27872 5302 27928
rect 5358 27872 5426 27928
rect 5482 27872 5550 27928
rect 5606 27872 5674 27928
rect 5730 27872 5798 27928
rect 5854 27872 5922 27928
rect 5978 27872 6046 27928
rect 6102 27872 6170 27928
rect 6226 27872 6294 27928
rect 6350 27872 6418 27928
rect 6474 27872 6542 27928
rect 6598 27872 6666 27928
rect 6722 27872 6790 27928
rect 6846 27872 6914 27928
rect 6970 27872 7038 27928
rect 7094 27872 7104 27928
rect 5168 27804 7104 27872
rect 5168 27748 5178 27804
rect 5234 27748 5302 27804
rect 5358 27748 5426 27804
rect 5482 27748 5550 27804
rect 5606 27748 5674 27804
rect 5730 27748 5798 27804
rect 5854 27748 5922 27804
rect 5978 27748 6046 27804
rect 6102 27748 6170 27804
rect 6226 27748 6294 27804
rect 6350 27748 6418 27804
rect 6474 27748 6542 27804
rect 6598 27748 6666 27804
rect 6722 27748 6790 27804
rect 6846 27748 6914 27804
rect 6970 27748 7038 27804
rect 7094 27748 7104 27804
rect 5168 27680 7104 27748
rect 5168 27624 5178 27680
rect 5234 27624 5302 27680
rect 5358 27624 5426 27680
rect 5482 27624 5550 27680
rect 5606 27624 5674 27680
rect 5730 27624 5798 27680
rect 5854 27624 5922 27680
rect 5978 27624 6046 27680
rect 6102 27624 6170 27680
rect 6226 27624 6294 27680
rect 6350 27624 6418 27680
rect 6474 27624 6542 27680
rect 6598 27624 6666 27680
rect 6722 27624 6790 27680
rect 6846 27624 6914 27680
rect 6970 27624 7038 27680
rect 7094 27624 7104 27680
rect 5168 27556 7104 27624
rect 5168 27500 5178 27556
rect 5234 27500 5302 27556
rect 5358 27500 5426 27556
rect 5482 27500 5550 27556
rect 5606 27500 5674 27556
rect 5730 27500 5798 27556
rect 5854 27500 5922 27556
rect 5978 27500 6046 27556
rect 6102 27500 6170 27556
rect 6226 27500 6294 27556
rect 6350 27500 6418 27556
rect 6474 27500 6542 27556
rect 6598 27500 6666 27556
rect 6722 27500 6790 27556
rect 6846 27500 6914 27556
rect 6970 27500 7038 27556
rect 7094 27500 7104 27556
rect 5168 27432 7104 27500
rect 5168 27376 5178 27432
rect 5234 27376 5302 27432
rect 5358 27376 5426 27432
rect 5482 27376 5550 27432
rect 5606 27376 5674 27432
rect 5730 27376 5798 27432
rect 5854 27376 5922 27432
rect 5978 27376 6046 27432
rect 6102 27376 6170 27432
rect 6226 27376 6294 27432
rect 6350 27376 6418 27432
rect 6474 27376 6542 27432
rect 6598 27376 6666 27432
rect 6722 27376 6790 27432
rect 6846 27376 6914 27432
rect 6970 27376 7038 27432
rect 7094 27376 7104 27432
rect 5168 27308 7104 27376
rect 5168 27252 5178 27308
rect 5234 27252 5302 27308
rect 5358 27252 5426 27308
rect 5482 27252 5550 27308
rect 5606 27252 5674 27308
rect 5730 27252 5798 27308
rect 5854 27252 5922 27308
rect 5978 27252 6046 27308
rect 6102 27252 6170 27308
rect 6226 27252 6294 27308
rect 6350 27252 6418 27308
rect 6474 27252 6542 27308
rect 6598 27252 6666 27308
rect 6722 27252 6790 27308
rect 6846 27252 6914 27308
rect 6970 27252 7038 27308
rect 7094 27252 7104 27308
rect 5168 27242 7104 27252
rect 7874 28548 9810 28558
rect 7874 28492 7884 28548
rect 7940 28492 8008 28548
rect 8064 28492 8132 28548
rect 8188 28492 8256 28548
rect 8312 28492 8380 28548
rect 8436 28492 8504 28548
rect 8560 28492 8628 28548
rect 8684 28492 8752 28548
rect 8808 28492 8876 28548
rect 8932 28492 9000 28548
rect 9056 28492 9124 28548
rect 9180 28492 9248 28548
rect 9304 28492 9372 28548
rect 9428 28492 9496 28548
rect 9552 28492 9620 28548
rect 9676 28492 9744 28548
rect 9800 28492 9810 28548
rect 7874 28424 9810 28492
rect 7874 28368 7884 28424
rect 7940 28368 8008 28424
rect 8064 28368 8132 28424
rect 8188 28368 8256 28424
rect 8312 28368 8380 28424
rect 8436 28368 8504 28424
rect 8560 28368 8628 28424
rect 8684 28368 8752 28424
rect 8808 28368 8876 28424
rect 8932 28368 9000 28424
rect 9056 28368 9124 28424
rect 9180 28368 9248 28424
rect 9304 28368 9372 28424
rect 9428 28368 9496 28424
rect 9552 28368 9620 28424
rect 9676 28368 9744 28424
rect 9800 28368 9810 28424
rect 7874 28300 9810 28368
rect 7874 28244 7884 28300
rect 7940 28244 8008 28300
rect 8064 28244 8132 28300
rect 8188 28244 8256 28300
rect 8312 28244 8380 28300
rect 8436 28244 8504 28300
rect 8560 28244 8628 28300
rect 8684 28244 8752 28300
rect 8808 28244 8876 28300
rect 8932 28244 9000 28300
rect 9056 28244 9124 28300
rect 9180 28244 9248 28300
rect 9304 28244 9372 28300
rect 9428 28244 9496 28300
rect 9552 28244 9620 28300
rect 9676 28244 9744 28300
rect 9800 28244 9810 28300
rect 7874 28176 9810 28244
rect 7874 28120 7884 28176
rect 7940 28120 8008 28176
rect 8064 28120 8132 28176
rect 8188 28120 8256 28176
rect 8312 28120 8380 28176
rect 8436 28120 8504 28176
rect 8560 28120 8628 28176
rect 8684 28120 8752 28176
rect 8808 28120 8876 28176
rect 8932 28120 9000 28176
rect 9056 28120 9124 28176
rect 9180 28120 9248 28176
rect 9304 28120 9372 28176
rect 9428 28120 9496 28176
rect 9552 28120 9620 28176
rect 9676 28120 9744 28176
rect 9800 28120 9810 28176
rect 7874 28052 9810 28120
rect 7874 27996 7884 28052
rect 7940 27996 8008 28052
rect 8064 27996 8132 28052
rect 8188 27996 8256 28052
rect 8312 27996 8380 28052
rect 8436 27996 8504 28052
rect 8560 27996 8628 28052
rect 8684 27996 8752 28052
rect 8808 27996 8876 28052
rect 8932 27996 9000 28052
rect 9056 27996 9124 28052
rect 9180 27996 9248 28052
rect 9304 27996 9372 28052
rect 9428 27996 9496 28052
rect 9552 27996 9620 28052
rect 9676 27996 9744 28052
rect 9800 27996 9810 28052
rect 7874 27928 9810 27996
rect 7874 27872 7884 27928
rect 7940 27872 8008 27928
rect 8064 27872 8132 27928
rect 8188 27872 8256 27928
rect 8312 27872 8380 27928
rect 8436 27872 8504 27928
rect 8560 27872 8628 27928
rect 8684 27872 8752 27928
rect 8808 27872 8876 27928
rect 8932 27872 9000 27928
rect 9056 27872 9124 27928
rect 9180 27872 9248 27928
rect 9304 27872 9372 27928
rect 9428 27872 9496 27928
rect 9552 27872 9620 27928
rect 9676 27872 9744 27928
rect 9800 27872 9810 27928
rect 7874 27804 9810 27872
rect 7874 27748 7884 27804
rect 7940 27748 8008 27804
rect 8064 27748 8132 27804
rect 8188 27748 8256 27804
rect 8312 27748 8380 27804
rect 8436 27748 8504 27804
rect 8560 27748 8628 27804
rect 8684 27748 8752 27804
rect 8808 27748 8876 27804
rect 8932 27748 9000 27804
rect 9056 27748 9124 27804
rect 9180 27748 9248 27804
rect 9304 27748 9372 27804
rect 9428 27748 9496 27804
rect 9552 27748 9620 27804
rect 9676 27748 9744 27804
rect 9800 27748 9810 27804
rect 7874 27680 9810 27748
rect 7874 27624 7884 27680
rect 7940 27624 8008 27680
rect 8064 27624 8132 27680
rect 8188 27624 8256 27680
rect 8312 27624 8380 27680
rect 8436 27624 8504 27680
rect 8560 27624 8628 27680
rect 8684 27624 8752 27680
rect 8808 27624 8876 27680
rect 8932 27624 9000 27680
rect 9056 27624 9124 27680
rect 9180 27624 9248 27680
rect 9304 27624 9372 27680
rect 9428 27624 9496 27680
rect 9552 27624 9620 27680
rect 9676 27624 9744 27680
rect 9800 27624 9810 27680
rect 7874 27556 9810 27624
rect 7874 27500 7884 27556
rect 7940 27500 8008 27556
rect 8064 27500 8132 27556
rect 8188 27500 8256 27556
rect 8312 27500 8380 27556
rect 8436 27500 8504 27556
rect 8560 27500 8628 27556
rect 8684 27500 8752 27556
rect 8808 27500 8876 27556
rect 8932 27500 9000 27556
rect 9056 27500 9124 27556
rect 9180 27500 9248 27556
rect 9304 27500 9372 27556
rect 9428 27500 9496 27556
rect 9552 27500 9620 27556
rect 9676 27500 9744 27556
rect 9800 27500 9810 27556
rect 7874 27432 9810 27500
rect 7874 27376 7884 27432
rect 7940 27376 8008 27432
rect 8064 27376 8132 27432
rect 8188 27376 8256 27432
rect 8312 27376 8380 27432
rect 8436 27376 8504 27432
rect 8560 27376 8628 27432
rect 8684 27376 8752 27432
rect 8808 27376 8876 27432
rect 8932 27376 9000 27432
rect 9056 27376 9124 27432
rect 9180 27376 9248 27432
rect 9304 27376 9372 27432
rect 9428 27376 9496 27432
rect 9552 27376 9620 27432
rect 9676 27376 9744 27432
rect 9800 27376 9810 27432
rect 7874 27308 9810 27376
rect 7874 27252 7884 27308
rect 7940 27252 8008 27308
rect 8064 27252 8132 27308
rect 8188 27252 8256 27308
rect 8312 27252 8380 27308
rect 8436 27252 8504 27308
rect 8560 27252 8628 27308
rect 8684 27252 8752 27308
rect 8808 27252 8876 27308
rect 8932 27252 9000 27308
rect 9056 27252 9124 27308
rect 9180 27252 9248 27308
rect 9304 27252 9372 27308
rect 9428 27252 9496 27308
rect 9552 27252 9620 27308
rect 9676 27252 9744 27308
rect 9800 27252 9810 27308
rect 7874 27242 9810 27252
rect 10244 28548 12180 28558
rect 10244 28492 10254 28548
rect 10310 28492 10378 28548
rect 10434 28492 10502 28548
rect 10558 28492 10626 28548
rect 10682 28492 10750 28548
rect 10806 28492 10874 28548
rect 10930 28492 10998 28548
rect 11054 28492 11122 28548
rect 11178 28492 11246 28548
rect 11302 28492 11370 28548
rect 11426 28492 11494 28548
rect 11550 28492 11618 28548
rect 11674 28492 11742 28548
rect 11798 28492 11866 28548
rect 11922 28492 11990 28548
rect 12046 28492 12114 28548
rect 12170 28492 12180 28548
rect 10244 28424 12180 28492
rect 10244 28368 10254 28424
rect 10310 28368 10378 28424
rect 10434 28368 10502 28424
rect 10558 28368 10626 28424
rect 10682 28368 10750 28424
rect 10806 28368 10874 28424
rect 10930 28368 10998 28424
rect 11054 28368 11122 28424
rect 11178 28368 11246 28424
rect 11302 28368 11370 28424
rect 11426 28368 11494 28424
rect 11550 28368 11618 28424
rect 11674 28368 11742 28424
rect 11798 28368 11866 28424
rect 11922 28368 11990 28424
rect 12046 28368 12114 28424
rect 12170 28368 12180 28424
rect 10244 28300 12180 28368
rect 10244 28244 10254 28300
rect 10310 28244 10378 28300
rect 10434 28244 10502 28300
rect 10558 28244 10626 28300
rect 10682 28244 10750 28300
rect 10806 28244 10874 28300
rect 10930 28244 10998 28300
rect 11054 28244 11122 28300
rect 11178 28244 11246 28300
rect 11302 28244 11370 28300
rect 11426 28244 11494 28300
rect 11550 28244 11618 28300
rect 11674 28244 11742 28300
rect 11798 28244 11866 28300
rect 11922 28244 11990 28300
rect 12046 28244 12114 28300
rect 12170 28244 12180 28300
rect 10244 28176 12180 28244
rect 10244 28120 10254 28176
rect 10310 28120 10378 28176
rect 10434 28120 10502 28176
rect 10558 28120 10626 28176
rect 10682 28120 10750 28176
rect 10806 28120 10874 28176
rect 10930 28120 10998 28176
rect 11054 28120 11122 28176
rect 11178 28120 11246 28176
rect 11302 28120 11370 28176
rect 11426 28120 11494 28176
rect 11550 28120 11618 28176
rect 11674 28120 11742 28176
rect 11798 28120 11866 28176
rect 11922 28120 11990 28176
rect 12046 28120 12114 28176
rect 12170 28120 12180 28176
rect 10244 28052 12180 28120
rect 10244 27996 10254 28052
rect 10310 27996 10378 28052
rect 10434 27996 10502 28052
rect 10558 27996 10626 28052
rect 10682 27996 10750 28052
rect 10806 27996 10874 28052
rect 10930 27996 10998 28052
rect 11054 27996 11122 28052
rect 11178 27996 11246 28052
rect 11302 27996 11370 28052
rect 11426 27996 11494 28052
rect 11550 27996 11618 28052
rect 11674 27996 11742 28052
rect 11798 27996 11866 28052
rect 11922 27996 11990 28052
rect 12046 27996 12114 28052
rect 12170 27996 12180 28052
rect 10244 27928 12180 27996
rect 10244 27872 10254 27928
rect 10310 27872 10378 27928
rect 10434 27872 10502 27928
rect 10558 27872 10626 27928
rect 10682 27872 10750 27928
rect 10806 27872 10874 27928
rect 10930 27872 10998 27928
rect 11054 27872 11122 27928
rect 11178 27872 11246 27928
rect 11302 27872 11370 27928
rect 11426 27872 11494 27928
rect 11550 27872 11618 27928
rect 11674 27872 11742 27928
rect 11798 27872 11866 27928
rect 11922 27872 11990 27928
rect 12046 27872 12114 27928
rect 12170 27872 12180 27928
rect 10244 27804 12180 27872
rect 10244 27748 10254 27804
rect 10310 27748 10378 27804
rect 10434 27748 10502 27804
rect 10558 27748 10626 27804
rect 10682 27748 10750 27804
rect 10806 27748 10874 27804
rect 10930 27748 10998 27804
rect 11054 27748 11122 27804
rect 11178 27748 11246 27804
rect 11302 27748 11370 27804
rect 11426 27748 11494 27804
rect 11550 27748 11618 27804
rect 11674 27748 11742 27804
rect 11798 27748 11866 27804
rect 11922 27748 11990 27804
rect 12046 27748 12114 27804
rect 12170 27748 12180 27804
rect 10244 27680 12180 27748
rect 10244 27624 10254 27680
rect 10310 27624 10378 27680
rect 10434 27624 10502 27680
rect 10558 27624 10626 27680
rect 10682 27624 10750 27680
rect 10806 27624 10874 27680
rect 10930 27624 10998 27680
rect 11054 27624 11122 27680
rect 11178 27624 11246 27680
rect 11302 27624 11370 27680
rect 11426 27624 11494 27680
rect 11550 27624 11618 27680
rect 11674 27624 11742 27680
rect 11798 27624 11866 27680
rect 11922 27624 11990 27680
rect 12046 27624 12114 27680
rect 12170 27624 12180 27680
rect 10244 27556 12180 27624
rect 10244 27500 10254 27556
rect 10310 27500 10378 27556
rect 10434 27500 10502 27556
rect 10558 27500 10626 27556
rect 10682 27500 10750 27556
rect 10806 27500 10874 27556
rect 10930 27500 10998 27556
rect 11054 27500 11122 27556
rect 11178 27500 11246 27556
rect 11302 27500 11370 27556
rect 11426 27500 11494 27556
rect 11550 27500 11618 27556
rect 11674 27500 11742 27556
rect 11798 27500 11866 27556
rect 11922 27500 11990 27556
rect 12046 27500 12114 27556
rect 12170 27500 12180 27556
rect 10244 27432 12180 27500
rect 10244 27376 10254 27432
rect 10310 27376 10378 27432
rect 10434 27376 10502 27432
rect 10558 27376 10626 27432
rect 10682 27376 10750 27432
rect 10806 27376 10874 27432
rect 10930 27376 10998 27432
rect 11054 27376 11122 27432
rect 11178 27376 11246 27432
rect 11302 27376 11370 27432
rect 11426 27376 11494 27432
rect 11550 27376 11618 27432
rect 11674 27376 11742 27432
rect 11798 27376 11866 27432
rect 11922 27376 11990 27432
rect 12046 27376 12114 27432
rect 12170 27376 12180 27432
rect 10244 27308 12180 27376
rect 10244 27252 10254 27308
rect 10310 27252 10378 27308
rect 10434 27252 10502 27308
rect 10558 27252 10626 27308
rect 10682 27252 10750 27308
rect 10806 27252 10874 27308
rect 10930 27252 10998 27308
rect 11054 27252 11122 27308
rect 11178 27252 11246 27308
rect 11302 27252 11370 27308
rect 11426 27252 11494 27308
rect 11550 27252 11618 27308
rect 11674 27252 11742 27308
rect 11798 27252 11866 27308
rect 11922 27252 11990 27308
rect 12046 27252 12114 27308
rect 12170 27252 12180 27308
rect 10244 27242 12180 27252
rect 12861 28548 14673 28558
rect 12861 28492 12871 28548
rect 12927 28492 12995 28548
rect 13051 28492 13119 28548
rect 13175 28492 13243 28548
rect 13299 28492 13367 28548
rect 13423 28492 13491 28548
rect 13547 28492 13615 28548
rect 13671 28492 13739 28548
rect 13795 28492 13863 28548
rect 13919 28492 13987 28548
rect 14043 28492 14111 28548
rect 14167 28492 14235 28548
rect 14291 28492 14359 28548
rect 14415 28492 14483 28548
rect 14539 28492 14607 28548
rect 14663 28492 14673 28548
rect 12861 28424 14673 28492
rect 12861 28368 12871 28424
rect 12927 28368 12995 28424
rect 13051 28368 13119 28424
rect 13175 28368 13243 28424
rect 13299 28368 13367 28424
rect 13423 28368 13491 28424
rect 13547 28368 13615 28424
rect 13671 28368 13739 28424
rect 13795 28368 13863 28424
rect 13919 28368 13987 28424
rect 14043 28368 14111 28424
rect 14167 28368 14235 28424
rect 14291 28368 14359 28424
rect 14415 28368 14483 28424
rect 14539 28368 14607 28424
rect 14663 28368 14673 28424
rect 12861 28300 14673 28368
rect 12861 28244 12871 28300
rect 12927 28244 12995 28300
rect 13051 28244 13119 28300
rect 13175 28244 13243 28300
rect 13299 28244 13367 28300
rect 13423 28244 13491 28300
rect 13547 28244 13615 28300
rect 13671 28244 13739 28300
rect 13795 28244 13863 28300
rect 13919 28244 13987 28300
rect 14043 28244 14111 28300
rect 14167 28244 14235 28300
rect 14291 28244 14359 28300
rect 14415 28244 14483 28300
rect 14539 28244 14607 28300
rect 14663 28244 14673 28300
rect 12861 28176 14673 28244
rect 12861 28120 12871 28176
rect 12927 28120 12995 28176
rect 13051 28120 13119 28176
rect 13175 28120 13243 28176
rect 13299 28120 13367 28176
rect 13423 28120 13491 28176
rect 13547 28120 13615 28176
rect 13671 28120 13739 28176
rect 13795 28120 13863 28176
rect 13919 28120 13987 28176
rect 14043 28120 14111 28176
rect 14167 28120 14235 28176
rect 14291 28120 14359 28176
rect 14415 28120 14483 28176
rect 14539 28120 14607 28176
rect 14663 28120 14673 28176
rect 12861 28052 14673 28120
rect 12861 27996 12871 28052
rect 12927 27996 12995 28052
rect 13051 27996 13119 28052
rect 13175 27996 13243 28052
rect 13299 27996 13367 28052
rect 13423 27996 13491 28052
rect 13547 27996 13615 28052
rect 13671 27996 13739 28052
rect 13795 27996 13863 28052
rect 13919 27996 13987 28052
rect 14043 27996 14111 28052
rect 14167 27996 14235 28052
rect 14291 27996 14359 28052
rect 14415 27996 14483 28052
rect 14539 27996 14607 28052
rect 14663 27996 14673 28052
rect 12861 27928 14673 27996
rect 12861 27872 12871 27928
rect 12927 27872 12995 27928
rect 13051 27872 13119 27928
rect 13175 27872 13243 27928
rect 13299 27872 13367 27928
rect 13423 27872 13491 27928
rect 13547 27872 13615 27928
rect 13671 27872 13739 27928
rect 13795 27872 13863 27928
rect 13919 27872 13987 27928
rect 14043 27872 14111 27928
rect 14167 27872 14235 27928
rect 14291 27872 14359 27928
rect 14415 27872 14483 27928
rect 14539 27872 14607 27928
rect 14663 27872 14673 27928
rect 12861 27804 14673 27872
rect 12861 27748 12871 27804
rect 12927 27748 12995 27804
rect 13051 27748 13119 27804
rect 13175 27748 13243 27804
rect 13299 27748 13367 27804
rect 13423 27748 13491 27804
rect 13547 27748 13615 27804
rect 13671 27748 13739 27804
rect 13795 27748 13863 27804
rect 13919 27748 13987 27804
rect 14043 27748 14111 27804
rect 14167 27748 14235 27804
rect 14291 27748 14359 27804
rect 14415 27748 14483 27804
rect 14539 27748 14607 27804
rect 14663 27748 14673 27804
rect 12861 27680 14673 27748
rect 12861 27624 12871 27680
rect 12927 27624 12995 27680
rect 13051 27624 13119 27680
rect 13175 27624 13243 27680
rect 13299 27624 13367 27680
rect 13423 27624 13491 27680
rect 13547 27624 13615 27680
rect 13671 27624 13739 27680
rect 13795 27624 13863 27680
rect 13919 27624 13987 27680
rect 14043 27624 14111 27680
rect 14167 27624 14235 27680
rect 14291 27624 14359 27680
rect 14415 27624 14483 27680
rect 14539 27624 14607 27680
rect 14663 27624 14673 27680
rect 12861 27556 14673 27624
rect 12861 27500 12871 27556
rect 12927 27500 12995 27556
rect 13051 27500 13119 27556
rect 13175 27500 13243 27556
rect 13299 27500 13367 27556
rect 13423 27500 13491 27556
rect 13547 27500 13615 27556
rect 13671 27500 13739 27556
rect 13795 27500 13863 27556
rect 13919 27500 13987 27556
rect 14043 27500 14111 27556
rect 14167 27500 14235 27556
rect 14291 27500 14359 27556
rect 14415 27500 14483 27556
rect 14539 27500 14607 27556
rect 14663 27500 14673 27556
rect 12861 27432 14673 27500
rect 12861 27376 12871 27432
rect 12927 27376 12995 27432
rect 13051 27376 13119 27432
rect 13175 27376 13243 27432
rect 13299 27376 13367 27432
rect 13423 27376 13491 27432
rect 13547 27376 13615 27432
rect 13671 27376 13739 27432
rect 13795 27376 13863 27432
rect 13919 27376 13987 27432
rect 14043 27376 14111 27432
rect 14167 27376 14235 27432
rect 14291 27376 14359 27432
rect 14415 27376 14483 27432
rect 14539 27376 14607 27432
rect 14663 27376 14673 27432
rect 12861 27308 14673 27376
rect 12861 27252 12871 27308
rect 12927 27252 12995 27308
rect 13051 27252 13119 27308
rect 13175 27252 13243 27308
rect 13299 27252 13367 27308
rect 13423 27252 13491 27308
rect 13547 27252 13615 27308
rect 13671 27252 13739 27308
rect 13795 27252 13863 27308
rect 13919 27252 13987 27308
rect 14043 27252 14111 27308
rect 14167 27252 14235 27308
rect 14291 27252 14359 27308
rect 14415 27252 14483 27308
rect 14539 27252 14607 27308
rect 14663 27252 14673 27308
rect 12861 27242 14673 27252
rect -11 27214 86 27224
rect 14892 27224 14902 28576
rect 14958 27224 14989 28576
rect 14892 27214 14989 27224
rect 2481 26954 2681 26964
rect 2481 26898 2491 26954
rect 2547 26898 2615 26954
rect 2671 26898 2681 26954
rect 2481 26830 2681 26898
rect 2481 26774 2491 26830
rect 2547 26774 2615 26830
rect 2671 26774 2681 26830
rect 2481 26706 2681 26774
rect 2481 26650 2491 26706
rect 2547 26650 2615 26706
rect 2671 26650 2681 26706
rect 2481 26582 2681 26650
rect 2481 26526 2491 26582
rect 2547 26526 2615 26582
rect 2671 26526 2681 26582
rect 2481 26458 2681 26526
rect 2481 26402 2491 26458
rect 2547 26402 2615 26458
rect 2671 26402 2681 26458
rect 2481 26334 2681 26402
rect 2481 26278 2491 26334
rect 2547 26278 2615 26334
rect 2671 26278 2681 26334
rect 2481 26210 2681 26278
rect 2481 26154 2491 26210
rect 2547 26154 2615 26210
rect 2671 26154 2681 26210
rect 2481 26086 2681 26154
rect 2481 26030 2491 26086
rect 2547 26030 2615 26086
rect 2671 26030 2681 26086
rect 2481 25962 2681 26030
rect 2481 25906 2491 25962
rect 2547 25906 2615 25962
rect 2671 25906 2681 25962
rect 2481 25838 2681 25906
rect 2481 25782 2491 25838
rect 2547 25782 2615 25838
rect 2671 25782 2681 25838
rect 2481 25714 2681 25782
rect 2481 25658 2491 25714
rect 2547 25658 2615 25714
rect 2671 25658 2681 25714
rect 2481 25590 2681 25658
rect 2481 25534 2491 25590
rect 2547 25534 2615 25590
rect 2671 25534 2681 25590
rect 2481 25466 2681 25534
rect 2481 25410 2491 25466
rect 2547 25410 2615 25466
rect 2671 25410 2681 25466
rect 2481 25342 2681 25410
rect 2481 25286 2491 25342
rect 2547 25286 2615 25342
rect 2671 25286 2681 25342
rect 2481 25218 2681 25286
rect 2481 25162 2491 25218
rect 2547 25162 2615 25218
rect 2671 25162 2681 25218
rect 2481 25094 2681 25162
rect 2481 25038 2491 25094
rect 2547 25038 2615 25094
rect 2671 25038 2681 25094
rect 2481 24970 2681 25038
rect 2481 24914 2491 24970
rect 2547 24914 2615 24970
rect 2671 24914 2681 24970
rect 2481 24846 2681 24914
rect 2481 24790 2491 24846
rect 2547 24790 2615 24846
rect 2671 24790 2681 24846
rect 2481 24722 2681 24790
rect 2481 24666 2491 24722
rect 2547 24666 2615 24722
rect 2671 24666 2681 24722
rect 2481 24598 2681 24666
rect 2481 24542 2491 24598
rect 2547 24542 2615 24598
rect 2671 24542 2681 24598
rect 2481 24474 2681 24542
rect 2481 24418 2491 24474
rect 2547 24418 2615 24474
rect 2671 24418 2681 24474
rect 2481 24350 2681 24418
rect 2481 24294 2491 24350
rect 2547 24294 2615 24350
rect 2671 24294 2681 24350
rect 2481 24226 2681 24294
rect 2481 24170 2491 24226
rect 2547 24170 2615 24226
rect 2671 24170 2681 24226
rect 2481 24102 2681 24170
rect 2481 24046 2491 24102
rect 2547 24046 2615 24102
rect 2671 24046 2681 24102
rect 2481 24036 2681 24046
rect 4851 26954 5051 26964
rect 4851 26898 4861 26954
rect 4917 26898 4985 26954
rect 5041 26898 5051 26954
rect 4851 26830 5051 26898
rect 4851 26774 4861 26830
rect 4917 26774 4985 26830
rect 5041 26774 5051 26830
rect 4851 26706 5051 26774
rect 4851 26650 4861 26706
rect 4917 26650 4985 26706
rect 5041 26650 5051 26706
rect 4851 26582 5051 26650
rect 4851 26526 4861 26582
rect 4917 26526 4985 26582
rect 5041 26526 5051 26582
rect 4851 26458 5051 26526
rect 4851 26402 4861 26458
rect 4917 26402 4985 26458
rect 5041 26402 5051 26458
rect 4851 26334 5051 26402
rect 4851 26278 4861 26334
rect 4917 26278 4985 26334
rect 5041 26278 5051 26334
rect 4851 26210 5051 26278
rect 4851 26154 4861 26210
rect 4917 26154 4985 26210
rect 5041 26154 5051 26210
rect 4851 26086 5051 26154
rect 4851 26030 4861 26086
rect 4917 26030 4985 26086
rect 5041 26030 5051 26086
rect 4851 25962 5051 26030
rect 4851 25906 4861 25962
rect 4917 25906 4985 25962
rect 5041 25906 5051 25962
rect 4851 25838 5051 25906
rect 4851 25782 4861 25838
rect 4917 25782 4985 25838
rect 5041 25782 5051 25838
rect 4851 25714 5051 25782
rect 4851 25658 4861 25714
rect 4917 25658 4985 25714
rect 5041 25658 5051 25714
rect 4851 25590 5051 25658
rect 4851 25534 4861 25590
rect 4917 25534 4985 25590
rect 5041 25534 5051 25590
rect 4851 25466 5051 25534
rect 4851 25410 4861 25466
rect 4917 25410 4985 25466
rect 5041 25410 5051 25466
rect 4851 25342 5051 25410
rect 4851 25286 4861 25342
rect 4917 25286 4985 25342
rect 5041 25286 5051 25342
rect 4851 25218 5051 25286
rect 4851 25162 4861 25218
rect 4917 25162 4985 25218
rect 5041 25162 5051 25218
rect 4851 25094 5051 25162
rect 4851 25038 4861 25094
rect 4917 25038 4985 25094
rect 5041 25038 5051 25094
rect 4851 24970 5051 25038
rect 4851 24914 4861 24970
rect 4917 24914 4985 24970
rect 5041 24914 5051 24970
rect 4851 24846 5051 24914
rect 4851 24790 4861 24846
rect 4917 24790 4985 24846
rect 5041 24790 5051 24846
rect 4851 24722 5051 24790
rect 4851 24666 4861 24722
rect 4917 24666 4985 24722
rect 5041 24666 5051 24722
rect 4851 24598 5051 24666
rect 4851 24542 4861 24598
rect 4917 24542 4985 24598
rect 5041 24542 5051 24598
rect 4851 24474 5051 24542
rect 4851 24418 4861 24474
rect 4917 24418 4985 24474
rect 5041 24418 5051 24474
rect 4851 24350 5051 24418
rect 4851 24294 4861 24350
rect 4917 24294 4985 24350
rect 5041 24294 5051 24350
rect 4851 24226 5051 24294
rect 4851 24170 4861 24226
rect 4917 24170 4985 24226
rect 5041 24170 5051 24226
rect 4851 24102 5051 24170
rect 4851 24046 4861 24102
rect 4917 24046 4985 24102
rect 5041 24046 5051 24102
rect 4851 24036 5051 24046
rect 7265 26954 7713 26964
rect 7265 26898 7275 26954
rect 7331 26898 7399 26954
rect 7455 26898 7523 26954
rect 7579 26898 7647 26954
rect 7703 26898 7713 26954
rect 7265 26830 7713 26898
rect 7265 26774 7275 26830
rect 7331 26774 7399 26830
rect 7455 26774 7523 26830
rect 7579 26774 7647 26830
rect 7703 26774 7713 26830
rect 7265 26706 7713 26774
rect 7265 26650 7275 26706
rect 7331 26650 7399 26706
rect 7455 26650 7523 26706
rect 7579 26650 7647 26706
rect 7703 26650 7713 26706
rect 7265 26582 7713 26650
rect 7265 26526 7275 26582
rect 7331 26526 7399 26582
rect 7455 26526 7523 26582
rect 7579 26526 7647 26582
rect 7703 26526 7713 26582
rect 7265 26458 7713 26526
rect 7265 26402 7275 26458
rect 7331 26402 7399 26458
rect 7455 26402 7523 26458
rect 7579 26402 7647 26458
rect 7703 26402 7713 26458
rect 7265 26334 7713 26402
rect 7265 26278 7275 26334
rect 7331 26278 7399 26334
rect 7455 26278 7523 26334
rect 7579 26278 7647 26334
rect 7703 26278 7713 26334
rect 7265 26210 7713 26278
rect 7265 26154 7275 26210
rect 7331 26154 7399 26210
rect 7455 26154 7523 26210
rect 7579 26154 7647 26210
rect 7703 26154 7713 26210
rect 7265 26086 7713 26154
rect 7265 26030 7275 26086
rect 7331 26030 7399 26086
rect 7455 26030 7523 26086
rect 7579 26030 7647 26086
rect 7703 26030 7713 26086
rect 7265 25962 7713 26030
rect 7265 25906 7275 25962
rect 7331 25906 7399 25962
rect 7455 25906 7523 25962
rect 7579 25906 7647 25962
rect 7703 25906 7713 25962
rect 7265 25838 7713 25906
rect 7265 25782 7275 25838
rect 7331 25782 7399 25838
rect 7455 25782 7523 25838
rect 7579 25782 7647 25838
rect 7703 25782 7713 25838
rect 7265 25714 7713 25782
rect 7265 25658 7275 25714
rect 7331 25658 7399 25714
rect 7455 25658 7523 25714
rect 7579 25658 7647 25714
rect 7703 25658 7713 25714
rect 7265 25590 7713 25658
rect 7265 25534 7275 25590
rect 7331 25534 7399 25590
rect 7455 25534 7523 25590
rect 7579 25534 7647 25590
rect 7703 25534 7713 25590
rect 7265 25466 7713 25534
rect 7265 25410 7275 25466
rect 7331 25410 7399 25466
rect 7455 25410 7523 25466
rect 7579 25410 7647 25466
rect 7703 25410 7713 25466
rect 7265 25342 7713 25410
rect 7265 25286 7275 25342
rect 7331 25286 7399 25342
rect 7455 25286 7523 25342
rect 7579 25286 7647 25342
rect 7703 25286 7713 25342
rect 7265 25218 7713 25286
rect 7265 25162 7275 25218
rect 7331 25162 7399 25218
rect 7455 25162 7523 25218
rect 7579 25162 7647 25218
rect 7703 25162 7713 25218
rect 7265 25094 7713 25162
rect 7265 25038 7275 25094
rect 7331 25038 7399 25094
rect 7455 25038 7523 25094
rect 7579 25038 7647 25094
rect 7703 25038 7713 25094
rect 7265 24970 7713 25038
rect 7265 24914 7275 24970
rect 7331 24914 7399 24970
rect 7455 24914 7523 24970
rect 7579 24914 7647 24970
rect 7703 24914 7713 24970
rect 7265 24846 7713 24914
rect 7265 24790 7275 24846
rect 7331 24790 7399 24846
rect 7455 24790 7523 24846
rect 7579 24790 7647 24846
rect 7703 24790 7713 24846
rect 7265 24722 7713 24790
rect 7265 24666 7275 24722
rect 7331 24666 7399 24722
rect 7455 24666 7523 24722
rect 7579 24666 7647 24722
rect 7703 24666 7713 24722
rect 7265 24598 7713 24666
rect 7265 24542 7275 24598
rect 7331 24542 7399 24598
rect 7455 24542 7523 24598
rect 7579 24542 7647 24598
rect 7703 24542 7713 24598
rect 7265 24474 7713 24542
rect 7265 24418 7275 24474
rect 7331 24418 7399 24474
rect 7455 24418 7523 24474
rect 7579 24418 7647 24474
rect 7703 24418 7713 24474
rect 7265 24350 7713 24418
rect 7265 24294 7275 24350
rect 7331 24294 7399 24350
rect 7455 24294 7523 24350
rect 7579 24294 7647 24350
rect 7703 24294 7713 24350
rect 7265 24226 7713 24294
rect 7265 24170 7275 24226
rect 7331 24170 7399 24226
rect 7455 24170 7523 24226
rect 7579 24170 7647 24226
rect 7703 24170 7713 24226
rect 7265 24102 7713 24170
rect 7265 24046 7275 24102
rect 7331 24046 7399 24102
rect 7455 24046 7523 24102
rect 7579 24046 7647 24102
rect 7703 24046 7713 24102
rect 7265 24036 7713 24046
rect 9927 26954 10127 26964
rect 9927 26898 9937 26954
rect 9993 26898 10061 26954
rect 10117 26898 10127 26954
rect 9927 26830 10127 26898
rect 9927 26774 9937 26830
rect 9993 26774 10061 26830
rect 10117 26774 10127 26830
rect 9927 26706 10127 26774
rect 9927 26650 9937 26706
rect 9993 26650 10061 26706
rect 10117 26650 10127 26706
rect 9927 26582 10127 26650
rect 9927 26526 9937 26582
rect 9993 26526 10061 26582
rect 10117 26526 10127 26582
rect 9927 26458 10127 26526
rect 9927 26402 9937 26458
rect 9993 26402 10061 26458
rect 10117 26402 10127 26458
rect 9927 26334 10127 26402
rect 9927 26278 9937 26334
rect 9993 26278 10061 26334
rect 10117 26278 10127 26334
rect 9927 26210 10127 26278
rect 9927 26154 9937 26210
rect 9993 26154 10061 26210
rect 10117 26154 10127 26210
rect 9927 26086 10127 26154
rect 9927 26030 9937 26086
rect 9993 26030 10061 26086
rect 10117 26030 10127 26086
rect 9927 25962 10127 26030
rect 9927 25906 9937 25962
rect 9993 25906 10061 25962
rect 10117 25906 10127 25962
rect 9927 25838 10127 25906
rect 9927 25782 9937 25838
rect 9993 25782 10061 25838
rect 10117 25782 10127 25838
rect 9927 25714 10127 25782
rect 9927 25658 9937 25714
rect 9993 25658 10061 25714
rect 10117 25658 10127 25714
rect 9927 25590 10127 25658
rect 9927 25534 9937 25590
rect 9993 25534 10061 25590
rect 10117 25534 10127 25590
rect 9927 25466 10127 25534
rect 9927 25410 9937 25466
rect 9993 25410 10061 25466
rect 10117 25410 10127 25466
rect 9927 25342 10127 25410
rect 9927 25286 9937 25342
rect 9993 25286 10061 25342
rect 10117 25286 10127 25342
rect 9927 25218 10127 25286
rect 9927 25162 9937 25218
rect 9993 25162 10061 25218
rect 10117 25162 10127 25218
rect 9927 25094 10127 25162
rect 9927 25038 9937 25094
rect 9993 25038 10061 25094
rect 10117 25038 10127 25094
rect 9927 24970 10127 25038
rect 9927 24914 9937 24970
rect 9993 24914 10061 24970
rect 10117 24914 10127 24970
rect 9927 24846 10127 24914
rect 9927 24790 9937 24846
rect 9993 24790 10061 24846
rect 10117 24790 10127 24846
rect 9927 24722 10127 24790
rect 9927 24666 9937 24722
rect 9993 24666 10061 24722
rect 10117 24666 10127 24722
rect 9927 24598 10127 24666
rect 9927 24542 9937 24598
rect 9993 24542 10061 24598
rect 10117 24542 10127 24598
rect 9927 24474 10127 24542
rect 9927 24418 9937 24474
rect 9993 24418 10061 24474
rect 10117 24418 10127 24474
rect 9927 24350 10127 24418
rect 9927 24294 9937 24350
rect 9993 24294 10061 24350
rect 10117 24294 10127 24350
rect 9927 24226 10127 24294
rect 9927 24170 9937 24226
rect 9993 24170 10061 24226
rect 10117 24170 10127 24226
rect 9927 24102 10127 24170
rect 9927 24046 9937 24102
rect 9993 24046 10061 24102
rect 10117 24046 10127 24102
rect 9927 24036 10127 24046
rect 12297 26954 12497 26964
rect 12297 26898 12307 26954
rect 12363 26898 12431 26954
rect 12487 26898 12497 26954
rect 12297 26830 12497 26898
rect 12297 26774 12307 26830
rect 12363 26774 12431 26830
rect 12487 26774 12497 26830
rect 12297 26706 12497 26774
rect 12297 26650 12307 26706
rect 12363 26650 12431 26706
rect 12487 26650 12497 26706
rect 12297 26582 12497 26650
rect 12297 26526 12307 26582
rect 12363 26526 12431 26582
rect 12487 26526 12497 26582
rect 12297 26458 12497 26526
rect 12297 26402 12307 26458
rect 12363 26402 12431 26458
rect 12487 26402 12497 26458
rect 12297 26334 12497 26402
rect 12297 26278 12307 26334
rect 12363 26278 12431 26334
rect 12487 26278 12497 26334
rect 12297 26210 12497 26278
rect 12297 26154 12307 26210
rect 12363 26154 12431 26210
rect 12487 26154 12497 26210
rect 12297 26086 12497 26154
rect 12297 26030 12307 26086
rect 12363 26030 12431 26086
rect 12487 26030 12497 26086
rect 12297 25962 12497 26030
rect 12297 25906 12307 25962
rect 12363 25906 12431 25962
rect 12487 25906 12497 25962
rect 12297 25838 12497 25906
rect 12297 25782 12307 25838
rect 12363 25782 12431 25838
rect 12487 25782 12497 25838
rect 12297 25714 12497 25782
rect 12297 25658 12307 25714
rect 12363 25658 12431 25714
rect 12487 25658 12497 25714
rect 12297 25590 12497 25658
rect 12297 25534 12307 25590
rect 12363 25534 12431 25590
rect 12487 25534 12497 25590
rect 12297 25466 12497 25534
rect 12297 25410 12307 25466
rect 12363 25410 12431 25466
rect 12487 25410 12497 25466
rect 12297 25342 12497 25410
rect 12297 25286 12307 25342
rect 12363 25286 12431 25342
rect 12487 25286 12497 25342
rect 12297 25218 12497 25286
rect 12297 25162 12307 25218
rect 12363 25162 12431 25218
rect 12487 25162 12497 25218
rect 12297 25094 12497 25162
rect 12297 25038 12307 25094
rect 12363 25038 12431 25094
rect 12487 25038 12497 25094
rect 12297 24970 12497 25038
rect 12297 24914 12307 24970
rect 12363 24914 12431 24970
rect 12487 24914 12497 24970
rect 12297 24846 12497 24914
rect 12297 24790 12307 24846
rect 12363 24790 12431 24846
rect 12487 24790 12497 24846
rect 12297 24722 12497 24790
rect 12297 24666 12307 24722
rect 12363 24666 12431 24722
rect 12487 24666 12497 24722
rect 12297 24598 12497 24666
rect 12297 24542 12307 24598
rect 12363 24542 12431 24598
rect 12487 24542 12497 24598
rect 12297 24474 12497 24542
rect 12297 24418 12307 24474
rect 12363 24418 12431 24474
rect 12487 24418 12497 24474
rect 12297 24350 12497 24418
rect 12297 24294 12307 24350
rect 12363 24294 12431 24350
rect 12487 24294 12497 24350
rect 12297 24226 12497 24294
rect 12297 24170 12307 24226
rect 12363 24170 12431 24226
rect 12487 24170 12497 24226
rect 12297 24102 12497 24170
rect 12297 24046 12307 24102
rect 12363 24046 12431 24102
rect 12487 24046 12497 24102
rect 12297 24036 12497 24046
rect 2481 23754 2681 23764
rect 2481 23698 2491 23754
rect 2547 23698 2615 23754
rect 2671 23698 2681 23754
rect 2481 23630 2681 23698
rect 2481 23574 2491 23630
rect 2547 23574 2615 23630
rect 2671 23574 2681 23630
rect 2481 23506 2681 23574
rect 2481 23450 2491 23506
rect 2547 23450 2615 23506
rect 2671 23450 2681 23506
rect 2481 23382 2681 23450
rect 2481 23326 2491 23382
rect 2547 23326 2615 23382
rect 2671 23326 2681 23382
rect 2481 23258 2681 23326
rect 2481 23202 2491 23258
rect 2547 23202 2615 23258
rect 2671 23202 2681 23258
rect 2481 23134 2681 23202
rect 2481 23078 2491 23134
rect 2547 23078 2615 23134
rect 2671 23078 2681 23134
rect 2481 23010 2681 23078
rect 2481 22954 2491 23010
rect 2547 22954 2615 23010
rect 2671 22954 2681 23010
rect 2481 22886 2681 22954
rect 2481 22830 2491 22886
rect 2547 22830 2615 22886
rect 2671 22830 2681 22886
rect 2481 22762 2681 22830
rect 2481 22706 2491 22762
rect 2547 22706 2615 22762
rect 2671 22706 2681 22762
rect 2481 22638 2681 22706
rect 2481 22582 2491 22638
rect 2547 22582 2615 22638
rect 2671 22582 2681 22638
rect 2481 22514 2681 22582
rect 2481 22458 2491 22514
rect 2547 22458 2615 22514
rect 2671 22458 2681 22514
rect 2481 22390 2681 22458
rect 2481 22334 2491 22390
rect 2547 22334 2615 22390
rect 2671 22334 2681 22390
rect 2481 22266 2681 22334
rect 2481 22210 2491 22266
rect 2547 22210 2615 22266
rect 2671 22210 2681 22266
rect 2481 22142 2681 22210
rect 2481 22086 2491 22142
rect 2547 22086 2615 22142
rect 2671 22086 2681 22142
rect 2481 22018 2681 22086
rect 2481 21962 2491 22018
rect 2547 21962 2615 22018
rect 2671 21962 2681 22018
rect 2481 21894 2681 21962
rect 2481 21838 2491 21894
rect 2547 21838 2615 21894
rect 2671 21838 2681 21894
rect 2481 21770 2681 21838
rect 2481 21714 2491 21770
rect 2547 21714 2615 21770
rect 2671 21714 2681 21770
rect 2481 21646 2681 21714
rect 2481 21590 2491 21646
rect 2547 21590 2615 21646
rect 2671 21590 2681 21646
rect 2481 21522 2681 21590
rect 2481 21466 2491 21522
rect 2547 21466 2615 21522
rect 2671 21466 2681 21522
rect 2481 21398 2681 21466
rect 2481 21342 2491 21398
rect 2547 21342 2615 21398
rect 2671 21342 2681 21398
rect 2481 21274 2681 21342
rect 2481 21218 2491 21274
rect 2547 21218 2615 21274
rect 2671 21218 2681 21274
rect 2481 21150 2681 21218
rect 2481 21094 2491 21150
rect 2547 21094 2615 21150
rect 2671 21094 2681 21150
rect 2481 21026 2681 21094
rect 2481 20970 2491 21026
rect 2547 20970 2615 21026
rect 2671 20970 2681 21026
rect 2481 20902 2681 20970
rect 2481 20846 2491 20902
rect 2547 20846 2615 20902
rect 2671 20846 2681 20902
rect 2481 20836 2681 20846
rect 4851 23754 5051 23764
rect 4851 23698 4861 23754
rect 4917 23698 4985 23754
rect 5041 23698 5051 23754
rect 4851 23630 5051 23698
rect 4851 23574 4861 23630
rect 4917 23574 4985 23630
rect 5041 23574 5051 23630
rect 4851 23506 5051 23574
rect 4851 23450 4861 23506
rect 4917 23450 4985 23506
rect 5041 23450 5051 23506
rect 4851 23382 5051 23450
rect 4851 23326 4861 23382
rect 4917 23326 4985 23382
rect 5041 23326 5051 23382
rect 4851 23258 5051 23326
rect 4851 23202 4861 23258
rect 4917 23202 4985 23258
rect 5041 23202 5051 23258
rect 4851 23134 5051 23202
rect 4851 23078 4861 23134
rect 4917 23078 4985 23134
rect 5041 23078 5051 23134
rect 4851 23010 5051 23078
rect 4851 22954 4861 23010
rect 4917 22954 4985 23010
rect 5041 22954 5051 23010
rect 4851 22886 5051 22954
rect 4851 22830 4861 22886
rect 4917 22830 4985 22886
rect 5041 22830 5051 22886
rect 4851 22762 5051 22830
rect 4851 22706 4861 22762
rect 4917 22706 4985 22762
rect 5041 22706 5051 22762
rect 4851 22638 5051 22706
rect 4851 22582 4861 22638
rect 4917 22582 4985 22638
rect 5041 22582 5051 22638
rect 4851 22514 5051 22582
rect 4851 22458 4861 22514
rect 4917 22458 4985 22514
rect 5041 22458 5051 22514
rect 4851 22390 5051 22458
rect 4851 22334 4861 22390
rect 4917 22334 4985 22390
rect 5041 22334 5051 22390
rect 4851 22266 5051 22334
rect 4851 22210 4861 22266
rect 4917 22210 4985 22266
rect 5041 22210 5051 22266
rect 4851 22142 5051 22210
rect 4851 22086 4861 22142
rect 4917 22086 4985 22142
rect 5041 22086 5051 22142
rect 4851 22018 5051 22086
rect 4851 21962 4861 22018
rect 4917 21962 4985 22018
rect 5041 21962 5051 22018
rect 4851 21894 5051 21962
rect 4851 21838 4861 21894
rect 4917 21838 4985 21894
rect 5041 21838 5051 21894
rect 4851 21770 5051 21838
rect 4851 21714 4861 21770
rect 4917 21714 4985 21770
rect 5041 21714 5051 21770
rect 4851 21646 5051 21714
rect 4851 21590 4861 21646
rect 4917 21590 4985 21646
rect 5041 21590 5051 21646
rect 4851 21522 5051 21590
rect 4851 21466 4861 21522
rect 4917 21466 4985 21522
rect 5041 21466 5051 21522
rect 4851 21398 5051 21466
rect 4851 21342 4861 21398
rect 4917 21342 4985 21398
rect 5041 21342 5051 21398
rect 4851 21274 5051 21342
rect 4851 21218 4861 21274
rect 4917 21218 4985 21274
rect 5041 21218 5051 21274
rect 4851 21150 5051 21218
rect 4851 21094 4861 21150
rect 4917 21094 4985 21150
rect 5041 21094 5051 21150
rect 4851 21026 5051 21094
rect 4851 20970 4861 21026
rect 4917 20970 4985 21026
rect 5041 20970 5051 21026
rect 4851 20902 5051 20970
rect 4851 20846 4861 20902
rect 4917 20846 4985 20902
rect 5041 20846 5051 20902
rect 4851 20836 5051 20846
rect 7265 23754 7713 23764
rect 7265 23698 7275 23754
rect 7331 23698 7399 23754
rect 7455 23698 7523 23754
rect 7579 23698 7647 23754
rect 7703 23698 7713 23754
rect 7265 23630 7713 23698
rect 7265 23574 7275 23630
rect 7331 23574 7399 23630
rect 7455 23574 7523 23630
rect 7579 23574 7647 23630
rect 7703 23574 7713 23630
rect 7265 23506 7713 23574
rect 7265 23450 7275 23506
rect 7331 23450 7399 23506
rect 7455 23450 7523 23506
rect 7579 23450 7647 23506
rect 7703 23450 7713 23506
rect 7265 23382 7713 23450
rect 7265 23326 7275 23382
rect 7331 23326 7399 23382
rect 7455 23326 7523 23382
rect 7579 23326 7647 23382
rect 7703 23326 7713 23382
rect 7265 23258 7713 23326
rect 7265 23202 7275 23258
rect 7331 23202 7399 23258
rect 7455 23202 7523 23258
rect 7579 23202 7647 23258
rect 7703 23202 7713 23258
rect 7265 23134 7713 23202
rect 7265 23078 7275 23134
rect 7331 23078 7399 23134
rect 7455 23078 7523 23134
rect 7579 23078 7647 23134
rect 7703 23078 7713 23134
rect 7265 23010 7713 23078
rect 7265 22954 7275 23010
rect 7331 22954 7399 23010
rect 7455 22954 7523 23010
rect 7579 22954 7647 23010
rect 7703 22954 7713 23010
rect 7265 22886 7713 22954
rect 7265 22830 7275 22886
rect 7331 22830 7399 22886
rect 7455 22830 7523 22886
rect 7579 22830 7647 22886
rect 7703 22830 7713 22886
rect 7265 22762 7713 22830
rect 7265 22706 7275 22762
rect 7331 22706 7399 22762
rect 7455 22706 7523 22762
rect 7579 22706 7647 22762
rect 7703 22706 7713 22762
rect 7265 22638 7713 22706
rect 7265 22582 7275 22638
rect 7331 22582 7399 22638
rect 7455 22582 7523 22638
rect 7579 22582 7647 22638
rect 7703 22582 7713 22638
rect 7265 22514 7713 22582
rect 7265 22458 7275 22514
rect 7331 22458 7399 22514
rect 7455 22458 7523 22514
rect 7579 22458 7647 22514
rect 7703 22458 7713 22514
rect 7265 22390 7713 22458
rect 7265 22334 7275 22390
rect 7331 22334 7399 22390
rect 7455 22334 7523 22390
rect 7579 22334 7647 22390
rect 7703 22334 7713 22390
rect 7265 22266 7713 22334
rect 7265 22210 7275 22266
rect 7331 22210 7399 22266
rect 7455 22210 7523 22266
rect 7579 22210 7647 22266
rect 7703 22210 7713 22266
rect 7265 22142 7713 22210
rect 7265 22086 7275 22142
rect 7331 22086 7399 22142
rect 7455 22086 7523 22142
rect 7579 22086 7647 22142
rect 7703 22086 7713 22142
rect 7265 22018 7713 22086
rect 7265 21962 7275 22018
rect 7331 21962 7399 22018
rect 7455 21962 7523 22018
rect 7579 21962 7647 22018
rect 7703 21962 7713 22018
rect 7265 21894 7713 21962
rect 7265 21838 7275 21894
rect 7331 21838 7399 21894
rect 7455 21838 7523 21894
rect 7579 21838 7647 21894
rect 7703 21838 7713 21894
rect 7265 21770 7713 21838
rect 7265 21714 7275 21770
rect 7331 21714 7399 21770
rect 7455 21714 7523 21770
rect 7579 21714 7647 21770
rect 7703 21714 7713 21770
rect 7265 21646 7713 21714
rect 7265 21590 7275 21646
rect 7331 21590 7399 21646
rect 7455 21590 7523 21646
rect 7579 21590 7647 21646
rect 7703 21590 7713 21646
rect 7265 21522 7713 21590
rect 7265 21466 7275 21522
rect 7331 21466 7399 21522
rect 7455 21466 7523 21522
rect 7579 21466 7647 21522
rect 7703 21466 7713 21522
rect 7265 21398 7713 21466
rect 7265 21342 7275 21398
rect 7331 21342 7399 21398
rect 7455 21342 7523 21398
rect 7579 21342 7647 21398
rect 7703 21342 7713 21398
rect 7265 21274 7713 21342
rect 7265 21218 7275 21274
rect 7331 21218 7399 21274
rect 7455 21218 7523 21274
rect 7579 21218 7647 21274
rect 7703 21218 7713 21274
rect 7265 21150 7713 21218
rect 7265 21094 7275 21150
rect 7331 21094 7399 21150
rect 7455 21094 7523 21150
rect 7579 21094 7647 21150
rect 7703 21094 7713 21150
rect 7265 21026 7713 21094
rect 7265 20970 7275 21026
rect 7331 20970 7399 21026
rect 7455 20970 7523 21026
rect 7579 20970 7647 21026
rect 7703 20970 7713 21026
rect 7265 20902 7713 20970
rect 7265 20846 7275 20902
rect 7331 20846 7399 20902
rect 7455 20846 7523 20902
rect 7579 20846 7647 20902
rect 7703 20846 7713 20902
rect 7265 20836 7713 20846
rect 9927 23754 10127 23764
rect 9927 23698 9937 23754
rect 9993 23698 10061 23754
rect 10117 23698 10127 23754
rect 9927 23630 10127 23698
rect 9927 23574 9937 23630
rect 9993 23574 10061 23630
rect 10117 23574 10127 23630
rect 9927 23506 10127 23574
rect 9927 23450 9937 23506
rect 9993 23450 10061 23506
rect 10117 23450 10127 23506
rect 9927 23382 10127 23450
rect 9927 23326 9937 23382
rect 9993 23326 10061 23382
rect 10117 23326 10127 23382
rect 9927 23258 10127 23326
rect 9927 23202 9937 23258
rect 9993 23202 10061 23258
rect 10117 23202 10127 23258
rect 9927 23134 10127 23202
rect 9927 23078 9937 23134
rect 9993 23078 10061 23134
rect 10117 23078 10127 23134
rect 9927 23010 10127 23078
rect 9927 22954 9937 23010
rect 9993 22954 10061 23010
rect 10117 22954 10127 23010
rect 9927 22886 10127 22954
rect 9927 22830 9937 22886
rect 9993 22830 10061 22886
rect 10117 22830 10127 22886
rect 9927 22762 10127 22830
rect 9927 22706 9937 22762
rect 9993 22706 10061 22762
rect 10117 22706 10127 22762
rect 9927 22638 10127 22706
rect 9927 22582 9937 22638
rect 9993 22582 10061 22638
rect 10117 22582 10127 22638
rect 9927 22514 10127 22582
rect 9927 22458 9937 22514
rect 9993 22458 10061 22514
rect 10117 22458 10127 22514
rect 9927 22390 10127 22458
rect 9927 22334 9937 22390
rect 9993 22334 10061 22390
rect 10117 22334 10127 22390
rect 9927 22266 10127 22334
rect 9927 22210 9937 22266
rect 9993 22210 10061 22266
rect 10117 22210 10127 22266
rect 9927 22142 10127 22210
rect 9927 22086 9937 22142
rect 9993 22086 10061 22142
rect 10117 22086 10127 22142
rect 9927 22018 10127 22086
rect 9927 21962 9937 22018
rect 9993 21962 10061 22018
rect 10117 21962 10127 22018
rect 9927 21894 10127 21962
rect 9927 21838 9937 21894
rect 9993 21838 10061 21894
rect 10117 21838 10127 21894
rect 9927 21770 10127 21838
rect 9927 21714 9937 21770
rect 9993 21714 10061 21770
rect 10117 21714 10127 21770
rect 9927 21646 10127 21714
rect 9927 21590 9937 21646
rect 9993 21590 10061 21646
rect 10117 21590 10127 21646
rect 9927 21522 10127 21590
rect 9927 21466 9937 21522
rect 9993 21466 10061 21522
rect 10117 21466 10127 21522
rect 9927 21398 10127 21466
rect 9927 21342 9937 21398
rect 9993 21342 10061 21398
rect 10117 21342 10127 21398
rect 9927 21274 10127 21342
rect 9927 21218 9937 21274
rect 9993 21218 10061 21274
rect 10117 21218 10127 21274
rect 9927 21150 10127 21218
rect 9927 21094 9937 21150
rect 9993 21094 10061 21150
rect 10117 21094 10127 21150
rect 9927 21026 10127 21094
rect 9927 20970 9937 21026
rect 9993 20970 10061 21026
rect 10117 20970 10127 21026
rect 9927 20902 10127 20970
rect 9927 20846 9937 20902
rect 9993 20846 10061 20902
rect 10117 20846 10127 20902
rect 9927 20836 10127 20846
rect 12297 23754 12497 23764
rect 12297 23698 12307 23754
rect 12363 23698 12431 23754
rect 12487 23698 12497 23754
rect 12297 23630 12497 23698
rect 12297 23574 12307 23630
rect 12363 23574 12431 23630
rect 12487 23574 12497 23630
rect 12297 23506 12497 23574
rect 12297 23450 12307 23506
rect 12363 23450 12431 23506
rect 12487 23450 12497 23506
rect 12297 23382 12497 23450
rect 12297 23326 12307 23382
rect 12363 23326 12431 23382
rect 12487 23326 12497 23382
rect 12297 23258 12497 23326
rect 12297 23202 12307 23258
rect 12363 23202 12431 23258
rect 12487 23202 12497 23258
rect 12297 23134 12497 23202
rect 12297 23078 12307 23134
rect 12363 23078 12431 23134
rect 12487 23078 12497 23134
rect 12297 23010 12497 23078
rect 12297 22954 12307 23010
rect 12363 22954 12431 23010
rect 12487 22954 12497 23010
rect 12297 22886 12497 22954
rect 12297 22830 12307 22886
rect 12363 22830 12431 22886
rect 12487 22830 12497 22886
rect 12297 22762 12497 22830
rect 12297 22706 12307 22762
rect 12363 22706 12431 22762
rect 12487 22706 12497 22762
rect 12297 22638 12497 22706
rect 12297 22582 12307 22638
rect 12363 22582 12431 22638
rect 12487 22582 12497 22638
rect 12297 22514 12497 22582
rect 12297 22458 12307 22514
rect 12363 22458 12431 22514
rect 12487 22458 12497 22514
rect 12297 22390 12497 22458
rect 12297 22334 12307 22390
rect 12363 22334 12431 22390
rect 12487 22334 12497 22390
rect 12297 22266 12497 22334
rect 12297 22210 12307 22266
rect 12363 22210 12431 22266
rect 12487 22210 12497 22266
rect 12297 22142 12497 22210
rect 12297 22086 12307 22142
rect 12363 22086 12431 22142
rect 12487 22086 12497 22142
rect 12297 22018 12497 22086
rect 12297 21962 12307 22018
rect 12363 21962 12431 22018
rect 12487 21962 12497 22018
rect 12297 21894 12497 21962
rect 12297 21838 12307 21894
rect 12363 21838 12431 21894
rect 12487 21838 12497 21894
rect 12297 21770 12497 21838
rect 12297 21714 12307 21770
rect 12363 21714 12431 21770
rect 12487 21714 12497 21770
rect 12297 21646 12497 21714
rect 12297 21590 12307 21646
rect 12363 21590 12431 21646
rect 12487 21590 12497 21646
rect 12297 21522 12497 21590
rect 12297 21466 12307 21522
rect 12363 21466 12431 21522
rect 12487 21466 12497 21522
rect 12297 21398 12497 21466
rect 12297 21342 12307 21398
rect 12363 21342 12431 21398
rect 12487 21342 12497 21398
rect 12297 21274 12497 21342
rect 12297 21218 12307 21274
rect 12363 21218 12431 21274
rect 12487 21218 12497 21274
rect 12297 21150 12497 21218
rect 12297 21094 12307 21150
rect 12363 21094 12431 21150
rect 12487 21094 12497 21150
rect 12297 21026 12497 21094
rect 12297 20970 12307 21026
rect 12363 20970 12431 21026
rect 12487 20970 12497 21026
rect 12297 20902 12497 20970
rect 12297 20846 12307 20902
rect 12363 20846 12431 20902
rect 12487 20846 12497 20902
rect 12297 20836 12497 20846
rect 2481 20554 2681 20564
rect 2481 20498 2491 20554
rect 2547 20498 2615 20554
rect 2671 20498 2681 20554
rect 2481 20430 2681 20498
rect 2481 20374 2491 20430
rect 2547 20374 2615 20430
rect 2671 20374 2681 20430
rect 2481 20306 2681 20374
rect 2481 20250 2491 20306
rect 2547 20250 2615 20306
rect 2671 20250 2681 20306
rect 2481 20182 2681 20250
rect 2481 20126 2491 20182
rect 2547 20126 2615 20182
rect 2671 20126 2681 20182
rect 2481 20058 2681 20126
rect 2481 20002 2491 20058
rect 2547 20002 2615 20058
rect 2671 20002 2681 20058
rect 2481 19934 2681 20002
rect 2481 19878 2491 19934
rect 2547 19878 2615 19934
rect 2671 19878 2681 19934
rect 2481 19810 2681 19878
rect 2481 19754 2491 19810
rect 2547 19754 2615 19810
rect 2671 19754 2681 19810
rect 2481 19686 2681 19754
rect 2481 19630 2491 19686
rect 2547 19630 2615 19686
rect 2671 19630 2681 19686
rect 2481 19562 2681 19630
rect 2481 19506 2491 19562
rect 2547 19506 2615 19562
rect 2671 19506 2681 19562
rect 2481 19438 2681 19506
rect 2481 19382 2491 19438
rect 2547 19382 2615 19438
rect 2671 19382 2681 19438
rect 2481 19314 2681 19382
rect 2481 19258 2491 19314
rect 2547 19258 2615 19314
rect 2671 19258 2681 19314
rect 2481 19190 2681 19258
rect 2481 19134 2491 19190
rect 2547 19134 2615 19190
rect 2671 19134 2681 19190
rect 2481 19066 2681 19134
rect 2481 19010 2491 19066
rect 2547 19010 2615 19066
rect 2671 19010 2681 19066
rect 2481 18942 2681 19010
rect 2481 18886 2491 18942
rect 2547 18886 2615 18942
rect 2671 18886 2681 18942
rect 2481 18818 2681 18886
rect 2481 18762 2491 18818
rect 2547 18762 2615 18818
rect 2671 18762 2681 18818
rect 2481 18694 2681 18762
rect 2481 18638 2491 18694
rect 2547 18638 2615 18694
rect 2671 18638 2681 18694
rect 2481 18570 2681 18638
rect 2481 18514 2491 18570
rect 2547 18514 2615 18570
rect 2671 18514 2681 18570
rect 2481 18446 2681 18514
rect 2481 18390 2491 18446
rect 2547 18390 2615 18446
rect 2671 18390 2681 18446
rect 2481 18322 2681 18390
rect 2481 18266 2491 18322
rect 2547 18266 2615 18322
rect 2671 18266 2681 18322
rect 2481 18198 2681 18266
rect 2481 18142 2491 18198
rect 2547 18142 2615 18198
rect 2671 18142 2681 18198
rect 2481 18074 2681 18142
rect 2481 18018 2491 18074
rect 2547 18018 2615 18074
rect 2671 18018 2681 18074
rect 2481 17950 2681 18018
rect 2481 17894 2491 17950
rect 2547 17894 2615 17950
rect 2671 17894 2681 17950
rect 2481 17826 2681 17894
rect 2481 17770 2491 17826
rect 2547 17770 2615 17826
rect 2671 17770 2681 17826
rect 2481 17702 2681 17770
rect 2481 17646 2491 17702
rect 2547 17646 2615 17702
rect 2671 17646 2681 17702
rect 2481 17636 2681 17646
rect 4851 20554 5051 20564
rect 4851 20498 4861 20554
rect 4917 20498 4985 20554
rect 5041 20498 5051 20554
rect 4851 20430 5051 20498
rect 4851 20374 4861 20430
rect 4917 20374 4985 20430
rect 5041 20374 5051 20430
rect 4851 20306 5051 20374
rect 4851 20250 4861 20306
rect 4917 20250 4985 20306
rect 5041 20250 5051 20306
rect 4851 20182 5051 20250
rect 4851 20126 4861 20182
rect 4917 20126 4985 20182
rect 5041 20126 5051 20182
rect 4851 20058 5051 20126
rect 4851 20002 4861 20058
rect 4917 20002 4985 20058
rect 5041 20002 5051 20058
rect 4851 19934 5051 20002
rect 4851 19878 4861 19934
rect 4917 19878 4985 19934
rect 5041 19878 5051 19934
rect 4851 19810 5051 19878
rect 4851 19754 4861 19810
rect 4917 19754 4985 19810
rect 5041 19754 5051 19810
rect 4851 19686 5051 19754
rect 4851 19630 4861 19686
rect 4917 19630 4985 19686
rect 5041 19630 5051 19686
rect 4851 19562 5051 19630
rect 4851 19506 4861 19562
rect 4917 19506 4985 19562
rect 5041 19506 5051 19562
rect 4851 19438 5051 19506
rect 4851 19382 4861 19438
rect 4917 19382 4985 19438
rect 5041 19382 5051 19438
rect 4851 19314 5051 19382
rect 4851 19258 4861 19314
rect 4917 19258 4985 19314
rect 5041 19258 5051 19314
rect 4851 19190 5051 19258
rect 4851 19134 4861 19190
rect 4917 19134 4985 19190
rect 5041 19134 5051 19190
rect 4851 19066 5051 19134
rect 4851 19010 4861 19066
rect 4917 19010 4985 19066
rect 5041 19010 5051 19066
rect 4851 18942 5051 19010
rect 4851 18886 4861 18942
rect 4917 18886 4985 18942
rect 5041 18886 5051 18942
rect 4851 18818 5051 18886
rect 4851 18762 4861 18818
rect 4917 18762 4985 18818
rect 5041 18762 5051 18818
rect 4851 18694 5051 18762
rect 4851 18638 4861 18694
rect 4917 18638 4985 18694
rect 5041 18638 5051 18694
rect 4851 18570 5051 18638
rect 4851 18514 4861 18570
rect 4917 18514 4985 18570
rect 5041 18514 5051 18570
rect 4851 18446 5051 18514
rect 4851 18390 4861 18446
rect 4917 18390 4985 18446
rect 5041 18390 5051 18446
rect 4851 18322 5051 18390
rect 4851 18266 4861 18322
rect 4917 18266 4985 18322
rect 5041 18266 5051 18322
rect 4851 18198 5051 18266
rect 4851 18142 4861 18198
rect 4917 18142 4985 18198
rect 5041 18142 5051 18198
rect 4851 18074 5051 18142
rect 4851 18018 4861 18074
rect 4917 18018 4985 18074
rect 5041 18018 5051 18074
rect 4851 17950 5051 18018
rect 4851 17894 4861 17950
rect 4917 17894 4985 17950
rect 5041 17894 5051 17950
rect 4851 17826 5051 17894
rect 4851 17770 4861 17826
rect 4917 17770 4985 17826
rect 5041 17770 5051 17826
rect 4851 17702 5051 17770
rect 4851 17646 4861 17702
rect 4917 17646 4985 17702
rect 5041 17646 5051 17702
rect 4851 17636 5051 17646
rect 7265 20554 7713 20564
rect 7265 20498 7275 20554
rect 7331 20498 7399 20554
rect 7455 20498 7523 20554
rect 7579 20498 7647 20554
rect 7703 20498 7713 20554
rect 7265 20430 7713 20498
rect 7265 20374 7275 20430
rect 7331 20374 7399 20430
rect 7455 20374 7523 20430
rect 7579 20374 7647 20430
rect 7703 20374 7713 20430
rect 7265 20306 7713 20374
rect 7265 20250 7275 20306
rect 7331 20250 7399 20306
rect 7455 20250 7523 20306
rect 7579 20250 7647 20306
rect 7703 20250 7713 20306
rect 7265 20182 7713 20250
rect 7265 20126 7275 20182
rect 7331 20126 7399 20182
rect 7455 20126 7523 20182
rect 7579 20126 7647 20182
rect 7703 20126 7713 20182
rect 7265 20058 7713 20126
rect 7265 20002 7275 20058
rect 7331 20002 7399 20058
rect 7455 20002 7523 20058
rect 7579 20002 7647 20058
rect 7703 20002 7713 20058
rect 7265 19934 7713 20002
rect 7265 19878 7275 19934
rect 7331 19878 7399 19934
rect 7455 19878 7523 19934
rect 7579 19878 7647 19934
rect 7703 19878 7713 19934
rect 7265 19810 7713 19878
rect 7265 19754 7275 19810
rect 7331 19754 7399 19810
rect 7455 19754 7523 19810
rect 7579 19754 7647 19810
rect 7703 19754 7713 19810
rect 7265 19686 7713 19754
rect 7265 19630 7275 19686
rect 7331 19630 7399 19686
rect 7455 19630 7523 19686
rect 7579 19630 7647 19686
rect 7703 19630 7713 19686
rect 7265 19562 7713 19630
rect 7265 19506 7275 19562
rect 7331 19506 7399 19562
rect 7455 19506 7523 19562
rect 7579 19506 7647 19562
rect 7703 19506 7713 19562
rect 7265 19438 7713 19506
rect 7265 19382 7275 19438
rect 7331 19382 7399 19438
rect 7455 19382 7523 19438
rect 7579 19382 7647 19438
rect 7703 19382 7713 19438
rect 7265 19314 7713 19382
rect 7265 19258 7275 19314
rect 7331 19258 7399 19314
rect 7455 19258 7523 19314
rect 7579 19258 7647 19314
rect 7703 19258 7713 19314
rect 7265 19190 7713 19258
rect 7265 19134 7275 19190
rect 7331 19134 7399 19190
rect 7455 19134 7523 19190
rect 7579 19134 7647 19190
rect 7703 19134 7713 19190
rect 7265 19066 7713 19134
rect 7265 19010 7275 19066
rect 7331 19010 7399 19066
rect 7455 19010 7523 19066
rect 7579 19010 7647 19066
rect 7703 19010 7713 19066
rect 7265 18942 7713 19010
rect 7265 18886 7275 18942
rect 7331 18886 7399 18942
rect 7455 18886 7523 18942
rect 7579 18886 7647 18942
rect 7703 18886 7713 18942
rect 7265 18818 7713 18886
rect 7265 18762 7275 18818
rect 7331 18762 7399 18818
rect 7455 18762 7523 18818
rect 7579 18762 7647 18818
rect 7703 18762 7713 18818
rect 7265 18694 7713 18762
rect 7265 18638 7275 18694
rect 7331 18638 7399 18694
rect 7455 18638 7523 18694
rect 7579 18638 7647 18694
rect 7703 18638 7713 18694
rect 7265 18570 7713 18638
rect 7265 18514 7275 18570
rect 7331 18514 7399 18570
rect 7455 18514 7523 18570
rect 7579 18514 7647 18570
rect 7703 18514 7713 18570
rect 7265 18446 7713 18514
rect 7265 18390 7275 18446
rect 7331 18390 7399 18446
rect 7455 18390 7523 18446
rect 7579 18390 7647 18446
rect 7703 18390 7713 18446
rect 7265 18322 7713 18390
rect 7265 18266 7275 18322
rect 7331 18266 7399 18322
rect 7455 18266 7523 18322
rect 7579 18266 7647 18322
rect 7703 18266 7713 18322
rect 7265 18198 7713 18266
rect 7265 18142 7275 18198
rect 7331 18142 7399 18198
rect 7455 18142 7523 18198
rect 7579 18142 7647 18198
rect 7703 18142 7713 18198
rect 7265 18074 7713 18142
rect 7265 18018 7275 18074
rect 7331 18018 7399 18074
rect 7455 18018 7523 18074
rect 7579 18018 7647 18074
rect 7703 18018 7713 18074
rect 7265 17950 7713 18018
rect 7265 17894 7275 17950
rect 7331 17894 7399 17950
rect 7455 17894 7523 17950
rect 7579 17894 7647 17950
rect 7703 17894 7713 17950
rect 7265 17826 7713 17894
rect 7265 17770 7275 17826
rect 7331 17770 7399 17826
rect 7455 17770 7523 17826
rect 7579 17770 7647 17826
rect 7703 17770 7713 17826
rect 7265 17702 7713 17770
rect 7265 17646 7275 17702
rect 7331 17646 7399 17702
rect 7455 17646 7523 17702
rect 7579 17646 7647 17702
rect 7703 17646 7713 17702
rect 7265 17636 7713 17646
rect 9927 20554 10127 20564
rect 9927 20498 9937 20554
rect 9993 20498 10061 20554
rect 10117 20498 10127 20554
rect 9927 20430 10127 20498
rect 9927 20374 9937 20430
rect 9993 20374 10061 20430
rect 10117 20374 10127 20430
rect 9927 20306 10127 20374
rect 9927 20250 9937 20306
rect 9993 20250 10061 20306
rect 10117 20250 10127 20306
rect 9927 20182 10127 20250
rect 9927 20126 9937 20182
rect 9993 20126 10061 20182
rect 10117 20126 10127 20182
rect 9927 20058 10127 20126
rect 9927 20002 9937 20058
rect 9993 20002 10061 20058
rect 10117 20002 10127 20058
rect 9927 19934 10127 20002
rect 9927 19878 9937 19934
rect 9993 19878 10061 19934
rect 10117 19878 10127 19934
rect 9927 19810 10127 19878
rect 9927 19754 9937 19810
rect 9993 19754 10061 19810
rect 10117 19754 10127 19810
rect 9927 19686 10127 19754
rect 9927 19630 9937 19686
rect 9993 19630 10061 19686
rect 10117 19630 10127 19686
rect 9927 19562 10127 19630
rect 9927 19506 9937 19562
rect 9993 19506 10061 19562
rect 10117 19506 10127 19562
rect 9927 19438 10127 19506
rect 9927 19382 9937 19438
rect 9993 19382 10061 19438
rect 10117 19382 10127 19438
rect 9927 19314 10127 19382
rect 9927 19258 9937 19314
rect 9993 19258 10061 19314
rect 10117 19258 10127 19314
rect 9927 19190 10127 19258
rect 9927 19134 9937 19190
rect 9993 19134 10061 19190
rect 10117 19134 10127 19190
rect 9927 19066 10127 19134
rect 9927 19010 9937 19066
rect 9993 19010 10061 19066
rect 10117 19010 10127 19066
rect 9927 18942 10127 19010
rect 9927 18886 9937 18942
rect 9993 18886 10061 18942
rect 10117 18886 10127 18942
rect 9927 18818 10127 18886
rect 9927 18762 9937 18818
rect 9993 18762 10061 18818
rect 10117 18762 10127 18818
rect 9927 18694 10127 18762
rect 9927 18638 9937 18694
rect 9993 18638 10061 18694
rect 10117 18638 10127 18694
rect 9927 18570 10127 18638
rect 9927 18514 9937 18570
rect 9993 18514 10061 18570
rect 10117 18514 10127 18570
rect 9927 18446 10127 18514
rect 9927 18390 9937 18446
rect 9993 18390 10061 18446
rect 10117 18390 10127 18446
rect 9927 18322 10127 18390
rect 9927 18266 9937 18322
rect 9993 18266 10061 18322
rect 10117 18266 10127 18322
rect 9927 18198 10127 18266
rect 9927 18142 9937 18198
rect 9993 18142 10061 18198
rect 10117 18142 10127 18198
rect 9927 18074 10127 18142
rect 9927 18018 9937 18074
rect 9993 18018 10061 18074
rect 10117 18018 10127 18074
rect 9927 17950 10127 18018
rect 9927 17894 9937 17950
rect 9993 17894 10061 17950
rect 10117 17894 10127 17950
rect 9927 17826 10127 17894
rect 9927 17770 9937 17826
rect 9993 17770 10061 17826
rect 10117 17770 10127 17826
rect 9927 17702 10127 17770
rect 9927 17646 9937 17702
rect 9993 17646 10061 17702
rect 10117 17646 10127 17702
rect 9927 17636 10127 17646
rect 12297 20554 12497 20564
rect 12297 20498 12307 20554
rect 12363 20498 12431 20554
rect 12487 20498 12497 20554
rect 12297 20430 12497 20498
rect 12297 20374 12307 20430
rect 12363 20374 12431 20430
rect 12487 20374 12497 20430
rect 12297 20306 12497 20374
rect 12297 20250 12307 20306
rect 12363 20250 12431 20306
rect 12487 20250 12497 20306
rect 12297 20182 12497 20250
rect 12297 20126 12307 20182
rect 12363 20126 12431 20182
rect 12487 20126 12497 20182
rect 12297 20058 12497 20126
rect 12297 20002 12307 20058
rect 12363 20002 12431 20058
rect 12487 20002 12497 20058
rect 12297 19934 12497 20002
rect 12297 19878 12307 19934
rect 12363 19878 12431 19934
rect 12487 19878 12497 19934
rect 12297 19810 12497 19878
rect 12297 19754 12307 19810
rect 12363 19754 12431 19810
rect 12487 19754 12497 19810
rect 12297 19686 12497 19754
rect 12297 19630 12307 19686
rect 12363 19630 12431 19686
rect 12487 19630 12497 19686
rect 12297 19562 12497 19630
rect 12297 19506 12307 19562
rect 12363 19506 12431 19562
rect 12487 19506 12497 19562
rect 12297 19438 12497 19506
rect 12297 19382 12307 19438
rect 12363 19382 12431 19438
rect 12487 19382 12497 19438
rect 12297 19314 12497 19382
rect 12297 19258 12307 19314
rect 12363 19258 12431 19314
rect 12487 19258 12497 19314
rect 12297 19190 12497 19258
rect 12297 19134 12307 19190
rect 12363 19134 12431 19190
rect 12487 19134 12497 19190
rect 12297 19066 12497 19134
rect 12297 19010 12307 19066
rect 12363 19010 12431 19066
rect 12487 19010 12497 19066
rect 12297 18942 12497 19010
rect 12297 18886 12307 18942
rect 12363 18886 12431 18942
rect 12487 18886 12497 18942
rect 12297 18818 12497 18886
rect 12297 18762 12307 18818
rect 12363 18762 12431 18818
rect 12487 18762 12497 18818
rect 12297 18694 12497 18762
rect 12297 18638 12307 18694
rect 12363 18638 12431 18694
rect 12487 18638 12497 18694
rect 12297 18570 12497 18638
rect 12297 18514 12307 18570
rect 12363 18514 12431 18570
rect 12487 18514 12497 18570
rect 12297 18446 12497 18514
rect 12297 18390 12307 18446
rect 12363 18390 12431 18446
rect 12487 18390 12497 18446
rect 12297 18322 12497 18390
rect 12297 18266 12307 18322
rect 12363 18266 12431 18322
rect 12487 18266 12497 18322
rect 12297 18198 12497 18266
rect 12297 18142 12307 18198
rect 12363 18142 12431 18198
rect 12487 18142 12497 18198
rect 12297 18074 12497 18142
rect 12297 18018 12307 18074
rect 12363 18018 12431 18074
rect 12487 18018 12497 18074
rect 12297 17950 12497 18018
rect 12297 17894 12307 17950
rect 12363 17894 12431 17950
rect 12487 17894 12497 17950
rect 12297 17826 12497 17894
rect 12297 17770 12307 17826
rect 12363 17770 12431 17826
rect 12487 17770 12497 17826
rect 12297 17702 12497 17770
rect 12297 17646 12307 17702
rect 12363 17646 12431 17702
rect 12487 17646 12497 17702
rect 12297 17636 12497 17646
rect 2481 17354 2681 17364
rect 2481 17298 2491 17354
rect 2547 17298 2615 17354
rect 2671 17298 2681 17354
rect 2481 17230 2681 17298
rect 2481 17174 2491 17230
rect 2547 17174 2615 17230
rect 2671 17174 2681 17230
rect 2481 17106 2681 17174
rect 2481 17050 2491 17106
rect 2547 17050 2615 17106
rect 2671 17050 2681 17106
rect 2481 16982 2681 17050
rect 2481 16926 2491 16982
rect 2547 16926 2615 16982
rect 2671 16926 2681 16982
rect 2481 16858 2681 16926
rect 2481 16802 2491 16858
rect 2547 16802 2615 16858
rect 2671 16802 2681 16858
rect 2481 16734 2681 16802
rect 2481 16678 2491 16734
rect 2547 16678 2615 16734
rect 2671 16678 2681 16734
rect 2481 16610 2681 16678
rect 2481 16554 2491 16610
rect 2547 16554 2615 16610
rect 2671 16554 2681 16610
rect 2481 16486 2681 16554
rect 2481 16430 2491 16486
rect 2547 16430 2615 16486
rect 2671 16430 2681 16486
rect 2481 16362 2681 16430
rect 2481 16306 2491 16362
rect 2547 16306 2615 16362
rect 2671 16306 2681 16362
rect 2481 16238 2681 16306
rect 2481 16182 2491 16238
rect 2547 16182 2615 16238
rect 2671 16182 2681 16238
rect 2481 16114 2681 16182
rect 2481 16058 2491 16114
rect 2547 16058 2615 16114
rect 2671 16058 2681 16114
rect 2481 15990 2681 16058
rect 2481 15934 2491 15990
rect 2547 15934 2615 15990
rect 2671 15934 2681 15990
rect 2481 15866 2681 15934
rect 2481 15810 2491 15866
rect 2547 15810 2615 15866
rect 2671 15810 2681 15866
rect 2481 15742 2681 15810
rect 2481 15686 2491 15742
rect 2547 15686 2615 15742
rect 2671 15686 2681 15742
rect 2481 15618 2681 15686
rect 2481 15562 2491 15618
rect 2547 15562 2615 15618
rect 2671 15562 2681 15618
rect 2481 15494 2681 15562
rect 2481 15438 2491 15494
rect 2547 15438 2615 15494
rect 2671 15438 2681 15494
rect 2481 15370 2681 15438
rect 2481 15314 2491 15370
rect 2547 15314 2615 15370
rect 2671 15314 2681 15370
rect 2481 15246 2681 15314
rect 2481 15190 2491 15246
rect 2547 15190 2615 15246
rect 2671 15190 2681 15246
rect 2481 15122 2681 15190
rect 2481 15066 2491 15122
rect 2547 15066 2615 15122
rect 2671 15066 2681 15122
rect 2481 14998 2681 15066
rect 2481 14942 2491 14998
rect 2547 14942 2615 14998
rect 2671 14942 2681 14998
rect 2481 14874 2681 14942
rect 2481 14818 2491 14874
rect 2547 14818 2615 14874
rect 2671 14818 2681 14874
rect 2481 14750 2681 14818
rect 2481 14694 2491 14750
rect 2547 14694 2615 14750
rect 2671 14694 2681 14750
rect 2481 14626 2681 14694
rect 2481 14570 2491 14626
rect 2547 14570 2615 14626
rect 2671 14570 2681 14626
rect 2481 14502 2681 14570
rect 2481 14446 2491 14502
rect 2547 14446 2615 14502
rect 2671 14446 2681 14502
rect 2481 14436 2681 14446
rect 4851 17354 5051 17364
rect 4851 17298 4861 17354
rect 4917 17298 4985 17354
rect 5041 17298 5051 17354
rect 4851 17230 5051 17298
rect 4851 17174 4861 17230
rect 4917 17174 4985 17230
rect 5041 17174 5051 17230
rect 4851 17106 5051 17174
rect 4851 17050 4861 17106
rect 4917 17050 4985 17106
rect 5041 17050 5051 17106
rect 4851 16982 5051 17050
rect 4851 16926 4861 16982
rect 4917 16926 4985 16982
rect 5041 16926 5051 16982
rect 4851 16858 5051 16926
rect 4851 16802 4861 16858
rect 4917 16802 4985 16858
rect 5041 16802 5051 16858
rect 4851 16734 5051 16802
rect 4851 16678 4861 16734
rect 4917 16678 4985 16734
rect 5041 16678 5051 16734
rect 4851 16610 5051 16678
rect 4851 16554 4861 16610
rect 4917 16554 4985 16610
rect 5041 16554 5051 16610
rect 4851 16486 5051 16554
rect 4851 16430 4861 16486
rect 4917 16430 4985 16486
rect 5041 16430 5051 16486
rect 4851 16362 5051 16430
rect 4851 16306 4861 16362
rect 4917 16306 4985 16362
rect 5041 16306 5051 16362
rect 4851 16238 5051 16306
rect 4851 16182 4861 16238
rect 4917 16182 4985 16238
rect 5041 16182 5051 16238
rect 4851 16114 5051 16182
rect 4851 16058 4861 16114
rect 4917 16058 4985 16114
rect 5041 16058 5051 16114
rect 4851 15990 5051 16058
rect 4851 15934 4861 15990
rect 4917 15934 4985 15990
rect 5041 15934 5051 15990
rect 4851 15866 5051 15934
rect 4851 15810 4861 15866
rect 4917 15810 4985 15866
rect 5041 15810 5051 15866
rect 4851 15742 5051 15810
rect 4851 15686 4861 15742
rect 4917 15686 4985 15742
rect 5041 15686 5051 15742
rect 4851 15618 5051 15686
rect 4851 15562 4861 15618
rect 4917 15562 4985 15618
rect 5041 15562 5051 15618
rect 4851 15494 5051 15562
rect 4851 15438 4861 15494
rect 4917 15438 4985 15494
rect 5041 15438 5051 15494
rect 4851 15370 5051 15438
rect 4851 15314 4861 15370
rect 4917 15314 4985 15370
rect 5041 15314 5051 15370
rect 4851 15246 5051 15314
rect 4851 15190 4861 15246
rect 4917 15190 4985 15246
rect 5041 15190 5051 15246
rect 4851 15122 5051 15190
rect 4851 15066 4861 15122
rect 4917 15066 4985 15122
rect 5041 15066 5051 15122
rect 4851 14998 5051 15066
rect 4851 14942 4861 14998
rect 4917 14942 4985 14998
rect 5041 14942 5051 14998
rect 4851 14874 5051 14942
rect 4851 14818 4861 14874
rect 4917 14818 4985 14874
rect 5041 14818 5051 14874
rect 4851 14750 5051 14818
rect 4851 14694 4861 14750
rect 4917 14694 4985 14750
rect 5041 14694 5051 14750
rect 4851 14626 5051 14694
rect 4851 14570 4861 14626
rect 4917 14570 4985 14626
rect 5041 14570 5051 14626
rect 4851 14502 5051 14570
rect 4851 14446 4861 14502
rect 4917 14446 4985 14502
rect 5041 14446 5051 14502
rect 4851 14436 5051 14446
rect 7265 17354 7713 17364
rect 7265 17298 7275 17354
rect 7331 17298 7399 17354
rect 7455 17298 7523 17354
rect 7579 17298 7647 17354
rect 7703 17298 7713 17354
rect 7265 17230 7713 17298
rect 7265 17174 7275 17230
rect 7331 17174 7399 17230
rect 7455 17174 7523 17230
rect 7579 17174 7647 17230
rect 7703 17174 7713 17230
rect 7265 17106 7713 17174
rect 7265 17050 7275 17106
rect 7331 17050 7399 17106
rect 7455 17050 7523 17106
rect 7579 17050 7647 17106
rect 7703 17050 7713 17106
rect 7265 16982 7713 17050
rect 7265 16926 7275 16982
rect 7331 16926 7399 16982
rect 7455 16926 7523 16982
rect 7579 16926 7647 16982
rect 7703 16926 7713 16982
rect 7265 16858 7713 16926
rect 7265 16802 7275 16858
rect 7331 16802 7399 16858
rect 7455 16802 7523 16858
rect 7579 16802 7647 16858
rect 7703 16802 7713 16858
rect 7265 16734 7713 16802
rect 7265 16678 7275 16734
rect 7331 16678 7399 16734
rect 7455 16678 7523 16734
rect 7579 16678 7647 16734
rect 7703 16678 7713 16734
rect 7265 16610 7713 16678
rect 7265 16554 7275 16610
rect 7331 16554 7399 16610
rect 7455 16554 7523 16610
rect 7579 16554 7647 16610
rect 7703 16554 7713 16610
rect 7265 16486 7713 16554
rect 7265 16430 7275 16486
rect 7331 16430 7399 16486
rect 7455 16430 7523 16486
rect 7579 16430 7647 16486
rect 7703 16430 7713 16486
rect 7265 16362 7713 16430
rect 7265 16306 7275 16362
rect 7331 16306 7399 16362
rect 7455 16306 7523 16362
rect 7579 16306 7647 16362
rect 7703 16306 7713 16362
rect 7265 16238 7713 16306
rect 7265 16182 7275 16238
rect 7331 16182 7399 16238
rect 7455 16182 7523 16238
rect 7579 16182 7647 16238
rect 7703 16182 7713 16238
rect 7265 16114 7713 16182
rect 7265 16058 7275 16114
rect 7331 16058 7399 16114
rect 7455 16058 7523 16114
rect 7579 16058 7647 16114
rect 7703 16058 7713 16114
rect 7265 15990 7713 16058
rect 7265 15934 7275 15990
rect 7331 15934 7399 15990
rect 7455 15934 7523 15990
rect 7579 15934 7647 15990
rect 7703 15934 7713 15990
rect 7265 15866 7713 15934
rect 7265 15810 7275 15866
rect 7331 15810 7399 15866
rect 7455 15810 7523 15866
rect 7579 15810 7647 15866
rect 7703 15810 7713 15866
rect 7265 15742 7713 15810
rect 7265 15686 7275 15742
rect 7331 15686 7399 15742
rect 7455 15686 7523 15742
rect 7579 15686 7647 15742
rect 7703 15686 7713 15742
rect 7265 15618 7713 15686
rect 7265 15562 7275 15618
rect 7331 15562 7399 15618
rect 7455 15562 7523 15618
rect 7579 15562 7647 15618
rect 7703 15562 7713 15618
rect 7265 15494 7713 15562
rect 7265 15438 7275 15494
rect 7331 15438 7399 15494
rect 7455 15438 7523 15494
rect 7579 15438 7647 15494
rect 7703 15438 7713 15494
rect 7265 15370 7713 15438
rect 7265 15314 7275 15370
rect 7331 15314 7399 15370
rect 7455 15314 7523 15370
rect 7579 15314 7647 15370
rect 7703 15314 7713 15370
rect 7265 15246 7713 15314
rect 7265 15190 7275 15246
rect 7331 15190 7399 15246
rect 7455 15190 7523 15246
rect 7579 15190 7647 15246
rect 7703 15190 7713 15246
rect 7265 15122 7713 15190
rect 7265 15066 7275 15122
rect 7331 15066 7399 15122
rect 7455 15066 7523 15122
rect 7579 15066 7647 15122
rect 7703 15066 7713 15122
rect 7265 14998 7713 15066
rect 7265 14942 7275 14998
rect 7331 14942 7399 14998
rect 7455 14942 7523 14998
rect 7579 14942 7647 14998
rect 7703 14942 7713 14998
rect 7265 14874 7713 14942
rect 7265 14818 7275 14874
rect 7331 14818 7399 14874
rect 7455 14818 7523 14874
rect 7579 14818 7647 14874
rect 7703 14818 7713 14874
rect 7265 14750 7713 14818
rect 7265 14694 7275 14750
rect 7331 14694 7399 14750
rect 7455 14694 7523 14750
rect 7579 14694 7647 14750
rect 7703 14694 7713 14750
rect 7265 14626 7713 14694
rect 7265 14570 7275 14626
rect 7331 14570 7399 14626
rect 7455 14570 7523 14626
rect 7579 14570 7647 14626
rect 7703 14570 7713 14626
rect 7265 14502 7713 14570
rect 7265 14446 7275 14502
rect 7331 14446 7399 14502
rect 7455 14446 7523 14502
rect 7579 14446 7647 14502
rect 7703 14446 7713 14502
rect 7265 14436 7713 14446
rect 9927 17354 10127 17364
rect 9927 17298 9937 17354
rect 9993 17298 10061 17354
rect 10117 17298 10127 17354
rect 9927 17230 10127 17298
rect 9927 17174 9937 17230
rect 9993 17174 10061 17230
rect 10117 17174 10127 17230
rect 9927 17106 10127 17174
rect 9927 17050 9937 17106
rect 9993 17050 10061 17106
rect 10117 17050 10127 17106
rect 9927 16982 10127 17050
rect 9927 16926 9937 16982
rect 9993 16926 10061 16982
rect 10117 16926 10127 16982
rect 9927 16858 10127 16926
rect 9927 16802 9937 16858
rect 9993 16802 10061 16858
rect 10117 16802 10127 16858
rect 9927 16734 10127 16802
rect 9927 16678 9937 16734
rect 9993 16678 10061 16734
rect 10117 16678 10127 16734
rect 9927 16610 10127 16678
rect 9927 16554 9937 16610
rect 9993 16554 10061 16610
rect 10117 16554 10127 16610
rect 9927 16486 10127 16554
rect 9927 16430 9937 16486
rect 9993 16430 10061 16486
rect 10117 16430 10127 16486
rect 9927 16362 10127 16430
rect 9927 16306 9937 16362
rect 9993 16306 10061 16362
rect 10117 16306 10127 16362
rect 9927 16238 10127 16306
rect 9927 16182 9937 16238
rect 9993 16182 10061 16238
rect 10117 16182 10127 16238
rect 9927 16114 10127 16182
rect 9927 16058 9937 16114
rect 9993 16058 10061 16114
rect 10117 16058 10127 16114
rect 9927 15990 10127 16058
rect 9927 15934 9937 15990
rect 9993 15934 10061 15990
rect 10117 15934 10127 15990
rect 9927 15866 10127 15934
rect 9927 15810 9937 15866
rect 9993 15810 10061 15866
rect 10117 15810 10127 15866
rect 9927 15742 10127 15810
rect 9927 15686 9937 15742
rect 9993 15686 10061 15742
rect 10117 15686 10127 15742
rect 9927 15618 10127 15686
rect 9927 15562 9937 15618
rect 9993 15562 10061 15618
rect 10117 15562 10127 15618
rect 9927 15494 10127 15562
rect 9927 15438 9937 15494
rect 9993 15438 10061 15494
rect 10117 15438 10127 15494
rect 9927 15370 10127 15438
rect 9927 15314 9937 15370
rect 9993 15314 10061 15370
rect 10117 15314 10127 15370
rect 9927 15246 10127 15314
rect 9927 15190 9937 15246
rect 9993 15190 10061 15246
rect 10117 15190 10127 15246
rect 9927 15122 10127 15190
rect 9927 15066 9937 15122
rect 9993 15066 10061 15122
rect 10117 15066 10127 15122
rect 9927 14998 10127 15066
rect 9927 14942 9937 14998
rect 9993 14942 10061 14998
rect 10117 14942 10127 14998
rect 9927 14874 10127 14942
rect 9927 14818 9937 14874
rect 9993 14818 10061 14874
rect 10117 14818 10127 14874
rect 9927 14750 10127 14818
rect 9927 14694 9937 14750
rect 9993 14694 10061 14750
rect 10117 14694 10127 14750
rect 9927 14626 10127 14694
rect 9927 14570 9937 14626
rect 9993 14570 10061 14626
rect 10117 14570 10127 14626
rect 9927 14502 10127 14570
rect 9927 14446 9937 14502
rect 9993 14446 10061 14502
rect 10117 14446 10127 14502
rect 9927 14436 10127 14446
rect 12297 17354 12497 17364
rect 12297 17298 12307 17354
rect 12363 17298 12431 17354
rect 12487 17298 12497 17354
rect 12297 17230 12497 17298
rect 12297 17174 12307 17230
rect 12363 17174 12431 17230
rect 12487 17174 12497 17230
rect 12297 17106 12497 17174
rect 12297 17050 12307 17106
rect 12363 17050 12431 17106
rect 12487 17050 12497 17106
rect 12297 16982 12497 17050
rect 12297 16926 12307 16982
rect 12363 16926 12431 16982
rect 12487 16926 12497 16982
rect 12297 16858 12497 16926
rect 12297 16802 12307 16858
rect 12363 16802 12431 16858
rect 12487 16802 12497 16858
rect 12297 16734 12497 16802
rect 12297 16678 12307 16734
rect 12363 16678 12431 16734
rect 12487 16678 12497 16734
rect 12297 16610 12497 16678
rect 12297 16554 12307 16610
rect 12363 16554 12431 16610
rect 12487 16554 12497 16610
rect 12297 16486 12497 16554
rect 12297 16430 12307 16486
rect 12363 16430 12431 16486
rect 12487 16430 12497 16486
rect 12297 16362 12497 16430
rect 12297 16306 12307 16362
rect 12363 16306 12431 16362
rect 12487 16306 12497 16362
rect 12297 16238 12497 16306
rect 12297 16182 12307 16238
rect 12363 16182 12431 16238
rect 12487 16182 12497 16238
rect 12297 16114 12497 16182
rect 12297 16058 12307 16114
rect 12363 16058 12431 16114
rect 12487 16058 12497 16114
rect 12297 15990 12497 16058
rect 12297 15934 12307 15990
rect 12363 15934 12431 15990
rect 12487 15934 12497 15990
rect 12297 15866 12497 15934
rect 12297 15810 12307 15866
rect 12363 15810 12431 15866
rect 12487 15810 12497 15866
rect 12297 15742 12497 15810
rect 12297 15686 12307 15742
rect 12363 15686 12431 15742
rect 12487 15686 12497 15742
rect 12297 15618 12497 15686
rect 12297 15562 12307 15618
rect 12363 15562 12431 15618
rect 12487 15562 12497 15618
rect 12297 15494 12497 15562
rect 12297 15438 12307 15494
rect 12363 15438 12431 15494
rect 12487 15438 12497 15494
rect 12297 15370 12497 15438
rect 12297 15314 12307 15370
rect 12363 15314 12431 15370
rect 12487 15314 12497 15370
rect 12297 15246 12497 15314
rect 12297 15190 12307 15246
rect 12363 15190 12431 15246
rect 12487 15190 12497 15246
rect 12297 15122 12497 15190
rect 12297 15066 12307 15122
rect 12363 15066 12431 15122
rect 12487 15066 12497 15122
rect 12297 14998 12497 15066
rect 12297 14942 12307 14998
rect 12363 14942 12431 14998
rect 12487 14942 12497 14998
rect 12297 14874 12497 14942
rect 12297 14818 12307 14874
rect 12363 14818 12431 14874
rect 12487 14818 12497 14874
rect 12297 14750 12497 14818
rect 12297 14694 12307 14750
rect 12363 14694 12431 14750
rect 12487 14694 12497 14750
rect 12297 14626 12497 14694
rect 12297 14570 12307 14626
rect 12363 14570 12431 14626
rect 12487 14570 12497 14626
rect 12297 14502 12497 14570
rect 12297 14446 12307 14502
rect 12363 14446 12431 14502
rect 12487 14446 12497 14502
rect 12297 14436 12497 14446
rect -11 14176 86 14186
rect -11 12824 20 14176
rect 76 12824 86 14176
rect 14892 14176 14989 14186
rect 305 14148 2117 14158
rect 305 14092 315 14148
rect 371 14092 439 14148
rect 495 14092 563 14148
rect 619 14092 687 14148
rect 743 14092 811 14148
rect 867 14092 935 14148
rect 991 14092 1059 14148
rect 1115 14092 1183 14148
rect 1239 14092 1307 14148
rect 1363 14092 1431 14148
rect 1487 14092 1555 14148
rect 1611 14092 1679 14148
rect 1735 14092 1803 14148
rect 1859 14092 1927 14148
rect 1983 14092 2051 14148
rect 2107 14092 2117 14148
rect 305 14024 2117 14092
rect 305 13968 315 14024
rect 371 13968 439 14024
rect 495 13968 563 14024
rect 619 13968 687 14024
rect 743 13968 811 14024
rect 867 13968 935 14024
rect 991 13968 1059 14024
rect 1115 13968 1183 14024
rect 1239 13968 1307 14024
rect 1363 13968 1431 14024
rect 1487 13968 1555 14024
rect 1611 13968 1679 14024
rect 1735 13968 1803 14024
rect 1859 13968 1927 14024
rect 1983 13968 2051 14024
rect 2107 13968 2117 14024
rect 305 13900 2117 13968
rect 305 13844 315 13900
rect 371 13844 439 13900
rect 495 13844 563 13900
rect 619 13844 687 13900
rect 743 13844 811 13900
rect 867 13844 935 13900
rect 991 13844 1059 13900
rect 1115 13844 1183 13900
rect 1239 13844 1307 13900
rect 1363 13844 1431 13900
rect 1487 13844 1555 13900
rect 1611 13844 1679 13900
rect 1735 13844 1803 13900
rect 1859 13844 1927 13900
rect 1983 13844 2051 13900
rect 2107 13844 2117 13900
rect 305 13776 2117 13844
rect 305 13720 315 13776
rect 371 13720 439 13776
rect 495 13720 563 13776
rect 619 13720 687 13776
rect 743 13720 811 13776
rect 867 13720 935 13776
rect 991 13720 1059 13776
rect 1115 13720 1183 13776
rect 1239 13720 1307 13776
rect 1363 13720 1431 13776
rect 1487 13720 1555 13776
rect 1611 13720 1679 13776
rect 1735 13720 1803 13776
rect 1859 13720 1927 13776
rect 1983 13720 2051 13776
rect 2107 13720 2117 13776
rect 305 13652 2117 13720
rect 305 13596 315 13652
rect 371 13596 439 13652
rect 495 13596 563 13652
rect 619 13596 687 13652
rect 743 13596 811 13652
rect 867 13596 935 13652
rect 991 13596 1059 13652
rect 1115 13596 1183 13652
rect 1239 13596 1307 13652
rect 1363 13596 1431 13652
rect 1487 13596 1555 13652
rect 1611 13596 1679 13652
rect 1735 13596 1803 13652
rect 1859 13596 1927 13652
rect 1983 13596 2051 13652
rect 2107 13596 2117 13652
rect 305 13528 2117 13596
rect 305 13472 315 13528
rect 371 13472 439 13528
rect 495 13472 563 13528
rect 619 13472 687 13528
rect 743 13472 811 13528
rect 867 13472 935 13528
rect 991 13472 1059 13528
rect 1115 13472 1183 13528
rect 1239 13472 1307 13528
rect 1363 13472 1431 13528
rect 1487 13472 1555 13528
rect 1611 13472 1679 13528
rect 1735 13472 1803 13528
rect 1859 13472 1927 13528
rect 1983 13472 2051 13528
rect 2107 13472 2117 13528
rect 305 13404 2117 13472
rect 305 13348 315 13404
rect 371 13348 439 13404
rect 495 13348 563 13404
rect 619 13348 687 13404
rect 743 13348 811 13404
rect 867 13348 935 13404
rect 991 13348 1059 13404
rect 1115 13348 1183 13404
rect 1239 13348 1307 13404
rect 1363 13348 1431 13404
rect 1487 13348 1555 13404
rect 1611 13348 1679 13404
rect 1735 13348 1803 13404
rect 1859 13348 1927 13404
rect 1983 13348 2051 13404
rect 2107 13348 2117 13404
rect 305 13280 2117 13348
rect 305 13224 315 13280
rect 371 13224 439 13280
rect 495 13224 563 13280
rect 619 13224 687 13280
rect 743 13224 811 13280
rect 867 13224 935 13280
rect 991 13224 1059 13280
rect 1115 13224 1183 13280
rect 1239 13224 1307 13280
rect 1363 13224 1431 13280
rect 1487 13224 1555 13280
rect 1611 13224 1679 13280
rect 1735 13224 1803 13280
rect 1859 13224 1927 13280
rect 1983 13224 2051 13280
rect 2107 13224 2117 13280
rect 305 13156 2117 13224
rect 305 13100 315 13156
rect 371 13100 439 13156
rect 495 13100 563 13156
rect 619 13100 687 13156
rect 743 13100 811 13156
rect 867 13100 935 13156
rect 991 13100 1059 13156
rect 1115 13100 1183 13156
rect 1239 13100 1307 13156
rect 1363 13100 1431 13156
rect 1487 13100 1555 13156
rect 1611 13100 1679 13156
rect 1735 13100 1803 13156
rect 1859 13100 1927 13156
rect 1983 13100 2051 13156
rect 2107 13100 2117 13156
rect 305 13032 2117 13100
rect 305 12976 315 13032
rect 371 12976 439 13032
rect 495 12976 563 13032
rect 619 12976 687 13032
rect 743 12976 811 13032
rect 867 12976 935 13032
rect 991 12976 1059 13032
rect 1115 12976 1183 13032
rect 1239 12976 1307 13032
rect 1363 12976 1431 13032
rect 1487 12976 1555 13032
rect 1611 12976 1679 13032
rect 1735 12976 1803 13032
rect 1859 12976 1927 13032
rect 1983 12976 2051 13032
rect 2107 12976 2117 13032
rect 305 12908 2117 12976
rect 305 12852 315 12908
rect 371 12852 439 12908
rect 495 12852 563 12908
rect 619 12852 687 12908
rect 743 12852 811 12908
rect 867 12852 935 12908
rect 991 12852 1059 12908
rect 1115 12852 1183 12908
rect 1239 12852 1307 12908
rect 1363 12852 1431 12908
rect 1487 12852 1555 12908
rect 1611 12852 1679 12908
rect 1735 12852 1803 12908
rect 1859 12852 1927 12908
rect 1983 12852 2051 12908
rect 2107 12852 2117 12908
rect 305 12842 2117 12852
rect 2798 14148 4734 14158
rect 2798 14092 2808 14148
rect 2864 14092 2932 14148
rect 2988 14092 3056 14148
rect 3112 14092 3180 14148
rect 3236 14092 3304 14148
rect 3360 14092 3428 14148
rect 3484 14092 3552 14148
rect 3608 14092 3676 14148
rect 3732 14092 3800 14148
rect 3856 14092 3924 14148
rect 3980 14092 4048 14148
rect 4104 14092 4172 14148
rect 4228 14092 4296 14148
rect 4352 14092 4420 14148
rect 4476 14092 4544 14148
rect 4600 14092 4668 14148
rect 4724 14092 4734 14148
rect 2798 14024 4734 14092
rect 2798 13968 2808 14024
rect 2864 13968 2932 14024
rect 2988 13968 3056 14024
rect 3112 13968 3180 14024
rect 3236 13968 3304 14024
rect 3360 13968 3428 14024
rect 3484 13968 3552 14024
rect 3608 13968 3676 14024
rect 3732 13968 3800 14024
rect 3856 13968 3924 14024
rect 3980 13968 4048 14024
rect 4104 13968 4172 14024
rect 4228 13968 4296 14024
rect 4352 13968 4420 14024
rect 4476 13968 4544 14024
rect 4600 13968 4668 14024
rect 4724 13968 4734 14024
rect 2798 13900 4734 13968
rect 2798 13844 2808 13900
rect 2864 13844 2932 13900
rect 2988 13844 3056 13900
rect 3112 13844 3180 13900
rect 3236 13844 3304 13900
rect 3360 13844 3428 13900
rect 3484 13844 3552 13900
rect 3608 13844 3676 13900
rect 3732 13844 3800 13900
rect 3856 13844 3924 13900
rect 3980 13844 4048 13900
rect 4104 13844 4172 13900
rect 4228 13844 4296 13900
rect 4352 13844 4420 13900
rect 4476 13844 4544 13900
rect 4600 13844 4668 13900
rect 4724 13844 4734 13900
rect 2798 13776 4734 13844
rect 2798 13720 2808 13776
rect 2864 13720 2932 13776
rect 2988 13720 3056 13776
rect 3112 13720 3180 13776
rect 3236 13720 3304 13776
rect 3360 13720 3428 13776
rect 3484 13720 3552 13776
rect 3608 13720 3676 13776
rect 3732 13720 3800 13776
rect 3856 13720 3924 13776
rect 3980 13720 4048 13776
rect 4104 13720 4172 13776
rect 4228 13720 4296 13776
rect 4352 13720 4420 13776
rect 4476 13720 4544 13776
rect 4600 13720 4668 13776
rect 4724 13720 4734 13776
rect 2798 13652 4734 13720
rect 2798 13596 2808 13652
rect 2864 13596 2932 13652
rect 2988 13596 3056 13652
rect 3112 13596 3180 13652
rect 3236 13596 3304 13652
rect 3360 13596 3428 13652
rect 3484 13596 3552 13652
rect 3608 13596 3676 13652
rect 3732 13596 3800 13652
rect 3856 13596 3924 13652
rect 3980 13596 4048 13652
rect 4104 13596 4172 13652
rect 4228 13596 4296 13652
rect 4352 13596 4420 13652
rect 4476 13596 4544 13652
rect 4600 13596 4668 13652
rect 4724 13596 4734 13652
rect 2798 13528 4734 13596
rect 2798 13472 2808 13528
rect 2864 13472 2932 13528
rect 2988 13472 3056 13528
rect 3112 13472 3180 13528
rect 3236 13472 3304 13528
rect 3360 13472 3428 13528
rect 3484 13472 3552 13528
rect 3608 13472 3676 13528
rect 3732 13472 3800 13528
rect 3856 13472 3924 13528
rect 3980 13472 4048 13528
rect 4104 13472 4172 13528
rect 4228 13472 4296 13528
rect 4352 13472 4420 13528
rect 4476 13472 4544 13528
rect 4600 13472 4668 13528
rect 4724 13472 4734 13528
rect 2798 13404 4734 13472
rect 2798 13348 2808 13404
rect 2864 13348 2932 13404
rect 2988 13348 3056 13404
rect 3112 13348 3180 13404
rect 3236 13348 3304 13404
rect 3360 13348 3428 13404
rect 3484 13348 3552 13404
rect 3608 13348 3676 13404
rect 3732 13348 3800 13404
rect 3856 13348 3924 13404
rect 3980 13348 4048 13404
rect 4104 13348 4172 13404
rect 4228 13348 4296 13404
rect 4352 13348 4420 13404
rect 4476 13348 4544 13404
rect 4600 13348 4668 13404
rect 4724 13348 4734 13404
rect 2798 13280 4734 13348
rect 2798 13224 2808 13280
rect 2864 13224 2932 13280
rect 2988 13224 3056 13280
rect 3112 13224 3180 13280
rect 3236 13224 3304 13280
rect 3360 13224 3428 13280
rect 3484 13224 3552 13280
rect 3608 13224 3676 13280
rect 3732 13224 3800 13280
rect 3856 13224 3924 13280
rect 3980 13224 4048 13280
rect 4104 13224 4172 13280
rect 4228 13224 4296 13280
rect 4352 13224 4420 13280
rect 4476 13224 4544 13280
rect 4600 13224 4668 13280
rect 4724 13224 4734 13280
rect 2798 13156 4734 13224
rect 2798 13100 2808 13156
rect 2864 13100 2932 13156
rect 2988 13100 3056 13156
rect 3112 13100 3180 13156
rect 3236 13100 3304 13156
rect 3360 13100 3428 13156
rect 3484 13100 3552 13156
rect 3608 13100 3676 13156
rect 3732 13100 3800 13156
rect 3856 13100 3924 13156
rect 3980 13100 4048 13156
rect 4104 13100 4172 13156
rect 4228 13100 4296 13156
rect 4352 13100 4420 13156
rect 4476 13100 4544 13156
rect 4600 13100 4668 13156
rect 4724 13100 4734 13156
rect 2798 13032 4734 13100
rect 2798 12976 2808 13032
rect 2864 12976 2932 13032
rect 2988 12976 3056 13032
rect 3112 12976 3180 13032
rect 3236 12976 3304 13032
rect 3360 12976 3428 13032
rect 3484 12976 3552 13032
rect 3608 12976 3676 13032
rect 3732 12976 3800 13032
rect 3856 12976 3924 13032
rect 3980 12976 4048 13032
rect 4104 12976 4172 13032
rect 4228 12976 4296 13032
rect 4352 12976 4420 13032
rect 4476 12976 4544 13032
rect 4600 12976 4668 13032
rect 4724 12976 4734 13032
rect 2798 12908 4734 12976
rect 2798 12852 2808 12908
rect 2864 12852 2932 12908
rect 2988 12852 3056 12908
rect 3112 12852 3180 12908
rect 3236 12852 3304 12908
rect 3360 12852 3428 12908
rect 3484 12852 3552 12908
rect 3608 12852 3676 12908
rect 3732 12852 3800 12908
rect 3856 12852 3924 12908
rect 3980 12852 4048 12908
rect 4104 12852 4172 12908
rect 4228 12852 4296 12908
rect 4352 12852 4420 12908
rect 4476 12852 4544 12908
rect 4600 12852 4668 12908
rect 4724 12852 4734 12908
rect 2798 12842 4734 12852
rect 5168 14148 7104 14158
rect 5168 14092 5178 14148
rect 5234 14092 5302 14148
rect 5358 14092 5426 14148
rect 5482 14092 5550 14148
rect 5606 14092 5674 14148
rect 5730 14092 5798 14148
rect 5854 14092 5922 14148
rect 5978 14092 6046 14148
rect 6102 14092 6170 14148
rect 6226 14092 6294 14148
rect 6350 14092 6418 14148
rect 6474 14092 6542 14148
rect 6598 14092 6666 14148
rect 6722 14092 6790 14148
rect 6846 14092 6914 14148
rect 6970 14092 7038 14148
rect 7094 14092 7104 14148
rect 5168 14024 7104 14092
rect 5168 13968 5178 14024
rect 5234 13968 5302 14024
rect 5358 13968 5426 14024
rect 5482 13968 5550 14024
rect 5606 13968 5674 14024
rect 5730 13968 5798 14024
rect 5854 13968 5922 14024
rect 5978 13968 6046 14024
rect 6102 13968 6170 14024
rect 6226 13968 6294 14024
rect 6350 13968 6418 14024
rect 6474 13968 6542 14024
rect 6598 13968 6666 14024
rect 6722 13968 6790 14024
rect 6846 13968 6914 14024
rect 6970 13968 7038 14024
rect 7094 13968 7104 14024
rect 5168 13900 7104 13968
rect 5168 13844 5178 13900
rect 5234 13844 5302 13900
rect 5358 13844 5426 13900
rect 5482 13844 5550 13900
rect 5606 13844 5674 13900
rect 5730 13844 5798 13900
rect 5854 13844 5922 13900
rect 5978 13844 6046 13900
rect 6102 13844 6170 13900
rect 6226 13844 6294 13900
rect 6350 13844 6418 13900
rect 6474 13844 6542 13900
rect 6598 13844 6666 13900
rect 6722 13844 6790 13900
rect 6846 13844 6914 13900
rect 6970 13844 7038 13900
rect 7094 13844 7104 13900
rect 5168 13776 7104 13844
rect 5168 13720 5178 13776
rect 5234 13720 5302 13776
rect 5358 13720 5426 13776
rect 5482 13720 5550 13776
rect 5606 13720 5674 13776
rect 5730 13720 5798 13776
rect 5854 13720 5922 13776
rect 5978 13720 6046 13776
rect 6102 13720 6170 13776
rect 6226 13720 6294 13776
rect 6350 13720 6418 13776
rect 6474 13720 6542 13776
rect 6598 13720 6666 13776
rect 6722 13720 6790 13776
rect 6846 13720 6914 13776
rect 6970 13720 7038 13776
rect 7094 13720 7104 13776
rect 5168 13652 7104 13720
rect 5168 13596 5178 13652
rect 5234 13596 5302 13652
rect 5358 13596 5426 13652
rect 5482 13596 5550 13652
rect 5606 13596 5674 13652
rect 5730 13596 5798 13652
rect 5854 13596 5922 13652
rect 5978 13596 6046 13652
rect 6102 13596 6170 13652
rect 6226 13596 6294 13652
rect 6350 13596 6418 13652
rect 6474 13596 6542 13652
rect 6598 13596 6666 13652
rect 6722 13596 6790 13652
rect 6846 13596 6914 13652
rect 6970 13596 7038 13652
rect 7094 13596 7104 13652
rect 5168 13528 7104 13596
rect 5168 13472 5178 13528
rect 5234 13472 5302 13528
rect 5358 13472 5426 13528
rect 5482 13472 5550 13528
rect 5606 13472 5674 13528
rect 5730 13472 5798 13528
rect 5854 13472 5922 13528
rect 5978 13472 6046 13528
rect 6102 13472 6170 13528
rect 6226 13472 6294 13528
rect 6350 13472 6418 13528
rect 6474 13472 6542 13528
rect 6598 13472 6666 13528
rect 6722 13472 6790 13528
rect 6846 13472 6914 13528
rect 6970 13472 7038 13528
rect 7094 13472 7104 13528
rect 5168 13404 7104 13472
rect 5168 13348 5178 13404
rect 5234 13348 5302 13404
rect 5358 13348 5426 13404
rect 5482 13348 5550 13404
rect 5606 13348 5674 13404
rect 5730 13348 5798 13404
rect 5854 13348 5922 13404
rect 5978 13348 6046 13404
rect 6102 13348 6170 13404
rect 6226 13348 6294 13404
rect 6350 13348 6418 13404
rect 6474 13348 6542 13404
rect 6598 13348 6666 13404
rect 6722 13348 6790 13404
rect 6846 13348 6914 13404
rect 6970 13348 7038 13404
rect 7094 13348 7104 13404
rect 5168 13280 7104 13348
rect 5168 13224 5178 13280
rect 5234 13224 5302 13280
rect 5358 13224 5426 13280
rect 5482 13224 5550 13280
rect 5606 13224 5674 13280
rect 5730 13224 5798 13280
rect 5854 13224 5922 13280
rect 5978 13224 6046 13280
rect 6102 13224 6170 13280
rect 6226 13224 6294 13280
rect 6350 13224 6418 13280
rect 6474 13224 6542 13280
rect 6598 13224 6666 13280
rect 6722 13224 6790 13280
rect 6846 13224 6914 13280
rect 6970 13224 7038 13280
rect 7094 13224 7104 13280
rect 5168 13156 7104 13224
rect 5168 13100 5178 13156
rect 5234 13100 5302 13156
rect 5358 13100 5426 13156
rect 5482 13100 5550 13156
rect 5606 13100 5674 13156
rect 5730 13100 5798 13156
rect 5854 13100 5922 13156
rect 5978 13100 6046 13156
rect 6102 13100 6170 13156
rect 6226 13100 6294 13156
rect 6350 13100 6418 13156
rect 6474 13100 6542 13156
rect 6598 13100 6666 13156
rect 6722 13100 6790 13156
rect 6846 13100 6914 13156
rect 6970 13100 7038 13156
rect 7094 13100 7104 13156
rect 5168 13032 7104 13100
rect 5168 12976 5178 13032
rect 5234 12976 5302 13032
rect 5358 12976 5426 13032
rect 5482 12976 5550 13032
rect 5606 12976 5674 13032
rect 5730 12976 5798 13032
rect 5854 12976 5922 13032
rect 5978 12976 6046 13032
rect 6102 12976 6170 13032
rect 6226 12976 6294 13032
rect 6350 12976 6418 13032
rect 6474 12976 6542 13032
rect 6598 12976 6666 13032
rect 6722 12976 6790 13032
rect 6846 12976 6914 13032
rect 6970 12976 7038 13032
rect 7094 12976 7104 13032
rect 5168 12908 7104 12976
rect 5168 12852 5178 12908
rect 5234 12852 5302 12908
rect 5358 12852 5426 12908
rect 5482 12852 5550 12908
rect 5606 12852 5674 12908
rect 5730 12852 5798 12908
rect 5854 12852 5922 12908
rect 5978 12852 6046 12908
rect 6102 12852 6170 12908
rect 6226 12852 6294 12908
rect 6350 12852 6418 12908
rect 6474 12852 6542 12908
rect 6598 12852 6666 12908
rect 6722 12852 6790 12908
rect 6846 12852 6914 12908
rect 6970 12852 7038 12908
rect 7094 12852 7104 12908
rect 5168 12842 7104 12852
rect 7874 14148 9810 14158
rect 7874 14092 7884 14148
rect 7940 14092 8008 14148
rect 8064 14092 8132 14148
rect 8188 14092 8256 14148
rect 8312 14092 8380 14148
rect 8436 14092 8504 14148
rect 8560 14092 8628 14148
rect 8684 14092 8752 14148
rect 8808 14092 8876 14148
rect 8932 14092 9000 14148
rect 9056 14092 9124 14148
rect 9180 14092 9248 14148
rect 9304 14092 9372 14148
rect 9428 14092 9496 14148
rect 9552 14092 9620 14148
rect 9676 14092 9744 14148
rect 9800 14092 9810 14148
rect 7874 14024 9810 14092
rect 7874 13968 7884 14024
rect 7940 13968 8008 14024
rect 8064 13968 8132 14024
rect 8188 13968 8256 14024
rect 8312 13968 8380 14024
rect 8436 13968 8504 14024
rect 8560 13968 8628 14024
rect 8684 13968 8752 14024
rect 8808 13968 8876 14024
rect 8932 13968 9000 14024
rect 9056 13968 9124 14024
rect 9180 13968 9248 14024
rect 9304 13968 9372 14024
rect 9428 13968 9496 14024
rect 9552 13968 9620 14024
rect 9676 13968 9744 14024
rect 9800 13968 9810 14024
rect 7874 13900 9810 13968
rect 7874 13844 7884 13900
rect 7940 13844 8008 13900
rect 8064 13844 8132 13900
rect 8188 13844 8256 13900
rect 8312 13844 8380 13900
rect 8436 13844 8504 13900
rect 8560 13844 8628 13900
rect 8684 13844 8752 13900
rect 8808 13844 8876 13900
rect 8932 13844 9000 13900
rect 9056 13844 9124 13900
rect 9180 13844 9248 13900
rect 9304 13844 9372 13900
rect 9428 13844 9496 13900
rect 9552 13844 9620 13900
rect 9676 13844 9744 13900
rect 9800 13844 9810 13900
rect 7874 13776 9810 13844
rect 7874 13720 7884 13776
rect 7940 13720 8008 13776
rect 8064 13720 8132 13776
rect 8188 13720 8256 13776
rect 8312 13720 8380 13776
rect 8436 13720 8504 13776
rect 8560 13720 8628 13776
rect 8684 13720 8752 13776
rect 8808 13720 8876 13776
rect 8932 13720 9000 13776
rect 9056 13720 9124 13776
rect 9180 13720 9248 13776
rect 9304 13720 9372 13776
rect 9428 13720 9496 13776
rect 9552 13720 9620 13776
rect 9676 13720 9744 13776
rect 9800 13720 9810 13776
rect 7874 13652 9810 13720
rect 7874 13596 7884 13652
rect 7940 13596 8008 13652
rect 8064 13596 8132 13652
rect 8188 13596 8256 13652
rect 8312 13596 8380 13652
rect 8436 13596 8504 13652
rect 8560 13596 8628 13652
rect 8684 13596 8752 13652
rect 8808 13596 8876 13652
rect 8932 13596 9000 13652
rect 9056 13596 9124 13652
rect 9180 13596 9248 13652
rect 9304 13596 9372 13652
rect 9428 13596 9496 13652
rect 9552 13596 9620 13652
rect 9676 13596 9744 13652
rect 9800 13596 9810 13652
rect 7874 13528 9810 13596
rect 7874 13472 7884 13528
rect 7940 13472 8008 13528
rect 8064 13472 8132 13528
rect 8188 13472 8256 13528
rect 8312 13472 8380 13528
rect 8436 13472 8504 13528
rect 8560 13472 8628 13528
rect 8684 13472 8752 13528
rect 8808 13472 8876 13528
rect 8932 13472 9000 13528
rect 9056 13472 9124 13528
rect 9180 13472 9248 13528
rect 9304 13472 9372 13528
rect 9428 13472 9496 13528
rect 9552 13472 9620 13528
rect 9676 13472 9744 13528
rect 9800 13472 9810 13528
rect 7874 13404 9810 13472
rect 7874 13348 7884 13404
rect 7940 13348 8008 13404
rect 8064 13348 8132 13404
rect 8188 13348 8256 13404
rect 8312 13348 8380 13404
rect 8436 13348 8504 13404
rect 8560 13348 8628 13404
rect 8684 13348 8752 13404
rect 8808 13348 8876 13404
rect 8932 13348 9000 13404
rect 9056 13348 9124 13404
rect 9180 13348 9248 13404
rect 9304 13348 9372 13404
rect 9428 13348 9496 13404
rect 9552 13348 9620 13404
rect 9676 13348 9744 13404
rect 9800 13348 9810 13404
rect 7874 13280 9810 13348
rect 7874 13224 7884 13280
rect 7940 13224 8008 13280
rect 8064 13224 8132 13280
rect 8188 13224 8256 13280
rect 8312 13224 8380 13280
rect 8436 13224 8504 13280
rect 8560 13224 8628 13280
rect 8684 13224 8752 13280
rect 8808 13224 8876 13280
rect 8932 13224 9000 13280
rect 9056 13224 9124 13280
rect 9180 13224 9248 13280
rect 9304 13224 9372 13280
rect 9428 13224 9496 13280
rect 9552 13224 9620 13280
rect 9676 13224 9744 13280
rect 9800 13224 9810 13280
rect 7874 13156 9810 13224
rect 7874 13100 7884 13156
rect 7940 13100 8008 13156
rect 8064 13100 8132 13156
rect 8188 13100 8256 13156
rect 8312 13100 8380 13156
rect 8436 13100 8504 13156
rect 8560 13100 8628 13156
rect 8684 13100 8752 13156
rect 8808 13100 8876 13156
rect 8932 13100 9000 13156
rect 9056 13100 9124 13156
rect 9180 13100 9248 13156
rect 9304 13100 9372 13156
rect 9428 13100 9496 13156
rect 9552 13100 9620 13156
rect 9676 13100 9744 13156
rect 9800 13100 9810 13156
rect 7874 13032 9810 13100
rect 7874 12976 7884 13032
rect 7940 12976 8008 13032
rect 8064 12976 8132 13032
rect 8188 12976 8256 13032
rect 8312 12976 8380 13032
rect 8436 12976 8504 13032
rect 8560 12976 8628 13032
rect 8684 12976 8752 13032
rect 8808 12976 8876 13032
rect 8932 12976 9000 13032
rect 9056 12976 9124 13032
rect 9180 12976 9248 13032
rect 9304 12976 9372 13032
rect 9428 12976 9496 13032
rect 9552 12976 9620 13032
rect 9676 12976 9744 13032
rect 9800 12976 9810 13032
rect 7874 12908 9810 12976
rect 7874 12852 7884 12908
rect 7940 12852 8008 12908
rect 8064 12852 8132 12908
rect 8188 12852 8256 12908
rect 8312 12852 8380 12908
rect 8436 12852 8504 12908
rect 8560 12852 8628 12908
rect 8684 12852 8752 12908
rect 8808 12852 8876 12908
rect 8932 12852 9000 12908
rect 9056 12852 9124 12908
rect 9180 12852 9248 12908
rect 9304 12852 9372 12908
rect 9428 12852 9496 12908
rect 9552 12852 9620 12908
rect 9676 12852 9744 12908
rect 9800 12852 9810 12908
rect 7874 12842 9810 12852
rect 10244 14148 12180 14158
rect 10244 14092 10254 14148
rect 10310 14092 10378 14148
rect 10434 14092 10502 14148
rect 10558 14092 10626 14148
rect 10682 14092 10750 14148
rect 10806 14092 10874 14148
rect 10930 14092 10998 14148
rect 11054 14092 11122 14148
rect 11178 14092 11246 14148
rect 11302 14092 11370 14148
rect 11426 14092 11494 14148
rect 11550 14092 11618 14148
rect 11674 14092 11742 14148
rect 11798 14092 11866 14148
rect 11922 14092 11990 14148
rect 12046 14092 12114 14148
rect 12170 14092 12180 14148
rect 10244 14024 12180 14092
rect 10244 13968 10254 14024
rect 10310 13968 10378 14024
rect 10434 13968 10502 14024
rect 10558 13968 10626 14024
rect 10682 13968 10750 14024
rect 10806 13968 10874 14024
rect 10930 13968 10998 14024
rect 11054 13968 11122 14024
rect 11178 13968 11246 14024
rect 11302 13968 11370 14024
rect 11426 13968 11494 14024
rect 11550 13968 11618 14024
rect 11674 13968 11742 14024
rect 11798 13968 11866 14024
rect 11922 13968 11990 14024
rect 12046 13968 12114 14024
rect 12170 13968 12180 14024
rect 10244 13900 12180 13968
rect 10244 13844 10254 13900
rect 10310 13844 10378 13900
rect 10434 13844 10502 13900
rect 10558 13844 10626 13900
rect 10682 13844 10750 13900
rect 10806 13844 10874 13900
rect 10930 13844 10998 13900
rect 11054 13844 11122 13900
rect 11178 13844 11246 13900
rect 11302 13844 11370 13900
rect 11426 13844 11494 13900
rect 11550 13844 11618 13900
rect 11674 13844 11742 13900
rect 11798 13844 11866 13900
rect 11922 13844 11990 13900
rect 12046 13844 12114 13900
rect 12170 13844 12180 13900
rect 10244 13776 12180 13844
rect 10244 13720 10254 13776
rect 10310 13720 10378 13776
rect 10434 13720 10502 13776
rect 10558 13720 10626 13776
rect 10682 13720 10750 13776
rect 10806 13720 10874 13776
rect 10930 13720 10998 13776
rect 11054 13720 11122 13776
rect 11178 13720 11246 13776
rect 11302 13720 11370 13776
rect 11426 13720 11494 13776
rect 11550 13720 11618 13776
rect 11674 13720 11742 13776
rect 11798 13720 11866 13776
rect 11922 13720 11990 13776
rect 12046 13720 12114 13776
rect 12170 13720 12180 13776
rect 10244 13652 12180 13720
rect 10244 13596 10254 13652
rect 10310 13596 10378 13652
rect 10434 13596 10502 13652
rect 10558 13596 10626 13652
rect 10682 13596 10750 13652
rect 10806 13596 10874 13652
rect 10930 13596 10998 13652
rect 11054 13596 11122 13652
rect 11178 13596 11246 13652
rect 11302 13596 11370 13652
rect 11426 13596 11494 13652
rect 11550 13596 11618 13652
rect 11674 13596 11742 13652
rect 11798 13596 11866 13652
rect 11922 13596 11990 13652
rect 12046 13596 12114 13652
rect 12170 13596 12180 13652
rect 10244 13528 12180 13596
rect 10244 13472 10254 13528
rect 10310 13472 10378 13528
rect 10434 13472 10502 13528
rect 10558 13472 10626 13528
rect 10682 13472 10750 13528
rect 10806 13472 10874 13528
rect 10930 13472 10998 13528
rect 11054 13472 11122 13528
rect 11178 13472 11246 13528
rect 11302 13472 11370 13528
rect 11426 13472 11494 13528
rect 11550 13472 11618 13528
rect 11674 13472 11742 13528
rect 11798 13472 11866 13528
rect 11922 13472 11990 13528
rect 12046 13472 12114 13528
rect 12170 13472 12180 13528
rect 10244 13404 12180 13472
rect 10244 13348 10254 13404
rect 10310 13348 10378 13404
rect 10434 13348 10502 13404
rect 10558 13348 10626 13404
rect 10682 13348 10750 13404
rect 10806 13348 10874 13404
rect 10930 13348 10998 13404
rect 11054 13348 11122 13404
rect 11178 13348 11246 13404
rect 11302 13348 11370 13404
rect 11426 13348 11494 13404
rect 11550 13348 11618 13404
rect 11674 13348 11742 13404
rect 11798 13348 11866 13404
rect 11922 13348 11990 13404
rect 12046 13348 12114 13404
rect 12170 13348 12180 13404
rect 10244 13280 12180 13348
rect 10244 13224 10254 13280
rect 10310 13224 10378 13280
rect 10434 13224 10502 13280
rect 10558 13224 10626 13280
rect 10682 13224 10750 13280
rect 10806 13224 10874 13280
rect 10930 13224 10998 13280
rect 11054 13224 11122 13280
rect 11178 13224 11246 13280
rect 11302 13224 11370 13280
rect 11426 13224 11494 13280
rect 11550 13224 11618 13280
rect 11674 13224 11742 13280
rect 11798 13224 11866 13280
rect 11922 13224 11990 13280
rect 12046 13224 12114 13280
rect 12170 13224 12180 13280
rect 10244 13156 12180 13224
rect 10244 13100 10254 13156
rect 10310 13100 10378 13156
rect 10434 13100 10502 13156
rect 10558 13100 10626 13156
rect 10682 13100 10750 13156
rect 10806 13100 10874 13156
rect 10930 13100 10998 13156
rect 11054 13100 11122 13156
rect 11178 13100 11246 13156
rect 11302 13100 11370 13156
rect 11426 13100 11494 13156
rect 11550 13100 11618 13156
rect 11674 13100 11742 13156
rect 11798 13100 11866 13156
rect 11922 13100 11990 13156
rect 12046 13100 12114 13156
rect 12170 13100 12180 13156
rect 10244 13032 12180 13100
rect 10244 12976 10254 13032
rect 10310 12976 10378 13032
rect 10434 12976 10502 13032
rect 10558 12976 10626 13032
rect 10682 12976 10750 13032
rect 10806 12976 10874 13032
rect 10930 12976 10998 13032
rect 11054 12976 11122 13032
rect 11178 12976 11246 13032
rect 11302 12976 11370 13032
rect 11426 12976 11494 13032
rect 11550 12976 11618 13032
rect 11674 12976 11742 13032
rect 11798 12976 11866 13032
rect 11922 12976 11990 13032
rect 12046 12976 12114 13032
rect 12170 12976 12180 13032
rect 10244 12908 12180 12976
rect 10244 12852 10254 12908
rect 10310 12852 10378 12908
rect 10434 12852 10502 12908
rect 10558 12852 10626 12908
rect 10682 12852 10750 12908
rect 10806 12852 10874 12908
rect 10930 12852 10998 12908
rect 11054 12852 11122 12908
rect 11178 12852 11246 12908
rect 11302 12852 11370 12908
rect 11426 12852 11494 12908
rect 11550 12852 11618 12908
rect 11674 12852 11742 12908
rect 11798 12852 11866 12908
rect 11922 12852 11990 12908
rect 12046 12852 12114 12908
rect 12170 12852 12180 12908
rect 10244 12842 12180 12852
rect 12861 14148 14673 14158
rect 12861 14092 12871 14148
rect 12927 14092 12995 14148
rect 13051 14092 13119 14148
rect 13175 14092 13243 14148
rect 13299 14092 13367 14148
rect 13423 14092 13491 14148
rect 13547 14092 13615 14148
rect 13671 14092 13739 14148
rect 13795 14092 13863 14148
rect 13919 14092 13987 14148
rect 14043 14092 14111 14148
rect 14167 14092 14235 14148
rect 14291 14092 14359 14148
rect 14415 14092 14483 14148
rect 14539 14092 14607 14148
rect 14663 14092 14673 14148
rect 12861 14024 14673 14092
rect 12861 13968 12871 14024
rect 12927 13968 12995 14024
rect 13051 13968 13119 14024
rect 13175 13968 13243 14024
rect 13299 13968 13367 14024
rect 13423 13968 13491 14024
rect 13547 13968 13615 14024
rect 13671 13968 13739 14024
rect 13795 13968 13863 14024
rect 13919 13968 13987 14024
rect 14043 13968 14111 14024
rect 14167 13968 14235 14024
rect 14291 13968 14359 14024
rect 14415 13968 14483 14024
rect 14539 13968 14607 14024
rect 14663 13968 14673 14024
rect 12861 13900 14673 13968
rect 12861 13844 12871 13900
rect 12927 13844 12995 13900
rect 13051 13844 13119 13900
rect 13175 13844 13243 13900
rect 13299 13844 13367 13900
rect 13423 13844 13491 13900
rect 13547 13844 13615 13900
rect 13671 13844 13739 13900
rect 13795 13844 13863 13900
rect 13919 13844 13987 13900
rect 14043 13844 14111 13900
rect 14167 13844 14235 13900
rect 14291 13844 14359 13900
rect 14415 13844 14483 13900
rect 14539 13844 14607 13900
rect 14663 13844 14673 13900
rect 12861 13776 14673 13844
rect 12861 13720 12871 13776
rect 12927 13720 12995 13776
rect 13051 13720 13119 13776
rect 13175 13720 13243 13776
rect 13299 13720 13367 13776
rect 13423 13720 13491 13776
rect 13547 13720 13615 13776
rect 13671 13720 13739 13776
rect 13795 13720 13863 13776
rect 13919 13720 13987 13776
rect 14043 13720 14111 13776
rect 14167 13720 14235 13776
rect 14291 13720 14359 13776
rect 14415 13720 14483 13776
rect 14539 13720 14607 13776
rect 14663 13720 14673 13776
rect 12861 13652 14673 13720
rect 12861 13596 12871 13652
rect 12927 13596 12995 13652
rect 13051 13596 13119 13652
rect 13175 13596 13243 13652
rect 13299 13596 13367 13652
rect 13423 13596 13491 13652
rect 13547 13596 13615 13652
rect 13671 13596 13739 13652
rect 13795 13596 13863 13652
rect 13919 13596 13987 13652
rect 14043 13596 14111 13652
rect 14167 13596 14235 13652
rect 14291 13596 14359 13652
rect 14415 13596 14483 13652
rect 14539 13596 14607 13652
rect 14663 13596 14673 13652
rect 12861 13528 14673 13596
rect 12861 13472 12871 13528
rect 12927 13472 12995 13528
rect 13051 13472 13119 13528
rect 13175 13472 13243 13528
rect 13299 13472 13367 13528
rect 13423 13472 13491 13528
rect 13547 13472 13615 13528
rect 13671 13472 13739 13528
rect 13795 13472 13863 13528
rect 13919 13472 13987 13528
rect 14043 13472 14111 13528
rect 14167 13472 14235 13528
rect 14291 13472 14359 13528
rect 14415 13472 14483 13528
rect 14539 13472 14607 13528
rect 14663 13472 14673 13528
rect 12861 13404 14673 13472
rect 12861 13348 12871 13404
rect 12927 13348 12995 13404
rect 13051 13348 13119 13404
rect 13175 13348 13243 13404
rect 13299 13348 13367 13404
rect 13423 13348 13491 13404
rect 13547 13348 13615 13404
rect 13671 13348 13739 13404
rect 13795 13348 13863 13404
rect 13919 13348 13987 13404
rect 14043 13348 14111 13404
rect 14167 13348 14235 13404
rect 14291 13348 14359 13404
rect 14415 13348 14483 13404
rect 14539 13348 14607 13404
rect 14663 13348 14673 13404
rect 12861 13280 14673 13348
rect 12861 13224 12871 13280
rect 12927 13224 12995 13280
rect 13051 13224 13119 13280
rect 13175 13224 13243 13280
rect 13299 13224 13367 13280
rect 13423 13224 13491 13280
rect 13547 13224 13615 13280
rect 13671 13224 13739 13280
rect 13795 13224 13863 13280
rect 13919 13224 13987 13280
rect 14043 13224 14111 13280
rect 14167 13224 14235 13280
rect 14291 13224 14359 13280
rect 14415 13224 14483 13280
rect 14539 13224 14607 13280
rect 14663 13224 14673 13280
rect 12861 13156 14673 13224
rect 12861 13100 12871 13156
rect 12927 13100 12995 13156
rect 13051 13100 13119 13156
rect 13175 13100 13243 13156
rect 13299 13100 13367 13156
rect 13423 13100 13491 13156
rect 13547 13100 13615 13156
rect 13671 13100 13739 13156
rect 13795 13100 13863 13156
rect 13919 13100 13987 13156
rect 14043 13100 14111 13156
rect 14167 13100 14235 13156
rect 14291 13100 14359 13156
rect 14415 13100 14483 13156
rect 14539 13100 14607 13156
rect 14663 13100 14673 13156
rect 12861 13032 14673 13100
rect 12861 12976 12871 13032
rect 12927 12976 12995 13032
rect 13051 12976 13119 13032
rect 13175 12976 13243 13032
rect 13299 12976 13367 13032
rect 13423 12976 13491 13032
rect 13547 12976 13615 13032
rect 13671 12976 13739 13032
rect 13795 12976 13863 13032
rect 13919 12976 13987 13032
rect 14043 12976 14111 13032
rect 14167 12976 14235 13032
rect 14291 12976 14359 13032
rect 14415 12976 14483 13032
rect 14539 12976 14607 13032
rect 14663 12976 14673 13032
rect 12861 12908 14673 12976
rect 12861 12852 12871 12908
rect 12927 12852 12995 12908
rect 13051 12852 13119 12908
rect 13175 12852 13243 12908
rect 13299 12852 13367 12908
rect 13423 12852 13491 12908
rect 13547 12852 13615 12908
rect 13671 12852 13739 12908
rect 13795 12852 13863 12908
rect 13919 12852 13987 12908
rect 14043 12852 14111 12908
rect 14167 12852 14235 12908
rect 14291 12852 14359 12908
rect 14415 12852 14483 12908
rect 14539 12852 14607 12908
rect 14663 12852 14673 12908
rect 12861 12842 14673 12852
rect -11 12814 86 12824
rect 14892 12824 14902 14176
rect 14958 12824 14989 14176
rect 14892 12814 14989 12824
rect 2481 12548 2681 12558
rect 2481 12492 2491 12548
rect 2547 12492 2615 12548
rect 2671 12492 2681 12548
rect 2481 12424 2681 12492
rect 2481 12368 2491 12424
rect 2547 12368 2615 12424
rect 2671 12368 2681 12424
rect 2481 12300 2681 12368
rect 2481 12244 2491 12300
rect 2547 12244 2615 12300
rect 2671 12244 2681 12300
rect 2481 12176 2681 12244
rect 2481 12120 2491 12176
rect 2547 12120 2615 12176
rect 2671 12120 2681 12176
rect 2481 12052 2681 12120
rect 2481 11996 2491 12052
rect 2547 11996 2615 12052
rect 2671 11996 2681 12052
rect 2481 11928 2681 11996
rect 2481 11872 2491 11928
rect 2547 11872 2615 11928
rect 2671 11872 2681 11928
rect 2481 11804 2681 11872
rect 2481 11748 2491 11804
rect 2547 11748 2615 11804
rect 2671 11748 2681 11804
rect 2481 11680 2681 11748
rect 2481 11624 2491 11680
rect 2547 11624 2615 11680
rect 2671 11624 2681 11680
rect 2481 11556 2681 11624
rect 2481 11500 2491 11556
rect 2547 11500 2615 11556
rect 2671 11500 2681 11556
rect 2481 11432 2681 11500
rect 2481 11376 2491 11432
rect 2547 11376 2615 11432
rect 2671 11376 2681 11432
rect 2481 11308 2681 11376
rect 2481 11252 2491 11308
rect 2547 11252 2615 11308
rect 2671 11252 2681 11308
rect 2481 11242 2681 11252
rect 4851 12548 5051 12558
rect 4851 12492 4861 12548
rect 4917 12492 4985 12548
rect 5041 12492 5051 12548
rect 4851 12424 5051 12492
rect 4851 12368 4861 12424
rect 4917 12368 4985 12424
rect 5041 12368 5051 12424
rect 4851 12300 5051 12368
rect 4851 12244 4861 12300
rect 4917 12244 4985 12300
rect 5041 12244 5051 12300
rect 4851 12176 5051 12244
rect 4851 12120 4861 12176
rect 4917 12120 4985 12176
rect 5041 12120 5051 12176
rect 4851 12052 5051 12120
rect 4851 11996 4861 12052
rect 4917 11996 4985 12052
rect 5041 11996 5051 12052
rect 4851 11928 5051 11996
rect 4851 11872 4861 11928
rect 4917 11872 4985 11928
rect 5041 11872 5051 11928
rect 4851 11804 5051 11872
rect 4851 11748 4861 11804
rect 4917 11748 4985 11804
rect 5041 11748 5051 11804
rect 4851 11680 5051 11748
rect 4851 11624 4861 11680
rect 4917 11624 4985 11680
rect 5041 11624 5051 11680
rect 4851 11556 5051 11624
rect 4851 11500 4861 11556
rect 4917 11500 4985 11556
rect 5041 11500 5051 11556
rect 4851 11432 5051 11500
rect 4851 11376 4861 11432
rect 4917 11376 4985 11432
rect 5041 11376 5051 11432
rect 4851 11308 5051 11376
rect 4851 11252 4861 11308
rect 4917 11252 4985 11308
rect 5041 11252 5051 11308
rect 4851 11242 5051 11252
rect 7265 12548 7713 12558
rect 7265 12492 7275 12548
rect 7331 12492 7399 12548
rect 7455 12492 7523 12548
rect 7579 12492 7647 12548
rect 7703 12492 7713 12548
rect 7265 12424 7713 12492
rect 7265 12368 7275 12424
rect 7331 12368 7399 12424
rect 7455 12368 7523 12424
rect 7579 12368 7647 12424
rect 7703 12368 7713 12424
rect 7265 12300 7713 12368
rect 7265 12244 7275 12300
rect 7331 12244 7399 12300
rect 7455 12244 7523 12300
rect 7579 12244 7647 12300
rect 7703 12244 7713 12300
rect 7265 12176 7713 12244
rect 7265 12120 7275 12176
rect 7331 12120 7399 12176
rect 7455 12120 7523 12176
rect 7579 12120 7647 12176
rect 7703 12120 7713 12176
rect 7265 12052 7713 12120
rect 7265 11996 7275 12052
rect 7331 11996 7399 12052
rect 7455 11996 7523 12052
rect 7579 11996 7647 12052
rect 7703 11996 7713 12052
rect 7265 11928 7713 11996
rect 7265 11872 7275 11928
rect 7331 11872 7399 11928
rect 7455 11872 7523 11928
rect 7579 11872 7647 11928
rect 7703 11872 7713 11928
rect 7265 11804 7713 11872
rect 7265 11748 7275 11804
rect 7331 11748 7399 11804
rect 7455 11748 7523 11804
rect 7579 11748 7647 11804
rect 7703 11748 7713 11804
rect 7265 11680 7713 11748
rect 7265 11624 7275 11680
rect 7331 11624 7399 11680
rect 7455 11624 7523 11680
rect 7579 11624 7647 11680
rect 7703 11624 7713 11680
rect 7265 11556 7713 11624
rect 7265 11500 7275 11556
rect 7331 11500 7399 11556
rect 7455 11500 7523 11556
rect 7579 11500 7647 11556
rect 7703 11500 7713 11556
rect 7265 11432 7713 11500
rect 7265 11376 7275 11432
rect 7331 11376 7399 11432
rect 7455 11376 7523 11432
rect 7579 11376 7647 11432
rect 7703 11376 7713 11432
rect 7265 11308 7713 11376
rect 7265 11252 7275 11308
rect 7331 11252 7399 11308
rect 7455 11252 7523 11308
rect 7579 11252 7647 11308
rect 7703 11252 7713 11308
rect 7265 11242 7713 11252
rect 9927 12548 10127 12558
rect 9927 12492 9937 12548
rect 9993 12492 10061 12548
rect 10117 12492 10127 12548
rect 9927 12424 10127 12492
rect 9927 12368 9937 12424
rect 9993 12368 10061 12424
rect 10117 12368 10127 12424
rect 9927 12300 10127 12368
rect 9927 12244 9937 12300
rect 9993 12244 10061 12300
rect 10117 12244 10127 12300
rect 9927 12176 10127 12244
rect 9927 12120 9937 12176
rect 9993 12120 10061 12176
rect 10117 12120 10127 12176
rect 9927 12052 10127 12120
rect 9927 11996 9937 12052
rect 9993 11996 10061 12052
rect 10117 11996 10127 12052
rect 9927 11928 10127 11996
rect 9927 11872 9937 11928
rect 9993 11872 10061 11928
rect 10117 11872 10127 11928
rect 9927 11804 10127 11872
rect 9927 11748 9937 11804
rect 9993 11748 10061 11804
rect 10117 11748 10127 11804
rect 9927 11680 10127 11748
rect 9927 11624 9937 11680
rect 9993 11624 10061 11680
rect 10117 11624 10127 11680
rect 9927 11556 10127 11624
rect 9927 11500 9937 11556
rect 9993 11500 10061 11556
rect 10117 11500 10127 11556
rect 9927 11432 10127 11500
rect 9927 11376 9937 11432
rect 9993 11376 10061 11432
rect 10117 11376 10127 11432
rect 9927 11308 10127 11376
rect 9927 11252 9937 11308
rect 9993 11252 10061 11308
rect 10117 11252 10127 11308
rect 9927 11242 10127 11252
rect 12297 12548 12497 12558
rect 12297 12492 12307 12548
rect 12363 12492 12431 12548
rect 12487 12492 12497 12548
rect 12297 12424 12497 12492
rect 12297 12368 12307 12424
rect 12363 12368 12431 12424
rect 12487 12368 12497 12424
rect 12297 12300 12497 12368
rect 12297 12244 12307 12300
rect 12363 12244 12431 12300
rect 12487 12244 12497 12300
rect 12297 12176 12497 12244
rect 12297 12120 12307 12176
rect 12363 12120 12431 12176
rect 12487 12120 12497 12176
rect 12297 12052 12497 12120
rect 12297 11996 12307 12052
rect 12363 11996 12431 12052
rect 12487 11996 12497 12052
rect 12297 11928 12497 11996
rect 12297 11872 12307 11928
rect 12363 11872 12431 11928
rect 12487 11872 12497 11928
rect 12297 11804 12497 11872
rect 12297 11748 12307 11804
rect 12363 11748 12431 11804
rect 12487 11748 12497 11804
rect 12297 11680 12497 11748
rect 12297 11624 12307 11680
rect 12363 11624 12431 11680
rect 12487 11624 12497 11680
rect 12297 11556 12497 11624
rect 12297 11500 12307 11556
rect 12363 11500 12431 11556
rect 12487 11500 12497 11556
rect 12297 11432 12497 11500
rect 12297 11376 12307 11432
rect 12363 11376 12431 11432
rect 12487 11376 12497 11432
rect 12297 11308 12497 11376
rect 12297 11252 12307 11308
rect 12363 11252 12431 11308
rect 12487 11252 12497 11308
rect 12297 11242 12497 11252
rect -11 10986 86 10996
rect -11 8014 20 10986
rect 76 8014 86 10986
rect 14892 10986 14989 10996
rect 305 10954 2117 10964
rect 305 10898 315 10954
rect 371 10898 439 10954
rect 495 10898 563 10954
rect 619 10898 687 10954
rect 743 10898 811 10954
rect 867 10898 935 10954
rect 991 10898 1059 10954
rect 1115 10898 1183 10954
rect 1239 10898 1307 10954
rect 1363 10898 1431 10954
rect 1487 10898 1555 10954
rect 1611 10898 1679 10954
rect 1735 10898 1803 10954
rect 1859 10898 1927 10954
rect 1983 10898 2051 10954
rect 2107 10898 2117 10954
rect 305 10830 2117 10898
rect 305 10774 315 10830
rect 371 10774 439 10830
rect 495 10774 563 10830
rect 619 10774 687 10830
rect 743 10774 811 10830
rect 867 10774 935 10830
rect 991 10774 1059 10830
rect 1115 10774 1183 10830
rect 1239 10774 1307 10830
rect 1363 10774 1431 10830
rect 1487 10774 1555 10830
rect 1611 10774 1679 10830
rect 1735 10774 1803 10830
rect 1859 10774 1927 10830
rect 1983 10774 2051 10830
rect 2107 10774 2117 10830
rect 305 10706 2117 10774
rect 305 10650 315 10706
rect 371 10650 439 10706
rect 495 10650 563 10706
rect 619 10650 687 10706
rect 743 10650 811 10706
rect 867 10650 935 10706
rect 991 10650 1059 10706
rect 1115 10650 1183 10706
rect 1239 10650 1307 10706
rect 1363 10650 1431 10706
rect 1487 10650 1555 10706
rect 1611 10650 1679 10706
rect 1735 10650 1803 10706
rect 1859 10650 1927 10706
rect 1983 10650 2051 10706
rect 2107 10650 2117 10706
rect 305 10582 2117 10650
rect 305 10526 315 10582
rect 371 10526 439 10582
rect 495 10526 563 10582
rect 619 10526 687 10582
rect 743 10526 811 10582
rect 867 10526 935 10582
rect 991 10526 1059 10582
rect 1115 10526 1183 10582
rect 1239 10526 1307 10582
rect 1363 10526 1431 10582
rect 1487 10526 1555 10582
rect 1611 10526 1679 10582
rect 1735 10526 1803 10582
rect 1859 10526 1927 10582
rect 1983 10526 2051 10582
rect 2107 10526 2117 10582
rect 305 10458 2117 10526
rect 305 10402 315 10458
rect 371 10402 439 10458
rect 495 10402 563 10458
rect 619 10402 687 10458
rect 743 10402 811 10458
rect 867 10402 935 10458
rect 991 10402 1059 10458
rect 1115 10402 1183 10458
rect 1239 10402 1307 10458
rect 1363 10402 1431 10458
rect 1487 10402 1555 10458
rect 1611 10402 1679 10458
rect 1735 10402 1803 10458
rect 1859 10402 1927 10458
rect 1983 10402 2051 10458
rect 2107 10402 2117 10458
rect 305 10334 2117 10402
rect 305 10278 315 10334
rect 371 10278 439 10334
rect 495 10278 563 10334
rect 619 10278 687 10334
rect 743 10278 811 10334
rect 867 10278 935 10334
rect 991 10278 1059 10334
rect 1115 10278 1183 10334
rect 1239 10278 1307 10334
rect 1363 10278 1431 10334
rect 1487 10278 1555 10334
rect 1611 10278 1679 10334
rect 1735 10278 1803 10334
rect 1859 10278 1927 10334
rect 1983 10278 2051 10334
rect 2107 10278 2117 10334
rect 305 10210 2117 10278
rect 305 10154 315 10210
rect 371 10154 439 10210
rect 495 10154 563 10210
rect 619 10154 687 10210
rect 743 10154 811 10210
rect 867 10154 935 10210
rect 991 10154 1059 10210
rect 1115 10154 1183 10210
rect 1239 10154 1307 10210
rect 1363 10154 1431 10210
rect 1487 10154 1555 10210
rect 1611 10154 1679 10210
rect 1735 10154 1803 10210
rect 1859 10154 1927 10210
rect 1983 10154 2051 10210
rect 2107 10154 2117 10210
rect 305 10086 2117 10154
rect 305 10030 315 10086
rect 371 10030 439 10086
rect 495 10030 563 10086
rect 619 10030 687 10086
rect 743 10030 811 10086
rect 867 10030 935 10086
rect 991 10030 1059 10086
rect 1115 10030 1183 10086
rect 1239 10030 1307 10086
rect 1363 10030 1431 10086
rect 1487 10030 1555 10086
rect 1611 10030 1679 10086
rect 1735 10030 1803 10086
rect 1859 10030 1927 10086
rect 1983 10030 2051 10086
rect 2107 10030 2117 10086
rect 305 9962 2117 10030
rect 305 9906 315 9962
rect 371 9906 439 9962
rect 495 9906 563 9962
rect 619 9906 687 9962
rect 743 9906 811 9962
rect 867 9906 935 9962
rect 991 9906 1059 9962
rect 1115 9906 1183 9962
rect 1239 9906 1307 9962
rect 1363 9906 1431 9962
rect 1487 9906 1555 9962
rect 1611 9906 1679 9962
rect 1735 9906 1803 9962
rect 1859 9906 1927 9962
rect 1983 9906 2051 9962
rect 2107 9906 2117 9962
rect 305 9838 2117 9906
rect 305 9782 315 9838
rect 371 9782 439 9838
rect 495 9782 563 9838
rect 619 9782 687 9838
rect 743 9782 811 9838
rect 867 9782 935 9838
rect 991 9782 1059 9838
rect 1115 9782 1183 9838
rect 1239 9782 1307 9838
rect 1363 9782 1431 9838
rect 1487 9782 1555 9838
rect 1611 9782 1679 9838
rect 1735 9782 1803 9838
rect 1859 9782 1927 9838
rect 1983 9782 2051 9838
rect 2107 9782 2117 9838
rect 305 9714 2117 9782
rect 305 9658 315 9714
rect 371 9658 439 9714
rect 495 9658 563 9714
rect 619 9658 687 9714
rect 743 9658 811 9714
rect 867 9658 935 9714
rect 991 9658 1059 9714
rect 1115 9658 1183 9714
rect 1239 9658 1307 9714
rect 1363 9658 1431 9714
rect 1487 9658 1555 9714
rect 1611 9658 1679 9714
rect 1735 9658 1803 9714
rect 1859 9658 1927 9714
rect 1983 9658 2051 9714
rect 2107 9658 2117 9714
rect 305 9590 2117 9658
rect 305 9534 315 9590
rect 371 9534 439 9590
rect 495 9534 563 9590
rect 619 9534 687 9590
rect 743 9534 811 9590
rect 867 9534 935 9590
rect 991 9534 1059 9590
rect 1115 9534 1183 9590
rect 1239 9534 1307 9590
rect 1363 9534 1431 9590
rect 1487 9534 1555 9590
rect 1611 9534 1679 9590
rect 1735 9534 1803 9590
rect 1859 9534 1927 9590
rect 1983 9534 2051 9590
rect 2107 9534 2117 9590
rect 305 9466 2117 9534
rect 305 9410 315 9466
rect 371 9410 439 9466
rect 495 9410 563 9466
rect 619 9410 687 9466
rect 743 9410 811 9466
rect 867 9410 935 9466
rect 991 9410 1059 9466
rect 1115 9410 1183 9466
rect 1239 9410 1307 9466
rect 1363 9410 1431 9466
rect 1487 9410 1555 9466
rect 1611 9410 1679 9466
rect 1735 9410 1803 9466
rect 1859 9410 1927 9466
rect 1983 9410 2051 9466
rect 2107 9410 2117 9466
rect 305 9342 2117 9410
rect 305 9286 315 9342
rect 371 9286 439 9342
rect 495 9286 563 9342
rect 619 9286 687 9342
rect 743 9286 811 9342
rect 867 9286 935 9342
rect 991 9286 1059 9342
rect 1115 9286 1183 9342
rect 1239 9286 1307 9342
rect 1363 9286 1431 9342
rect 1487 9286 1555 9342
rect 1611 9286 1679 9342
rect 1735 9286 1803 9342
rect 1859 9286 1927 9342
rect 1983 9286 2051 9342
rect 2107 9286 2117 9342
rect 305 9218 2117 9286
rect 305 9162 315 9218
rect 371 9162 439 9218
rect 495 9162 563 9218
rect 619 9162 687 9218
rect 743 9162 811 9218
rect 867 9162 935 9218
rect 991 9162 1059 9218
rect 1115 9162 1183 9218
rect 1239 9162 1307 9218
rect 1363 9162 1431 9218
rect 1487 9162 1555 9218
rect 1611 9162 1679 9218
rect 1735 9162 1803 9218
rect 1859 9162 1927 9218
rect 1983 9162 2051 9218
rect 2107 9162 2117 9218
rect 305 9094 2117 9162
rect 305 9038 315 9094
rect 371 9038 439 9094
rect 495 9038 563 9094
rect 619 9038 687 9094
rect 743 9038 811 9094
rect 867 9038 935 9094
rect 991 9038 1059 9094
rect 1115 9038 1183 9094
rect 1239 9038 1307 9094
rect 1363 9038 1431 9094
rect 1487 9038 1555 9094
rect 1611 9038 1679 9094
rect 1735 9038 1803 9094
rect 1859 9038 1927 9094
rect 1983 9038 2051 9094
rect 2107 9038 2117 9094
rect 305 8970 2117 9038
rect 305 8914 315 8970
rect 371 8914 439 8970
rect 495 8914 563 8970
rect 619 8914 687 8970
rect 743 8914 811 8970
rect 867 8914 935 8970
rect 991 8914 1059 8970
rect 1115 8914 1183 8970
rect 1239 8914 1307 8970
rect 1363 8914 1431 8970
rect 1487 8914 1555 8970
rect 1611 8914 1679 8970
rect 1735 8914 1803 8970
rect 1859 8914 1927 8970
rect 1983 8914 2051 8970
rect 2107 8914 2117 8970
rect 305 8846 2117 8914
rect 305 8790 315 8846
rect 371 8790 439 8846
rect 495 8790 563 8846
rect 619 8790 687 8846
rect 743 8790 811 8846
rect 867 8790 935 8846
rect 991 8790 1059 8846
rect 1115 8790 1183 8846
rect 1239 8790 1307 8846
rect 1363 8790 1431 8846
rect 1487 8790 1555 8846
rect 1611 8790 1679 8846
rect 1735 8790 1803 8846
rect 1859 8790 1927 8846
rect 1983 8790 2051 8846
rect 2107 8790 2117 8846
rect 305 8722 2117 8790
rect 305 8666 315 8722
rect 371 8666 439 8722
rect 495 8666 563 8722
rect 619 8666 687 8722
rect 743 8666 811 8722
rect 867 8666 935 8722
rect 991 8666 1059 8722
rect 1115 8666 1183 8722
rect 1239 8666 1307 8722
rect 1363 8666 1431 8722
rect 1487 8666 1555 8722
rect 1611 8666 1679 8722
rect 1735 8666 1803 8722
rect 1859 8666 1927 8722
rect 1983 8666 2051 8722
rect 2107 8666 2117 8722
rect 305 8598 2117 8666
rect 305 8542 315 8598
rect 371 8542 439 8598
rect 495 8542 563 8598
rect 619 8542 687 8598
rect 743 8542 811 8598
rect 867 8542 935 8598
rect 991 8542 1059 8598
rect 1115 8542 1183 8598
rect 1239 8542 1307 8598
rect 1363 8542 1431 8598
rect 1487 8542 1555 8598
rect 1611 8542 1679 8598
rect 1735 8542 1803 8598
rect 1859 8542 1927 8598
rect 1983 8542 2051 8598
rect 2107 8542 2117 8598
rect 305 8474 2117 8542
rect 305 8418 315 8474
rect 371 8418 439 8474
rect 495 8418 563 8474
rect 619 8418 687 8474
rect 743 8418 811 8474
rect 867 8418 935 8474
rect 991 8418 1059 8474
rect 1115 8418 1183 8474
rect 1239 8418 1307 8474
rect 1363 8418 1431 8474
rect 1487 8418 1555 8474
rect 1611 8418 1679 8474
rect 1735 8418 1803 8474
rect 1859 8418 1927 8474
rect 1983 8418 2051 8474
rect 2107 8418 2117 8474
rect 305 8350 2117 8418
rect 305 8294 315 8350
rect 371 8294 439 8350
rect 495 8294 563 8350
rect 619 8294 687 8350
rect 743 8294 811 8350
rect 867 8294 935 8350
rect 991 8294 1059 8350
rect 1115 8294 1183 8350
rect 1239 8294 1307 8350
rect 1363 8294 1431 8350
rect 1487 8294 1555 8350
rect 1611 8294 1679 8350
rect 1735 8294 1803 8350
rect 1859 8294 1927 8350
rect 1983 8294 2051 8350
rect 2107 8294 2117 8350
rect 305 8226 2117 8294
rect 305 8170 315 8226
rect 371 8170 439 8226
rect 495 8170 563 8226
rect 619 8170 687 8226
rect 743 8170 811 8226
rect 867 8170 935 8226
rect 991 8170 1059 8226
rect 1115 8170 1183 8226
rect 1239 8170 1307 8226
rect 1363 8170 1431 8226
rect 1487 8170 1555 8226
rect 1611 8170 1679 8226
rect 1735 8170 1803 8226
rect 1859 8170 1927 8226
rect 1983 8170 2051 8226
rect 2107 8170 2117 8226
rect 305 8102 2117 8170
rect 305 8046 315 8102
rect 371 8046 439 8102
rect 495 8046 563 8102
rect 619 8046 687 8102
rect 743 8046 811 8102
rect 867 8046 935 8102
rect 991 8046 1059 8102
rect 1115 8046 1183 8102
rect 1239 8046 1307 8102
rect 1363 8046 1431 8102
rect 1487 8046 1555 8102
rect 1611 8046 1679 8102
rect 1735 8046 1803 8102
rect 1859 8046 1927 8102
rect 1983 8046 2051 8102
rect 2107 8046 2117 8102
rect 305 8036 2117 8046
rect 2798 10954 4734 10964
rect 2798 10898 2808 10954
rect 2864 10898 2932 10954
rect 2988 10898 3056 10954
rect 3112 10898 3180 10954
rect 3236 10898 3304 10954
rect 3360 10898 3428 10954
rect 3484 10898 3552 10954
rect 3608 10898 3676 10954
rect 3732 10898 3800 10954
rect 3856 10898 3924 10954
rect 3980 10898 4048 10954
rect 4104 10898 4172 10954
rect 4228 10898 4296 10954
rect 4352 10898 4420 10954
rect 4476 10898 4544 10954
rect 4600 10898 4668 10954
rect 4724 10898 4734 10954
rect 2798 10830 4734 10898
rect 2798 10774 2808 10830
rect 2864 10774 2932 10830
rect 2988 10774 3056 10830
rect 3112 10774 3180 10830
rect 3236 10774 3304 10830
rect 3360 10774 3428 10830
rect 3484 10774 3552 10830
rect 3608 10774 3676 10830
rect 3732 10774 3800 10830
rect 3856 10774 3924 10830
rect 3980 10774 4048 10830
rect 4104 10774 4172 10830
rect 4228 10774 4296 10830
rect 4352 10774 4420 10830
rect 4476 10774 4544 10830
rect 4600 10774 4668 10830
rect 4724 10774 4734 10830
rect 2798 10706 4734 10774
rect 2798 10650 2808 10706
rect 2864 10650 2932 10706
rect 2988 10650 3056 10706
rect 3112 10650 3180 10706
rect 3236 10650 3304 10706
rect 3360 10650 3428 10706
rect 3484 10650 3552 10706
rect 3608 10650 3676 10706
rect 3732 10650 3800 10706
rect 3856 10650 3924 10706
rect 3980 10650 4048 10706
rect 4104 10650 4172 10706
rect 4228 10650 4296 10706
rect 4352 10650 4420 10706
rect 4476 10650 4544 10706
rect 4600 10650 4668 10706
rect 4724 10650 4734 10706
rect 2798 10582 4734 10650
rect 2798 10526 2808 10582
rect 2864 10526 2932 10582
rect 2988 10526 3056 10582
rect 3112 10526 3180 10582
rect 3236 10526 3304 10582
rect 3360 10526 3428 10582
rect 3484 10526 3552 10582
rect 3608 10526 3676 10582
rect 3732 10526 3800 10582
rect 3856 10526 3924 10582
rect 3980 10526 4048 10582
rect 4104 10526 4172 10582
rect 4228 10526 4296 10582
rect 4352 10526 4420 10582
rect 4476 10526 4544 10582
rect 4600 10526 4668 10582
rect 4724 10526 4734 10582
rect 2798 10458 4734 10526
rect 2798 10402 2808 10458
rect 2864 10402 2932 10458
rect 2988 10402 3056 10458
rect 3112 10402 3180 10458
rect 3236 10402 3304 10458
rect 3360 10402 3428 10458
rect 3484 10402 3552 10458
rect 3608 10402 3676 10458
rect 3732 10402 3800 10458
rect 3856 10402 3924 10458
rect 3980 10402 4048 10458
rect 4104 10402 4172 10458
rect 4228 10402 4296 10458
rect 4352 10402 4420 10458
rect 4476 10402 4544 10458
rect 4600 10402 4668 10458
rect 4724 10402 4734 10458
rect 2798 10334 4734 10402
rect 2798 10278 2808 10334
rect 2864 10278 2932 10334
rect 2988 10278 3056 10334
rect 3112 10278 3180 10334
rect 3236 10278 3304 10334
rect 3360 10278 3428 10334
rect 3484 10278 3552 10334
rect 3608 10278 3676 10334
rect 3732 10278 3800 10334
rect 3856 10278 3924 10334
rect 3980 10278 4048 10334
rect 4104 10278 4172 10334
rect 4228 10278 4296 10334
rect 4352 10278 4420 10334
rect 4476 10278 4544 10334
rect 4600 10278 4668 10334
rect 4724 10278 4734 10334
rect 2798 10210 4734 10278
rect 2798 10154 2808 10210
rect 2864 10154 2932 10210
rect 2988 10154 3056 10210
rect 3112 10154 3180 10210
rect 3236 10154 3304 10210
rect 3360 10154 3428 10210
rect 3484 10154 3552 10210
rect 3608 10154 3676 10210
rect 3732 10154 3800 10210
rect 3856 10154 3924 10210
rect 3980 10154 4048 10210
rect 4104 10154 4172 10210
rect 4228 10154 4296 10210
rect 4352 10154 4420 10210
rect 4476 10154 4544 10210
rect 4600 10154 4668 10210
rect 4724 10154 4734 10210
rect 2798 10086 4734 10154
rect 2798 10030 2808 10086
rect 2864 10030 2932 10086
rect 2988 10030 3056 10086
rect 3112 10030 3180 10086
rect 3236 10030 3304 10086
rect 3360 10030 3428 10086
rect 3484 10030 3552 10086
rect 3608 10030 3676 10086
rect 3732 10030 3800 10086
rect 3856 10030 3924 10086
rect 3980 10030 4048 10086
rect 4104 10030 4172 10086
rect 4228 10030 4296 10086
rect 4352 10030 4420 10086
rect 4476 10030 4544 10086
rect 4600 10030 4668 10086
rect 4724 10030 4734 10086
rect 2798 9962 4734 10030
rect 2798 9906 2808 9962
rect 2864 9906 2932 9962
rect 2988 9906 3056 9962
rect 3112 9906 3180 9962
rect 3236 9906 3304 9962
rect 3360 9906 3428 9962
rect 3484 9906 3552 9962
rect 3608 9906 3676 9962
rect 3732 9906 3800 9962
rect 3856 9906 3924 9962
rect 3980 9906 4048 9962
rect 4104 9906 4172 9962
rect 4228 9906 4296 9962
rect 4352 9906 4420 9962
rect 4476 9906 4544 9962
rect 4600 9906 4668 9962
rect 4724 9906 4734 9962
rect 2798 9838 4734 9906
rect 2798 9782 2808 9838
rect 2864 9782 2932 9838
rect 2988 9782 3056 9838
rect 3112 9782 3180 9838
rect 3236 9782 3304 9838
rect 3360 9782 3428 9838
rect 3484 9782 3552 9838
rect 3608 9782 3676 9838
rect 3732 9782 3800 9838
rect 3856 9782 3924 9838
rect 3980 9782 4048 9838
rect 4104 9782 4172 9838
rect 4228 9782 4296 9838
rect 4352 9782 4420 9838
rect 4476 9782 4544 9838
rect 4600 9782 4668 9838
rect 4724 9782 4734 9838
rect 2798 9714 4734 9782
rect 2798 9658 2808 9714
rect 2864 9658 2932 9714
rect 2988 9658 3056 9714
rect 3112 9658 3180 9714
rect 3236 9658 3304 9714
rect 3360 9658 3428 9714
rect 3484 9658 3552 9714
rect 3608 9658 3676 9714
rect 3732 9658 3800 9714
rect 3856 9658 3924 9714
rect 3980 9658 4048 9714
rect 4104 9658 4172 9714
rect 4228 9658 4296 9714
rect 4352 9658 4420 9714
rect 4476 9658 4544 9714
rect 4600 9658 4668 9714
rect 4724 9658 4734 9714
rect 2798 9590 4734 9658
rect 2798 9534 2808 9590
rect 2864 9534 2932 9590
rect 2988 9534 3056 9590
rect 3112 9534 3180 9590
rect 3236 9534 3304 9590
rect 3360 9534 3428 9590
rect 3484 9534 3552 9590
rect 3608 9534 3676 9590
rect 3732 9534 3800 9590
rect 3856 9534 3924 9590
rect 3980 9534 4048 9590
rect 4104 9534 4172 9590
rect 4228 9534 4296 9590
rect 4352 9534 4420 9590
rect 4476 9534 4544 9590
rect 4600 9534 4668 9590
rect 4724 9534 4734 9590
rect 2798 9466 4734 9534
rect 2798 9410 2808 9466
rect 2864 9410 2932 9466
rect 2988 9410 3056 9466
rect 3112 9410 3180 9466
rect 3236 9410 3304 9466
rect 3360 9410 3428 9466
rect 3484 9410 3552 9466
rect 3608 9410 3676 9466
rect 3732 9410 3800 9466
rect 3856 9410 3924 9466
rect 3980 9410 4048 9466
rect 4104 9410 4172 9466
rect 4228 9410 4296 9466
rect 4352 9410 4420 9466
rect 4476 9410 4544 9466
rect 4600 9410 4668 9466
rect 4724 9410 4734 9466
rect 2798 9342 4734 9410
rect 2798 9286 2808 9342
rect 2864 9286 2932 9342
rect 2988 9286 3056 9342
rect 3112 9286 3180 9342
rect 3236 9286 3304 9342
rect 3360 9286 3428 9342
rect 3484 9286 3552 9342
rect 3608 9286 3676 9342
rect 3732 9286 3800 9342
rect 3856 9286 3924 9342
rect 3980 9286 4048 9342
rect 4104 9286 4172 9342
rect 4228 9286 4296 9342
rect 4352 9286 4420 9342
rect 4476 9286 4544 9342
rect 4600 9286 4668 9342
rect 4724 9286 4734 9342
rect 2798 9218 4734 9286
rect 2798 9162 2808 9218
rect 2864 9162 2932 9218
rect 2988 9162 3056 9218
rect 3112 9162 3180 9218
rect 3236 9162 3304 9218
rect 3360 9162 3428 9218
rect 3484 9162 3552 9218
rect 3608 9162 3676 9218
rect 3732 9162 3800 9218
rect 3856 9162 3924 9218
rect 3980 9162 4048 9218
rect 4104 9162 4172 9218
rect 4228 9162 4296 9218
rect 4352 9162 4420 9218
rect 4476 9162 4544 9218
rect 4600 9162 4668 9218
rect 4724 9162 4734 9218
rect 2798 9094 4734 9162
rect 2798 9038 2808 9094
rect 2864 9038 2932 9094
rect 2988 9038 3056 9094
rect 3112 9038 3180 9094
rect 3236 9038 3304 9094
rect 3360 9038 3428 9094
rect 3484 9038 3552 9094
rect 3608 9038 3676 9094
rect 3732 9038 3800 9094
rect 3856 9038 3924 9094
rect 3980 9038 4048 9094
rect 4104 9038 4172 9094
rect 4228 9038 4296 9094
rect 4352 9038 4420 9094
rect 4476 9038 4544 9094
rect 4600 9038 4668 9094
rect 4724 9038 4734 9094
rect 2798 8970 4734 9038
rect 2798 8914 2808 8970
rect 2864 8914 2932 8970
rect 2988 8914 3056 8970
rect 3112 8914 3180 8970
rect 3236 8914 3304 8970
rect 3360 8914 3428 8970
rect 3484 8914 3552 8970
rect 3608 8914 3676 8970
rect 3732 8914 3800 8970
rect 3856 8914 3924 8970
rect 3980 8914 4048 8970
rect 4104 8914 4172 8970
rect 4228 8914 4296 8970
rect 4352 8914 4420 8970
rect 4476 8914 4544 8970
rect 4600 8914 4668 8970
rect 4724 8914 4734 8970
rect 2798 8846 4734 8914
rect 2798 8790 2808 8846
rect 2864 8790 2932 8846
rect 2988 8790 3056 8846
rect 3112 8790 3180 8846
rect 3236 8790 3304 8846
rect 3360 8790 3428 8846
rect 3484 8790 3552 8846
rect 3608 8790 3676 8846
rect 3732 8790 3800 8846
rect 3856 8790 3924 8846
rect 3980 8790 4048 8846
rect 4104 8790 4172 8846
rect 4228 8790 4296 8846
rect 4352 8790 4420 8846
rect 4476 8790 4544 8846
rect 4600 8790 4668 8846
rect 4724 8790 4734 8846
rect 2798 8722 4734 8790
rect 2798 8666 2808 8722
rect 2864 8666 2932 8722
rect 2988 8666 3056 8722
rect 3112 8666 3180 8722
rect 3236 8666 3304 8722
rect 3360 8666 3428 8722
rect 3484 8666 3552 8722
rect 3608 8666 3676 8722
rect 3732 8666 3800 8722
rect 3856 8666 3924 8722
rect 3980 8666 4048 8722
rect 4104 8666 4172 8722
rect 4228 8666 4296 8722
rect 4352 8666 4420 8722
rect 4476 8666 4544 8722
rect 4600 8666 4668 8722
rect 4724 8666 4734 8722
rect 2798 8598 4734 8666
rect 2798 8542 2808 8598
rect 2864 8542 2932 8598
rect 2988 8542 3056 8598
rect 3112 8542 3180 8598
rect 3236 8542 3304 8598
rect 3360 8542 3428 8598
rect 3484 8542 3552 8598
rect 3608 8542 3676 8598
rect 3732 8542 3800 8598
rect 3856 8542 3924 8598
rect 3980 8542 4048 8598
rect 4104 8542 4172 8598
rect 4228 8542 4296 8598
rect 4352 8542 4420 8598
rect 4476 8542 4544 8598
rect 4600 8542 4668 8598
rect 4724 8542 4734 8598
rect 2798 8474 4734 8542
rect 2798 8418 2808 8474
rect 2864 8418 2932 8474
rect 2988 8418 3056 8474
rect 3112 8418 3180 8474
rect 3236 8418 3304 8474
rect 3360 8418 3428 8474
rect 3484 8418 3552 8474
rect 3608 8418 3676 8474
rect 3732 8418 3800 8474
rect 3856 8418 3924 8474
rect 3980 8418 4048 8474
rect 4104 8418 4172 8474
rect 4228 8418 4296 8474
rect 4352 8418 4420 8474
rect 4476 8418 4544 8474
rect 4600 8418 4668 8474
rect 4724 8418 4734 8474
rect 2798 8350 4734 8418
rect 2798 8294 2808 8350
rect 2864 8294 2932 8350
rect 2988 8294 3056 8350
rect 3112 8294 3180 8350
rect 3236 8294 3304 8350
rect 3360 8294 3428 8350
rect 3484 8294 3552 8350
rect 3608 8294 3676 8350
rect 3732 8294 3800 8350
rect 3856 8294 3924 8350
rect 3980 8294 4048 8350
rect 4104 8294 4172 8350
rect 4228 8294 4296 8350
rect 4352 8294 4420 8350
rect 4476 8294 4544 8350
rect 4600 8294 4668 8350
rect 4724 8294 4734 8350
rect 2798 8226 4734 8294
rect 2798 8170 2808 8226
rect 2864 8170 2932 8226
rect 2988 8170 3056 8226
rect 3112 8170 3180 8226
rect 3236 8170 3304 8226
rect 3360 8170 3428 8226
rect 3484 8170 3552 8226
rect 3608 8170 3676 8226
rect 3732 8170 3800 8226
rect 3856 8170 3924 8226
rect 3980 8170 4048 8226
rect 4104 8170 4172 8226
rect 4228 8170 4296 8226
rect 4352 8170 4420 8226
rect 4476 8170 4544 8226
rect 4600 8170 4668 8226
rect 4724 8170 4734 8226
rect 2798 8102 4734 8170
rect 2798 8046 2808 8102
rect 2864 8046 2932 8102
rect 2988 8046 3056 8102
rect 3112 8046 3180 8102
rect 3236 8046 3304 8102
rect 3360 8046 3428 8102
rect 3484 8046 3552 8102
rect 3608 8046 3676 8102
rect 3732 8046 3800 8102
rect 3856 8046 3924 8102
rect 3980 8046 4048 8102
rect 4104 8046 4172 8102
rect 4228 8046 4296 8102
rect 4352 8046 4420 8102
rect 4476 8046 4544 8102
rect 4600 8046 4668 8102
rect 4724 8046 4734 8102
rect 2798 8036 4734 8046
rect 5168 10954 7104 10964
rect 5168 10898 5178 10954
rect 5234 10898 5302 10954
rect 5358 10898 5426 10954
rect 5482 10898 5550 10954
rect 5606 10898 5674 10954
rect 5730 10898 5798 10954
rect 5854 10898 5922 10954
rect 5978 10898 6046 10954
rect 6102 10898 6170 10954
rect 6226 10898 6294 10954
rect 6350 10898 6418 10954
rect 6474 10898 6542 10954
rect 6598 10898 6666 10954
rect 6722 10898 6790 10954
rect 6846 10898 6914 10954
rect 6970 10898 7038 10954
rect 7094 10898 7104 10954
rect 5168 10830 7104 10898
rect 5168 10774 5178 10830
rect 5234 10774 5302 10830
rect 5358 10774 5426 10830
rect 5482 10774 5550 10830
rect 5606 10774 5674 10830
rect 5730 10774 5798 10830
rect 5854 10774 5922 10830
rect 5978 10774 6046 10830
rect 6102 10774 6170 10830
rect 6226 10774 6294 10830
rect 6350 10774 6418 10830
rect 6474 10774 6542 10830
rect 6598 10774 6666 10830
rect 6722 10774 6790 10830
rect 6846 10774 6914 10830
rect 6970 10774 7038 10830
rect 7094 10774 7104 10830
rect 5168 10706 7104 10774
rect 5168 10650 5178 10706
rect 5234 10650 5302 10706
rect 5358 10650 5426 10706
rect 5482 10650 5550 10706
rect 5606 10650 5674 10706
rect 5730 10650 5798 10706
rect 5854 10650 5922 10706
rect 5978 10650 6046 10706
rect 6102 10650 6170 10706
rect 6226 10650 6294 10706
rect 6350 10650 6418 10706
rect 6474 10650 6542 10706
rect 6598 10650 6666 10706
rect 6722 10650 6790 10706
rect 6846 10650 6914 10706
rect 6970 10650 7038 10706
rect 7094 10650 7104 10706
rect 5168 10582 7104 10650
rect 5168 10526 5178 10582
rect 5234 10526 5302 10582
rect 5358 10526 5426 10582
rect 5482 10526 5550 10582
rect 5606 10526 5674 10582
rect 5730 10526 5798 10582
rect 5854 10526 5922 10582
rect 5978 10526 6046 10582
rect 6102 10526 6170 10582
rect 6226 10526 6294 10582
rect 6350 10526 6418 10582
rect 6474 10526 6542 10582
rect 6598 10526 6666 10582
rect 6722 10526 6790 10582
rect 6846 10526 6914 10582
rect 6970 10526 7038 10582
rect 7094 10526 7104 10582
rect 5168 10458 7104 10526
rect 5168 10402 5178 10458
rect 5234 10402 5302 10458
rect 5358 10402 5426 10458
rect 5482 10402 5550 10458
rect 5606 10402 5674 10458
rect 5730 10402 5798 10458
rect 5854 10402 5922 10458
rect 5978 10402 6046 10458
rect 6102 10402 6170 10458
rect 6226 10402 6294 10458
rect 6350 10402 6418 10458
rect 6474 10402 6542 10458
rect 6598 10402 6666 10458
rect 6722 10402 6790 10458
rect 6846 10402 6914 10458
rect 6970 10402 7038 10458
rect 7094 10402 7104 10458
rect 5168 10334 7104 10402
rect 5168 10278 5178 10334
rect 5234 10278 5302 10334
rect 5358 10278 5426 10334
rect 5482 10278 5550 10334
rect 5606 10278 5674 10334
rect 5730 10278 5798 10334
rect 5854 10278 5922 10334
rect 5978 10278 6046 10334
rect 6102 10278 6170 10334
rect 6226 10278 6294 10334
rect 6350 10278 6418 10334
rect 6474 10278 6542 10334
rect 6598 10278 6666 10334
rect 6722 10278 6790 10334
rect 6846 10278 6914 10334
rect 6970 10278 7038 10334
rect 7094 10278 7104 10334
rect 5168 10210 7104 10278
rect 5168 10154 5178 10210
rect 5234 10154 5302 10210
rect 5358 10154 5426 10210
rect 5482 10154 5550 10210
rect 5606 10154 5674 10210
rect 5730 10154 5798 10210
rect 5854 10154 5922 10210
rect 5978 10154 6046 10210
rect 6102 10154 6170 10210
rect 6226 10154 6294 10210
rect 6350 10154 6418 10210
rect 6474 10154 6542 10210
rect 6598 10154 6666 10210
rect 6722 10154 6790 10210
rect 6846 10154 6914 10210
rect 6970 10154 7038 10210
rect 7094 10154 7104 10210
rect 5168 10086 7104 10154
rect 5168 10030 5178 10086
rect 5234 10030 5302 10086
rect 5358 10030 5426 10086
rect 5482 10030 5550 10086
rect 5606 10030 5674 10086
rect 5730 10030 5798 10086
rect 5854 10030 5922 10086
rect 5978 10030 6046 10086
rect 6102 10030 6170 10086
rect 6226 10030 6294 10086
rect 6350 10030 6418 10086
rect 6474 10030 6542 10086
rect 6598 10030 6666 10086
rect 6722 10030 6790 10086
rect 6846 10030 6914 10086
rect 6970 10030 7038 10086
rect 7094 10030 7104 10086
rect 5168 9962 7104 10030
rect 5168 9906 5178 9962
rect 5234 9906 5302 9962
rect 5358 9906 5426 9962
rect 5482 9906 5550 9962
rect 5606 9906 5674 9962
rect 5730 9906 5798 9962
rect 5854 9906 5922 9962
rect 5978 9906 6046 9962
rect 6102 9906 6170 9962
rect 6226 9906 6294 9962
rect 6350 9906 6418 9962
rect 6474 9906 6542 9962
rect 6598 9906 6666 9962
rect 6722 9906 6790 9962
rect 6846 9906 6914 9962
rect 6970 9906 7038 9962
rect 7094 9906 7104 9962
rect 5168 9838 7104 9906
rect 5168 9782 5178 9838
rect 5234 9782 5302 9838
rect 5358 9782 5426 9838
rect 5482 9782 5550 9838
rect 5606 9782 5674 9838
rect 5730 9782 5798 9838
rect 5854 9782 5922 9838
rect 5978 9782 6046 9838
rect 6102 9782 6170 9838
rect 6226 9782 6294 9838
rect 6350 9782 6418 9838
rect 6474 9782 6542 9838
rect 6598 9782 6666 9838
rect 6722 9782 6790 9838
rect 6846 9782 6914 9838
rect 6970 9782 7038 9838
rect 7094 9782 7104 9838
rect 5168 9714 7104 9782
rect 5168 9658 5178 9714
rect 5234 9658 5302 9714
rect 5358 9658 5426 9714
rect 5482 9658 5550 9714
rect 5606 9658 5674 9714
rect 5730 9658 5798 9714
rect 5854 9658 5922 9714
rect 5978 9658 6046 9714
rect 6102 9658 6170 9714
rect 6226 9658 6294 9714
rect 6350 9658 6418 9714
rect 6474 9658 6542 9714
rect 6598 9658 6666 9714
rect 6722 9658 6790 9714
rect 6846 9658 6914 9714
rect 6970 9658 7038 9714
rect 7094 9658 7104 9714
rect 5168 9590 7104 9658
rect 5168 9534 5178 9590
rect 5234 9534 5302 9590
rect 5358 9534 5426 9590
rect 5482 9534 5550 9590
rect 5606 9534 5674 9590
rect 5730 9534 5798 9590
rect 5854 9534 5922 9590
rect 5978 9534 6046 9590
rect 6102 9534 6170 9590
rect 6226 9534 6294 9590
rect 6350 9534 6418 9590
rect 6474 9534 6542 9590
rect 6598 9534 6666 9590
rect 6722 9534 6790 9590
rect 6846 9534 6914 9590
rect 6970 9534 7038 9590
rect 7094 9534 7104 9590
rect 5168 9466 7104 9534
rect 5168 9410 5178 9466
rect 5234 9410 5302 9466
rect 5358 9410 5426 9466
rect 5482 9410 5550 9466
rect 5606 9410 5674 9466
rect 5730 9410 5798 9466
rect 5854 9410 5922 9466
rect 5978 9410 6046 9466
rect 6102 9410 6170 9466
rect 6226 9410 6294 9466
rect 6350 9410 6418 9466
rect 6474 9410 6542 9466
rect 6598 9410 6666 9466
rect 6722 9410 6790 9466
rect 6846 9410 6914 9466
rect 6970 9410 7038 9466
rect 7094 9410 7104 9466
rect 5168 9342 7104 9410
rect 5168 9286 5178 9342
rect 5234 9286 5302 9342
rect 5358 9286 5426 9342
rect 5482 9286 5550 9342
rect 5606 9286 5674 9342
rect 5730 9286 5798 9342
rect 5854 9286 5922 9342
rect 5978 9286 6046 9342
rect 6102 9286 6170 9342
rect 6226 9286 6294 9342
rect 6350 9286 6418 9342
rect 6474 9286 6542 9342
rect 6598 9286 6666 9342
rect 6722 9286 6790 9342
rect 6846 9286 6914 9342
rect 6970 9286 7038 9342
rect 7094 9286 7104 9342
rect 5168 9218 7104 9286
rect 5168 9162 5178 9218
rect 5234 9162 5302 9218
rect 5358 9162 5426 9218
rect 5482 9162 5550 9218
rect 5606 9162 5674 9218
rect 5730 9162 5798 9218
rect 5854 9162 5922 9218
rect 5978 9162 6046 9218
rect 6102 9162 6170 9218
rect 6226 9162 6294 9218
rect 6350 9162 6418 9218
rect 6474 9162 6542 9218
rect 6598 9162 6666 9218
rect 6722 9162 6790 9218
rect 6846 9162 6914 9218
rect 6970 9162 7038 9218
rect 7094 9162 7104 9218
rect 5168 9094 7104 9162
rect 5168 9038 5178 9094
rect 5234 9038 5302 9094
rect 5358 9038 5426 9094
rect 5482 9038 5550 9094
rect 5606 9038 5674 9094
rect 5730 9038 5798 9094
rect 5854 9038 5922 9094
rect 5978 9038 6046 9094
rect 6102 9038 6170 9094
rect 6226 9038 6294 9094
rect 6350 9038 6418 9094
rect 6474 9038 6542 9094
rect 6598 9038 6666 9094
rect 6722 9038 6790 9094
rect 6846 9038 6914 9094
rect 6970 9038 7038 9094
rect 7094 9038 7104 9094
rect 5168 8970 7104 9038
rect 5168 8914 5178 8970
rect 5234 8914 5302 8970
rect 5358 8914 5426 8970
rect 5482 8914 5550 8970
rect 5606 8914 5674 8970
rect 5730 8914 5798 8970
rect 5854 8914 5922 8970
rect 5978 8914 6046 8970
rect 6102 8914 6170 8970
rect 6226 8914 6294 8970
rect 6350 8914 6418 8970
rect 6474 8914 6542 8970
rect 6598 8914 6666 8970
rect 6722 8914 6790 8970
rect 6846 8914 6914 8970
rect 6970 8914 7038 8970
rect 7094 8914 7104 8970
rect 5168 8846 7104 8914
rect 5168 8790 5178 8846
rect 5234 8790 5302 8846
rect 5358 8790 5426 8846
rect 5482 8790 5550 8846
rect 5606 8790 5674 8846
rect 5730 8790 5798 8846
rect 5854 8790 5922 8846
rect 5978 8790 6046 8846
rect 6102 8790 6170 8846
rect 6226 8790 6294 8846
rect 6350 8790 6418 8846
rect 6474 8790 6542 8846
rect 6598 8790 6666 8846
rect 6722 8790 6790 8846
rect 6846 8790 6914 8846
rect 6970 8790 7038 8846
rect 7094 8790 7104 8846
rect 5168 8722 7104 8790
rect 5168 8666 5178 8722
rect 5234 8666 5302 8722
rect 5358 8666 5426 8722
rect 5482 8666 5550 8722
rect 5606 8666 5674 8722
rect 5730 8666 5798 8722
rect 5854 8666 5922 8722
rect 5978 8666 6046 8722
rect 6102 8666 6170 8722
rect 6226 8666 6294 8722
rect 6350 8666 6418 8722
rect 6474 8666 6542 8722
rect 6598 8666 6666 8722
rect 6722 8666 6790 8722
rect 6846 8666 6914 8722
rect 6970 8666 7038 8722
rect 7094 8666 7104 8722
rect 5168 8598 7104 8666
rect 5168 8542 5178 8598
rect 5234 8542 5302 8598
rect 5358 8542 5426 8598
rect 5482 8542 5550 8598
rect 5606 8542 5674 8598
rect 5730 8542 5798 8598
rect 5854 8542 5922 8598
rect 5978 8542 6046 8598
rect 6102 8542 6170 8598
rect 6226 8542 6294 8598
rect 6350 8542 6418 8598
rect 6474 8542 6542 8598
rect 6598 8542 6666 8598
rect 6722 8542 6790 8598
rect 6846 8542 6914 8598
rect 6970 8542 7038 8598
rect 7094 8542 7104 8598
rect 5168 8474 7104 8542
rect 5168 8418 5178 8474
rect 5234 8418 5302 8474
rect 5358 8418 5426 8474
rect 5482 8418 5550 8474
rect 5606 8418 5674 8474
rect 5730 8418 5798 8474
rect 5854 8418 5922 8474
rect 5978 8418 6046 8474
rect 6102 8418 6170 8474
rect 6226 8418 6294 8474
rect 6350 8418 6418 8474
rect 6474 8418 6542 8474
rect 6598 8418 6666 8474
rect 6722 8418 6790 8474
rect 6846 8418 6914 8474
rect 6970 8418 7038 8474
rect 7094 8418 7104 8474
rect 5168 8350 7104 8418
rect 5168 8294 5178 8350
rect 5234 8294 5302 8350
rect 5358 8294 5426 8350
rect 5482 8294 5550 8350
rect 5606 8294 5674 8350
rect 5730 8294 5798 8350
rect 5854 8294 5922 8350
rect 5978 8294 6046 8350
rect 6102 8294 6170 8350
rect 6226 8294 6294 8350
rect 6350 8294 6418 8350
rect 6474 8294 6542 8350
rect 6598 8294 6666 8350
rect 6722 8294 6790 8350
rect 6846 8294 6914 8350
rect 6970 8294 7038 8350
rect 7094 8294 7104 8350
rect 5168 8226 7104 8294
rect 5168 8170 5178 8226
rect 5234 8170 5302 8226
rect 5358 8170 5426 8226
rect 5482 8170 5550 8226
rect 5606 8170 5674 8226
rect 5730 8170 5798 8226
rect 5854 8170 5922 8226
rect 5978 8170 6046 8226
rect 6102 8170 6170 8226
rect 6226 8170 6294 8226
rect 6350 8170 6418 8226
rect 6474 8170 6542 8226
rect 6598 8170 6666 8226
rect 6722 8170 6790 8226
rect 6846 8170 6914 8226
rect 6970 8170 7038 8226
rect 7094 8170 7104 8226
rect 5168 8102 7104 8170
rect 5168 8046 5178 8102
rect 5234 8046 5302 8102
rect 5358 8046 5426 8102
rect 5482 8046 5550 8102
rect 5606 8046 5674 8102
rect 5730 8046 5798 8102
rect 5854 8046 5922 8102
rect 5978 8046 6046 8102
rect 6102 8046 6170 8102
rect 6226 8046 6294 8102
rect 6350 8046 6418 8102
rect 6474 8046 6542 8102
rect 6598 8046 6666 8102
rect 6722 8046 6790 8102
rect 6846 8046 6914 8102
rect 6970 8046 7038 8102
rect 7094 8046 7104 8102
rect 5168 8036 7104 8046
rect 7874 10954 9810 10964
rect 7874 10898 7884 10954
rect 7940 10898 8008 10954
rect 8064 10898 8132 10954
rect 8188 10898 8256 10954
rect 8312 10898 8380 10954
rect 8436 10898 8504 10954
rect 8560 10898 8628 10954
rect 8684 10898 8752 10954
rect 8808 10898 8876 10954
rect 8932 10898 9000 10954
rect 9056 10898 9124 10954
rect 9180 10898 9248 10954
rect 9304 10898 9372 10954
rect 9428 10898 9496 10954
rect 9552 10898 9620 10954
rect 9676 10898 9744 10954
rect 9800 10898 9810 10954
rect 7874 10830 9810 10898
rect 7874 10774 7884 10830
rect 7940 10774 8008 10830
rect 8064 10774 8132 10830
rect 8188 10774 8256 10830
rect 8312 10774 8380 10830
rect 8436 10774 8504 10830
rect 8560 10774 8628 10830
rect 8684 10774 8752 10830
rect 8808 10774 8876 10830
rect 8932 10774 9000 10830
rect 9056 10774 9124 10830
rect 9180 10774 9248 10830
rect 9304 10774 9372 10830
rect 9428 10774 9496 10830
rect 9552 10774 9620 10830
rect 9676 10774 9744 10830
rect 9800 10774 9810 10830
rect 7874 10706 9810 10774
rect 7874 10650 7884 10706
rect 7940 10650 8008 10706
rect 8064 10650 8132 10706
rect 8188 10650 8256 10706
rect 8312 10650 8380 10706
rect 8436 10650 8504 10706
rect 8560 10650 8628 10706
rect 8684 10650 8752 10706
rect 8808 10650 8876 10706
rect 8932 10650 9000 10706
rect 9056 10650 9124 10706
rect 9180 10650 9248 10706
rect 9304 10650 9372 10706
rect 9428 10650 9496 10706
rect 9552 10650 9620 10706
rect 9676 10650 9744 10706
rect 9800 10650 9810 10706
rect 7874 10582 9810 10650
rect 7874 10526 7884 10582
rect 7940 10526 8008 10582
rect 8064 10526 8132 10582
rect 8188 10526 8256 10582
rect 8312 10526 8380 10582
rect 8436 10526 8504 10582
rect 8560 10526 8628 10582
rect 8684 10526 8752 10582
rect 8808 10526 8876 10582
rect 8932 10526 9000 10582
rect 9056 10526 9124 10582
rect 9180 10526 9248 10582
rect 9304 10526 9372 10582
rect 9428 10526 9496 10582
rect 9552 10526 9620 10582
rect 9676 10526 9744 10582
rect 9800 10526 9810 10582
rect 7874 10458 9810 10526
rect 7874 10402 7884 10458
rect 7940 10402 8008 10458
rect 8064 10402 8132 10458
rect 8188 10402 8256 10458
rect 8312 10402 8380 10458
rect 8436 10402 8504 10458
rect 8560 10402 8628 10458
rect 8684 10402 8752 10458
rect 8808 10402 8876 10458
rect 8932 10402 9000 10458
rect 9056 10402 9124 10458
rect 9180 10402 9248 10458
rect 9304 10402 9372 10458
rect 9428 10402 9496 10458
rect 9552 10402 9620 10458
rect 9676 10402 9744 10458
rect 9800 10402 9810 10458
rect 7874 10334 9810 10402
rect 7874 10278 7884 10334
rect 7940 10278 8008 10334
rect 8064 10278 8132 10334
rect 8188 10278 8256 10334
rect 8312 10278 8380 10334
rect 8436 10278 8504 10334
rect 8560 10278 8628 10334
rect 8684 10278 8752 10334
rect 8808 10278 8876 10334
rect 8932 10278 9000 10334
rect 9056 10278 9124 10334
rect 9180 10278 9248 10334
rect 9304 10278 9372 10334
rect 9428 10278 9496 10334
rect 9552 10278 9620 10334
rect 9676 10278 9744 10334
rect 9800 10278 9810 10334
rect 7874 10210 9810 10278
rect 7874 10154 7884 10210
rect 7940 10154 8008 10210
rect 8064 10154 8132 10210
rect 8188 10154 8256 10210
rect 8312 10154 8380 10210
rect 8436 10154 8504 10210
rect 8560 10154 8628 10210
rect 8684 10154 8752 10210
rect 8808 10154 8876 10210
rect 8932 10154 9000 10210
rect 9056 10154 9124 10210
rect 9180 10154 9248 10210
rect 9304 10154 9372 10210
rect 9428 10154 9496 10210
rect 9552 10154 9620 10210
rect 9676 10154 9744 10210
rect 9800 10154 9810 10210
rect 7874 10086 9810 10154
rect 7874 10030 7884 10086
rect 7940 10030 8008 10086
rect 8064 10030 8132 10086
rect 8188 10030 8256 10086
rect 8312 10030 8380 10086
rect 8436 10030 8504 10086
rect 8560 10030 8628 10086
rect 8684 10030 8752 10086
rect 8808 10030 8876 10086
rect 8932 10030 9000 10086
rect 9056 10030 9124 10086
rect 9180 10030 9248 10086
rect 9304 10030 9372 10086
rect 9428 10030 9496 10086
rect 9552 10030 9620 10086
rect 9676 10030 9744 10086
rect 9800 10030 9810 10086
rect 7874 9962 9810 10030
rect 7874 9906 7884 9962
rect 7940 9906 8008 9962
rect 8064 9906 8132 9962
rect 8188 9906 8256 9962
rect 8312 9906 8380 9962
rect 8436 9906 8504 9962
rect 8560 9906 8628 9962
rect 8684 9906 8752 9962
rect 8808 9906 8876 9962
rect 8932 9906 9000 9962
rect 9056 9906 9124 9962
rect 9180 9906 9248 9962
rect 9304 9906 9372 9962
rect 9428 9906 9496 9962
rect 9552 9906 9620 9962
rect 9676 9906 9744 9962
rect 9800 9906 9810 9962
rect 7874 9838 9810 9906
rect 7874 9782 7884 9838
rect 7940 9782 8008 9838
rect 8064 9782 8132 9838
rect 8188 9782 8256 9838
rect 8312 9782 8380 9838
rect 8436 9782 8504 9838
rect 8560 9782 8628 9838
rect 8684 9782 8752 9838
rect 8808 9782 8876 9838
rect 8932 9782 9000 9838
rect 9056 9782 9124 9838
rect 9180 9782 9248 9838
rect 9304 9782 9372 9838
rect 9428 9782 9496 9838
rect 9552 9782 9620 9838
rect 9676 9782 9744 9838
rect 9800 9782 9810 9838
rect 7874 9714 9810 9782
rect 7874 9658 7884 9714
rect 7940 9658 8008 9714
rect 8064 9658 8132 9714
rect 8188 9658 8256 9714
rect 8312 9658 8380 9714
rect 8436 9658 8504 9714
rect 8560 9658 8628 9714
rect 8684 9658 8752 9714
rect 8808 9658 8876 9714
rect 8932 9658 9000 9714
rect 9056 9658 9124 9714
rect 9180 9658 9248 9714
rect 9304 9658 9372 9714
rect 9428 9658 9496 9714
rect 9552 9658 9620 9714
rect 9676 9658 9744 9714
rect 9800 9658 9810 9714
rect 7874 9590 9810 9658
rect 7874 9534 7884 9590
rect 7940 9534 8008 9590
rect 8064 9534 8132 9590
rect 8188 9534 8256 9590
rect 8312 9534 8380 9590
rect 8436 9534 8504 9590
rect 8560 9534 8628 9590
rect 8684 9534 8752 9590
rect 8808 9534 8876 9590
rect 8932 9534 9000 9590
rect 9056 9534 9124 9590
rect 9180 9534 9248 9590
rect 9304 9534 9372 9590
rect 9428 9534 9496 9590
rect 9552 9534 9620 9590
rect 9676 9534 9744 9590
rect 9800 9534 9810 9590
rect 7874 9466 9810 9534
rect 7874 9410 7884 9466
rect 7940 9410 8008 9466
rect 8064 9410 8132 9466
rect 8188 9410 8256 9466
rect 8312 9410 8380 9466
rect 8436 9410 8504 9466
rect 8560 9410 8628 9466
rect 8684 9410 8752 9466
rect 8808 9410 8876 9466
rect 8932 9410 9000 9466
rect 9056 9410 9124 9466
rect 9180 9410 9248 9466
rect 9304 9410 9372 9466
rect 9428 9410 9496 9466
rect 9552 9410 9620 9466
rect 9676 9410 9744 9466
rect 9800 9410 9810 9466
rect 7874 9342 9810 9410
rect 7874 9286 7884 9342
rect 7940 9286 8008 9342
rect 8064 9286 8132 9342
rect 8188 9286 8256 9342
rect 8312 9286 8380 9342
rect 8436 9286 8504 9342
rect 8560 9286 8628 9342
rect 8684 9286 8752 9342
rect 8808 9286 8876 9342
rect 8932 9286 9000 9342
rect 9056 9286 9124 9342
rect 9180 9286 9248 9342
rect 9304 9286 9372 9342
rect 9428 9286 9496 9342
rect 9552 9286 9620 9342
rect 9676 9286 9744 9342
rect 9800 9286 9810 9342
rect 7874 9218 9810 9286
rect 7874 9162 7884 9218
rect 7940 9162 8008 9218
rect 8064 9162 8132 9218
rect 8188 9162 8256 9218
rect 8312 9162 8380 9218
rect 8436 9162 8504 9218
rect 8560 9162 8628 9218
rect 8684 9162 8752 9218
rect 8808 9162 8876 9218
rect 8932 9162 9000 9218
rect 9056 9162 9124 9218
rect 9180 9162 9248 9218
rect 9304 9162 9372 9218
rect 9428 9162 9496 9218
rect 9552 9162 9620 9218
rect 9676 9162 9744 9218
rect 9800 9162 9810 9218
rect 7874 9094 9810 9162
rect 7874 9038 7884 9094
rect 7940 9038 8008 9094
rect 8064 9038 8132 9094
rect 8188 9038 8256 9094
rect 8312 9038 8380 9094
rect 8436 9038 8504 9094
rect 8560 9038 8628 9094
rect 8684 9038 8752 9094
rect 8808 9038 8876 9094
rect 8932 9038 9000 9094
rect 9056 9038 9124 9094
rect 9180 9038 9248 9094
rect 9304 9038 9372 9094
rect 9428 9038 9496 9094
rect 9552 9038 9620 9094
rect 9676 9038 9744 9094
rect 9800 9038 9810 9094
rect 7874 8970 9810 9038
rect 7874 8914 7884 8970
rect 7940 8914 8008 8970
rect 8064 8914 8132 8970
rect 8188 8914 8256 8970
rect 8312 8914 8380 8970
rect 8436 8914 8504 8970
rect 8560 8914 8628 8970
rect 8684 8914 8752 8970
rect 8808 8914 8876 8970
rect 8932 8914 9000 8970
rect 9056 8914 9124 8970
rect 9180 8914 9248 8970
rect 9304 8914 9372 8970
rect 9428 8914 9496 8970
rect 9552 8914 9620 8970
rect 9676 8914 9744 8970
rect 9800 8914 9810 8970
rect 7874 8846 9810 8914
rect 7874 8790 7884 8846
rect 7940 8790 8008 8846
rect 8064 8790 8132 8846
rect 8188 8790 8256 8846
rect 8312 8790 8380 8846
rect 8436 8790 8504 8846
rect 8560 8790 8628 8846
rect 8684 8790 8752 8846
rect 8808 8790 8876 8846
rect 8932 8790 9000 8846
rect 9056 8790 9124 8846
rect 9180 8790 9248 8846
rect 9304 8790 9372 8846
rect 9428 8790 9496 8846
rect 9552 8790 9620 8846
rect 9676 8790 9744 8846
rect 9800 8790 9810 8846
rect 7874 8722 9810 8790
rect 7874 8666 7884 8722
rect 7940 8666 8008 8722
rect 8064 8666 8132 8722
rect 8188 8666 8256 8722
rect 8312 8666 8380 8722
rect 8436 8666 8504 8722
rect 8560 8666 8628 8722
rect 8684 8666 8752 8722
rect 8808 8666 8876 8722
rect 8932 8666 9000 8722
rect 9056 8666 9124 8722
rect 9180 8666 9248 8722
rect 9304 8666 9372 8722
rect 9428 8666 9496 8722
rect 9552 8666 9620 8722
rect 9676 8666 9744 8722
rect 9800 8666 9810 8722
rect 7874 8598 9810 8666
rect 7874 8542 7884 8598
rect 7940 8542 8008 8598
rect 8064 8542 8132 8598
rect 8188 8542 8256 8598
rect 8312 8542 8380 8598
rect 8436 8542 8504 8598
rect 8560 8542 8628 8598
rect 8684 8542 8752 8598
rect 8808 8542 8876 8598
rect 8932 8542 9000 8598
rect 9056 8542 9124 8598
rect 9180 8542 9248 8598
rect 9304 8542 9372 8598
rect 9428 8542 9496 8598
rect 9552 8542 9620 8598
rect 9676 8542 9744 8598
rect 9800 8542 9810 8598
rect 7874 8474 9810 8542
rect 7874 8418 7884 8474
rect 7940 8418 8008 8474
rect 8064 8418 8132 8474
rect 8188 8418 8256 8474
rect 8312 8418 8380 8474
rect 8436 8418 8504 8474
rect 8560 8418 8628 8474
rect 8684 8418 8752 8474
rect 8808 8418 8876 8474
rect 8932 8418 9000 8474
rect 9056 8418 9124 8474
rect 9180 8418 9248 8474
rect 9304 8418 9372 8474
rect 9428 8418 9496 8474
rect 9552 8418 9620 8474
rect 9676 8418 9744 8474
rect 9800 8418 9810 8474
rect 7874 8350 9810 8418
rect 7874 8294 7884 8350
rect 7940 8294 8008 8350
rect 8064 8294 8132 8350
rect 8188 8294 8256 8350
rect 8312 8294 8380 8350
rect 8436 8294 8504 8350
rect 8560 8294 8628 8350
rect 8684 8294 8752 8350
rect 8808 8294 8876 8350
rect 8932 8294 9000 8350
rect 9056 8294 9124 8350
rect 9180 8294 9248 8350
rect 9304 8294 9372 8350
rect 9428 8294 9496 8350
rect 9552 8294 9620 8350
rect 9676 8294 9744 8350
rect 9800 8294 9810 8350
rect 7874 8226 9810 8294
rect 7874 8170 7884 8226
rect 7940 8170 8008 8226
rect 8064 8170 8132 8226
rect 8188 8170 8256 8226
rect 8312 8170 8380 8226
rect 8436 8170 8504 8226
rect 8560 8170 8628 8226
rect 8684 8170 8752 8226
rect 8808 8170 8876 8226
rect 8932 8170 9000 8226
rect 9056 8170 9124 8226
rect 9180 8170 9248 8226
rect 9304 8170 9372 8226
rect 9428 8170 9496 8226
rect 9552 8170 9620 8226
rect 9676 8170 9744 8226
rect 9800 8170 9810 8226
rect 7874 8102 9810 8170
rect 7874 8046 7884 8102
rect 7940 8046 8008 8102
rect 8064 8046 8132 8102
rect 8188 8046 8256 8102
rect 8312 8046 8380 8102
rect 8436 8046 8504 8102
rect 8560 8046 8628 8102
rect 8684 8046 8752 8102
rect 8808 8046 8876 8102
rect 8932 8046 9000 8102
rect 9056 8046 9124 8102
rect 9180 8046 9248 8102
rect 9304 8046 9372 8102
rect 9428 8046 9496 8102
rect 9552 8046 9620 8102
rect 9676 8046 9744 8102
rect 9800 8046 9810 8102
rect 7874 8036 9810 8046
rect 10244 10954 12180 10964
rect 10244 10898 10254 10954
rect 10310 10898 10378 10954
rect 10434 10898 10502 10954
rect 10558 10898 10626 10954
rect 10682 10898 10750 10954
rect 10806 10898 10874 10954
rect 10930 10898 10998 10954
rect 11054 10898 11122 10954
rect 11178 10898 11246 10954
rect 11302 10898 11370 10954
rect 11426 10898 11494 10954
rect 11550 10898 11618 10954
rect 11674 10898 11742 10954
rect 11798 10898 11866 10954
rect 11922 10898 11990 10954
rect 12046 10898 12114 10954
rect 12170 10898 12180 10954
rect 10244 10830 12180 10898
rect 10244 10774 10254 10830
rect 10310 10774 10378 10830
rect 10434 10774 10502 10830
rect 10558 10774 10626 10830
rect 10682 10774 10750 10830
rect 10806 10774 10874 10830
rect 10930 10774 10998 10830
rect 11054 10774 11122 10830
rect 11178 10774 11246 10830
rect 11302 10774 11370 10830
rect 11426 10774 11494 10830
rect 11550 10774 11618 10830
rect 11674 10774 11742 10830
rect 11798 10774 11866 10830
rect 11922 10774 11990 10830
rect 12046 10774 12114 10830
rect 12170 10774 12180 10830
rect 10244 10706 12180 10774
rect 10244 10650 10254 10706
rect 10310 10650 10378 10706
rect 10434 10650 10502 10706
rect 10558 10650 10626 10706
rect 10682 10650 10750 10706
rect 10806 10650 10874 10706
rect 10930 10650 10998 10706
rect 11054 10650 11122 10706
rect 11178 10650 11246 10706
rect 11302 10650 11370 10706
rect 11426 10650 11494 10706
rect 11550 10650 11618 10706
rect 11674 10650 11742 10706
rect 11798 10650 11866 10706
rect 11922 10650 11990 10706
rect 12046 10650 12114 10706
rect 12170 10650 12180 10706
rect 10244 10582 12180 10650
rect 10244 10526 10254 10582
rect 10310 10526 10378 10582
rect 10434 10526 10502 10582
rect 10558 10526 10626 10582
rect 10682 10526 10750 10582
rect 10806 10526 10874 10582
rect 10930 10526 10998 10582
rect 11054 10526 11122 10582
rect 11178 10526 11246 10582
rect 11302 10526 11370 10582
rect 11426 10526 11494 10582
rect 11550 10526 11618 10582
rect 11674 10526 11742 10582
rect 11798 10526 11866 10582
rect 11922 10526 11990 10582
rect 12046 10526 12114 10582
rect 12170 10526 12180 10582
rect 10244 10458 12180 10526
rect 10244 10402 10254 10458
rect 10310 10402 10378 10458
rect 10434 10402 10502 10458
rect 10558 10402 10626 10458
rect 10682 10402 10750 10458
rect 10806 10402 10874 10458
rect 10930 10402 10998 10458
rect 11054 10402 11122 10458
rect 11178 10402 11246 10458
rect 11302 10402 11370 10458
rect 11426 10402 11494 10458
rect 11550 10402 11618 10458
rect 11674 10402 11742 10458
rect 11798 10402 11866 10458
rect 11922 10402 11990 10458
rect 12046 10402 12114 10458
rect 12170 10402 12180 10458
rect 10244 10334 12180 10402
rect 10244 10278 10254 10334
rect 10310 10278 10378 10334
rect 10434 10278 10502 10334
rect 10558 10278 10626 10334
rect 10682 10278 10750 10334
rect 10806 10278 10874 10334
rect 10930 10278 10998 10334
rect 11054 10278 11122 10334
rect 11178 10278 11246 10334
rect 11302 10278 11370 10334
rect 11426 10278 11494 10334
rect 11550 10278 11618 10334
rect 11674 10278 11742 10334
rect 11798 10278 11866 10334
rect 11922 10278 11990 10334
rect 12046 10278 12114 10334
rect 12170 10278 12180 10334
rect 10244 10210 12180 10278
rect 10244 10154 10254 10210
rect 10310 10154 10378 10210
rect 10434 10154 10502 10210
rect 10558 10154 10626 10210
rect 10682 10154 10750 10210
rect 10806 10154 10874 10210
rect 10930 10154 10998 10210
rect 11054 10154 11122 10210
rect 11178 10154 11246 10210
rect 11302 10154 11370 10210
rect 11426 10154 11494 10210
rect 11550 10154 11618 10210
rect 11674 10154 11742 10210
rect 11798 10154 11866 10210
rect 11922 10154 11990 10210
rect 12046 10154 12114 10210
rect 12170 10154 12180 10210
rect 10244 10086 12180 10154
rect 10244 10030 10254 10086
rect 10310 10030 10378 10086
rect 10434 10030 10502 10086
rect 10558 10030 10626 10086
rect 10682 10030 10750 10086
rect 10806 10030 10874 10086
rect 10930 10030 10998 10086
rect 11054 10030 11122 10086
rect 11178 10030 11246 10086
rect 11302 10030 11370 10086
rect 11426 10030 11494 10086
rect 11550 10030 11618 10086
rect 11674 10030 11742 10086
rect 11798 10030 11866 10086
rect 11922 10030 11990 10086
rect 12046 10030 12114 10086
rect 12170 10030 12180 10086
rect 10244 9962 12180 10030
rect 10244 9906 10254 9962
rect 10310 9906 10378 9962
rect 10434 9906 10502 9962
rect 10558 9906 10626 9962
rect 10682 9906 10750 9962
rect 10806 9906 10874 9962
rect 10930 9906 10998 9962
rect 11054 9906 11122 9962
rect 11178 9906 11246 9962
rect 11302 9906 11370 9962
rect 11426 9906 11494 9962
rect 11550 9906 11618 9962
rect 11674 9906 11742 9962
rect 11798 9906 11866 9962
rect 11922 9906 11990 9962
rect 12046 9906 12114 9962
rect 12170 9906 12180 9962
rect 10244 9838 12180 9906
rect 10244 9782 10254 9838
rect 10310 9782 10378 9838
rect 10434 9782 10502 9838
rect 10558 9782 10626 9838
rect 10682 9782 10750 9838
rect 10806 9782 10874 9838
rect 10930 9782 10998 9838
rect 11054 9782 11122 9838
rect 11178 9782 11246 9838
rect 11302 9782 11370 9838
rect 11426 9782 11494 9838
rect 11550 9782 11618 9838
rect 11674 9782 11742 9838
rect 11798 9782 11866 9838
rect 11922 9782 11990 9838
rect 12046 9782 12114 9838
rect 12170 9782 12180 9838
rect 10244 9714 12180 9782
rect 10244 9658 10254 9714
rect 10310 9658 10378 9714
rect 10434 9658 10502 9714
rect 10558 9658 10626 9714
rect 10682 9658 10750 9714
rect 10806 9658 10874 9714
rect 10930 9658 10998 9714
rect 11054 9658 11122 9714
rect 11178 9658 11246 9714
rect 11302 9658 11370 9714
rect 11426 9658 11494 9714
rect 11550 9658 11618 9714
rect 11674 9658 11742 9714
rect 11798 9658 11866 9714
rect 11922 9658 11990 9714
rect 12046 9658 12114 9714
rect 12170 9658 12180 9714
rect 10244 9590 12180 9658
rect 10244 9534 10254 9590
rect 10310 9534 10378 9590
rect 10434 9534 10502 9590
rect 10558 9534 10626 9590
rect 10682 9534 10750 9590
rect 10806 9534 10874 9590
rect 10930 9534 10998 9590
rect 11054 9534 11122 9590
rect 11178 9534 11246 9590
rect 11302 9534 11370 9590
rect 11426 9534 11494 9590
rect 11550 9534 11618 9590
rect 11674 9534 11742 9590
rect 11798 9534 11866 9590
rect 11922 9534 11990 9590
rect 12046 9534 12114 9590
rect 12170 9534 12180 9590
rect 10244 9466 12180 9534
rect 10244 9410 10254 9466
rect 10310 9410 10378 9466
rect 10434 9410 10502 9466
rect 10558 9410 10626 9466
rect 10682 9410 10750 9466
rect 10806 9410 10874 9466
rect 10930 9410 10998 9466
rect 11054 9410 11122 9466
rect 11178 9410 11246 9466
rect 11302 9410 11370 9466
rect 11426 9410 11494 9466
rect 11550 9410 11618 9466
rect 11674 9410 11742 9466
rect 11798 9410 11866 9466
rect 11922 9410 11990 9466
rect 12046 9410 12114 9466
rect 12170 9410 12180 9466
rect 10244 9342 12180 9410
rect 10244 9286 10254 9342
rect 10310 9286 10378 9342
rect 10434 9286 10502 9342
rect 10558 9286 10626 9342
rect 10682 9286 10750 9342
rect 10806 9286 10874 9342
rect 10930 9286 10998 9342
rect 11054 9286 11122 9342
rect 11178 9286 11246 9342
rect 11302 9286 11370 9342
rect 11426 9286 11494 9342
rect 11550 9286 11618 9342
rect 11674 9286 11742 9342
rect 11798 9286 11866 9342
rect 11922 9286 11990 9342
rect 12046 9286 12114 9342
rect 12170 9286 12180 9342
rect 10244 9218 12180 9286
rect 10244 9162 10254 9218
rect 10310 9162 10378 9218
rect 10434 9162 10502 9218
rect 10558 9162 10626 9218
rect 10682 9162 10750 9218
rect 10806 9162 10874 9218
rect 10930 9162 10998 9218
rect 11054 9162 11122 9218
rect 11178 9162 11246 9218
rect 11302 9162 11370 9218
rect 11426 9162 11494 9218
rect 11550 9162 11618 9218
rect 11674 9162 11742 9218
rect 11798 9162 11866 9218
rect 11922 9162 11990 9218
rect 12046 9162 12114 9218
rect 12170 9162 12180 9218
rect 10244 9094 12180 9162
rect 10244 9038 10254 9094
rect 10310 9038 10378 9094
rect 10434 9038 10502 9094
rect 10558 9038 10626 9094
rect 10682 9038 10750 9094
rect 10806 9038 10874 9094
rect 10930 9038 10998 9094
rect 11054 9038 11122 9094
rect 11178 9038 11246 9094
rect 11302 9038 11370 9094
rect 11426 9038 11494 9094
rect 11550 9038 11618 9094
rect 11674 9038 11742 9094
rect 11798 9038 11866 9094
rect 11922 9038 11990 9094
rect 12046 9038 12114 9094
rect 12170 9038 12180 9094
rect 10244 8970 12180 9038
rect 10244 8914 10254 8970
rect 10310 8914 10378 8970
rect 10434 8914 10502 8970
rect 10558 8914 10626 8970
rect 10682 8914 10750 8970
rect 10806 8914 10874 8970
rect 10930 8914 10998 8970
rect 11054 8914 11122 8970
rect 11178 8914 11246 8970
rect 11302 8914 11370 8970
rect 11426 8914 11494 8970
rect 11550 8914 11618 8970
rect 11674 8914 11742 8970
rect 11798 8914 11866 8970
rect 11922 8914 11990 8970
rect 12046 8914 12114 8970
rect 12170 8914 12180 8970
rect 10244 8846 12180 8914
rect 10244 8790 10254 8846
rect 10310 8790 10378 8846
rect 10434 8790 10502 8846
rect 10558 8790 10626 8846
rect 10682 8790 10750 8846
rect 10806 8790 10874 8846
rect 10930 8790 10998 8846
rect 11054 8790 11122 8846
rect 11178 8790 11246 8846
rect 11302 8790 11370 8846
rect 11426 8790 11494 8846
rect 11550 8790 11618 8846
rect 11674 8790 11742 8846
rect 11798 8790 11866 8846
rect 11922 8790 11990 8846
rect 12046 8790 12114 8846
rect 12170 8790 12180 8846
rect 10244 8722 12180 8790
rect 10244 8666 10254 8722
rect 10310 8666 10378 8722
rect 10434 8666 10502 8722
rect 10558 8666 10626 8722
rect 10682 8666 10750 8722
rect 10806 8666 10874 8722
rect 10930 8666 10998 8722
rect 11054 8666 11122 8722
rect 11178 8666 11246 8722
rect 11302 8666 11370 8722
rect 11426 8666 11494 8722
rect 11550 8666 11618 8722
rect 11674 8666 11742 8722
rect 11798 8666 11866 8722
rect 11922 8666 11990 8722
rect 12046 8666 12114 8722
rect 12170 8666 12180 8722
rect 10244 8598 12180 8666
rect 10244 8542 10254 8598
rect 10310 8542 10378 8598
rect 10434 8542 10502 8598
rect 10558 8542 10626 8598
rect 10682 8542 10750 8598
rect 10806 8542 10874 8598
rect 10930 8542 10998 8598
rect 11054 8542 11122 8598
rect 11178 8542 11246 8598
rect 11302 8542 11370 8598
rect 11426 8542 11494 8598
rect 11550 8542 11618 8598
rect 11674 8542 11742 8598
rect 11798 8542 11866 8598
rect 11922 8542 11990 8598
rect 12046 8542 12114 8598
rect 12170 8542 12180 8598
rect 10244 8474 12180 8542
rect 10244 8418 10254 8474
rect 10310 8418 10378 8474
rect 10434 8418 10502 8474
rect 10558 8418 10626 8474
rect 10682 8418 10750 8474
rect 10806 8418 10874 8474
rect 10930 8418 10998 8474
rect 11054 8418 11122 8474
rect 11178 8418 11246 8474
rect 11302 8418 11370 8474
rect 11426 8418 11494 8474
rect 11550 8418 11618 8474
rect 11674 8418 11742 8474
rect 11798 8418 11866 8474
rect 11922 8418 11990 8474
rect 12046 8418 12114 8474
rect 12170 8418 12180 8474
rect 10244 8350 12180 8418
rect 10244 8294 10254 8350
rect 10310 8294 10378 8350
rect 10434 8294 10502 8350
rect 10558 8294 10626 8350
rect 10682 8294 10750 8350
rect 10806 8294 10874 8350
rect 10930 8294 10998 8350
rect 11054 8294 11122 8350
rect 11178 8294 11246 8350
rect 11302 8294 11370 8350
rect 11426 8294 11494 8350
rect 11550 8294 11618 8350
rect 11674 8294 11742 8350
rect 11798 8294 11866 8350
rect 11922 8294 11990 8350
rect 12046 8294 12114 8350
rect 12170 8294 12180 8350
rect 10244 8226 12180 8294
rect 10244 8170 10254 8226
rect 10310 8170 10378 8226
rect 10434 8170 10502 8226
rect 10558 8170 10626 8226
rect 10682 8170 10750 8226
rect 10806 8170 10874 8226
rect 10930 8170 10998 8226
rect 11054 8170 11122 8226
rect 11178 8170 11246 8226
rect 11302 8170 11370 8226
rect 11426 8170 11494 8226
rect 11550 8170 11618 8226
rect 11674 8170 11742 8226
rect 11798 8170 11866 8226
rect 11922 8170 11990 8226
rect 12046 8170 12114 8226
rect 12170 8170 12180 8226
rect 10244 8102 12180 8170
rect 10244 8046 10254 8102
rect 10310 8046 10378 8102
rect 10434 8046 10502 8102
rect 10558 8046 10626 8102
rect 10682 8046 10750 8102
rect 10806 8046 10874 8102
rect 10930 8046 10998 8102
rect 11054 8046 11122 8102
rect 11178 8046 11246 8102
rect 11302 8046 11370 8102
rect 11426 8046 11494 8102
rect 11550 8046 11618 8102
rect 11674 8046 11742 8102
rect 11798 8046 11866 8102
rect 11922 8046 11990 8102
rect 12046 8046 12114 8102
rect 12170 8046 12180 8102
rect 10244 8036 12180 8046
rect 12861 10954 14673 10964
rect 12861 10898 12871 10954
rect 12927 10898 12995 10954
rect 13051 10898 13119 10954
rect 13175 10898 13243 10954
rect 13299 10898 13367 10954
rect 13423 10898 13491 10954
rect 13547 10898 13615 10954
rect 13671 10898 13739 10954
rect 13795 10898 13863 10954
rect 13919 10898 13987 10954
rect 14043 10898 14111 10954
rect 14167 10898 14235 10954
rect 14291 10898 14359 10954
rect 14415 10898 14483 10954
rect 14539 10898 14607 10954
rect 14663 10898 14673 10954
rect 12861 10830 14673 10898
rect 12861 10774 12871 10830
rect 12927 10774 12995 10830
rect 13051 10774 13119 10830
rect 13175 10774 13243 10830
rect 13299 10774 13367 10830
rect 13423 10774 13491 10830
rect 13547 10774 13615 10830
rect 13671 10774 13739 10830
rect 13795 10774 13863 10830
rect 13919 10774 13987 10830
rect 14043 10774 14111 10830
rect 14167 10774 14235 10830
rect 14291 10774 14359 10830
rect 14415 10774 14483 10830
rect 14539 10774 14607 10830
rect 14663 10774 14673 10830
rect 12861 10706 14673 10774
rect 12861 10650 12871 10706
rect 12927 10650 12995 10706
rect 13051 10650 13119 10706
rect 13175 10650 13243 10706
rect 13299 10650 13367 10706
rect 13423 10650 13491 10706
rect 13547 10650 13615 10706
rect 13671 10650 13739 10706
rect 13795 10650 13863 10706
rect 13919 10650 13987 10706
rect 14043 10650 14111 10706
rect 14167 10650 14235 10706
rect 14291 10650 14359 10706
rect 14415 10650 14483 10706
rect 14539 10650 14607 10706
rect 14663 10650 14673 10706
rect 12861 10582 14673 10650
rect 12861 10526 12871 10582
rect 12927 10526 12995 10582
rect 13051 10526 13119 10582
rect 13175 10526 13243 10582
rect 13299 10526 13367 10582
rect 13423 10526 13491 10582
rect 13547 10526 13615 10582
rect 13671 10526 13739 10582
rect 13795 10526 13863 10582
rect 13919 10526 13987 10582
rect 14043 10526 14111 10582
rect 14167 10526 14235 10582
rect 14291 10526 14359 10582
rect 14415 10526 14483 10582
rect 14539 10526 14607 10582
rect 14663 10526 14673 10582
rect 12861 10458 14673 10526
rect 12861 10402 12871 10458
rect 12927 10402 12995 10458
rect 13051 10402 13119 10458
rect 13175 10402 13243 10458
rect 13299 10402 13367 10458
rect 13423 10402 13491 10458
rect 13547 10402 13615 10458
rect 13671 10402 13739 10458
rect 13795 10402 13863 10458
rect 13919 10402 13987 10458
rect 14043 10402 14111 10458
rect 14167 10402 14235 10458
rect 14291 10402 14359 10458
rect 14415 10402 14483 10458
rect 14539 10402 14607 10458
rect 14663 10402 14673 10458
rect 12861 10334 14673 10402
rect 12861 10278 12871 10334
rect 12927 10278 12995 10334
rect 13051 10278 13119 10334
rect 13175 10278 13243 10334
rect 13299 10278 13367 10334
rect 13423 10278 13491 10334
rect 13547 10278 13615 10334
rect 13671 10278 13739 10334
rect 13795 10278 13863 10334
rect 13919 10278 13987 10334
rect 14043 10278 14111 10334
rect 14167 10278 14235 10334
rect 14291 10278 14359 10334
rect 14415 10278 14483 10334
rect 14539 10278 14607 10334
rect 14663 10278 14673 10334
rect 12861 10210 14673 10278
rect 12861 10154 12871 10210
rect 12927 10154 12995 10210
rect 13051 10154 13119 10210
rect 13175 10154 13243 10210
rect 13299 10154 13367 10210
rect 13423 10154 13491 10210
rect 13547 10154 13615 10210
rect 13671 10154 13739 10210
rect 13795 10154 13863 10210
rect 13919 10154 13987 10210
rect 14043 10154 14111 10210
rect 14167 10154 14235 10210
rect 14291 10154 14359 10210
rect 14415 10154 14483 10210
rect 14539 10154 14607 10210
rect 14663 10154 14673 10210
rect 12861 10086 14673 10154
rect 12861 10030 12871 10086
rect 12927 10030 12995 10086
rect 13051 10030 13119 10086
rect 13175 10030 13243 10086
rect 13299 10030 13367 10086
rect 13423 10030 13491 10086
rect 13547 10030 13615 10086
rect 13671 10030 13739 10086
rect 13795 10030 13863 10086
rect 13919 10030 13987 10086
rect 14043 10030 14111 10086
rect 14167 10030 14235 10086
rect 14291 10030 14359 10086
rect 14415 10030 14483 10086
rect 14539 10030 14607 10086
rect 14663 10030 14673 10086
rect 12861 9962 14673 10030
rect 12861 9906 12871 9962
rect 12927 9906 12995 9962
rect 13051 9906 13119 9962
rect 13175 9906 13243 9962
rect 13299 9906 13367 9962
rect 13423 9906 13491 9962
rect 13547 9906 13615 9962
rect 13671 9906 13739 9962
rect 13795 9906 13863 9962
rect 13919 9906 13987 9962
rect 14043 9906 14111 9962
rect 14167 9906 14235 9962
rect 14291 9906 14359 9962
rect 14415 9906 14483 9962
rect 14539 9906 14607 9962
rect 14663 9906 14673 9962
rect 12861 9838 14673 9906
rect 12861 9782 12871 9838
rect 12927 9782 12995 9838
rect 13051 9782 13119 9838
rect 13175 9782 13243 9838
rect 13299 9782 13367 9838
rect 13423 9782 13491 9838
rect 13547 9782 13615 9838
rect 13671 9782 13739 9838
rect 13795 9782 13863 9838
rect 13919 9782 13987 9838
rect 14043 9782 14111 9838
rect 14167 9782 14235 9838
rect 14291 9782 14359 9838
rect 14415 9782 14483 9838
rect 14539 9782 14607 9838
rect 14663 9782 14673 9838
rect 12861 9714 14673 9782
rect 12861 9658 12871 9714
rect 12927 9658 12995 9714
rect 13051 9658 13119 9714
rect 13175 9658 13243 9714
rect 13299 9658 13367 9714
rect 13423 9658 13491 9714
rect 13547 9658 13615 9714
rect 13671 9658 13739 9714
rect 13795 9658 13863 9714
rect 13919 9658 13987 9714
rect 14043 9658 14111 9714
rect 14167 9658 14235 9714
rect 14291 9658 14359 9714
rect 14415 9658 14483 9714
rect 14539 9658 14607 9714
rect 14663 9658 14673 9714
rect 12861 9590 14673 9658
rect 12861 9534 12871 9590
rect 12927 9534 12995 9590
rect 13051 9534 13119 9590
rect 13175 9534 13243 9590
rect 13299 9534 13367 9590
rect 13423 9534 13491 9590
rect 13547 9534 13615 9590
rect 13671 9534 13739 9590
rect 13795 9534 13863 9590
rect 13919 9534 13987 9590
rect 14043 9534 14111 9590
rect 14167 9534 14235 9590
rect 14291 9534 14359 9590
rect 14415 9534 14483 9590
rect 14539 9534 14607 9590
rect 14663 9534 14673 9590
rect 12861 9466 14673 9534
rect 12861 9410 12871 9466
rect 12927 9410 12995 9466
rect 13051 9410 13119 9466
rect 13175 9410 13243 9466
rect 13299 9410 13367 9466
rect 13423 9410 13491 9466
rect 13547 9410 13615 9466
rect 13671 9410 13739 9466
rect 13795 9410 13863 9466
rect 13919 9410 13987 9466
rect 14043 9410 14111 9466
rect 14167 9410 14235 9466
rect 14291 9410 14359 9466
rect 14415 9410 14483 9466
rect 14539 9410 14607 9466
rect 14663 9410 14673 9466
rect 12861 9342 14673 9410
rect 12861 9286 12871 9342
rect 12927 9286 12995 9342
rect 13051 9286 13119 9342
rect 13175 9286 13243 9342
rect 13299 9286 13367 9342
rect 13423 9286 13491 9342
rect 13547 9286 13615 9342
rect 13671 9286 13739 9342
rect 13795 9286 13863 9342
rect 13919 9286 13987 9342
rect 14043 9286 14111 9342
rect 14167 9286 14235 9342
rect 14291 9286 14359 9342
rect 14415 9286 14483 9342
rect 14539 9286 14607 9342
rect 14663 9286 14673 9342
rect 12861 9218 14673 9286
rect 12861 9162 12871 9218
rect 12927 9162 12995 9218
rect 13051 9162 13119 9218
rect 13175 9162 13243 9218
rect 13299 9162 13367 9218
rect 13423 9162 13491 9218
rect 13547 9162 13615 9218
rect 13671 9162 13739 9218
rect 13795 9162 13863 9218
rect 13919 9162 13987 9218
rect 14043 9162 14111 9218
rect 14167 9162 14235 9218
rect 14291 9162 14359 9218
rect 14415 9162 14483 9218
rect 14539 9162 14607 9218
rect 14663 9162 14673 9218
rect 12861 9094 14673 9162
rect 12861 9038 12871 9094
rect 12927 9038 12995 9094
rect 13051 9038 13119 9094
rect 13175 9038 13243 9094
rect 13299 9038 13367 9094
rect 13423 9038 13491 9094
rect 13547 9038 13615 9094
rect 13671 9038 13739 9094
rect 13795 9038 13863 9094
rect 13919 9038 13987 9094
rect 14043 9038 14111 9094
rect 14167 9038 14235 9094
rect 14291 9038 14359 9094
rect 14415 9038 14483 9094
rect 14539 9038 14607 9094
rect 14663 9038 14673 9094
rect 12861 8970 14673 9038
rect 12861 8914 12871 8970
rect 12927 8914 12995 8970
rect 13051 8914 13119 8970
rect 13175 8914 13243 8970
rect 13299 8914 13367 8970
rect 13423 8914 13491 8970
rect 13547 8914 13615 8970
rect 13671 8914 13739 8970
rect 13795 8914 13863 8970
rect 13919 8914 13987 8970
rect 14043 8914 14111 8970
rect 14167 8914 14235 8970
rect 14291 8914 14359 8970
rect 14415 8914 14483 8970
rect 14539 8914 14607 8970
rect 14663 8914 14673 8970
rect 12861 8846 14673 8914
rect 12861 8790 12871 8846
rect 12927 8790 12995 8846
rect 13051 8790 13119 8846
rect 13175 8790 13243 8846
rect 13299 8790 13367 8846
rect 13423 8790 13491 8846
rect 13547 8790 13615 8846
rect 13671 8790 13739 8846
rect 13795 8790 13863 8846
rect 13919 8790 13987 8846
rect 14043 8790 14111 8846
rect 14167 8790 14235 8846
rect 14291 8790 14359 8846
rect 14415 8790 14483 8846
rect 14539 8790 14607 8846
rect 14663 8790 14673 8846
rect 12861 8722 14673 8790
rect 12861 8666 12871 8722
rect 12927 8666 12995 8722
rect 13051 8666 13119 8722
rect 13175 8666 13243 8722
rect 13299 8666 13367 8722
rect 13423 8666 13491 8722
rect 13547 8666 13615 8722
rect 13671 8666 13739 8722
rect 13795 8666 13863 8722
rect 13919 8666 13987 8722
rect 14043 8666 14111 8722
rect 14167 8666 14235 8722
rect 14291 8666 14359 8722
rect 14415 8666 14483 8722
rect 14539 8666 14607 8722
rect 14663 8666 14673 8722
rect 12861 8598 14673 8666
rect 12861 8542 12871 8598
rect 12927 8542 12995 8598
rect 13051 8542 13119 8598
rect 13175 8542 13243 8598
rect 13299 8542 13367 8598
rect 13423 8542 13491 8598
rect 13547 8542 13615 8598
rect 13671 8542 13739 8598
rect 13795 8542 13863 8598
rect 13919 8542 13987 8598
rect 14043 8542 14111 8598
rect 14167 8542 14235 8598
rect 14291 8542 14359 8598
rect 14415 8542 14483 8598
rect 14539 8542 14607 8598
rect 14663 8542 14673 8598
rect 12861 8474 14673 8542
rect 12861 8418 12871 8474
rect 12927 8418 12995 8474
rect 13051 8418 13119 8474
rect 13175 8418 13243 8474
rect 13299 8418 13367 8474
rect 13423 8418 13491 8474
rect 13547 8418 13615 8474
rect 13671 8418 13739 8474
rect 13795 8418 13863 8474
rect 13919 8418 13987 8474
rect 14043 8418 14111 8474
rect 14167 8418 14235 8474
rect 14291 8418 14359 8474
rect 14415 8418 14483 8474
rect 14539 8418 14607 8474
rect 14663 8418 14673 8474
rect 12861 8350 14673 8418
rect 12861 8294 12871 8350
rect 12927 8294 12995 8350
rect 13051 8294 13119 8350
rect 13175 8294 13243 8350
rect 13299 8294 13367 8350
rect 13423 8294 13491 8350
rect 13547 8294 13615 8350
rect 13671 8294 13739 8350
rect 13795 8294 13863 8350
rect 13919 8294 13987 8350
rect 14043 8294 14111 8350
rect 14167 8294 14235 8350
rect 14291 8294 14359 8350
rect 14415 8294 14483 8350
rect 14539 8294 14607 8350
rect 14663 8294 14673 8350
rect 12861 8226 14673 8294
rect 12861 8170 12871 8226
rect 12927 8170 12995 8226
rect 13051 8170 13119 8226
rect 13175 8170 13243 8226
rect 13299 8170 13367 8226
rect 13423 8170 13491 8226
rect 13547 8170 13615 8226
rect 13671 8170 13739 8226
rect 13795 8170 13863 8226
rect 13919 8170 13987 8226
rect 14043 8170 14111 8226
rect 14167 8170 14235 8226
rect 14291 8170 14359 8226
rect 14415 8170 14483 8226
rect 14539 8170 14607 8226
rect 14663 8170 14673 8226
rect 12861 8102 14673 8170
rect 12861 8046 12871 8102
rect 12927 8046 12995 8102
rect 13051 8046 13119 8102
rect 13175 8046 13243 8102
rect 13299 8046 13367 8102
rect 13423 8046 13491 8102
rect 13547 8046 13615 8102
rect 13671 8046 13739 8102
rect 13795 8046 13863 8102
rect 13919 8046 13987 8102
rect 14043 8046 14111 8102
rect 14167 8046 14235 8102
rect 14291 8046 14359 8102
rect 14415 8046 14483 8102
rect 14539 8046 14607 8102
rect 14663 8046 14673 8102
rect 12861 8036 14673 8046
rect -11 8004 86 8014
rect 14892 8014 14902 10986
rect 14958 8014 14989 10986
rect 14892 8004 14989 8014
rect -11 7786 86 7796
rect -11 4814 20 7786
rect 76 4814 86 7786
rect 14892 7786 14989 7796
rect 305 7754 2117 7764
rect 305 7698 315 7754
rect 371 7698 439 7754
rect 495 7698 563 7754
rect 619 7698 687 7754
rect 743 7698 811 7754
rect 867 7698 935 7754
rect 991 7698 1059 7754
rect 1115 7698 1183 7754
rect 1239 7698 1307 7754
rect 1363 7698 1431 7754
rect 1487 7698 1555 7754
rect 1611 7698 1679 7754
rect 1735 7698 1803 7754
rect 1859 7698 1927 7754
rect 1983 7698 2051 7754
rect 2107 7698 2117 7754
rect 305 7630 2117 7698
rect 305 7574 315 7630
rect 371 7574 439 7630
rect 495 7574 563 7630
rect 619 7574 687 7630
rect 743 7574 811 7630
rect 867 7574 935 7630
rect 991 7574 1059 7630
rect 1115 7574 1183 7630
rect 1239 7574 1307 7630
rect 1363 7574 1431 7630
rect 1487 7574 1555 7630
rect 1611 7574 1679 7630
rect 1735 7574 1803 7630
rect 1859 7574 1927 7630
rect 1983 7574 2051 7630
rect 2107 7574 2117 7630
rect 305 7506 2117 7574
rect 305 7450 315 7506
rect 371 7450 439 7506
rect 495 7450 563 7506
rect 619 7450 687 7506
rect 743 7450 811 7506
rect 867 7450 935 7506
rect 991 7450 1059 7506
rect 1115 7450 1183 7506
rect 1239 7450 1307 7506
rect 1363 7450 1431 7506
rect 1487 7450 1555 7506
rect 1611 7450 1679 7506
rect 1735 7450 1803 7506
rect 1859 7450 1927 7506
rect 1983 7450 2051 7506
rect 2107 7450 2117 7506
rect 305 7382 2117 7450
rect 305 7326 315 7382
rect 371 7326 439 7382
rect 495 7326 563 7382
rect 619 7326 687 7382
rect 743 7326 811 7382
rect 867 7326 935 7382
rect 991 7326 1059 7382
rect 1115 7326 1183 7382
rect 1239 7326 1307 7382
rect 1363 7326 1431 7382
rect 1487 7326 1555 7382
rect 1611 7326 1679 7382
rect 1735 7326 1803 7382
rect 1859 7326 1927 7382
rect 1983 7326 2051 7382
rect 2107 7326 2117 7382
rect 305 7258 2117 7326
rect 305 7202 315 7258
rect 371 7202 439 7258
rect 495 7202 563 7258
rect 619 7202 687 7258
rect 743 7202 811 7258
rect 867 7202 935 7258
rect 991 7202 1059 7258
rect 1115 7202 1183 7258
rect 1239 7202 1307 7258
rect 1363 7202 1431 7258
rect 1487 7202 1555 7258
rect 1611 7202 1679 7258
rect 1735 7202 1803 7258
rect 1859 7202 1927 7258
rect 1983 7202 2051 7258
rect 2107 7202 2117 7258
rect 305 7134 2117 7202
rect 305 7078 315 7134
rect 371 7078 439 7134
rect 495 7078 563 7134
rect 619 7078 687 7134
rect 743 7078 811 7134
rect 867 7078 935 7134
rect 991 7078 1059 7134
rect 1115 7078 1183 7134
rect 1239 7078 1307 7134
rect 1363 7078 1431 7134
rect 1487 7078 1555 7134
rect 1611 7078 1679 7134
rect 1735 7078 1803 7134
rect 1859 7078 1927 7134
rect 1983 7078 2051 7134
rect 2107 7078 2117 7134
rect 305 7010 2117 7078
rect 305 6954 315 7010
rect 371 6954 439 7010
rect 495 6954 563 7010
rect 619 6954 687 7010
rect 743 6954 811 7010
rect 867 6954 935 7010
rect 991 6954 1059 7010
rect 1115 6954 1183 7010
rect 1239 6954 1307 7010
rect 1363 6954 1431 7010
rect 1487 6954 1555 7010
rect 1611 6954 1679 7010
rect 1735 6954 1803 7010
rect 1859 6954 1927 7010
rect 1983 6954 2051 7010
rect 2107 6954 2117 7010
rect 305 6886 2117 6954
rect 305 6830 315 6886
rect 371 6830 439 6886
rect 495 6830 563 6886
rect 619 6830 687 6886
rect 743 6830 811 6886
rect 867 6830 935 6886
rect 991 6830 1059 6886
rect 1115 6830 1183 6886
rect 1239 6830 1307 6886
rect 1363 6830 1431 6886
rect 1487 6830 1555 6886
rect 1611 6830 1679 6886
rect 1735 6830 1803 6886
rect 1859 6830 1927 6886
rect 1983 6830 2051 6886
rect 2107 6830 2117 6886
rect 305 6762 2117 6830
rect 305 6706 315 6762
rect 371 6706 439 6762
rect 495 6706 563 6762
rect 619 6706 687 6762
rect 743 6706 811 6762
rect 867 6706 935 6762
rect 991 6706 1059 6762
rect 1115 6706 1183 6762
rect 1239 6706 1307 6762
rect 1363 6706 1431 6762
rect 1487 6706 1555 6762
rect 1611 6706 1679 6762
rect 1735 6706 1803 6762
rect 1859 6706 1927 6762
rect 1983 6706 2051 6762
rect 2107 6706 2117 6762
rect 305 6638 2117 6706
rect 305 6582 315 6638
rect 371 6582 439 6638
rect 495 6582 563 6638
rect 619 6582 687 6638
rect 743 6582 811 6638
rect 867 6582 935 6638
rect 991 6582 1059 6638
rect 1115 6582 1183 6638
rect 1239 6582 1307 6638
rect 1363 6582 1431 6638
rect 1487 6582 1555 6638
rect 1611 6582 1679 6638
rect 1735 6582 1803 6638
rect 1859 6582 1927 6638
rect 1983 6582 2051 6638
rect 2107 6582 2117 6638
rect 305 6514 2117 6582
rect 305 6458 315 6514
rect 371 6458 439 6514
rect 495 6458 563 6514
rect 619 6458 687 6514
rect 743 6458 811 6514
rect 867 6458 935 6514
rect 991 6458 1059 6514
rect 1115 6458 1183 6514
rect 1239 6458 1307 6514
rect 1363 6458 1431 6514
rect 1487 6458 1555 6514
rect 1611 6458 1679 6514
rect 1735 6458 1803 6514
rect 1859 6458 1927 6514
rect 1983 6458 2051 6514
rect 2107 6458 2117 6514
rect 305 6390 2117 6458
rect 305 6334 315 6390
rect 371 6334 439 6390
rect 495 6334 563 6390
rect 619 6334 687 6390
rect 743 6334 811 6390
rect 867 6334 935 6390
rect 991 6334 1059 6390
rect 1115 6334 1183 6390
rect 1239 6334 1307 6390
rect 1363 6334 1431 6390
rect 1487 6334 1555 6390
rect 1611 6334 1679 6390
rect 1735 6334 1803 6390
rect 1859 6334 1927 6390
rect 1983 6334 2051 6390
rect 2107 6334 2117 6390
rect 305 6266 2117 6334
rect 305 6210 315 6266
rect 371 6210 439 6266
rect 495 6210 563 6266
rect 619 6210 687 6266
rect 743 6210 811 6266
rect 867 6210 935 6266
rect 991 6210 1059 6266
rect 1115 6210 1183 6266
rect 1239 6210 1307 6266
rect 1363 6210 1431 6266
rect 1487 6210 1555 6266
rect 1611 6210 1679 6266
rect 1735 6210 1803 6266
rect 1859 6210 1927 6266
rect 1983 6210 2051 6266
rect 2107 6210 2117 6266
rect 305 6142 2117 6210
rect 305 6086 315 6142
rect 371 6086 439 6142
rect 495 6086 563 6142
rect 619 6086 687 6142
rect 743 6086 811 6142
rect 867 6086 935 6142
rect 991 6086 1059 6142
rect 1115 6086 1183 6142
rect 1239 6086 1307 6142
rect 1363 6086 1431 6142
rect 1487 6086 1555 6142
rect 1611 6086 1679 6142
rect 1735 6086 1803 6142
rect 1859 6086 1927 6142
rect 1983 6086 2051 6142
rect 2107 6086 2117 6142
rect 305 6018 2117 6086
rect 305 5962 315 6018
rect 371 5962 439 6018
rect 495 5962 563 6018
rect 619 5962 687 6018
rect 743 5962 811 6018
rect 867 5962 935 6018
rect 991 5962 1059 6018
rect 1115 5962 1183 6018
rect 1239 5962 1307 6018
rect 1363 5962 1431 6018
rect 1487 5962 1555 6018
rect 1611 5962 1679 6018
rect 1735 5962 1803 6018
rect 1859 5962 1927 6018
rect 1983 5962 2051 6018
rect 2107 5962 2117 6018
rect 305 5894 2117 5962
rect 305 5838 315 5894
rect 371 5838 439 5894
rect 495 5838 563 5894
rect 619 5838 687 5894
rect 743 5838 811 5894
rect 867 5838 935 5894
rect 991 5838 1059 5894
rect 1115 5838 1183 5894
rect 1239 5838 1307 5894
rect 1363 5838 1431 5894
rect 1487 5838 1555 5894
rect 1611 5838 1679 5894
rect 1735 5838 1803 5894
rect 1859 5838 1927 5894
rect 1983 5838 2051 5894
rect 2107 5838 2117 5894
rect 305 5770 2117 5838
rect 305 5714 315 5770
rect 371 5714 439 5770
rect 495 5714 563 5770
rect 619 5714 687 5770
rect 743 5714 811 5770
rect 867 5714 935 5770
rect 991 5714 1059 5770
rect 1115 5714 1183 5770
rect 1239 5714 1307 5770
rect 1363 5714 1431 5770
rect 1487 5714 1555 5770
rect 1611 5714 1679 5770
rect 1735 5714 1803 5770
rect 1859 5714 1927 5770
rect 1983 5714 2051 5770
rect 2107 5714 2117 5770
rect 305 5646 2117 5714
rect 305 5590 315 5646
rect 371 5590 439 5646
rect 495 5590 563 5646
rect 619 5590 687 5646
rect 743 5590 811 5646
rect 867 5590 935 5646
rect 991 5590 1059 5646
rect 1115 5590 1183 5646
rect 1239 5590 1307 5646
rect 1363 5590 1431 5646
rect 1487 5590 1555 5646
rect 1611 5590 1679 5646
rect 1735 5590 1803 5646
rect 1859 5590 1927 5646
rect 1983 5590 2051 5646
rect 2107 5590 2117 5646
rect 305 5522 2117 5590
rect 305 5466 315 5522
rect 371 5466 439 5522
rect 495 5466 563 5522
rect 619 5466 687 5522
rect 743 5466 811 5522
rect 867 5466 935 5522
rect 991 5466 1059 5522
rect 1115 5466 1183 5522
rect 1239 5466 1307 5522
rect 1363 5466 1431 5522
rect 1487 5466 1555 5522
rect 1611 5466 1679 5522
rect 1735 5466 1803 5522
rect 1859 5466 1927 5522
rect 1983 5466 2051 5522
rect 2107 5466 2117 5522
rect 305 5398 2117 5466
rect 305 5342 315 5398
rect 371 5342 439 5398
rect 495 5342 563 5398
rect 619 5342 687 5398
rect 743 5342 811 5398
rect 867 5342 935 5398
rect 991 5342 1059 5398
rect 1115 5342 1183 5398
rect 1239 5342 1307 5398
rect 1363 5342 1431 5398
rect 1487 5342 1555 5398
rect 1611 5342 1679 5398
rect 1735 5342 1803 5398
rect 1859 5342 1927 5398
rect 1983 5342 2051 5398
rect 2107 5342 2117 5398
rect 305 5274 2117 5342
rect 305 5218 315 5274
rect 371 5218 439 5274
rect 495 5218 563 5274
rect 619 5218 687 5274
rect 743 5218 811 5274
rect 867 5218 935 5274
rect 991 5218 1059 5274
rect 1115 5218 1183 5274
rect 1239 5218 1307 5274
rect 1363 5218 1431 5274
rect 1487 5218 1555 5274
rect 1611 5218 1679 5274
rect 1735 5218 1803 5274
rect 1859 5218 1927 5274
rect 1983 5218 2051 5274
rect 2107 5218 2117 5274
rect 305 5150 2117 5218
rect 305 5094 315 5150
rect 371 5094 439 5150
rect 495 5094 563 5150
rect 619 5094 687 5150
rect 743 5094 811 5150
rect 867 5094 935 5150
rect 991 5094 1059 5150
rect 1115 5094 1183 5150
rect 1239 5094 1307 5150
rect 1363 5094 1431 5150
rect 1487 5094 1555 5150
rect 1611 5094 1679 5150
rect 1735 5094 1803 5150
rect 1859 5094 1927 5150
rect 1983 5094 2051 5150
rect 2107 5094 2117 5150
rect 305 5026 2117 5094
rect 305 4970 315 5026
rect 371 4970 439 5026
rect 495 4970 563 5026
rect 619 4970 687 5026
rect 743 4970 811 5026
rect 867 4970 935 5026
rect 991 4970 1059 5026
rect 1115 4970 1183 5026
rect 1239 4970 1307 5026
rect 1363 4970 1431 5026
rect 1487 4970 1555 5026
rect 1611 4970 1679 5026
rect 1735 4970 1803 5026
rect 1859 4970 1927 5026
rect 1983 4970 2051 5026
rect 2107 4970 2117 5026
rect 305 4902 2117 4970
rect 305 4846 315 4902
rect 371 4846 439 4902
rect 495 4846 563 4902
rect 619 4846 687 4902
rect 743 4846 811 4902
rect 867 4846 935 4902
rect 991 4846 1059 4902
rect 1115 4846 1183 4902
rect 1239 4846 1307 4902
rect 1363 4846 1431 4902
rect 1487 4846 1555 4902
rect 1611 4846 1679 4902
rect 1735 4846 1803 4902
rect 1859 4846 1927 4902
rect 1983 4846 2051 4902
rect 2107 4846 2117 4902
rect 305 4836 2117 4846
rect 2798 7754 4734 7764
rect 2798 7698 2808 7754
rect 2864 7698 2932 7754
rect 2988 7698 3056 7754
rect 3112 7698 3180 7754
rect 3236 7698 3304 7754
rect 3360 7698 3428 7754
rect 3484 7698 3552 7754
rect 3608 7698 3676 7754
rect 3732 7698 3800 7754
rect 3856 7698 3924 7754
rect 3980 7698 4048 7754
rect 4104 7698 4172 7754
rect 4228 7698 4296 7754
rect 4352 7698 4420 7754
rect 4476 7698 4544 7754
rect 4600 7698 4668 7754
rect 4724 7698 4734 7754
rect 2798 7630 4734 7698
rect 2798 7574 2808 7630
rect 2864 7574 2932 7630
rect 2988 7574 3056 7630
rect 3112 7574 3180 7630
rect 3236 7574 3304 7630
rect 3360 7574 3428 7630
rect 3484 7574 3552 7630
rect 3608 7574 3676 7630
rect 3732 7574 3800 7630
rect 3856 7574 3924 7630
rect 3980 7574 4048 7630
rect 4104 7574 4172 7630
rect 4228 7574 4296 7630
rect 4352 7574 4420 7630
rect 4476 7574 4544 7630
rect 4600 7574 4668 7630
rect 4724 7574 4734 7630
rect 2798 7506 4734 7574
rect 2798 7450 2808 7506
rect 2864 7450 2932 7506
rect 2988 7450 3056 7506
rect 3112 7450 3180 7506
rect 3236 7450 3304 7506
rect 3360 7450 3428 7506
rect 3484 7450 3552 7506
rect 3608 7450 3676 7506
rect 3732 7450 3800 7506
rect 3856 7450 3924 7506
rect 3980 7450 4048 7506
rect 4104 7450 4172 7506
rect 4228 7450 4296 7506
rect 4352 7450 4420 7506
rect 4476 7450 4544 7506
rect 4600 7450 4668 7506
rect 4724 7450 4734 7506
rect 2798 7382 4734 7450
rect 2798 7326 2808 7382
rect 2864 7326 2932 7382
rect 2988 7326 3056 7382
rect 3112 7326 3180 7382
rect 3236 7326 3304 7382
rect 3360 7326 3428 7382
rect 3484 7326 3552 7382
rect 3608 7326 3676 7382
rect 3732 7326 3800 7382
rect 3856 7326 3924 7382
rect 3980 7326 4048 7382
rect 4104 7326 4172 7382
rect 4228 7326 4296 7382
rect 4352 7326 4420 7382
rect 4476 7326 4544 7382
rect 4600 7326 4668 7382
rect 4724 7326 4734 7382
rect 2798 7258 4734 7326
rect 2798 7202 2808 7258
rect 2864 7202 2932 7258
rect 2988 7202 3056 7258
rect 3112 7202 3180 7258
rect 3236 7202 3304 7258
rect 3360 7202 3428 7258
rect 3484 7202 3552 7258
rect 3608 7202 3676 7258
rect 3732 7202 3800 7258
rect 3856 7202 3924 7258
rect 3980 7202 4048 7258
rect 4104 7202 4172 7258
rect 4228 7202 4296 7258
rect 4352 7202 4420 7258
rect 4476 7202 4544 7258
rect 4600 7202 4668 7258
rect 4724 7202 4734 7258
rect 2798 7134 4734 7202
rect 2798 7078 2808 7134
rect 2864 7078 2932 7134
rect 2988 7078 3056 7134
rect 3112 7078 3180 7134
rect 3236 7078 3304 7134
rect 3360 7078 3428 7134
rect 3484 7078 3552 7134
rect 3608 7078 3676 7134
rect 3732 7078 3800 7134
rect 3856 7078 3924 7134
rect 3980 7078 4048 7134
rect 4104 7078 4172 7134
rect 4228 7078 4296 7134
rect 4352 7078 4420 7134
rect 4476 7078 4544 7134
rect 4600 7078 4668 7134
rect 4724 7078 4734 7134
rect 2798 7010 4734 7078
rect 2798 6954 2808 7010
rect 2864 6954 2932 7010
rect 2988 6954 3056 7010
rect 3112 6954 3180 7010
rect 3236 6954 3304 7010
rect 3360 6954 3428 7010
rect 3484 6954 3552 7010
rect 3608 6954 3676 7010
rect 3732 6954 3800 7010
rect 3856 6954 3924 7010
rect 3980 6954 4048 7010
rect 4104 6954 4172 7010
rect 4228 6954 4296 7010
rect 4352 6954 4420 7010
rect 4476 6954 4544 7010
rect 4600 6954 4668 7010
rect 4724 6954 4734 7010
rect 2798 6886 4734 6954
rect 2798 6830 2808 6886
rect 2864 6830 2932 6886
rect 2988 6830 3056 6886
rect 3112 6830 3180 6886
rect 3236 6830 3304 6886
rect 3360 6830 3428 6886
rect 3484 6830 3552 6886
rect 3608 6830 3676 6886
rect 3732 6830 3800 6886
rect 3856 6830 3924 6886
rect 3980 6830 4048 6886
rect 4104 6830 4172 6886
rect 4228 6830 4296 6886
rect 4352 6830 4420 6886
rect 4476 6830 4544 6886
rect 4600 6830 4668 6886
rect 4724 6830 4734 6886
rect 2798 6762 4734 6830
rect 2798 6706 2808 6762
rect 2864 6706 2932 6762
rect 2988 6706 3056 6762
rect 3112 6706 3180 6762
rect 3236 6706 3304 6762
rect 3360 6706 3428 6762
rect 3484 6706 3552 6762
rect 3608 6706 3676 6762
rect 3732 6706 3800 6762
rect 3856 6706 3924 6762
rect 3980 6706 4048 6762
rect 4104 6706 4172 6762
rect 4228 6706 4296 6762
rect 4352 6706 4420 6762
rect 4476 6706 4544 6762
rect 4600 6706 4668 6762
rect 4724 6706 4734 6762
rect 2798 6638 4734 6706
rect 2798 6582 2808 6638
rect 2864 6582 2932 6638
rect 2988 6582 3056 6638
rect 3112 6582 3180 6638
rect 3236 6582 3304 6638
rect 3360 6582 3428 6638
rect 3484 6582 3552 6638
rect 3608 6582 3676 6638
rect 3732 6582 3800 6638
rect 3856 6582 3924 6638
rect 3980 6582 4048 6638
rect 4104 6582 4172 6638
rect 4228 6582 4296 6638
rect 4352 6582 4420 6638
rect 4476 6582 4544 6638
rect 4600 6582 4668 6638
rect 4724 6582 4734 6638
rect 2798 6514 4734 6582
rect 2798 6458 2808 6514
rect 2864 6458 2932 6514
rect 2988 6458 3056 6514
rect 3112 6458 3180 6514
rect 3236 6458 3304 6514
rect 3360 6458 3428 6514
rect 3484 6458 3552 6514
rect 3608 6458 3676 6514
rect 3732 6458 3800 6514
rect 3856 6458 3924 6514
rect 3980 6458 4048 6514
rect 4104 6458 4172 6514
rect 4228 6458 4296 6514
rect 4352 6458 4420 6514
rect 4476 6458 4544 6514
rect 4600 6458 4668 6514
rect 4724 6458 4734 6514
rect 2798 6390 4734 6458
rect 2798 6334 2808 6390
rect 2864 6334 2932 6390
rect 2988 6334 3056 6390
rect 3112 6334 3180 6390
rect 3236 6334 3304 6390
rect 3360 6334 3428 6390
rect 3484 6334 3552 6390
rect 3608 6334 3676 6390
rect 3732 6334 3800 6390
rect 3856 6334 3924 6390
rect 3980 6334 4048 6390
rect 4104 6334 4172 6390
rect 4228 6334 4296 6390
rect 4352 6334 4420 6390
rect 4476 6334 4544 6390
rect 4600 6334 4668 6390
rect 4724 6334 4734 6390
rect 2798 6266 4734 6334
rect 2798 6210 2808 6266
rect 2864 6210 2932 6266
rect 2988 6210 3056 6266
rect 3112 6210 3180 6266
rect 3236 6210 3304 6266
rect 3360 6210 3428 6266
rect 3484 6210 3552 6266
rect 3608 6210 3676 6266
rect 3732 6210 3800 6266
rect 3856 6210 3924 6266
rect 3980 6210 4048 6266
rect 4104 6210 4172 6266
rect 4228 6210 4296 6266
rect 4352 6210 4420 6266
rect 4476 6210 4544 6266
rect 4600 6210 4668 6266
rect 4724 6210 4734 6266
rect 2798 6142 4734 6210
rect 2798 6086 2808 6142
rect 2864 6086 2932 6142
rect 2988 6086 3056 6142
rect 3112 6086 3180 6142
rect 3236 6086 3304 6142
rect 3360 6086 3428 6142
rect 3484 6086 3552 6142
rect 3608 6086 3676 6142
rect 3732 6086 3800 6142
rect 3856 6086 3924 6142
rect 3980 6086 4048 6142
rect 4104 6086 4172 6142
rect 4228 6086 4296 6142
rect 4352 6086 4420 6142
rect 4476 6086 4544 6142
rect 4600 6086 4668 6142
rect 4724 6086 4734 6142
rect 2798 6018 4734 6086
rect 2798 5962 2808 6018
rect 2864 5962 2932 6018
rect 2988 5962 3056 6018
rect 3112 5962 3180 6018
rect 3236 5962 3304 6018
rect 3360 5962 3428 6018
rect 3484 5962 3552 6018
rect 3608 5962 3676 6018
rect 3732 5962 3800 6018
rect 3856 5962 3924 6018
rect 3980 5962 4048 6018
rect 4104 5962 4172 6018
rect 4228 5962 4296 6018
rect 4352 5962 4420 6018
rect 4476 5962 4544 6018
rect 4600 5962 4668 6018
rect 4724 5962 4734 6018
rect 2798 5894 4734 5962
rect 2798 5838 2808 5894
rect 2864 5838 2932 5894
rect 2988 5838 3056 5894
rect 3112 5838 3180 5894
rect 3236 5838 3304 5894
rect 3360 5838 3428 5894
rect 3484 5838 3552 5894
rect 3608 5838 3676 5894
rect 3732 5838 3800 5894
rect 3856 5838 3924 5894
rect 3980 5838 4048 5894
rect 4104 5838 4172 5894
rect 4228 5838 4296 5894
rect 4352 5838 4420 5894
rect 4476 5838 4544 5894
rect 4600 5838 4668 5894
rect 4724 5838 4734 5894
rect 2798 5770 4734 5838
rect 2798 5714 2808 5770
rect 2864 5714 2932 5770
rect 2988 5714 3056 5770
rect 3112 5714 3180 5770
rect 3236 5714 3304 5770
rect 3360 5714 3428 5770
rect 3484 5714 3552 5770
rect 3608 5714 3676 5770
rect 3732 5714 3800 5770
rect 3856 5714 3924 5770
rect 3980 5714 4048 5770
rect 4104 5714 4172 5770
rect 4228 5714 4296 5770
rect 4352 5714 4420 5770
rect 4476 5714 4544 5770
rect 4600 5714 4668 5770
rect 4724 5714 4734 5770
rect 2798 5646 4734 5714
rect 2798 5590 2808 5646
rect 2864 5590 2932 5646
rect 2988 5590 3056 5646
rect 3112 5590 3180 5646
rect 3236 5590 3304 5646
rect 3360 5590 3428 5646
rect 3484 5590 3552 5646
rect 3608 5590 3676 5646
rect 3732 5590 3800 5646
rect 3856 5590 3924 5646
rect 3980 5590 4048 5646
rect 4104 5590 4172 5646
rect 4228 5590 4296 5646
rect 4352 5590 4420 5646
rect 4476 5590 4544 5646
rect 4600 5590 4668 5646
rect 4724 5590 4734 5646
rect 2798 5522 4734 5590
rect 2798 5466 2808 5522
rect 2864 5466 2932 5522
rect 2988 5466 3056 5522
rect 3112 5466 3180 5522
rect 3236 5466 3304 5522
rect 3360 5466 3428 5522
rect 3484 5466 3552 5522
rect 3608 5466 3676 5522
rect 3732 5466 3800 5522
rect 3856 5466 3924 5522
rect 3980 5466 4048 5522
rect 4104 5466 4172 5522
rect 4228 5466 4296 5522
rect 4352 5466 4420 5522
rect 4476 5466 4544 5522
rect 4600 5466 4668 5522
rect 4724 5466 4734 5522
rect 2798 5398 4734 5466
rect 2798 5342 2808 5398
rect 2864 5342 2932 5398
rect 2988 5342 3056 5398
rect 3112 5342 3180 5398
rect 3236 5342 3304 5398
rect 3360 5342 3428 5398
rect 3484 5342 3552 5398
rect 3608 5342 3676 5398
rect 3732 5342 3800 5398
rect 3856 5342 3924 5398
rect 3980 5342 4048 5398
rect 4104 5342 4172 5398
rect 4228 5342 4296 5398
rect 4352 5342 4420 5398
rect 4476 5342 4544 5398
rect 4600 5342 4668 5398
rect 4724 5342 4734 5398
rect 2798 5274 4734 5342
rect 2798 5218 2808 5274
rect 2864 5218 2932 5274
rect 2988 5218 3056 5274
rect 3112 5218 3180 5274
rect 3236 5218 3304 5274
rect 3360 5218 3428 5274
rect 3484 5218 3552 5274
rect 3608 5218 3676 5274
rect 3732 5218 3800 5274
rect 3856 5218 3924 5274
rect 3980 5218 4048 5274
rect 4104 5218 4172 5274
rect 4228 5218 4296 5274
rect 4352 5218 4420 5274
rect 4476 5218 4544 5274
rect 4600 5218 4668 5274
rect 4724 5218 4734 5274
rect 2798 5150 4734 5218
rect 2798 5094 2808 5150
rect 2864 5094 2932 5150
rect 2988 5094 3056 5150
rect 3112 5094 3180 5150
rect 3236 5094 3304 5150
rect 3360 5094 3428 5150
rect 3484 5094 3552 5150
rect 3608 5094 3676 5150
rect 3732 5094 3800 5150
rect 3856 5094 3924 5150
rect 3980 5094 4048 5150
rect 4104 5094 4172 5150
rect 4228 5094 4296 5150
rect 4352 5094 4420 5150
rect 4476 5094 4544 5150
rect 4600 5094 4668 5150
rect 4724 5094 4734 5150
rect 2798 5026 4734 5094
rect 2798 4970 2808 5026
rect 2864 4970 2932 5026
rect 2988 4970 3056 5026
rect 3112 4970 3180 5026
rect 3236 4970 3304 5026
rect 3360 4970 3428 5026
rect 3484 4970 3552 5026
rect 3608 4970 3676 5026
rect 3732 4970 3800 5026
rect 3856 4970 3924 5026
rect 3980 4970 4048 5026
rect 4104 4970 4172 5026
rect 4228 4970 4296 5026
rect 4352 4970 4420 5026
rect 4476 4970 4544 5026
rect 4600 4970 4668 5026
rect 4724 4970 4734 5026
rect 2798 4902 4734 4970
rect 2798 4846 2808 4902
rect 2864 4846 2932 4902
rect 2988 4846 3056 4902
rect 3112 4846 3180 4902
rect 3236 4846 3304 4902
rect 3360 4846 3428 4902
rect 3484 4846 3552 4902
rect 3608 4846 3676 4902
rect 3732 4846 3800 4902
rect 3856 4846 3924 4902
rect 3980 4846 4048 4902
rect 4104 4846 4172 4902
rect 4228 4846 4296 4902
rect 4352 4846 4420 4902
rect 4476 4846 4544 4902
rect 4600 4846 4668 4902
rect 4724 4846 4734 4902
rect 2798 4836 4734 4846
rect 5168 7754 7104 7764
rect 5168 7698 5178 7754
rect 5234 7698 5302 7754
rect 5358 7698 5426 7754
rect 5482 7698 5550 7754
rect 5606 7698 5674 7754
rect 5730 7698 5798 7754
rect 5854 7698 5922 7754
rect 5978 7698 6046 7754
rect 6102 7698 6170 7754
rect 6226 7698 6294 7754
rect 6350 7698 6418 7754
rect 6474 7698 6542 7754
rect 6598 7698 6666 7754
rect 6722 7698 6790 7754
rect 6846 7698 6914 7754
rect 6970 7698 7038 7754
rect 7094 7698 7104 7754
rect 5168 7630 7104 7698
rect 5168 7574 5178 7630
rect 5234 7574 5302 7630
rect 5358 7574 5426 7630
rect 5482 7574 5550 7630
rect 5606 7574 5674 7630
rect 5730 7574 5798 7630
rect 5854 7574 5922 7630
rect 5978 7574 6046 7630
rect 6102 7574 6170 7630
rect 6226 7574 6294 7630
rect 6350 7574 6418 7630
rect 6474 7574 6542 7630
rect 6598 7574 6666 7630
rect 6722 7574 6790 7630
rect 6846 7574 6914 7630
rect 6970 7574 7038 7630
rect 7094 7574 7104 7630
rect 5168 7506 7104 7574
rect 5168 7450 5178 7506
rect 5234 7450 5302 7506
rect 5358 7450 5426 7506
rect 5482 7450 5550 7506
rect 5606 7450 5674 7506
rect 5730 7450 5798 7506
rect 5854 7450 5922 7506
rect 5978 7450 6046 7506
rect 6102 7450 6170 7506
rect 6226 7450 6294 7506
rect 6350 7450 6418 7506
rect 6474 7450 6542 7506
rect 6598 7450 6666 7506
rect 6722 7450 6790 7506
rect 6846 7450 6914 7506
rect 6970 7450 7038 7506
rect 7094 7450 7104 7506
rect 5168 7382 7104 7450
rect 5168 7326 5178 7382
rect 5234 7326 5302 7382
rect 5358 7326 5426 7382
rect 5482 7326 5550 7382
rect 5606 7326 5674 7382
rect 5730 7326 5798 7382
rect 5854 7326 5922 7382
rect 5978 7326 6046 7382
rect 6102 7326 6170 7382
rect 6226 7326 6294 7382
rect 6350 7326 6418 7382
rect 6474 7326 6542 7382
rect 6598 7326 6666 7382
rect 6722 7326 6790 7382
rect 6846 7326 6914 7382
rect 6970 7326 7038 7382
rect 7094 7326 7104 7382
rect 5168 7258 7104 7326
rect 5168 7202 5178 7258
rect 5234 7202 5302 7258
rect 5358 7202 5426 7258
rect 5482 7202 5550 7258
rect 5606 7202 5674 7258
rect 5730 7202 5798 7258
rect 5854 7202 5922 7258
rect 5978 7202 6046 7258
rect 6102 7202 6170 7258
rect 6226 7202 6294 7258
rect 6350 7202 6418 7258
rect 6474 7202 6542 7258
rect 6598 7202 6666 7258
rect 6722 7202 6790 7258
rect 6846 7202 6914 7258
rect 6970 7202 7038 7258
rect 7094 7202 7104 7258
rect 5168 7134 7104 7202
rect 5168 7078 5178 7134
rect 5234 7078 5302 7134
rect 5358 7078 5426 7134
rect 5482 7078 5550 7134
rect 5606 7078 5674 7134
rect 5730 7078 5798 7134
rect 5854 7078 5922 7134
rect 5978 7078 6046 7134
rect 6102 7078 6170 7134
rect 6226 7078 6294 7134
rect 6350 7078 6418 7134
rect 6474 7078 6542 7134
rect 6598 7078 6666 7134
rect 6722 7078 6790 7134
rect 6846 7078 6914 7134
rect 6970 7078 7038 7134
rect 7094 7078 7104 7134
rect 5168 7010 7104 7078
rect 5168 6954 5178 7010
rect 5234 6954 5302 7010
rect 5358 6954 5426 7010
rect 5482 6954 5550 7010
rect 5606 6954 5674 7010
rect 5730 6954 5798 7010
rect 5854 6954 5922 7010
rect 5978 6954 6046 7010
rect 6102 6954 6170 7010
rect 6226 6954 6294 7010
rect 6350 6954 6418 7010
rect 6474 6954 6542 7010
rect 6598 6954 6666 7010
rect 6722 6954 6790 7010
rect 6846 6954 6914 7010
rect 6970 6954 7038 7010
rect 7094 6954 7104 7010
rect 5168 6886 7104 6954
rect 5168 6830 5178 6886
rect 5234 6830 5302 6886
rect 5358 6830 5426 6886
rect 5482 6830 5550 6886
rect 5606 6830 5674 6886
rect 5730 6830 5798 6886
rect 5854 6830 5922 6886
rect 5978 6830 6046 6886
rect 6102 6830 6170 6886
rect 6226 6830 6294 6886
rect 6350 6830 6418 6886
rect 6474 6830 6542 6886
rect 6598 6830 6666 6886
rect 6722 6830 6790 6886
rect 6846 6830 6914 6886
rect 6970 6830 7038 6886
rect 7094 6830 7104 6886
rect 5168 6762 7104 6830
rect 5168 6706 5178 6762
rect 5234 6706 5302 6762
rect 5358 6706 5426 6762
rect 5482 6706 5550 6762
rect 5606 6706 5674 6762
rect 5730 6706 5798 6762
rect 5854 6706 5922 6762
rect 5978 6706 6046 6762
rect 6102 6706 6170 6762
rect 6226 6706 6294 6762
rect 6350 6706 6418 6762
rect 6474 6706 6542 6762
rect 6598 6706 6666 6762
rect 6722 6706 6790 6762
rect 6846 6706 6914 6762
rect 6970 6706 7038 6762
rect 7094 6706 7104 6762
rect 5168 6638 7104 6706
rect 5168 6582 5178 6638
rect 5234 6582 5302 6638
rect 5358 6582 5426 6638
rect 5482 6582 5550 6638
rect 5606 6582 5674 6638
rect 5730 6582 5798 6638
rect 5854 6582 5922 6638
rect 5978 6582 6046 6638
rect 6102 6582 6170 6638
rect 6226 6582 6294 6638
rect 6350 6582 6418 6638
rect 6474 6582 6542 6638
rect 6598 6582 6666 6638
rect 6722 6582 6790 6638
rect 6846 6582 6914 6638
rect 6970 6582 7038 6638
rect 7094 6582 7104 6638
rect 5168 6514 7104 6582
rect 5168 6458 5178 6514
rect 5234 6458 5302 6514
rect 5358 6458 5426 6514
rect 5482 6458 5550 6514
rect 5606 6458 5674 6514
rect 5730 6458 5798 6514
rect 5854 6458 5922 6514
rect 5978 6458 6046 6514
rect 6102 6458 6170 6514
rect 6226 6458 6294 6514
rect 6350 6458 6418 6514
rect 6474 6458 6542 6514
rect 6598 6458 6666 6514
rect 6722 6458 6790 6514
rect 6846 6458 6914 6514
rect 6970 6458 7038 6514
rect 7094 6458 7104 6514
rect 5168 6390 7104 6458
rect 5168 6334 5178 6390
rect 5234 6334 5302 6390
rect 5358 6334 5426 6390
rect 5482 6334 5550 6390
rect 5606 6334 5674 6390
rect 5730 6334 5798 6390
rect 5854 6334 5922 6390
rect 5978 6334 6046 6390
rect 6102 6334 6170 6390
rect 6226 6334 6294 6390
rect 6350 6334 6418 6390
rect 6474 6334 6542 6390
rect 6598 6334 6666 6390
rect 6722 6334 6790 6390
rect 6846 6334 6914 6390
rect 6970 6334 7038 6390
rect 7094 6334 7104 6390
rect 5168 6266 7104 6334
rect 5168 6210 5178 6266
rect 5234 6210 5302 6266
rect 5358 6210 5426 6266
rect 5482 6210 5550 6266
rect 5606 6210 5674 6266
rect 5730 6210 5798 6266
rect 5854 6210 5922 6266
rect 5978 6210 6046 6266
rect 6102 6210 6170 6266
rect 6226 6210 6294 6266
rect 6350 6210 6418 6266
rect 6474 6210 6542 6266
rect 6598 6210 6666 6266
rect 6722 6210 6790 6266
rect 6846 6210 6914 6266
rect 6970 6210 7038 6266
rect 7094 6210 7104 6266
rect 5168 6142 7104 6210
rect 5168 6086 5178 6142
rect 5234 6086 5302 6142
rect 5358 6086 5426 6142
rect 5482 6086 5550 6142
rect 5606 6086 5674 6142
rect 5730 6086 5798 6142
rect 5854 6086 5922 6142
rect 5978 6086 6046 6142
rect 6102 6086 6170 6142
rect 6226 6086 6294 6142
rect 6350 6086 6418 6142
rect 6474 6086 6542 6142
rect 6598 6086 6666 6142
rect 6722 6086 6790 6142
rect 6846 6086 6914 6142
rect 6970 6086 7038 6142
rect 7094 6086 7104 6142
rect 5168 6018 7104 6086
rect 5168 5962 5178 6018
rect 5234 5962 5302 6018
rect 5358 5962 5426 6018
rect 5482 5962 5550 6018
rect 5606 5962 5674 6018
rect 5730 5962 5798 6018
rect 5854 5962 5922 6018
rect 5978 5962 6046 6018
rect 6102 5962 6170 6018
rect 6226 5962 6294 6018
rect 6350 5962 6418 6018
rect 6474 5962 6542 6018
rect 6598 5962 6666 6018
rect 6722 5962 6790 6018
rect 6846 5962 6914 6018
rect 6970 5962 7038 6018
rect 7094 5962 7104 6018
rect 5168 5894 7104 5962
rect 5168 5838 5178 5894
rect 5234 5838 5302 5894
rect 5358 5838 5426 5894
rect 5482 5838 5550 5894
rect 5606 5838 5674 5894
rect 5730 5838 5798 5894
rect 5854 5838 5922 5894
rect 5978 5838 6046 5894
rect 6102 5838 6170 5894
rect 6226 5838 6294 5894
rect 6350 5838 6418 5894
rect 6474 5838 6542 5894
rect 6598 5838 6666 5894
rect 6722 5838 6790 5894
rect 6846 5838 6914 5894
rect 6970 5838 7038 5894
rect 7094 5838 7104 5894
rect 5168 5770 7104 5838
rect 5168 5714 5178 5770
rect 5234 5714 5302 5770
rect 5358 5714 5426 5770
rect 5482 5714 5550 5770
rect 5606 5714 5674 5770
rect 5730 5714 5798 5770
rect 5854 5714 5922 5770
rect 5978 5714 6046 5770
rect 6102 5714 6170 5770
rect 6226 5714 6294 5770
rect 6350 5714 6418 5770
rect 6474 5714 6542 5770
rect 6598 5714 6666 5770
rect 6722 5714 6790 5770
rect 6846 5714 6914 5770
rect 6970 5714 7038 5770
rect 7094 5714 7104 5770
rect 5168 5646 7104 5714
rect 5168 5590 5178 5646
rect 5234 5590 5302 5646
rect 5358 5590 5426 5646
rect 5482 5590 5550 5646
rect 5606 5590 5674 5646
rect 5730 5590 5798 5646
rect 5854 5590 5922 5646
rect 5978 5590 6046 5646
rect 6102 5590 6170 5646
rect 6226 5590 6294 5646
rect 6350 5590 6418 5646
rect 6474 5590 6542 5646
rect 6598 5590 6666 5646
rect 6722 5590 6790 5646
rect 6846 5590 6914 5646
rect 6970 5590 7038 5646
rect 7094 5590 7104 5646
rect 5168 5522 7104 5590
rect 5168 5466 5178 5522
rect 5234 5466 5302 5522
rect 5358 5466 5426 5522
rect 5482 5466 5550 5522
rect 5606 5466 5674 5522
rect 5730 5466 5798 5522
rect 5854 5466 5922 5522
rect 5978 5466 6046 5522
rect 6102 5466 6170 5522
rect 6226 5466 6294 5522
rect 6350 5466 6418 5522
rect 6474 5466 6542 5522
rect 6598 5466 6666 5522
rect 6722 5466 6790 5522
rect 6846 5466 6914 5522
rect 6970 5466 7038 5522
rect 7094 5466 7104 5522
rect 5168 5398 7104 5466
rect 5168 5342 5178 5398
rect 5234 5342 5302 5398
rect 5358 5342 5426 5398
rect 5482 5342 5550 5398
rect 5606 5342 5674 5398
rect 5730 5342 5798 5398
rect 5854 5342 5922 5398
rect 5978 5342 6046 5398
rect 6102 5342 6170 5398
rect 6226 5342 6294 5398
rect 6350 5342 6418 5398
rect 6474 5342 6542 5398
rect 6598 5342 6666 5398
rect 6722 5342 6790 5398
rect 6846 5342 6914 5398
rect 6970 5342 7038 5398
rect 7094 5342 7104 5398
rect 5168 5274 7104 5342
rect 5168 5218 5178 5274
rect 5234 5218 5302 5274
rect 5358 5218 5426 5274
rect 5482 5218 5550 5274
rect 5606 5218 5674 5274
rect 5730 5218 5798 5274
rect 5854 5218 5922 5274
rect 5978 5218 6046 5274
rect 6102 5218 6170 5274
rect 6226 5218 6294 5274
rect 6350 5218 6418 5274
rect 6474 5218 6542 5274
rect 6598 5218 6666 5274
rect 6722 5218 6790 5274
rect 6846 5218 6914 5274
rect 6970 5218 7038 5274
rect 7094 5218 7104 5274
rect 5168 5150 7104 5218
rect 5168 5094 5178 5150
rect 5234 5094 5302 5150
rect 5358 5094 5426 5150
rect 5482 5094 5550 5150
rect 5606 5094 5674 5150
rect 5730 5094 5798 5150
rect 5854 5094 5922 5150
rect 5978 5094 6046 5150
rect 6102 5094 6170 5150
rect 6226 5094 6294 5150
rect 6350 5094 6418 5150
rect 6474 5094 6542 5150
rect 6598 5094 6666 5150
rect 6722 5094 6790 5150
rect 6846 5094 6914 5150
rect 6970 5094 7038 5150
rect 7094 5094 7104 5150
rect 5168 5026 7104 5094
rect 5168 4970 5178 5026
rect 5234 4970 5302 5026
rect 5358 4970 5426 5026
rect 5482 4970 5550 5026
rect 5606 4970 5674 5026
rect 5730 4970 5798 5026
rect 5854 4970 5922 5026
rect 5978 4970 6046 5026
rect 6102 4970 6170 5026
rect 6226 4970 6294 5026
rect 6350 4970 6418 5026
rect 6474 4970 6542 5026
rect 6598 4970 6666 5026
rect 6722 4970 6790 5026
rect 6846 4970 6914 5026
rect 6970 4970 7038 5026
rect 7094 4970 7104 5026
rect 5168 4902 7104 4970
rect 5168 4846 5178 4902
rect 5234 4846 5302 4902
rect 5358 4846 5426 4902
rect 5482 4846 5550 4902
rect 5606 4846 5674 4902
rect 5730 4846 5798 4902
rect 5854 4846 5922 4902
rect 5978 4846 6046 4902
rect 6102 4846 6170 4902
rect 6226 4846 6294 4902
rect 6350 4846 6418 4902
rect 6474 4846 6542 4902
rect 6598 4846 6666 4902
rect 6722 4846 6790 4902
rect 6846 4846 6914 4902
rect 6970 4846 7038 4902
rect 7094 4846 7104 4902
rect 5168 4836 7104 4846
rect 7874 7754 9810 7764
rect 7874 7698 7884 7754
rect 7940 7698 8008 7754
rect 8064 7698 8132 7754
rect 8188 7698 8256 7754
rect 8312 7698 8380 7754
rect 8436 7698 8504 7754
rect 8560 7698 8628 7754
rect 8684 7698 8752 7754
rect 8808 7698 8876 7754
rect 8932 7698 9000 7754
rect 9056 7698 9124 7754
rect 9180 7698 9248 7754
rect 9304 7698 9372 7754
rect 9428 7698 9496 7754
rect 9552 7698 9620 7754
rect 9676 7698 9744 7754
rect 9800 7698 9810 7754
rect 7874 7630 9810 7698
rect 7874 7574 7884 7630
rect 7940 7574 8008 7630
rect 8064 7574 8132 7630
rect 8188 7574 8256 7630
rect 8312 7574 8380 7630
rect 8436 7574 8504 7630
rect 8560 7574 8628 7630
rect 8684 7574 8752 7630
rect 8808 7574 8876 7630
rect 8932 7574 9000 7630
rect 9056 7574 9124 7630
rect 9180 7574 9248 7630
rect 9304 7574 9372 7630
rect 9428 7574 9496 7630
rect 9552 7574 9620 7630
rect 9676 7574 9744 7630
rect 9800 7574 9810 7630
rect 7874 7506 9810 7574
rect 7874 7450 7884 7506
rect 7940 7450 8008 7506
rect 8064 7450 8132 7506
rect 8188 7450 8256 7506
rect 8312 7450 8380 7506
rect 8436 7450 8504 7506
rect 8560 7450 8628 7506
rect 8684 7450 8752 7506
rect 8808 7450 8876 7506
rect 8932 7450 9000 7506
rect 9056 7450 9124 7506
rect 9180 7450 9248 7506
rect 9304 7450 9372 7506
rect 9428 7450 9496 7506
rect 9552 7450 9620 7506
rect 9676 7450 9744 7506
rect 9800 7450 9810 7506
rect 7874 7382 9810 7450
rect 7874 7326 7884 7382
rect 7940 7326 8008 7382
rect 8064 7326 8132 7382
rect 8188 7326 8256 7382
rect 8312 7326 8380 7382
rect 8436 7326 8504 7382
rect 8560 7326 8628 7382
rect 8684 7326 8752 7382
rect 8808 7326 8876 7382
rect 8932 7326 9000 7382
rect 9056 7326 9124 7382
rect 9180 7326 9248 7382
rect 9304 7326 9372 7382
rect 9428 7326 9496 7382
rect 9552 7326 9620 7382
rect 9676 7326 9744 7382
rect 9800 7326 9810 7382
rect 7874 7258 9810 7326
rect 7874 7202 7884 7258
rect 7940 7202 8008 7258
rect 8064 7202 8132 7258
rect 8188 7202 8256 7258
rect 8312 7202 8380 7258
rect 8436 7202 8504 7258
rect 8560 7202 8628 7258
rect 8684 7202 8752 7258
rect 8808 7202 8876 7258
rect 8932 7202 9000 7258
rect 9056 7202 9124 7258
rect 9180 7202 9248 7258
rect 9304 7202 9372 7258
rect 9428 7202 9496 7258
rect 9552 7202 9620 7258
rect 9676 7202 9744 7258
rect 9800 7202 9810 7258
rect 7874 7134 9810 7202
rect 7874 7078 7884 7134
rect 7940 7078 8008 7134
rect 8064 7078 8132 7134
rect 8188 7078 8256 7134
rect 8312 7078 8380 7134
rect 8436 7078 8504 7134
rect 8560 7078 8628 7134
rect 8684 7078 8752 7134
rect 8808 7078 8876 7134
rect 8932 7078 9000 7134
rect 9056 7078 9124 7134
rect 9180 7078 9248 7134
rect 9304 7078 9372 7134
rect 9428 7078 9496 7134
rect 9552 7078 9620 7134
rect 9676 7078 9744 7134
rect 9800 7078 9810 7134
rect 7874 7010 9810 7078
rect 7874 6954 7884 7010
rect 7940 6954 8008 7010
rect 8064 6954 8132 7010
rect 8188 6954 8256 7010
rect 8312 6954 8380 7010
rect 8436 6954 8504 7010
rect 8560 6954 8628 7010
rect 8684 6954 8752 7010
rect 8808 6954 8876 7010
rect 8932 6954 9000 7010
rect 9056 6954 9124 7010
rect 9180 6954 9248 7010
rect 9304 6954 9372 7010
rect 9428 6954 9496 7010
rect 9552 6954 9620 7010
rect 9676 6954 9744 7010
rect 9800 6954 9810 7010
rect 7874 6886 9810 6954
rect 7874 6830 7884 6886
rect 7940 6830 8008 6886
rect 8064 6830 8132 6886
rect 8188 6830 8256 6886
rect 8312 6830 8380 6886
rect 8436 6830 8504 6886
rect 8560 6830 8628 6886
rect 8684 6830 8752 6886
rect 8808 6830 8876 6886
rect 8932 6830 9000 6886
rect 9056 6830 9124 6886
rect 9180 6830 9248 6886
rect 9304 6830 9372 6886
rect 9428 6830 9496 6886
rect 9552 6830 9620 6886
rect 9676 6830 9744 6886
rect 9800 6830 9810 6886
rect 7874 6762 9810 6830
rect 7874 6706 7884 6762
rect 7940 6706 8008 6762
rect 8064 6706 8132 6762
rect 8188 6706 8256 6762
rect 8312 6706 8380 6762
rect 8436 6706 8504 6762
rect 8560 6706 8628 6762
rect 8684 6706 8752 6762
rect 8808 6706 8876 6762
rect 8932 6706 9000 6762
rect 9056 6706 9124 6762
rect 9180 6706 9248 6762
rect 9304 6706 9372 6762
rect 9428 6706 9496 6762
rect 9552 6706 9620 6762
rect 9676 6706 9744 6762
rect 9800 6706 9810 6762
rect 7874 6638 9810 6706
rect 7874 6582 7884 6638
rect 7940 6582 8008 6638
rect 8064 6582 8132 6638
rect 8188 6582 8256 6638
rect 8312 6582 8380 6638
rect 8436 6582 8504 6638
rect 8560 6582 8628 6638
rect 8684 6582 8752 6638
rect 8808 6582 8876 6638
rect 8932 6582 9000 6638
rect 9056 6582 9124 6638
rect 9180 6582 9248 6638
rect 9304 6582 9372 6638
rect 9428 6582 9496 6638
rect 9552 6582 9620 6638
rect 9676 6582 9744 6638
rect 9800 6582 9810 6638
rect 7874 6514 9810 6582
rect 7874 6458 7884 6514
rect 7940 6458 8008 6514
rect 8064 6458 8132 6514
rect 8188 6458 8256 6514
rect 8312 6458 8380 6514
rect 8436 6458 8504 6514
rect 8560 6458 8628 6514
rect 8684 6458 8752 6514
rect 8808 6458 8876 6514
rect 8932 6458 9000 6514
rect 9056 6458 9124 6514
rect 9180 6458 9248 6514
rect 9304 6458 9372 6514
rect 9428 6458 9496 6514
rect 9552 6458 9620 6514
rect 9676 6458 9744 6514
rect 9800 6458 9810 6514
rect 7874 6390 9810 6458
rect 7874 6334 7884 6390
rect 7940 6334 8008 6390
rect 8064 6334 8132 6390
rect 8188 6334 8256 6390
rect 8312 6334 8380 6390
rect 8436 6334 8504 6390
rect 8560 6334 8628 6390
rect 8684 6334 8752 6390
rect 8808 6334 8876 6390
rect 8932 6334 9000 6390
rect 9056 6334 9124 6390
rect 9180 6334 9248 6390
rect 9304 6334 9372 6390
rect 9428 6334 9496 6390
rect 9552 6334 9620 6390
rect 9676 6334 9744 6390
rect 9800 6334 9810 6390
rect 7874 6266 9810 6334
rect 7874 6210 7884 6266
rect 7940 6210 8008 6266
rect 8064 6210 8132 6266
rect 8188 6210 8256 6266
rect 8312 6210 8380 6266
rect 8436 6210 8504 6266
rect 8560 6210 8628 6266
rect 8684 6210 8752 6266
rect 8808 6210 8876 6266
rect 8932 6210 9000 6266
rect 9056 6210 9124 6266
rect 9180 6210 9248 6266
rect 9304 6210 9372 6266
rect 9428 6210 9496 6266
rect 9552 6210 9620 6266
rect 9676 6210 9744 6266
rect 9800 6210 9810 6266
rect 7874 6142 9810 6210
rect 7874 6086 7884 6142
rect 7940 6086 8008 6142
rect 8064 6086 8132 6142
rect 8188 6086 8256 6142
rect 8312 6086 8380 6142
rect 8436 6086 8504 6142
rect 8560 6086 8628 6142
rect 8684 6086 8752 6142
rect 8808 6086 8876 6142
rect 8932 6086 9000 6142
rect 9056 6086 9124 6142
rect 9180 6086 9248 6142
rect 9304 6086 9372 6142
rect 9428 6086 9496 6142
rect 9552 6086 9620 6142
rect 9676 6086 9744 6142
rect 9800 6086 9810 6142
rect 7874 6018 9810 6086
rect 7874 5962 7884 6018
rect 7940 5962 8008 6018
rect 8064 5962 8132 6018
rect 8188 5962 8256 6018
rect 8312 5962 8380 6018
rect 8436 5962 8504 6018
rect 8560 5962 8628 6018
rect 8684 5962 8752 6018
rect 8808 5962 8876 6018
rect 8932 5962 9000 6018
rect 9056 5962 9124 6018
rect 9180 5962 9248 6018
rect 9304 5962 9372 6018
rect 9428 5962 9496 6018
rect 9552 5962 9620 6018
rect 9676 5962 9744 6018
rect 9800 5962 9810 6018
rect 7874 5894 9810 5962
rect 7874 5838 7884 5894
rect 7940 5838 8008 5894
rect 8064 5838 8132 5894
rect 8188 5838 8256 5894
rect 8312 5838 8380 5894
rect 8436 5838 8504 5894
rect 8560 5838 8628 5894
rect 8684 5838 8752 5894
rect 8808 5838 8876 5894
rect 8932 5838 9000 5894
rect 9056 5838 9124 5894
rect 9180 5838 9248 5894
rect 9304 5838 9372 5894
rect 9428 5838 9496 5894
rect 9552 5838 9620 5894
rect 9676 5838 9744 5894
rect 9800 5838 9810 5894
rect 7874 5770 9810 5838
rect 7874 5714 7884 5770
rect 7940 5714 8008 5770
rect 8064 5714 8132 5770
rect 8188 5714 8256 5770
rect 8312 5714 8380 5770
rect 8436 5714 8504 5770
rect 8560 5714 8628 5770
rect 8684 5714 8752 5770
rect 8808 5714 8876 5770
rect 8932 5714 9000 5770
rect 9056 5714 9124 5770
rect 9180 5714 9248 5770
rect 9304 5714 9372 5770
rect 9428 5714 9496 5770
rect 9552 5714 9620 5770
rect 9676 5714 9744 5770
rect 9800 5714 9810 5770
rect 7874 5646 9810 5714
rect 7874 5590 7884 5646
rect 7940 5590 8008 5646
rect 8064 5590 8132 5646
rect 8188 5590 8256 5646
rect 8312 5590 8380 5646
rect 8436 5590 8504 5646
rect 8560 5590 8628 5646
rect 8684 5590 8752 5646
rect 8808 5590 8876 5646
rect 8932 5590 9000 5646
rect 9056 5590 9124 5646
rect 9180 5590 9248 5646
rect 9304 5590 9372 5646
rect 9428 5590 9496 5646
rect 9552 5590 9620 5646
rect 9676 5590 9744 5646
rect 9800 5590 9810 5646
rect 7874 5522 9810 5590
rect 7874 5466 7884 5522
rect 7940 5466 8008 5522
rect 8064 5466 8132 5522
rect 8188 5466 8256 5522
rect 8312 5466 8380 5522
rect 8436 5466 8504 5522
rect 8560 5466 8628 5522
rect 8684 5466 8752 5522
rect 8808 5466 8876 5522
rect 8932 5466 9000 5522
rect 9056 5466 9124 5522
rect 9180 5466 9248 5522
rect 9304 5466 9372 5522
rect 9428 5466 9496 5522
rect 9552 5466 9620 5522
rect 9676 5466 9744 5522
rect 9800 5466 9810 5522
rect 7874 5398 9810 5466
rect 7874 5342 7884 5398
rect 7940 5342 8008 5398
rect 8064 5342 8132 5398
rect 8188 5342 8256 5398
rect 8312 5342 8380 5398
rect 8436 5342 8504 5398
rect 8560 5342 8628 5398
rect 8684 5342 8752 5398
rect 8808 5342 8876 5398
rect 8932 5342 9000 5398
rect 9056 5342 9124 5398
rect 9180 5342 9248 5398
rect 9304 5342 9372 5398
rect 9428 5342 9496 5398
rect 9552 5342 9620 5398
rect 9676 5342 9744 5398
rect 9800 5342 9810 5398
rect 7874 5274 9810 5342
rect 7874 5218 7884 5274
rect 7940 5218 8008 5274
rect 8064 5218 8132 5274
rect 8188 5218 8256 5274
rect 8312 5218 8380 5274
rect 8436 5218 8504 5274
rect 8560 5218 8628 5274
rect 8684 5218 8752 5274
rect 8808 5218 8876 5274
rect 8932 5218 9000 5274
rect 9056 5218 9124 5274
rect 9180 5218 9248 5274
rect 9304 5218 9372 5274
rect 9428 5218 9496 5274
rect 9552 5218 9620 5274
rect 9676 5218 9744 5274
rect 9800 5218 9810 5274
rect 7874 5150 9810 5218
rect 7874 5094 7884 5150
rect 7940 5094 8008 5150
rect 8064 5094 8132 5150
rect 8188 5094 8256 5150
rect 8312 5094 8380 5150
rect 8436 5094 8504 5150
rect 8560 5094 8628 5150
rect 8684 5094 8752 5150
rect 8808 5094 8876 5150
rect 8932 5094 9000 5150
rect 9056 5094 9124 5150
rect 9180 5094 9248 5150
rect 9304 5094 9372 5150
rect 9428 5094 9496 5150
rect 9552 5094 9620 5150
rect 9676 5094 9744 5150
rect 9800 5094 9810 5150
rect 7874 5026 9810 5094
rect 7874 4970 7884 5026
rect 7940 4970 8008 5026
rect 8064 4970 8132 5026
rect 8188 4970 8256 5026
rect 8312 4970 8380 5026
rect 8436 4970 8504 5026
rect 8560 4970 8628 5026
rect 8684 4970 8752 5026
rect 8808 4970 8876 5026
rect 8932 4970 9000 5026
rect 9056 4970 9124 5026
rect 9180 4970 9248 5026
rect 9304 4970 9372 5026
rect 9428 4970 9496 5026
rect 9552 4970 9620 5026
rect 9676 4970 9744 5026
rect 9800 4970 9810 5026
rect 7874 4902 9810 4970
rect 7874 4846 7884 4902
rect 7940 4846 8008 4902
rect 8064 4846 8132 4902
rect 8188 4846 8256 4902
rect 8312 4846 8380 4902
rect 8436 4846 8504 4902
rect 8560 4846 8628 4902
rect 8684 4846 8752 4902
rect 8808 4846 8876 4902
rect 8932 4846 9000 4902
rect 9056 4846 9124 4902
rect 9180 4846 9248 4902
rect 9304 4846 9372 4902
rect 9428 4846 9496 4902
rect 9552 4846 9620 4902
rect 9676 4846 9744 4902
rect 9800 4846 9810 4902
rect 7874 4836 9810 4846
rect 10244 7754 12180 7764
rect 10244 7698 10254 7754
rect 10310 7698 10378 7754
rect 10434 7698 10502 7754
rect 10558 7698 10626 7754
rect 10682 7698 10750 7754
rect 10806 7698 10874 7754
rect 10930 7698 10998 7754
rect 11054 7698 11122 7754
rect 11178 7698 11246 7754
rect 11302 7698 11370 7754
rect 11426 7698 11494 7754
rect 11550 7698 11618 7754
rect 11674 7698 11742 7754
rect 11798 7698 11866 7754
rect 11922 7698 11990 7754
rect 12046 7698 12114 7754
rect 12170 7698 12180 7754
rect 10244 7630 12180 7698
rect 10244 7574 10254 7630
rect 10310 7574 10378 7630
rect 10434 7574 10502 7630
rect 10558 7574 10626 7630
rect 10682 7574 10750 7630
rect 10806 7574 10874 7630
rect 10930 7574 10998 7630
rect 11054 7574 11122 7630
rect 11178 7574 11246 7630
rect 11302 7574 11370 7630
rect 11426 7574 11494 7630
rect 11550 7574 11618 7630
rect 11674 7574 11742 7630
rect 11798 7574 11866 7630
rect 11922 7574 11990 7630
rect 12046 7574 12114 7630
rect 12170 7574 12180 7630
rect 10244 7506 12180 7574
rect 10244 7450 10254 7506
rect 10310 7450 10378 7506
rect 10434 7450 10502 7506
rect 10558 7450 10626 7506
rect 10682 7450 10750 7506
rect 10806 7450 10874 7506
rect 10930 7450 10998 7506
rect 11054 7450 11122 7506
rect 11178 7450 11246 7506
rect 11302 7450 11370 7506
rect 11426 7450 11494 7506
rect 11550 7450 11618 7506
rect 11674 7450 11742 7506
rect 11798 7450 11866 7506
rect 11922 7450 11990 7506
rect 12046 7450 12114 7506
rect 12170 7450 12180 7506
rect 10244 7382 12180 7450
rect 10244 7326 10254 7382
rect 10310 7326 10378 7382
rect 10434 7326 10502 7382
rect 10558 7326 10626 7382
rect 10682 7326 10750 7382
rect 10806 7326 10874 7382
rect 10930 7326 10998 7382
rect 11054 7326 11122 7382
rect 11178 7326 11246 7382
rect 11302 7326 11370 7382
rect 11426 7326 11494 7382
rect 11550 7326 11618 7382
rect 11674 7326 11742 7382
rect 11798 7326 11866 7382
rect 11922 7326 11990 7382
rect 12046 7326 12114 7382
rect 12170 7326 12180 7382
rect 10244 7258 12180 7326
rect 10244 7202 10254 7258
rect 10310 7202 10378 7258
rect 10434 7202 10502 7258
rect 10558 7202 10626 7258
rect 10682 7202 10750 7258
rect 10806 7202 10874 7258
rect 10930 7202 10998 7258
rect 11054 7202 11122 7258
rect 11178 7202 11246 7258
rect 11302 7202 11370 7258
rect 11426 7202 11494 7258
rect 11550 7202 11618 7258
rect 11674 7202 11742 7258
rect 11798 7202 11866 7258
rect 11922 7202 11990 7258
rect 12046 7202 12114 7258
rect 12170 7202 12180 7258
rect 10244 7134 12180 7202
rect 10244 7078 10254 7134
rect 10310 7078 10378 7134
rect 10434 7078 10502 7134
rect 10558 7078 10626 7134
rect 10682 7078 10750 7134
rect 10806 7078 10874 7134
rect 10930 7078 10998 7134
rect 11054 7078 11122 7134
rect 11178 7078 11246 7134
rect 11302 7078 11370 7134
rect 11426 7078 11494 7134
rect 11550 7078 11618 7134
rect 11674 7078 11742 7134
rect 11798 7078 11866 7134
rect 11922 7078 11990 7134
rect 12046 7078 12114 7134
rect 12170 7078 12180 7134
rect 10244 7010 12180 7078
rect 10244 6954 10254 7010
rect 10310 6954 10378 7010
rect 10434 6954 10502 7010
rect 10558 6954 10626 7010
rect 10682 6954 10750 7010
rect 10806 6954 10874 7010
rect 10930 6954 10998 7010
rect 11054 6954 11122 7010
rect 11178 6954 11246 7010
rect 11302 6954 11370 7010
rect 11426 6954 11494 7010
rect 11550 6954 11618 7010
rect 11674 6954 11742 7010
rect 11798 6954 11866 7010
rect 11922 6954 11990 7010
rect 12046 6954 12114 7010
rect 12170 6954 12180 7010
rect 10244 6886 12180 6954
rect 10244 6830 10254 6886
rect 10310 6830 10378 6886
rect 10434 6830 10502 6886
rect 10558 6830 10626 6886
rect 10682 6830 10750 6886
rect 10806 6830 10874 6886
rect 10930 6830 10998 6886
rect 11054 6830 11122 6886
rect 11178 6830 11246 6886
rect 11302 6830 11370 6886
rect 11426 6830 11494 6886
rect 11550 6830 11618 6886
rect 11674 6830 11742 6886
rect 11798 6830 11866 6886
rect 11922 6830 11990 6886
rect 12046 6830 12114 6886
rect 12170 6830 12180 6886
rect 10244 6762 12180 6830
rect 10244 6706 10254 6762
rect 10310 6706 10378 6762
rect 10434 6706 10502 6762
rect 10558 6706 10626 6762
rect 10682 6706 10750 6762
rect 10806 6706 10874 6762
rect 10930 6706 10998 6762
rect 11054 6706 11122 6762
rect 11178 6706 11246 6762
rect 11302 6706 11370 6762
rect 11426 6706 11494 6762
rect 11550 6706 11618 6762
rect 11674 6706 11742 6762
rect 11798 6706 11866 6762
rect 11922 6706 11990 6762
rect 12046 6706 12114 6762
rect 12170 6706 12180 6762
rect 10244 6638 12180 6706
rect 10244 6582 10254 6638
rect 10310 6582 10378 6638
rect 10434 6582 10502 6638
rect 10558 6582 10626 6638
rect 10682 6582 10750 6638
rect 10806 6582 10874 6638
rect 10930 6582 10998 6638
rect 11054 6582 11122 6638
rect 11178 6582 11246 6638
rect 11302 6582 11370 6638
rect 11426 6582 11494 6638
rect 11550 6582 11618 6638
rect 11674 6582 11742 6638
rect 11798 6582 11866 6638
rect 11922 6582 11990 6638
rect 12046 6582 12114 6638
rect 12170 6582 12180 6638
rect 10244 6514 12180 6582
rect 10244 6458 10254 6514
rect 10310 6458 10378 6514
rect 10434 6458 10502 6514
rect 10558 6458 10626 6514
rect 10682 6458 10750 6514
rect 10806 6458 10874 6514
rect 10930 6458 10998 6514
rect 11054 6458 11122 6514
rect 11178 6458 11246 6514
rect 11302 6458 11370 6514
rect 11426 6458 11494 6514
rect 11550 6458 11618 6514
rect 11674 6458 11742 6514
rect 11798 6458 11866 6514
rect 11922 6458 11990 6514
rect 12046 6458 12114 6514
rect 12170 6458 12180 6514
rect 10244 6390 12180 6458
rect 10244 6334 10254 6390
rect 10310 6334 10378 6390
rect 10434 6334 10502 6390
rect 10558 6334 10626 6390
rect 10682 6334 10750 6390
rect 10806 6334 10874 6390
rect 10930 6334 10998 6390
rect 11054 6334 11122 6390
rect 11178 6334 11246 6390
rect 11302 6334 11370 6390
rect 11426 6334 11494 6390
rect 11550 6334 11618 6390
rect 11674 6334 11742 6390
rect 11798 6334 11866 6390
rect 11922 6334 11990 6390
rect 12046 6334 12114 6390
rect 12170 6334 12180 6390
rect 10244 6266 12180 6334
rect 10244 6210 10254 6266
rect 10310 6210 10378 6266
rect 10434 6210 10502 6266
rect 10558 6210 10626 6266
rect 10682 6210 10750 6266
rect 10806 6210 10874 6266
rect 10930 6210 10998 6266
rect 11054 6210 11122 6266
rect 11178 6210 11246 6266
rect 11302 6210 11370 6266
rect 11426 6210 11494 6266
rect 11550 6210 11618 6266
rect 11674 6210 11742 6266
rect 11798 6210 11866 6266
rect 11922 6210 11990 6266
rect 12046 6210 12114 6266
rect 12170 6210 12180 6266
rect 10244 6142 12180 6210
rect 10244 6086 10254 6142
rect 10310 6086 10378 6142
rect 10434 6086 10502 6142
rect 10558 6086 10626 6142
rect 10682 6086 10750 6142
rect 10806 6086 10874 6142
rect 10930 6086 10998 6142
rect 11054 6086 11122 6142
rect 11178 6086 11246 6142
rect 11302 6086 11370 6142
rect 11426 6086 11494 6142
rect 11550 6086 11618 6142
rect 11674 6086 11742 6142
rect 11798 6086 11866 6142
rect 11922 6086 11990 6142
rect 12046 6086 12114 6142
rect 12170 6086 12180 6142
rect 10244 6018 12180 6086
rect 10244 5962 10254 6018
rect 10310 5962 10378 6018
rect 10434 5962 10502 6018
rect 10558 5962 10626 6018
rect 10682 5962 10750 6018
rect 10806 5962 10874 6018
rect 10930 5962 10998 6018
rect 11054 5962 11122 6018
rect 11178 5962 11246 6018
rect 11302 5962 11370 6018
rect 11426 5962 11494 6018
rect 11550 5962 11618 6018
rect 11674 5962 11742 6018
rect 11798 5962 11866 6018
rect 11922 5962 11990 6018
rect 12046 5962 12114 6018
rect 12170 5962 12180 6018
rect 10244 5894 12180 5962
rect 10244 5838 10254 5894
rect 10310 5838 10378 5894
rect 10434 5838 10502 5894
rect 10558 5838 10626 5894
rect 10682 5838 10750 5894
rect 10806 5838 10874 5894
rect 10930 5838 10998 5894
rect 11054 5838 11122 5894
rect 11178 5838 11246 5894
rect 11302 5838 11370 5894
rect 11426 5838 11494 5894
rect 11550 5838 11618 5894
rect 11674 5838 11742 5894
rect 11798 5838 11866 5894
rect 11922 5838 11990 5894
rect 12046 5838 12114 5894
rect 12170 5838 12180 5894
rect 10244 5770 12180 5838
rect 10244 5714 10254 5770
rect 10310 5714 10378 5770
rect 10434 5714 10502 5770
rect 10558 5714 10626 5770
rect 10682 5714 10750 5770
rect 10806 5714 10874 5770
rect 10930 5714 10998 5770
rect 11054 5714 11122 5770
rect 11178 5714 11246 5770
rect 11302 5714 11370 5770
rect 11426 5714 11494 5770
rect 11550 5714 11618 5770
rect 11674 5714 11742 5770
rect 11798 5714 11866 5770
rect 11922 5714 11990 5770
rect 12046 5714 12114 5770
rect 12170 5714 12180 5770
rect 10244 5646 12180 5714
rect 10244 5590 10254 5646
rect 10310 5590 10378 5646
rect 10434 5590 10502 5646
rect 10558 5590 10626 5646
rect 10682 5590 10750 5646
rect 10806 5590 10874 5646
rect 10930 5590 10998 5646
rect 11054 5590 11122 5646
rect 11178 5590 11246 5646
rect 11302 5590 11370 5646
rect 11426 5590 11494 5646
rect 11550 5590 11618 5646
rect 11674 5590 11742 5646
rect 11798 5590 11866 5646
rect 11922 5590 11990 5646
rect 12046 5590 12114 5646
rect 12170 5590 12180 5646
rect 10244 5522 12180 5590
rect 10244 5466 10254 5522
rect 10310 5466 10378 5522
rect 10434 5466 10502 5522
rect 10558 5466 10626 5522
rect 10682 5466 10750 5522
rect 10806 5466 10874 5522
rect 10930 5466 10998 5522
rect 11054 5466 11122 5522
rect 11178 5466 11246 5522
rect 11302 5466 11370 5522
rect 11426 5466 11494 5522
rect 11550 5466 11618 5522
rect 11674 5466 11742 5522
rect 11798 5466 11866 5522
rect 11922 5466 11990 5522
rect 12046 5466 12114 5522
rect 12170 5466 12180 5522
rect 10244 5398 12180 5466
rect 10244 5342 10254 5398
rect 10310 5342 10378 5398
rect 10434 5342 10502 5398
rect 10558 5342 10626 5398
rect 10682 5342 10750 5398
rect 10806 5342 10874 5398
rect 10930 5342 10998 5398
rect 11054 5342 11122 5398
rect 11178 5342 11246 5398
rect 11302 5342 11370 5398
rect 11426 5342 11494 5398
rect 11550 5342 11618 5398
rect 11674 5342 11742 5398
rect 11798 5342 11866 5398
rect 11922 5342 11990 5398
rect 12046 5342 12114 5398
rect 12170 5342 12180 5398
rect 10244 5274 12180 5342
rect 10244 5218 10254 5274
rect 10310 5218 10378 5274
rect 10434 5218 10502 5274
rect 10558 5218 10626 5274
rect 10682 5218 10750 5274
rect 10806 5218 10874 5274
rect 10930 5218 10998 5274
rect 11054 5218 11122 5274
rect 11178 5218 11246 5274
rect 11302 5218 11370 5274
rect 11426 5218 11494 5274
rect 11550 5218 11618 5274
rect 11674 5218 11742 5274
rect 11798 5218 11866 5274
rect 11922 5218 11990 5274
rect 12046 5218 12114 5274
rect 12170 5218 12180 5274
rect 10244 5150 12180 5218
rect 10244 5094 10254 5150
rect 10310 5094 10378 5150
rect 10434 5094 10502 5150
rect 10558 5094 10626 5150
rect 10682 5094 10750 5150
rect 10806 5094 10874 5150
rect 10930 5094 10998 5150
rect 11054 5094 11122 5150
rect 11178 5094 11246 5150
rect 11302 5094 11370 5150
rect 11426 5094 11494 5150
rect 11550 5094 11618 5150
rect 11674 5094 11742 5150
rect 11798 5094 11866 5150
rect 11922 5094 11990 5150
rect 12046 5094 12114 5150
rect 12170 5094 12180 5150
rect 10244 5026 12180 5094
rect 10244 4970 10254 5026
rect 10310 4970 10378 5026
rect 10434 4970 10502 5026
rect 10558 4970 10626 5026
rect 10682 4970 10750 5026
rect 10806 4970 10874 5026
rect 10930 4970 10998 5026
rect 11054 4970 11122 5026
rect 11178 4970 11246 5026
rect 11302 4970 11370 5026
rect 11426 4970 11494 5026
rect 11550 4970 11618 5026
rect 11674 4970 11742 5026
rect 11798 4970 11866 5026
rect 11922 4970 11990 5026
rect 12046 4970 12114 5026
rect 12170 4970 12180 5026
rect 10244 4902 12180 4970
rect 10244 4846 10254 4902
rect 10310 4846 10378 4902
rect 10434 4846 10502 4902
rect 10558 4846 10626 4902
rect 10682 4846 10750 4902
rect 10806 4846 10874 4902
rect 10930 4846 10998 4902
rect 11054 4846 11122 4902
rect 11178 4846 11246 4902
rect 11302 4846 11370 4902
rect 11426 4846 11494 4902
rect 11550 4846 11618 4902
rect 11674 4846 11742 4902
rect 11798 4846 11866 4902
rect 11922 4846 11990 4902
rect 12046 4846 12114 4902
rect 12170 4846 12180 4902
rect 10244 4836 12180 4846
rect 12861 7754 14673 7764
rect 12861 7698 12871 7754
rect 12927 7698 12995 7754
rect 13051 7698 13119 7754
rect 13175 7698 13243 7754
rect 13299 7698 13367 7754
rect 13423 7698 13491 7754
rect 13547 7698 13615 7754
rect 13671 7698 13739 7754
rect 13795 7698 13863 7754
rect 13919 7698 13987 7754
rect 14043 7698 14111 7754
rect 14167 7698 14235 7754
rect 14291 7698 14359 7754
rect 14415 7698 14483 7754
rect 14539 7698 14607 7754
rect 14663 7698 14673 7754
rect 12861 7630 14673 7698
rect 12861 7574 12871 7630
rect 12927 7574 12995 7630
rect 13051 7574 13119 7630
rect 13175 7574 13243 7630
rect 13299 7574 13367 7630
rect 13423 7574 13491 7630
rect 13547 7574 13615 7630
rect 13671 7574 13739 7630
rect 13795 7574 13863 7630
rect 13919 7574 13987 7630
rect 14043 7574 14111 7630
rect 14167 7574 14235 7630
rect 14291 7574 14359 7630
rect 14415 7574 14483 7630
rect 14539 7574 14607 7630
rect 14663 7574 14673 7630
rect 12861 7506 14673 7574
rect 12861 7450 12871 7506
rect 12927 7450 12995 7506
rect 13051 7450 13119 7506
rect 13175 7450 13243 7506
rect 13299 7450 13367 7506
rect 13423 7450 13491 7506
rect 13547 7450 13615 7506
rect 13671 7450 13739 7506
rect 13795 7450 13863 7506
rect 13919 7450 13987 7506
rect 14043 7450 14111 7506
rect 14167 7450 14235 7506
rect 14291 7450 14359 7506
rect 14415 7450 14483 7506
rect 14539 7450 14607 7506
rect 14663 7450 14673 7506
rect 12861 7382 14673 7450
rect 12861 7326 12871 7382
rect 12927 7326 12995 7382
rect 13051 7326 13119 7382
rect 13175 7326 13243 7382
rect 13299 7326 13367 7382
rect 13423 7326 13491 7382
rect 13547 7326 13615 7382
rect 13671 7326 13739 7382
rect 13795 7326 13863 7382
rect 13919 7326 13987 7382
rect 14043 7326 14111 7382
rect 14167 7326 14235 7382
rect 14291 7326 14359 7382
rect 14415 7326 14483 7382
rect 14539 7326 14607 7382
rect 14663 7326 14673 7382
rect 12861 7258 14673 7326
rect 12861 7202 12871 7258
rect 12927 7202 12995 7258
rect 13051 7202 13119 7258
rect 13175 7202 13243 7258
rect 13299 7202 13367 7258
rect 13423 7202 13491 7258
rect 13547 7202 13615 7258
rect 13671 7202 13739 7258
rect 13795 7202 13863 7258
rect 13919 7202 13987 7258
rect 14043 7202 14111 7258
rect 14167 7202 14235 7258
rect 14291 7202 14359 7258
rect 14415 7202 14483 7258
rect 14539 7202 14607 7258
rect 14663 7202 14673 7258
rect 12861 7134 14673 7202
rect 12861 7078 12871 7134
rect 12927 7078 12995 7134
rect 13051 7078 13119 7134
rect 13175 7078 13243 7134
rect 13299 7078 13367 7134
rect 13423 7078 13491 7134
rect 13547 7078 13615 7134
rect 13671 7078 13739 7134
rect 13795 7078 13863 7134
rect 13919 7078 13987 7134
rect 14043 7078 14111 7134
rect 14167 7078 14235 7134
rect 14291 7078 14359 7134
rect 14415 7078 14483 7134
rect 14539 7078 14607 7134
rect 14663 7078 14673 7134
rect 12861 7010 14673 7078
rect 12861 6954 12871 7010
rect 12927 6954 12995 7010
rect 13051 6954 13119 7010
rect 13175 6954 13243 7010
rect 13299 6954 13367 7010
rect 13423 6954 13491 7010
rect 13547 6954 13615 7010
rect 13671 6954 13739 7010
rect 13795 6954 13863 7010
rect 13919 6954 13987 7010
rect 14043 6954 14111 7010
rect 14167 6954 14235 7010
rect 14291 6954 14359 7010
rect 14415 6954 14483 7010
rect 14539 6954 14607 7010
rect 14663 6954 14673 7010
rect 12861 6886 14673 6954
rect 12861 6830 12871 6886
rect 12927 6830 12995 6886
rect 13051 6830 13119 6886
rect 13175 6830 13243 6886
rect 13299 6830 13367 6886
rect 13423 6830 13491 6886
rect 13547 6830 13615 6886
rect 13671 6830 13739 6886
rect 13795 6830 13863 6886
rect 13919 6830 13987 6886
rect 14043 6830 14111 6886
rect 14167 6830 14235 6886
rect 14291 6830 14359 6886
rect 14415 6830 14483 6886
rect 14539 6830 14607 6886
rect 14663 6830 14673 6886
rect 12861 6762 14673 6830
rect 12861 6706 12871 6762
rect 12927 6706 12995 6762
rect 13051 6706 13119 6762
rect 13175 6706 13243 6762
rect 13299 6706 13367 6762
rect 13423 6706 13491 6762
rect 13547 6706 13615 6762
rect 13671 6706 13739 6762
rect 13795 6706 13863 6762
rect 13919 6706 13987 6762
rect 14043 6706 14111 6762
rect 14167 6706 14235 6762
rect 14291 6706 14359 6762
rect 14415 6706 14483 6762
rect 14539 6706 14607 6762
rect 14663 6706 14673 6762
rect 12861 6638 14673 6706
rect 12861 6582 12871 6638
rect 12927 6582 12995 6638
rect 13051 6582 13119 6638
rect 13175 6582 13243 6638
rect 13299 6582 13367 6638
rect 13423 6582 13491 6638
rect 13547 6582 13615 6638
rect 13671 6582 13739 6638
rect 13795 6582 13863 6638
rect 13919 6582 13987 6638
rect 14043 6582 14111 6638
rect 14167 6582 14235 6638
rect 14291 6582 14359 6638
rect 14415 6582 14483 6638
rect 14539 6582 14607 6638
rect 14663 6582 14673 6638
rect 12861 6514 14673 6582
rect 12861 6458 12871 6514
rect 12927 6458 12995 6514
rect 13051 6458 13119 6514
rect 13175 6458 13243 6514
rect 13299 6458 13367 6514
rect 13423 6458 13491 6514
rect 13547 6458 13615 6514
rect 13671 6458 13739 6514
rect 13795 6458 13863 6514
rect 13919 6458 13987 6514
rect 14043 6458 14111 6514
rect 14167 6458 14235 6514
rect 14291 6458 14359 6514
rect 14415 6458 14483 6514
rect 14539 6458 14607 6514
rect 14663 6458 14673 6514
rect 12861 6390 14673 6458
rect 12861 6334 12871 6390
rect 12927 6334 12995 6390
rect 13051 6334 13119 6390
rect 13175 6334 13243 6390
rect 13299 6334 13367 6390
rect 13423 6334 13491 6390
rect 13547 6334 13615 6390
rect 13671 6334 13739 6390
rect 13795 6334 13863 6390
rect 13919 6334 13987 6390
rect 14043 6334 14111 6390
rect 14167 6334 14235 6390
rect 14291 6334 14359 6390
rect 14415 6334 14483 6390
rect 14539 6334 14607 6390
rect 14663 6334 14673 6390
rect 12861 6266 14673 6334
rect 12861 6210 12871 6266
rect 12927 6210 12995 6266
rect 13051 6210 13119 6266
rect 13175 6210 13243 6266
rect 13299 6210 13367 6266
rect 13423 6210 13491 6266
rect 13547 6210 13615 6266
rect 13671 6210 13739 6266
rect 13795 6210 13863 6266
rect 13919 6210 13987 6266
rect 14043 6210 14111 6266
rect 14167 6210 14235 6266
rect 14291 6210 14359 6266
rect 14415 6210 14483 6266
rect 14539 6210 14607 6266
rect 14663 6210 14673 6266
rect 12861 6142 14673 6210
rect 12861 6086 12871 6142
rect 12927 6086 12995 6142
rect 13051 6086 13119 6142
rect 13175 6086 13243 6142
rect 13299 6086 13367 6142
rect 13423 6086 13491 6142
rect 13547 6086 13615 6142
rect 13671 6086 13739 6142
rect 13795 6086 13863 6142
rect 13919 6086 13987 6142
rect 14043 6086 14111 6142
rect 14167 6086 14235 6142
rect 14291 6086 14359 6142
rect 14415 6086 14483 6142
rect 14539 6086 14607 6142
rect 14663 6086 14673 6142
rect 12861 6018 14673 6086
rect 12861 5962 12871 6018
rect 12927 5962 12995 6018
rect 13051 5962 13119 6018
rect 13175 5962 13243 6018
rect 13299 5962 13367 6018
rect 13423 5962 13491 6018
rect 13547 5962 13615 6018
rect 13671 5962 13739 6018
rect 13795 5962 13863 6018
rect 13919 5962 13987 6018
rect 14043 5962 14111 6018
rect 14167 5962 14235 6018
rect 14291 5962 14359 6018
rect 14415 5962 14483 6018
rect 14539 5962 14607 6018
rect 14663 5962 14673 6018
rect 12861 5894 14673 5962
rect 12861 5838 12871 5894
rect 12927 5838 12995 5894
rect 13051 5838 13119 5894
rect 13175 5838 13243 5894
rect 13299 5838 13367 5894
rect 13423 5838 13491 5894
rect 13547 5838 13615 5894
rect 13671 5838 13739 5894
rect 13795 5838 13863 5894
rect 13919 5838 13987 5894
rect 14043 5838 14111 5894
rect 14167 5838 14235 5894
rect 14291 5838 14359 5894
rect 14415 5838 14483 5894
rect 14539 5838 14607 5894
rect 14663 5838 14673 5894
rect 12861 5770 14673 5838
rect 12861 5714 12871 5770
rect 12927 5714 12995 5770
rect 13051 5714 13119 5770
rect 13175 5714 13243 5770
rect 13299 5714 13367 5770
rect 13423 5714 13491 5770
rect 13547 5714 13615 5770
rect 13671 5714 13739 5770
rect 13795 5714 13863 5770
rect 13919 5714 13987 5770
rect 14043 5714 14111 5770
rect 14167 5714 14235 5770
rect 14291 5714 14359 5770
rect 14415 5714 14483 5770
rect 14539 5714 14607 5770
rect 14663 5714 14673 5770
rect 12861 5646 14673 5714
rect 12861 5590 12871 5646
rect 12927 5590 12995 5646
rect 13051 5590 13119 5646
rect 13175 5590 13243 5646
rect 13299 5590 13367 5646
rect 13423 5590 13491 5646
rect 13547 5590 13615 5646
rect 13671 5590 13739 5646
rect 13795 5590 13863 5646
rect 13919 5590 13987 5646
rect 14043 5590 14111 5646
rect 14167 5590 14235 5646
rect 14291 5590 14359 5646
rect 14415 5590 14483 5646
rect 14539 5590 14607 5646
rect 14663 5590 14673 5646
rect 12861 5522 14673 5590
rect 12861 5466 12871 5522
rect 12927 5466 12995 5522
rect 13051 5466 13119 5522
rect 13175 5466 13243 5522
rect 13299 5466 13367 5522
rect 13423 5466 13491 5522
rect 13547 5466 13615 5522
rect 13671 5466 13739 5522
rect 13795 5466 13863 5522
rect 13919 5466 13987 5522
rect 14043 5466 14111 5522
rect 14167 5466 14235 5522
rect 14291 5466 14359 5522
rect 14415 5466 14483 5522
rect 14539 5466 14607 5522
rect 14663 5466 14673 5522
rect 12861 5398 14673 5466
rect 12861 5342 12871 5398
rect 12927 5342 12995 5398
rect 13051 5342 13119 5398
rect 13175 5342 13243 5398
rect 13299 5342 13367 5398
rect 13423 5342 13491 5398
rect 13547 5342 13615 5398
rect 13671 5342 13739 5398
rect 13795 5342 13863 5398
rect 13919 5342 13987 5398
rect 14043 5342 14111 5398
rect 14167 5342 14235 5398
rect 14291 5342 14359 5398
rect 14415 5342 14483 5398
rect 14539 5342 14607 5398
rect 14663 5342 14673 5398
rect 12861 5274 14673 5342
rect 12861 5218 12871 5274
rect 12927 5218 12995 5274
rect 13051 5218 13119 5274
rect 13175 5218 13243 5274
rect 13299 5218 13367 5274
rect 13423 5218 13491 5274
rect 13547 5218 13615 5274
rect 13671 5218 13739 5274
rect 13795 5218 13863 5274
rect 13919 5218 13987 5274
rect 14043 5218 14111 5274
rect 14167 5218 14235 5274
rect 14291 5218 14359 5274
rect 14415 5218 14483 5274
rect 14539 5218 14607 5274
rect 14663 5218 14673 5274
rect 12861 5150 14673 5218
rect 12861 5094 12871 5150
rect 12927 5094 12995 5150
rect 13051 5094 13119 5150
rect 13175 5094 13243 5150
rect 13299 5094 13367 5150
rect 13423 5094 13491 5150
rect 13547 5094 13615 5150
rect 13671 5094 13739 5150
rect 13795 5094 13863 5150
rect 13919 5094 13987 5150
rect 14043 5094 14111 5150
rect 14167 5094 14235 5150
rect 14291 5094 14359 5150
rect 14415 5094 14483 5150
rect 14539 5094 14607 5150
rect 14663 5094 14673 5150
rect 12861 5026 14673 5094
rect 12861 4970 12871 5026
rect 12927 4970 12995 5026
rect 13051 4970 13119 5026
rect 13175 4970 13243 5026
rect 13299 4970 13367 5026
rect 13423 4970 13491 5026
rect 13547 4970 13615 5026
rect 13671 4970 13739 5026
rect 13795 4970 13863 5026
rect 13919 4970 13987 5026
rect 14043 4970 14111 5026
rect 14167 4970 14235 5026
rect 14291 4970 14359 5026
rect 14415 4970 14483 5026
rect 14539 4970 14607 5026
rect 14663 4970 14673 5026
rect 12861 4902 14673 4970
rect 12861 4846 12871 4902
rect 12927 4846 12995 4902
rect 13051 4846 13119 4902
rect 13175 4846 13243 4902
rect 13299 4846 13367 4902
rect 13423 4846 13491 4902
rect 13547 4846 13615 4902
rect 13671 4846 13739 4902
rect 13795 4846 13863 4902
rect 13919 4846 13987 4902
rect 14043 4846 14111 4902
rect 14167 4846 14235 4902
rect 14291 4846 14359 4902
rect 14415 4846 14483 4902
rect 14539 4846 14607 4902
rect 14663 4846 14673 4902
rect 12861 4836 14673 4846
rect -11 4804 86 4814
rect 14892 4814 14902 7786
rect 14958 4814 14989 7786
rect 14892 4804 14989 4814
rect -11 4586 86 4596
rect -11 1614 20 4586
rect 76 1614 86 4586
rect 14892 4586 14989 4596
rect 305 4554 2117 4564
rect 305 4498 315 4554
rect 371 4498 439 4554
rect 495 4498 563 4554
rect 619 4498 687 4554
rect 743 4498 811 4554
rect 867 4498 935 4554
rect 991 4498 1059 4554
rect 1115 4498 1183 4554
rect 1239 4498 1307 4554
rect 1363 4498 1431 4554
rect 1487 4498 1555 4554
rect 1611 4498 1679 4554
rect 1735 4498 1803 4554
rect 1859 4498 1927 4554
rect 1983 4498 2051 4554
rect 2107 4498 2117 4554
rect 305 4430 2117 4498
rect 305 4374 315 4430
rect 371 4374 439 4430
rect 495 4374 563 4430
rect 619 4374 687 4430
rect 743 4374 811 4430
rect 867 4374 935 4430
rect 991 4374 1059 4430
rect 1115 4374 1183 4430
rect 1239 4374 1307 4430
rect 1363 4374 1431 4430
rect 1487 4374 1555 4430
rect 1611 4374 1679 4430
rect 1735 4374 1803 4430
rect 1859 4374 1927 4430
rect 1983 4374 2051 4430
rect 2107 4374 2117 4430
rect 305 4306 2117 4374
rect 305 4250 315 4306
rect 371 4250 439 4306
rect 495 4250 563 4306
rect 619 4250 687 4306
rect 743 4250 811 4306
rect 867 4250 935 4306
rect 991 4250 1059 4306
rect 1115 4250 1183 4306
rect 1239 4250 1307 4306
rect 1363 4250 1431 4306
rect 1487 4250 1555 4306
rect 1611 4250 1679 4306
rect 1735 4250 1803 4306
rect 1859 4250 1927 4306
rect 1983 4250 2051 4306
rect 2107 4250 2117 4306
rect 305 4182 2117 4250
rect 305 4126 315 4182
rect 371 4126 439 4182
rect 495 4126 563 4182
rect 619 4126 687 4182
rect 743 4126 811 4182
rect 867 4126 935 4182
rect 991 4126 1059 4182
rect 1115 4126 1183 4182
rect 1239 4126 1307 4182
rect 1363 4126 1431 4182
rect 1487 4126 1555 4182
rect 1611 4126 1679 4182
rect 1735 4126 1803 4182
rect 1859 4126 1927 4182
rect 1983 4126 2051 4182
rect 2107 4126 2117 4182
rect 305 4058 2117 4126
rect 305 4002 315 4058
rect 371 4002 439 4058
rect 495 4002 563 4058
rect 619 4002 687 4058
rect 743 4002 811 4058
rect 867 4002 935 4058
rect 991 4002 1059 4058
rect 1115 4002 1183 4058
rect 1239 4002 1307 4058
rect 1363 4002 1431 4058
rect 1487 4002 1555 4058
rect 1611 4002 1679 4058
rect 1735 4002 1803 4058
rect 1859 4002 1927 4058
rect 1983 4002 2051 4058
rect 2107 4002 2117 4058
rect 305 3934 2117 4002
rect 305 3878 315 3934
rect 371 3878 439 3934
rect 495 3878 563 3934
rect 619 3878 687 3934
rect 743 3878 811 3934
rect 867 3878 935 3934
rect 991 3878 1059 3934
rect 1115 3878 1183 3934
rect 1239 3878 1307 3934
rect 1363 3878 1431 3934
rect 1487 3878 1555 3934
rect 1611 3878 1679 3934
rect 1735 3878 1803 3934
rect 1859 3878 1927 3934
rect 1983 3878 2051 3934
rect 2107 3878 2117 3934
rect 305 3810 2117 3878
rect 305 3754 315 3810
rect 371 3754 439 3810
rect 495 3754 563 3810
rect 619 3754 687 3810
rect 743 3754 811 3810
rect 867 3754 935 3810
rect 991 3754 1059 3810
rect 1115 3754 1183 3810
rect 1239 3754 1307 3810
rect 1363 3754 1431 3810
rect 1487 3754 1555 3810
rect 1611 3754 1679 3810
rect 1735 3754 1803 3810
rect 1859 3754 1927 3810
rect 1983 3754 2051 3810
rect 2107 3754 2117 3810
rect 305 3686 2117 3754
rect 305 3630 315 3686
rect 371 3630 439 3686
rect 495 3630 563 3686
rect 619 3630 687 3686
rect 743 3630 811 3686
rect 867 3630 935 3686
rect 991 3630 1059 3686
rect 1115 3630 1183 3686
rect 1239 3630 1307 3686
rect 1363 3630 1431 3686
rect 1487 3630 1555 3686
rect 1611 3630 1679 3686
rect 1735 3630 1803 3686
rect 1859 3630 1927 3686
rect 1983 3630 2051 3686
rect 2107 3630 2117 3686
rect 305 3562 2117 3630
rect 305 3506 315 3562
rect 371 3506 439 3562
rect 495 3506 563 3562
rect 619 3506 687 3562
rect 743 3506 811 3562
rect 867 3506 935 3562
rect 991 3506 1059 3562
rect 1115 3506 1183 3562
rect 1239 3506 1307 3562
rect 1363 3506 1431 3562
rect 1487 3506 1555 3562
rect 1611 3506 1679 3562
rect 1735 3506 1803 3562
rect 1859 3506 1927 3562
rect 1983 3506 2051 3562
rect 2107 3506 2117 3562
rect 305 3438 2117 3506
rect 305 3382 315 3438
rect 371 3382 439 3438
rect 495 3382 563 3438
rect 619 3382 687 3438
rect 743 3382 811 3438
rect 867 3382 935 3438
rect 991 3382 1059 3438
rect 1115 3382 1183 3438
rect 1239 3382 1307 3438
rect 1363 3382 1431 3438
rect 1487 3382 1555 3438
rect 1611 3382 1679 3438
rect 1735 3382 1803 3438
rect 1859 3382 1927 3438
rect 1983 3382 2051 3438
rect 2107 3382 2117 3438
rect 305 3314 2117 3382
rect 305 3258 315 3314
rect 371 3258 439 3314
rect 495 3258 563 3314
rect 619 3258 687 3314
rect 743 3258 811 3314
rect 867 3258 935 3314
rect 991 3258 1059 3314
rect 1115 3258 1183 3314
rect 1239 3258 1307 3314
rect 1363 3258 1431 3314
rect 1487 3258 1555 3314
rect 1611 3258 1679 3314
rect 1735 3258 1803 3314
rect 1859 3258 1927 3314
rect 1983 3258 2051 3314
rect 2107 3258 2117 3314
rect 305 3190 2117 3258
rect 305 3134 315 3190
rect 371 3134 439 3190
rect 495 3134 563 3190
rect 619 3134 687 3190
rect 743 3134 811 3190
rect 867 3134 935 3190
rect 991 3134 1059 3190
rect 1115 3134 1183 3190
rect 1239 3134 1307 3190
rect 1363 3134 1431 3190
rect 1487 3134 1555 3190
rect 1611 3134 1679 3190
rect 1735 3134 1803 3190
rect 1859 3134 1927 3190
rect 1983 3134 2051 3190
rect 2107 3134 2117 3190
rect 305 3066 2117 3134
rect 305 3010 315 3066
rect 371 3010 439 3066
rect 495 3010 563 3066
rect 619 3010 687 3066
rect 743 3010 811 3066
rect 867 3010 935 3066
rect 991 3010 1059 3066
rect 1115 3010 1183 3066
rect 1239 3010 1307 3066
rect 1363 3010 1431 3066
rect 1487 3010 1555 3066
rect 1611 3010 1679 3066
rect 1735 3010 1803 3066
rect 1859 3010 1927 3066
rect 1983 3010 2051 3066
rect 2107 3010 2117 3066
rect 305 2942 2117 3010
rect 305 2886 315 2942
rect 371 2886 439 2942
rect 495 2886 563 2942
rect 619 2886 687 2942
rect 743 2886 811 2942
rect 867 2886 935 2942
rect 991 2886 1059 2942
rect 1115 2886 1183 2942
rect 1239 2886 1307 2942
rect 1363 2886 1431 2942
rect 1487 2886 1555 2942
rect 1611 2886 1679 2942
rect 1735 2886 1803 2942
rect 1859 2886 1927 2942
rect 1983 2886 2051 2942
rect 2107 2886 2117 2942
rect 305 2818 2117 2886
rect 305 2762 315 2818
rect 371 2762 439 2818
rect 495 2762 563 2818
rect 619 2762 687 2818
rect 743 2762 811 2818
rect 867 2762 935 2818
rect 991 2762 1059 2818
rect 1115 2762 1183 2818
rect 1239 2762 1307 2818
rect 1363 2762 1431 2818
rect 1487 2762 1555 2818
rect 1611 2762 1679 2818
rect 1735 2762 1803 2818
rect 1859 2762 1927 2818
rect 1983 2762 2051 2818
rect 2107 2762 2117 2818
rect 305 2694 2117 2762
rect 305 2638 315 2694
rect 371 2638 439 2694
rect 495 2638 563 2694
rect 619 2638 687 2694
rect 743 2638 811 2694
rect 867 2638 935 2694
rect 991 2638 1059 2694
rect 1115 2638 1183 2694
rect 1239 2638 1307 2694
rect 1363 2638 1431 2694
rect 1487 2638 1555 2694
rect 1611 2638 1679 2694
rect 1735 2638 1803 2694
rect 1859 2638 1927 2694
rect 1983 2638 2051 2694
rect 2107 2638 2117 2694
rect 305 2570 2117 2638
rect 305 2514 315 2570
rect 371 2514 439 2570
rect 495 2514 563 2570
rect 619 2514 687 2570
rect 743 2514 811 2570
rect 867 2514 935 2570
rect 991 2514 1059 2570
rect 1115 2514 1183 2570
rect 1239 2514 1307 2570
rect 1363 2514 1431 2570
rect 1487 2514 1555 2570
rect 1611 2514 1679 2570
rect 1735 2514 1803 2570
rect 1859 2514 1927 2570
rect 1983 2514 2051 2570
rect 2107 2514 2117 2570
rect 305 2446 2117 2514
rect 305 2390 315 2446
rect 371 2390 439 2446
rect 495 2390 563 2446
rect 619 2390 687 2446
rect 743 2390 811 2446
rect 867 2390 935 2446
rect 991 2390 1059 2446
rect 1115 2390 1183 2446
rect 1239 2390 1307 2446
rect 1363 2390 1431 2446
rect 1487 2390 1555 2446
rect 1611 2390 1679 2446
rect 1735 2390 1803 2446
rect 1859 2390 1927 2446
rect 1983 2390 2051 2446
rect 2107 2390 2117 2446
rect 305 2322 2117 2390
rect 305 2266 315 2322
rect 371 2266 439 2322
rect 495 2266 563 2322
rect 619 2266 687 2322
rect 743 2266 811 2322
rect 867 2266 935 2322
rect 991 2266 1059 2322
rect 1115 2266 1183 2322
rect 1239 2266 1307 2322
rect 1363 2266 1431 2322
rect 1487 2266 1555 2322
rect 1611 2266 1679 2322
rect 1735 2266 1803 2322
rect 1859 2266 1927 2322
rect 1983 2266 2051 2322
rect 2107 2266 2117 2322
rect 305 2198 2117 2266
rect 305 2142 315 2198
rect 371 2142 439 2198
rect 495 2142 563 2198
rect 619 2142 687 2198
rect 743 2142 811 2198
rect 867 2142 935 2198
rect 991 2142 1059 2198
rect 1115 2142 1183 2198
rect 1239 2142 1307 2198
rect 1363 2142 1431 2198
rect 1487 2142 1555 2198
rect 1611 2142 1679 2198
rect 1735 2142 1803 2198
rect 1859 2142 1927 2198
rect 1983 2142 2051 2198
rect 2107 2142 2117 2198
rect 305 2074 2117 2142
rect 305 2018 315 2074
rect 371 2018 439 2074
rect 495 2018 563 2074
rect 619 2018 687 2074
rect 743 2018 811 2074
rect 867 2018 935 2074
rect 991 2018 1059 2074
rect 1115 2018 1183 2074
rect 1239 2018 1307 2074
rect 1363 2018 1431 2074
rect 1487 2018 1555 2074
rect 1611 2018 1679 2074
rect 1735 2018 1803 2074
rect 1859 2018 1927 2074
rect 1983 2018 2051 2074
rect 2107 2018 2117 2074
rect 305 1950 2117 2018
rect 305 1894 315 1950
rect 371 1894 439 1950
rect 495 1894 563 1950
rect 619 1894 687 1950
rect 743 1894 811 1950
rect 867 1894 935 1950
rect 991 1894 1059 1950
rect 1115 1894 1183 1950
rect 1239 1894 1307 1950
rect 1363 1894 1431 1950
rect 1487 1894 1555 1950
rect 1611 1894 1679 1950
rect 1735 1894 1803 1950
rect 1859 1894 1927 1950
rect 1983 1894 2051 1950
rect 2107 1894 2117 1950
rect 305 1826 2117 1894
rect 305 1770 315 1826
rect 371 1770 439 1826
rect 495 1770 563 1826
rect 619 1770 687 1826
rect 743 1770 811 1826
rect 867 1770 935 1826
rect 991 1770 1059 1826
rect 1115 1770 1183 1826
rect 1239 1770 1307 1826
rect 1363 1770 1431 1826
rect 1487 1770 1555 1826
rect 1611 1770 1679 1826
rect 1735 1770 1803 1826
rect 1859 1770 1927 1826
rect 1983 1770 2051 1826
rect 2107 1770 2117 1826
rect 305 1702 2117 1770
rect 305 1646 315 1702
rect 371 1646 439 1702
rect 495 1646 563 1702
rect 619 1646 687 1702
rect 743 1646 811 1702
rect 867 1646 935 1702
rect 991 1646 1059 1702
rect 1115 1646 1183 1702
rect 1239 1646 1307 1702
rect 1363 1646 1431 1702
rect 1487 1646 1555 1702
rect 1611 1646 1679 1702
rect 1735 1646 1803 1702
rect 1859 1646 1927 1702
rect 1983 1646 2051 1702
rect 2107 1646 2117 1702
rect 305 1636 2117 1646
rect 2798 4554 4734 4564
rect 2798 4498 2808 4554
rect 2864 4498 2932 4554
rect 2988 4498 3056 4554
rect 3112 4498 3180 4554
rect 3236 4498 3304 4554
rect 3360 4498 3428 4554
rect 3484 4498 3552 4554
rect 3608 4498 3676 4554
rect 3732 4498 3800 4554
rect 3856 4498 3924 4554
rect 3980 4498 4048 4554
rect 4104 4498 4172 4554
rect 4228 4498 4296 4554
rect 4352 4498 4420 4554
rect 4476 4498 4544 4554
rect 4600 4498 4668 4554
rect 4724 4498 4734 4554
rect 2798 4430 4734 4498
rect 2798 4374 2808 4430
rect 2864 4374 2932 4430
rect 2988 4374 3056 4430
rect 3112 4374 3180 4430
rect 3236 4374 3304 4430
rect 3360 4374 3428 4430
rect 3484 4374 3552 4430
rect 3608 4374 3676 4430
rect 3732 4374 3800 4430
rect 3856 4374 3924 4430
rect 3980 4374 4048 4430
rect 4104 4374 4172 4430
rect 4228 4374 4296 4430
rect 4352 4374 4420 4430
rect 4476 4374 4544 4430
rect 4600 4374 4668 4430
rect 4724 4374 4734 4430
rect 2798 4306 4734 4374
rect 2798 4250 2808 4306
rect 2864 4250 2932 4306
rect 2988 4250 3056 4306
rect 3112 4250 3180 4306
rect 3236 4250 3304 4306
rect 3360 4250 3428 4306
rect 3484 4250 3552 4306
rect 3608 4250 3676 4306
rect 3732 4250 3800 4306
rect 3856 4250 3924 4306
rect 3980 4250 4048 4306
rect 4104 4250 4172 4306
rect 4228 4250 4296 4306
rect 4352 4250 4420 4306
rect 4476 4250 4544 4306
rect 4600 4250 4668 4306
rect 4724 4250 4734 4306
rect 2798 4182 4734 4250
rect 2798 4126 2808 4182
rect 2864 4126 2932 4182
rect 2988 4126 3056 4182
rect 3112 4126 3180 4182
rect 3236 4126 3304 4182
rect 3360 4126 3428 4182
rect 3484 4126 3552 4182
rect 3608 4126 3676 4182
rect 3732 4126 3800 4182
rect 3856 4126 3924 4182
rect 3980 4126 4048 4182
rect 4104 4126 4172 4182
rect 4228 4126 4296 4182
rect 4352 4126 4420 4182
rect 4476 4126 4544 4182
rect 4600 4126 4668 4182
rect 4724 4126 4734 4182
rect 2798 4058 4734 4126
rect 2798 4002 2808 4058
rect 2864 4002 2932 4058
rect 2988 4002 3056 4058
rect 3112 4002 3180 4058
rect 3236 4002 3304 4058
rect 3360 4002 3428 4058
rect 3484 4002 3552 4058
rect 3608 4002 3676 4058
rect 3732 4002 3800 4058
rect 3856 4002 3924 4058
rect 3980 4002 4048 4058
rect 4104 4002 4172 4058
rect 4228 4002 4296 4058
rect 4352 4002 4420 4058
rect 4476 4002 4544 4058
rect 4600 4002 4668 4058
rect 4724 4002 4734 4058
rect 2798 3934 4734 4002
rect 2798 3878 2808 3934
rect 2864 3878 2932 3934
rect 2988 3878 3056 3934
rect 3112 3878 3180 3934
rect 3236 3878 3304 3934
rect 3360 3878 3428 3934
rect 3484 3878 3552 3934
rect 3608 3878 3676 3934
rect 3732 3878 3800 3934
rect 3856 3878 3924 3934
rect 3980 3878 4048 3934
rect 4104 3878 4172 3934
rect 4228 3878 4296 3934
rect 4352 3878 4420 3934
rect 4476 3878 4544 3934
rect 4600 3878 4668 3934
rect 4724 3878 4734 3934
rect 2798 3810 4734 3878
rect 2798 3754 2808 3810
rect 2864 3754 2932 3810
rect 2988 3754 3056 3810
rect 3112 3754 3180 3810
rect 3236 3754 3304 3810
rect 3360 3754 3428 3810
rect 3484 3754 3552 3810
rect 3608 3754 3676 3810
rect 3732 3754 3800 3810
rect 3856 3754 3924 3810
rect 3980 3754 4048 3810
rect 4104 3754 4172 3810
rect 4228 3754 4296 3810
rect 4352 3754 4420 3810
rect 4476 3754 4544 3810
rect 4600 3754 4668 3810
rect 4724 3754 4734 3810
rect 2798 3686 4734 3754
rect 2798 3630 2808 3686
rect 2864 3630 2932 3686
rect 2988 3630 3056 3686
rect 3112 3630 3180 3686
rect 3236 3630 3304 3686
rect 3360 3630 3428 3686
rect 3484 3630 3552 3686
rect 3608 3630 3676 3686
rect 3732 3630 3800 3686
rect 3856 3630 3924 3686
rect 3980 3630 4048 3686
rect 4104 3630 4172 3686
rect 4228 3630 4296 3686
rect 4352 3630 4420 3686
rect 4476 3630 4544 3686
rect 4600 3630 4668 3686
rect 4724 3630 4734 3686
rect 2798 3562 4734 3630
rect 2798 3506 2808 3562
rect 2864 3506 2932 3562
rect 2988 3506 3056 3562
rect 3112 3506 3180 3562
rect 3236 3506 3304 3562
rect 3360 3506 3428 3562
rect 3484 3506 3552 3562
rect 3608 3506 3676 3562
rect 3732 3506 3800 3562
rect 3856 3506 3924 3562
rect 3980 3506 4048 3562
rect 4104 3506 4172 3562
rect 4228 3506 4296 3562
rect 4352 3506 4420 3562
rect 4476 3506 4544 3562
rect 4600 3506 4668 3562
rect 4724 3506 4734 3562
rect 2798 3438 4734 3506
rect 2798 3382 2808 3438
rect 2864 3382 2932 3438
rect 2988 3382 3056 3438
rect 3112 3382 3180 3438
rect 3236 3382 3304 3438
rect 3360 3382 3428 3438
rect 3484 3382 3552 3438
rect 3608 3382 3676 3438
rect 3732 3382 3800 3438
rect 3856 3382 3924 3438
rect 3980 3382 4048 3438
rect 4104 3382 4172 3438
rect 4228 3382 4296 3438
rect 4352 3382 4420 3438
rect 4476 3382 4544 3438
rect 4600 3382 4668 3438
rect 4724 3382 4734 3438
rect 2798 3314 4734 3382
rect 2798 3258 2808 3314
rect 2864 3258 2932 3314
rect 2988 3258 3056 3314
rect 3112 3258 3180 3314
rect 3236 3258 3304 3314
rect 3360 3258 3428 3314
rect 3484 3258 3552 3314
rect 3608 3258 3676 3314
rect 3732 3258 3800 3314
rect 3856 3258 3924 3314
rect 3980 3258 4048 3314
rect 4104 3258 4172 3314
rect 4228 3258 4296 3314
rect 4352 3258 4420 3314
rect 4476 3258 4544 3314
rect 4600 3258 4668 3314
rect 4724 3258 4734 3314
rect 2798 3190 4734 3258
rect 2798 3134 2808 3190
rect 2864 3134 2932 3190
rect 2988 3134 3056 3190
rect 3112 3134 3180 3190
rect 3236 3134 3304 3190
rect 3360 3134 3428 3190
rect 3484 3134 3552 3190
rect 3608 3134 3676 3190
rect 3732 3134 3800 3190
rect 3856 3134 3924 3190
rect 3980 3134 4048 3190
rect 4104 3134 4172 3190
rect 4228 3134 4296 3190
rect 4352 3134 4420 3190
rect 4476 3134 4544 3190
rect 4600 3134 4668 3190
rect 4724 3134 4734 3190
rect 2798 3066 4734 3134
rect 2798 3010 2808 3066
rect 2864 3010 2932 3066
rect 2988 3010 3056 3066
rect 3112 3010 3180 3066
rect 3236 3010 3304 3066
rect 3360 3010 3428 3066
rect 3484 3010 3552 3066
rect 3608 3010 3676 3066
rect 3732 3010 3800 3066
rect 3856 3010 3924 3066
rect 3980 3010 4048 3066
rect 4104 3010 4172 3066
rect 4228 3010 4296 3066
rect 4352 3010 4420 3066
rect 4476 3010 4544 3066
rect 4600 3010 4668 3066
rect 4724 3010 4734 3066
rect 2798 2942 4734 3010
rect 2798 2886 2808 2942
rect 2864 2886 2932 2942
rect 2988 2886 3056 2942
rect 3112 2886 3180 2942
rect 3236 2886 3304 2942
rect 3360 2886 3428 2942
rect 3484 2886 3552 2942
rect 3608 2886 3676 2942
rect 3732 2886 3800 2942
rect 3856 2886 3924 2942
rect 3980 2886 4048 2942
rect 4104 2886 4172 2942
rect 4228 2886 4296 2942
rect 4352 2886 4420 2942
rect 4476 2886 4544 2942
rect 4600 2886 4668 2942
rect 4724 2886 4734 2942
rect 2798 2818 4734 2886
rect 2798 2762 2808 2818
rect 2864 2762 2932 2818
rect 2988 2762 3056 2818
rect 3112 2762 3180 2818
rect 3236 2762 3304 2818
rect 3360 2762 3428 2818
rect 3484 2762 3552 2818
rect 3608 2762 3676 2818
rect 3732 2762 3800 2818
rect 3856 2762 3924 2818
rect 3980 2762 4048 2818
rect 4104 2762 4172 2818
rect 4228 2762 4296 2818
rect 4352 2762 4420 2818
rect 4476 2762 4544 2818
rect 4600 2762 4668 2818
rect 4724 2762 4734 2818
rect 2798 2694 4734 2762
rect 2798 2638 2808 2694
rect 2864 2638 2932 2694
rect 2988 2638 3056 2694
rect 3112 2638 3180 2694
rect 3236 2638 3304 2694
rect 3360 2638 3428 2694
rect 3484 2638 3552 2694
rect 3608 2638 3676 2694
rect 3732 2638 3800 2694
rect 3856 2638 3924 2694
rect 3980 2638 4048 2694
rect 4104 2638 4172 2694
rect 4228 2638 4296 2694
rect 4352 2638 4420 2694
rect 4476 2638 4544 2694
rect 4600 2638 4668 2694
rect 4724 2638 4734 2694
rect 2798 2570 4734 2638
rect 2798 2514 2808 2570
rect 2864 2514 2932 2570
rect 2988 2514 3056 2570
rect 3112 2514 3180 2570
rect 3236 2514 3304 2570
rect 3360 2514 3428 2570
rect 3484 2514 3552 2570
rect 3608 2514 3676 2570
rect 3732 2514 3800 2570
rect 3856 2514 3924 2570
rect 3980 2514 4048 2570
rect 4104 2514 4172 2570
rect 4228 2514 4296 2570
rect 4352 2514 4420 2570
rect 4476 2514 4544 2570
rect 4600 2514 4668 2570
rect 4724 2514 4734 2570
rect 2798 2446 4734 2514
rect 2798 2390 2808 2446
rect 2864 2390 2932 2446
rect 2988 2390 3056 2446
rect 3112 2390 3180 2446
rect 3236 2390 3304 2446
rect 3360 2390 3428 2446
rect 3484 2390 3552 2446
rect 3608 2390 3676 2446
rect 3732 2390 3800 2446
rect 3856 2390 3924 2446
rect 3980 2390 4048 2446
rect 4104 2390 4172 2446
rect 4228 2390 4296 2446
rect 4352 2390 4420 2446
rect 4476 2390 4544 2446
rect 4600 2390 4668 2446
rect 4724 2390 4734 2446
rect 2798 2322 4734 2390
rect 2798 2266 2808 2322
rect 2864 2266 2932 2322
rect 2988 2266 3056 2322
rect 3112 2266 3180 2322
rect 3236 2266 3304 2322
rect 3360 2266 3428 2322
rect 3484 2266 3552 2322
rect 3608 2266 3676 2322
rect 3732 2266 3800 2322
rect 3856 2266 3924 2322
rect 3980 2266 4048 2322
rect 4104 2266 4172 2322
rect 4228 2266 4296 2322
rect 4352 2266 4420 2322
rect 4476 2266 4544 2322
rect 4600 2266 4668 2322
rect 4724 2266 4734 2322
rect 2798 2198 4734 2266
rect 2798 2142 2808 2198
rect 2864 2142 2932 2198
rect 2988 2142 3056 2198
rect 3112 2142 3180 2198
rect 3236 2142 3304 2198
rect 3360 2142 3428 2198
rect 3484 2142 3552 2198
rect 3608 2142 3676 2198
rect 3732 2142 3800 2198
rect 3856 2142 3924 2198
rect 3980 2142 4048 2198
rect 4104 2142 4172 2198
rect 4228 2142 4296 2198
rect 4352 2142 4420 2198
rect 4476 2142 4544 2198
rect 4600 2142 4668 2198
rect 4724 2142 4734 2198
rect 2798 2074 4734 2142
rect 2798 2018 2808 2074
rect 2864 2018 2932 2074
rect 2988 2018 3056 2074
rect 3112 2018 3180 2074
rect 3236 2018 3304 2074
rect 3360 2018 3428 2074
rect 3484 2018 3552 2074
rect 3608 2018 3676 2074
rect 3732 2018 3800 2074
rect 3856 2018 3924 2074
rect 3980 2018 4048 2074
rect 4104 2018 4172 2074
rect 4228 2018 4296 2074
rect 4352 2018 4420 2074
rect 4476 2018 4544 2074
rect 4600 2018 4668 2074
rect 4724 2018 4734 2074
rect 2798 1950 4734 2018
rect 2798 1894 2808 1950
rect 2864 1894 2932 1950
rect 2988 1894 3056 1950
rect 3112 1894 3180 1950
rect 3236 1894 3304 1950
rect 3360 1894 3428 1950
rect 3484 1894 3552 1950
rect 3608 1894 3676 1950
rect 3732 1894 3800 1950
rect 3856 1894 3924 1950
rect 3980 1894 4048 1950
rect 4104 1894 4172 1950
rect 4228 1894 4296 1950
rect 4352 1894 4420 1950
rect 4476 1894 4544 1950
rect 4600 1894 4668 1950
rect 4724 1894 4734 1950
rect 2798 1826 4734 1894
rect 2798 1770 2808 1826
rect 2864 1770 2932 1826
rect 2988 1770 3056 1826
rect 3112 1770 3180 1826
rect 3236 1770 3304 1826
rect 3360 1770 3428 1826
rect 3484 1770 3552 1826
rect 3608 1770 3676 1826
rect 3732 1770 3800 1826
rect 3856 1770 3924 1826
rect 3980 1770 4048 1826
rect 4104 1770 4172 1826
rect 4228 1770 4296 1826
rect 4352 1770 4420 1826
rect 4476 1770 4544 1826
rect 4600 1770 4668 1826
rect 4724 1770 4734 1826
rect 2798 1702 4734 1770
rect 2798 1646 2808 1702
rect 2864 1646 2932 1702
rect 2988 1646 3056 1702
rect 3112 1646 3180 1702
rect 3236 1646 3304 1702
rect 3360 1646 3428 1702
rect 3484 1646 3552 1702
rect 3608 1646 3676 1702
rect 3732 1646 3800 1702
rect 3856 1646 3924 1702
rect 3980 1646 4048 1702
rect 4104 1646 4172 1702
rect 4228 1646 4296 1702
rect 4352 1646 4420 1702
rect 4476 1646 4544 1702
rect 4600 1646 4668 1702
rect 4724 1646 4734 1702
rect 2798 1636 4734 1646
rect 5168 4554 7104 4564
rect 5168 4498 5178 4554
rect 5234 4498 5302 4554
rect 5358 4498 5426 4554
rect 5482 4498 5550 4554
rect 5606 4498 5674 4554
rect 5730 4498 5798 4554
rect 5854 4498 5922 4554
rect 5978 4498 6046 4554
rect 6102 4498 6170 4554
rect 6226 4498 6294 4554
rect 6350 4498 6418 4554
rect 6474 4498 6542 4554
rect 6598 4498 6666 4554
rect 6722 4498 6790 4554
rect 6846 4498 6914 4554
rect 6970 4498 7038 4554
rect 7094 4498 7104 4554
rect 5168 4430 7104 4498
rect 5168 4374 5178 4430
rect 5234 4374 5302 4430
rect 5358 4374 5426 4430
rect 5482 4374 5550 4430
rect 5606 4374 5674 4430
rect 5730 4374 5798 4430
rect 5854 4374 5922 4430
rect 5978 4374 6046 4430
rect 6102 4374 6170 4430
rect 6226 4374 6294 4430
rect 6350 4374 6418 4430
rect 6474 4374 6542 4430
rect 6598 4374 6666 4430
rect 6722 4374 6790 4430
rect 6846 4374 6914 4430
rect 6970 4374 7038 4430
rect 7094 4374 7104 4430
rect 5168 4306 7104 4374
rect 5168 4250 5178 4306
rect 5234 4250 5302 4306
rect 5358 4250 5426 4306
rect 5482 4250 5550 4306
rect 5606 4250 5674 4306
rect 5730 4250 5798 4306
rect 5854 4250 5922 4306
rect 5978 4250 6046 4306
rect 6102 4250 6170 4306
rect 6226 4250 6294 4306
rect 6350 4250 6418 4306
rect 6474 4250 6542 4306
rect 6598 4250 6666 4306
rect 6722 4250 6790 4306
rect 6846 4250 6914 4306
rect 6970 4250 7038 4306
rect 7094 4250 7104 4306
rect 5168 4182 7104 4250
rect 5168 4126 5178 4182
rect 5234 4126 5302 4182
rect 5358 4126 5426 4182
rect 5482 4126 5550 4182
rect 5606 4126 5674 4182
rect 5730 4126 5798 4182
rect 5854 4126 5922 4182
rect 5978 4126 6046 4182
rect 6102 4126 6170 4182
rect 6226 4126 6294 4182
rect 6350 4126 6418 4182
rect 6474 4126 6542 4182
rect 6598 4126 6666 4182
rect 6722 4126 6790 4182
rect 6846 4126 6914 4182
rect 6970 4126 7038 4182
rect 7094 4126 7104 4182
rect 5168 4058 7104 4126
rect 5168 4002 5178 4058
rect 5234 4002 5302 4058
rect 5358 4002 5426 4058
rect 5482 4002 5550 4058
rect 5606 4002 5674 4058
rect 5730 4002 5798 4058
rect 5854 4002 5922 4058
rect 5978 4002 6046 4058
rect 6102 4002 6170 4058
rect 6226 4002 6294 4058
rect 6350 4002 6418 4058
rect 6474 4002 6542 4058
rect 6598 4002 6666 4058
rect 6722 4002 6790 4058
rect 6846 4002 6914 4058
rect 6970 4002 7038 4058
rect 7094 4002 7104 4058
rect 5168 3934 7104 4002
rect 5168 3878 5178 3934
rect 5234 3878 5302 3934
rect 5358 3878 5426 3934
rect 5482 3878 5550 3934
rect 5606 3878 5674 3934
rect 5730 3878 5798 3934
rect 5854 3878 5922 3934
rect 5978 3878 6046 3934
rect 6102 3878 6170 3934
rect 6226 3878 6294 3934
rect 6350 3878 6418 3934
rect 6474 3878 6542 3934
rect 6598 3878 6666 3934
rect 6722 3878 6790 3934
rect 6846 3878 6914 3934
rect 6970 3878 7038 3934
rect 7094 3878 7104 3934
rect 5168 3810 7104 3878
rect 5168 3754 5178 3810
rect 5234 3754 5302 3810
rect 5358 3754 5426 3810
rect 5482 3754 5550 3810
rect 5606 3754 5674 3810
rect 5730 3754 5798 3810
rect 5854 3754 5922 3810
rect 5978 3754 6046 3810
rect 6102 3754 6170 3810
rect 6226 3754 6294 3810
rect 6350 3754 6418 3810
rect 6474 3754 6542 3810
rect 6598 3754 6666 3810
rect 6722 3754 6790 3810
rect 6846 3754 6914 3810
rect 6970 3754 7038 3810
rect 7094 3754 7104 3810
rect 5168 3686 7104 3754
rect 5168 3630 5178 3686
rect 5234 3630 5302 3686
rect 5358 3630 5426 3686
rect 5482 3630 5550 3686
rect 5606 3630 5674 3686
rect 5730 3630 5798 3686
rect 5854 3630 5922 3686
rect 5978 3630 6046 3686
rect 6102 3630 6170 3686
rect 6226 3630 6294 3686
rect 6350 3630 6418 3686
rect 6474 3630 6542 3686
rect 6598 3630 6666 3686
rect 6722 3630 6790 3686
rect 6846 3630 6914 3686
rect 6970 3630 7038 3686
rect 7094 3630 7104 3686
rect 5168 3562 7104 3630
rect 5168 3506 5178 3562
rect 5234 3506 5302 3562
rect 5358 3506 5426 3562
rect 5482 3506 5550 3562
rect 5606 3506 5674 3562
rect 5730 3506 5798 3562
rect 5854 3506 5922 3562
rect 5978 3506 6046 3562
rect 6102 3506 6170 3562
rect 6226 3506 6294 3562
rect 6350 3506 6418 3562
rect 6474 3506 6542 3562
rect 6598 3506 6666 3562
rect 6722 3506 6790 3562
rect 6846 3506 6914 3562
rect 6970 3506 7038 3562
rect 7094 3506 7104 3562
rect 5168 3438 7104 3506
rect 5168 3382 5178 3438
rect 5234 3382 5302 3438
rect 5358 3382 5426 3438
rect 5482 3382 5550 3438
rect 5606 3382 5674 3438
rect 5730 3382 5798 3438
rect 5854 3382 5922 3438
rect 5978 3382 6046 3438
rect 6102 3382 6170 3438
rect 6226 3382 6294 3438
rect 6350 3382 6418 3438
rect 6474 3382 6542 3438
rect 6598 3382 6666 3438
rect 6722 3382 6790 3438
rect 6846 3382 6914 3438
rect 6970 3382 7038 3438
rect 7094 3382 7104 3438
rect 5168 3314 7104 3382
rect 5168 3258 5178 3314
rect 5234 3258 5302 3314
rect 5358 3258 5426 3314
rect 5482 3258 5550 3314
rect 5606 3258 5674 3314
rect 5730 3258 5798 3314
rect 5854 3258 5922 3314
rect 5978 3258 6046 3314
rect 6102 3258 6170 3314
rect 6226 3258 6294 3314
rect 6350 3258 6418 3314
rect 6474 3258 6542 3314
rect 6598 3258 6666 3314
rect 6722 3258 6790 3314
rect 6846 3258 6914 3314
rect 6970 3258 7038 3314
rect 7094 3258 7104 3314
rect 5168 3190 7104 3258
rect 5168 3134 5178 3190
rect 5234 3134 5302 3190
rect 5358 3134 5426 3190
rect 5482 3134 5550 3190
rect 5606 3134 5674 3190
rect 5730 3134 5798 3190
rect 5854 3134 5922 3190
rect 5978 3134 6046 3190
rect 6102 3134 6170 3190
rect 6226 3134 6294 3190
rect 6350 3134 6418 3190
rect 6474 3134 6542 3190
rect 6598 3134 6666 3190
rect 6722 3134 6790 3190
rect 6846 3134 6914 3190
rect 6970 3134 7038 3190
rect 7094 3134 7104 3190
rect 5168 3066 7104 3134
rect 5168 3010 5178 3066
rect 5234 3010 5302 3066
rect 5358 3010 5426 3066
rect 5482 3010 5550 3066
rect 5606 3010 5674 3066
rect 5730 3010 5798 3066
rect 5854 3010 5922 3066
rect 5978 3010 6046 3066
rect 6102 3010 6170 3066
rect 6226 3010 6294 3066
rect 6350 3010 6418 3066
rect 6474 3010 6542 3066
rect 6598 3010 6666 3066
rect 6722 3010 6790 3066
rect 6846 3010 6914 3066
rect 6970 3010 7038 3066
rect 7094 3010 7104 3066
rect 5168 2942 7104 3010
rect 5168 2886 5178 2942
rect 5234 2886 5302 2942
rect 5358 2886 5426 2942
rect 5482 2886 5550 2942
rect 5606 2886 5674 2942
rect 5730 2886 5798 2942
rect 5854 2886 5922 2942
rect 5978 2886 6046 2942
rect 6102 2886 6170 2942
rect 6226 2886 6294 2942
rect 6350 2886 6418 2942
rect 6474 2886 6542 2942
rect 6598 2886 6666 2942
rect 6722 2886 6790 2942
rect 6846 2886 6914 2942
rect 6970 2886 7038 2942
rect 7094 2886 7104 2942
rect 5168 2818 7104 2886
rect 5168 2762 5178 2818
rect 5234 2762 5302 2818
rect 5358 2762 5426 2818
rect 5482 2762 5550 2818
rect 5606 2762 5674 2818
rect 5730 2762 5798 2818
rect 5854 2762 5922 2818
rect 5978 2762 6046 2818
rect 6102 2762 6170 2818
rect 6226 2762 6294 2818
rect 6350 2762 6418 2818
rect 6474 2762 6542 2818
rect 6598 2762 6666 2818
rect 6722 2762 6790 2818
rect 6846 2762 6914 2818
rect 6970 2762 7038 2818
rect 7094 2762 7104 2818
rect 5168 2694 7104 2762
rect 5168 2638 5178 2694
rect 5234 2638 5302 2694
rect 5358 2638 5426 2694
rect 5482 2638 5550 2694
rect 5606 2638 5674 2694
rect 5730 2638 5798 2694
rect 5854 2638 5922 2694
rect 5978 2638 6046 2694
rect 6102 2638 6170 2694
rect 6226 2638 6294 2694
rect 6350 2638 6418 2694
rect 6474 2638 6542 2694
rect 6598 2638 6666 2694
rect 6722 2638 6790 2694
rect 6846 2638 6914 2694
rect 6970 2638 7038 2694
rect 7094 2638 7104 2694
rect 5168 2570 7104 2638
rect 5168 2514 5178 2570
rect 5234 2514 5302 2570
rect 5358 2514 5426 2570
rect 5482 2514 5550 2570
rect 5606 2514 5674 2570
rect 5730 2514 5798 2570
rect 5854 2514 5922 2570
rect 5978 2514 6046 2570
rect 6102 2514 6170 2570
rect 6226 2514 6294 2570
rect 6350 2514 6418 2570
rect 6474 2514 6542 2570
rect 6598 2514 6666 2570
rect 6722 2514 6790 2570
rect 6846 2514 6914 2570
rect 6970 2514 7038 2570
rect 7094 2514 7104 2570
rect 5168 2446 7104 2514
rect 5168 2390 5178 2446
rect 5234 2390 5302 2446
rect 5358 2390 5426 2446
rect 5482 2390 5550 2446
rect 5606 2390 5674 2446
rect 5730 2390 5798 2446
rect 5854 2390 5922 2446
rect 5978 2390 6046 2446
rect 6102 2390 6170 2446
rect 6226 2390 6294 2446
rect 6350 2390 6418 2446
rect 6474 2390 6542 2446
rect 6598 2390 6666 2446
rect 6722 2390 6790 2446
rect 6846 2390 6914 2446
rect 6970 2390 7038 2446
rect 7094 2390 7104 2446
rect 5168 2322 7104 2390
rect 5168 2266 5178 2322
rect 5234 2266 5302 2322
rect 5358 2266 5426 2322
rect 5482 2266 5550 2322
rect 5606 2266 5674 2322
rect 5730 2266 5798 2322
rect 5854 2266 5922 2322
rect 5978 2266 6046 2322
rect 6102 2266 6170 2322
rect 6226 2266 6294 2322
rect 6350 2266 6418 2322
rect 6474 2266 6542 2322
rect 6598 2266 6666 2322
rect 6722 2266 6790 2322
rect 6846 2266 6914 2322
rect 6970 2266 7038 2322
rect 7094 2266 7104 2322
rect 5168 2198 7104 2266
rect 5168 2142 5178 2198
rect 5234 2142 5302 2198
rect 5358 2142 5426 2198
rect 5482 2142 5550 2198
rect 5606 2142 5674 2198
rect 5730 2142 5798 2198
rect 5854 2142 5922 2198
rect 5978 2142 6046 2198
rect 6102 2142 6170 2198
rect 6226 2142 6294 2198
rect 6350 2142 6418 2198
rect 6474 2142 6542 2198
rect 6598 2142 6666 2198
rect 6722 2142 6790 2198
rect 6846 2142 6914 2198
rect 6970 2142 7038 2198
rect 7094 2142 7104 2198
rect 5168 2074 7104 2142
rect 5168 2018 5178 2074
rect 5234 2018 5302 2074
rect 5358 2018 5426 2074
rect 5482 2018 5550 2074
rect 5606 2018 5674 2074
rect 5730 2018 5798 2074
rect 5854 2018 5922 2074
rect 5978 2018 6046 2074
rect 6102 2018 6170 2074
rect 6226 2018 6294 2074
rect 6350 2018 6418 2074
rect 6474 2018 6542 2074
rect 6598 2018 6666 2074
rect 6722 2018 6790 2074
rect 6846 2018 6914 2074
rect 6970 2018 7038 2074
rect 7094 2018 7104 2074
rect 5168 1950 7104 2018
rect 5168 1894 5178 1950
rect 5234 1894 5302 1950
rect 5358 1894 5426 1950
rect 5482 1894 5550 1950
rect 5606 1894 5674 1950
rect 5730 1894 5798 1950
rect 5854 1894 5922 1950
rect 5978 1894 6046 1950
rect 6102 1894 6170 1950
rect 6226 1894 6294 1950
rect 6350 1894 6418 1950
rect 6474 1894 6542 1950
rect 6598 1894 6666 1950
rect 6722 1894 6790 1950
rect 6846 1894 6914 1950
rect 6970 1894 7038 1950
rect 7094 1894 7104 1950
rect 5168 1826 7104 1894
rect 5168 1770 5178 1826
rect 5234 1770 5302 1826
rect 5358 1770 5426 1826
rect 5482 1770 5550 1826
rect 5606 1770 5674 1826
rect 5730 1770 5798 1826
rect 5854 1770 5922 1826
rect 5978 1770 6046 1826
rect 6102 1770 6170 1826
rect 6226 1770 6294 1826
rect 6350 1770 6418 1826
rect 6474 1770 6542 1826
rect 6598 1770 6666 1826
rect 6722 1770 6790 1826
rect 6846 1770 6914 1826
rect 6970 1770 7038 1826
rect 7094 1770 7104 1826
rect 5168 1702 7104 1770
rect 5168 1646 5178 1702
rect 5234 1646 5302 1702
rect 5358 1646 5426 1702
rect 5482 1646 5550 1702
rect 5606 1646 5674 1702
rect 5730 1646 5798 1702
rect 5854 1646 5922 1702
rect 5978 1646 6046 1702
rect 6102 1646 6170 1702
rect 6226 1646 6294 1702
rect 6350 1646 6418 1702
rect 6474 1646 6542 1702
rect 6598 1646 6666 1702
rect 6722 1646 6790 1702
rect 6846 1646 6914 1702
rect 6970 1646 7038 1702
rect 7094 1646 7104 1702
rect 5168 1636 7104 1646
rect 7874 4554 9810 4564
rect 7874 4498 7884 4554
rect 7940 4498 8008 4554
rect 8064 4498 8132 4554
rect 8188 4498 8256 4554
rect 8312 4498 8380 4554
rect 8436 4498 8504 4554
rect 8560 4498 8628 4554
rect 8684 4498 8752 4554
rect 8808 4498 8876 4554
rect 8932 4498 9000 4554
rect 9056 4498 9124 4554
rect 9180 4498 9248 4554
rect 9304 4498 9372 4554
rect 9428 4498 9496 4554
rect 9552 4498 9620 4554
rect 9676 4498 9744 4554
rect 9800 4498 9810 4554
rect 7874 4430 9810 4498
rect 7874 4374 7884 4430
rect 7940 4374 8008 4430
rect 8064 4374 8132 4430
rect 8188 4374 8256 4430
rect 8312 4374 8380 4430
rect 8436 4374 8504 4430
rect 8560 4374 8628 4430
rect 8684 4374 8752 4430
rect 8808 4374 8876 4430
rect 8932 4374 9000 4430
rect 9056 4374 9124 4430
rect 9180 4374 9248 4430
rect 9304 4374 9372 4430
rect 9428 4374 9496 4430
rect 9552 4374 9620 4430
rect 9676 4374 9744 4430
rect 9800 4374 9810 4430
rect 7874 4306 9810 4374
rect 7874 4250 7884 4306
rect 7940 4250 8008 4306
rect 8064 4250 8132 4306
rect 8188 4250 8256 4306
rect 8312 4250 8380 4306
rect 8436 4250 8504 4306
rect 8560 4250 8628 4306
rect 8684 4250 8752 4306
rect 8808 4250 8876 4306
rect 8932 4250 9000 4306
rect 9056 4250 9124 4306
rect 9180 4250 9248 4306
rect 9304 4250 9372 4306
rect 9428 4250 9496 4306
rect 9552 4250 9620 4306
rect 9676 4250 9744 4306
rect 9800 4250 9810 4306
rect 7874 4182 9810 4250
rect 7874 4126 7884 4182
rect 7940 4126 8008 4182
rect 8064 4126 8132 4182
rect 8188 4126 8256 4182
rect 8312 4126 8380 4182
rect 8436 4126 8504 4182
rect 8560 4126 8628 4182
rect 8684 4126 8752 4182
rect 8808 4126 8876 4182
rect 8932 4126 9000 4182
rect 9056 4126 9124 4182
rect 9180 4126 9248 4182
rect 9304 4126 9372 4182
rect 9428 4126 9496 4182
rect 9552 4126 9620 4182
rect 9676 4126 9744 4182
rect 9800 4126 9810 4182
rect 7874 4058 9810 4126
rect 7874 4002 7884 4058
rect 7940 4002 8008 4058
rect 8064 4002 8132 4058
rect 8188 4002 8256 4058
rect 8312 4002 8380 4058
rect 8436 4002 8504 4058
rect 8560 4002 8628 4058
rect 8684 4002 8752 4058
rect 8808 4002 8876 4058
rect 8932 4002 9000 4058
rect 9056 4002 9124 4058
rect 9180 4002 9248 4058
rect 9304 4002 9372 4058
rect 9428 4002 9496 4058
rect 9552 4002 9620 4058
rect 9676 4002 9744 4058
rect 9800 4002 9810 4058
rect 7874 3934 9810 4002
rect 7874 3878 7884 3934
rect 7940 3878 8008 3934
rect 8064 3878 8132 3934
rect 8188 3878 8256 3934
rect 8312 3878 8380 3934
rect 8436 3878 8504 3934
rect 8560 3878 8628 3934
rect 8684 3878 8752 3934
rect 8808 3878 8876 3934
rect 8932 3878 9000 3934
rect 9056 3878 9124 3934
rect 9180 3878 9248 3934
rect 9304 3878 9372 3934
rect 9428 3878 9496 3934
rect 9552 3878 9620 3934
rect 9676 3878 9744 3934
rect 9800 3878 9810 3934
rect 7874 3810 9810 3878
rect 7874 3754 7884 3810
rect 7940 3754 8008 3810
rect 8064 3754 8132 3810
rect 8188 3754 8256 3810
rect 8312 3754 8380 3810
rect 8436 3754 8504 3810
rect 8560 3754 8628 3810
rect 8684 3754 8752 3810
rect 8808 3754 8876 3810
rect 8932 3754 9000 3810
rect 9056 3754 9124 3810
rect 9180 3754 9248 3810
rect 9304 3754 9372 3810
rect 9428 3754 9496 3810
rect 9552 3754 9620 3810
rect 9676 3754 9744 3810
rect 9800 3754 9810 3810
rect 7874 3686 9810 3754
rect 7874 3630 7884 3686
rect 7940 3630 8008 3686
rect 8064 3630 8132 3686
rect 8188 3630 8256 3686
rect 8312 3630 8380 3686
rect 8436 3630 8504 3686
rect 8560 3630 8628 3686
rect 8684 3630 8752 3686
rect 8808 3630 8876 3686
rect 8932 3630 9000 3686
rect 9056 3630 9124 3686
rect 9180 3630 9248 3686
rect 9304 3630 9372 3686
rect 9428 3630 9496 3686
rect 9552 3630 9620 3686
rect 9676 3630 9744 3686
rect 9800 3630 9810 3686
rect 7874 3562 9810 3630
rect 7874 3506 7884 3562
rect 7940 3506 8008 3562
rect 8064 3506 8132 3562
rect 8188 3506 8256 3562
rect 8312 3506 8380 3562
rect 8436 3506 8504 3562
rect 8560 3506 8628 3562
rect 8684 3506 8752 3562
rect 8808 3506 8876 3562
rect 8932 3506 9000 3562
rect 9056 3506 9124 3562
rect 9180 3506 9248 3562
rect 9304 3506 9372 3562
rect 9428 3506 9496 3562
rect 9552 3506 9620 3562
rect 9676 3506 9744 3562
rect 9800 3506 9810 3562
rect 7874 3438 9810 3506
rect 7874 3382 7884 3438
rect 7940 3382 8008 3438
rect 8064 3382 8132 3438
rect 8188 3382 8256 3438
rect 8312 3382 8380 3438
rect 8436 3382 8504 3438
rect 8560 3382 8628 3438
rect 8684 3382 8752 3438
rect 8808 3382 8876 3438
rect 8932 3382 9000 3438
rect 9056 3382 9124 3438
rect 9180 3382 9248 3438
rect 9304 3382 9372 3438
rect 9428 3382 9496 3438
rect 9552 3382 9620 3438
rect 9676 3382 9744 3438
rect 9800 3382 9810 3438
rect 7874 3314 9810 3382
rect 7874 3258 7884 3314
rect 7940 3258 8008 3314
rect 8064 3258 8132 3314
rect 8188 3258 8256 3314
rect 8312 3258 8380 3314
rect 8436 3258 8504 3314
rect 8560 3258 8628 3314
rect 8684 3258 8752 3314
rect 8808 3258 8876 3314
rect 8932 3258 9000 3314
rect 9056 3258 9124 3314
rect 9180 3258 9248 3314
rect 9304 3258 9372 3314
rect 9428 3258 9496 3314
rect 9552 3258 9620 3314
rect 9676 3258 9744 3314
rect 9800 3258 9810 3314
rect 7874 3190 9810 3258
rect 7874 3134 7884 3190
rect 7940 3134 8008 3190
rect 8064 3134 8132 3190
rect 8188 3134 8256 3190
rect 8312 3134 8380 3190
rect 8436 3134 8504 3190
rect 8560 3134 8628 3190
rect 8684 3134 8752 3190
rect 8808 3134 8876 3190
rect 8932 3134 9000 3190
rect 9056 3134 9124 3190
rect 9180 3134 9248 3190
rect 9304 3134 9372 3190
rect 9428 3134 9496 3190
rect 9552 3134 9620 3190
rect 9676 3134 9744 3190
rect 9800 3134 9810 3190
rect 7874 3066 9810 3134
rect 7874 3010 7884 3066
rect 7940 3010 8008 3066
rect 8064 3010 8132 3066
rect 8188 3010 8256 3066
rect 8312 3010 8380 3066
rect 8436 3010 8504 3066
rect 8560 3010 8628 3066
rect 8684 3010 8752 3066
rect 8808 3010 8876 3066
rect 8932 3010 9000 3066
rect 9056 3010 9124 3066
rect 9180 3010 9248 3066
rect 9304 3010 9372 3066
rect 9428 3010 9496 3066
rect 9552 3010 9620 3066
rect 9676 3010 9744 3066
rect 9800 3010 9810 3066
rect 7874 2942 9810 3010
rect 7874 2886 7884 2942
rect 7940 2886 8008 2942
rect 8064 2886 8132 2942
rect 8188 2886 8256 2942
rect 8312 2886 8380 2942
rect 8436 2886 8504 2942
rect 8560 2886 8628 2942
rect 8684 2886 8752 2942
rect 8808 2886 8876 2942
rect 8932 2886 9000 2942
rect 9056 2886 9124 2942
rect 9180 2886 9248 2942
rect 9304 2886 9372 2942
rect 9428 2886 9496 2942
rect 9552 2886 9620 2942
rect 9676 2886 9744 2942
rect 9800 2886 9810 2942
rect 7874 2818 9810 2886
rect 7874 2762 7884 2818
rect 7940 2762 8008 2818
rect 8064 2762 8132 2818
rect 8188 2762 8256 2818
rect 8312 2762 8380 2818
rect 8436 2762 8504 2818
rect 8560 2762 8628 2818
rect 8684 2762 8752 2818
rect 8808 2762 8876 2818
rect 8932 2762 9000 2818
rect 9056 2762 9124 2818
rect 9180 2762 9248 2818
rect 9304 2762 9372 2818
rect 9428 2762 9496 2818
rect 9552 2762 9620 2818
rect 9676 2762 9744 2818
rect 9800 2762 9810 2818
rect 7874 2694 9810 2762
rect 7874 2638 7884 2694
rect 7940 2638 8008 2694
rect 8064 2638 8132 2694
rect 8188 2638 8256 2694
rect 8312 2638 8380 2694
rect 8436 2638 8504 2694
rect 8560 2638 8628 2694
rect 8684 2638 8752 2694
rect 8808 2638 8876 2694
rect 8932 2638 9000 2694
rect 9056 2638 9124 2694
rect 9180 2638 9248 2694
rect 9304 2638 9372 2694
rect 9428 2638 9496 2694
rect 9552 2638 9620 2694
rect 9676 2638 9744 2694
rect 9800 2638 9810 2694
rect 7874 2570 9810 2638
rect 7874 2514 7884 2570
rect 7940 2514 8008 2570
rect 8064 2514 8132 2570
rect 8188 2514 8256 2570
rect 8312 2514 8380 2570
rect 8436 2514 8504 2570
rect 8560 2514 8628 2570
rect 8684 2514 8752 2570
rect 8808 2514 8876 2570
rect 8932 2514 9000 2570
rect 9056 2514 9124 2570
rect 9180 2514 9248 2570
rect 9304 2514 9372 2570
rect 9428 2514 9496 2570
rect 9552 2514 9620 2570
rect 9676 2514 9744 2570
rect 9800 2514 9810 2570
rect 7874 2446 9810 2514
rect 7874 2390 7884 2446
rect 7940 2390 8008 2446
rect 8064 2390 8132 2446
rect 8188 2390 8256 2446
rect 8312 2390 8380 2446
rect 8436 2390 8504 2446
rect 8560 2390 8628 2446
rect 8684 2390 8752 2446
rect 8808 2390 8876 2446
rect 8932 2390 9000 2446
rect 9056 2390 9124 2446
rect 9180 2390 9248 2446
rect 9304 2390 9372 2446
rect 9428 2390 9496 2446
rect 9552 2390 9620 2446
rect 9676 2390 9744 2446
rect 9800 2390 9810 2446
rect 7874 2322 9810 2390
rect 7874 2266 7884 2322
rect 7940 2266 8008 2322
rect 8064 2266 8132 2322
rect 8188 2266 8256 2322
rect 8312 2266 8380 2322
rect 8436 2266 8504 2322
rect 8560 2266 8628 2322
rect 8684 2266 8752 2322
rect 8808 2266 8876 2322
rect 8932 2266 9000 2322
rect 9056 2266 9124 2322
rect 9180 2266 9248 2322
rect 9304 2266 9372 2322
rect 9428 2266 9496 2322
rect 9552 2266 9620 2322
rect 9676 2266 9744 2322
rect 9800 2266 9810 2322
rect 7874 2198 9810 2266
rect 7874 2142 7884 2198
rect 7940 2142 8008 2198
rect 8064 2142 8132 2198
rect 8188 2142 8256 2198
rect 8312 2142 8380 2198
rect 8436 2142 8504 2198
rect 8560 2142 8628 2198
rect 8684 2142 8752 2198
rect 8808 2142 8876 2198
rect 8932 2142 9000 2198
rect 9056 2142 9124 2198
rect 9180 2142 9248 2198
rect 9304 2142 9372 2198
rect 9428 2142 9496 2198
rect 9552 2142 9620 2198
rect 9676 2142 9744 2198
rect 9800 2142 9810 2198
rect 7874 2074 9810 2142
rect 7874 2018 7884 2074
rect 7940 2018 8008 2074
rect 8064 2018 8132 2074
rect 8188 2018 8256 2074
rect 8312 2018 8380 2074
rect 8436 2018 8504 2074
rect 8560 2018 8628 2074
rect 8684 2018 8752 2074
rect 8808 2018 8876 2074
rect 8932 2018 9000 2074
rect 9056 2018 9124 2074
rect 9180 2018 9248 2074
rect 9304 2018 9372 2074
rect 9428 2018 9496 2074
rect 9552 2018 9620 2074
rect 9676 2018 9744 2074
rect 9800 2018 9810 2074
rect 7874 1950 9810 2018
rect 7874 1894 7884 1950
rect 7940 1894 8008 1950
rect 8064 1894 8132 1950
rect 8188 1894 8256 1950
rect 8312 1894 8380 1950
rect 8436 1894 8504 1950
rect 8560 1894 8628 1950
rect 8684 1894 8752 1950
rect 8808 1894 8876 1950
rect 8932 1894 9000 1950
rect 9056 1894 9124 1950
rect 9180 1894 9248 1950
rect 9304 1894 9372 1950
rect 9428 1894 9496 1950
rect 9552 1894 9620 1950
rect 9676 1894 9744 1950
rect 9800 1894 9810 1950
rect 7874 1826 9810 1894
rect 7874 1770 7884 1826
rect 7940 1770 8008 1826
rect 8064 1770 8132 1826
rect 8188 1770 8256 1826
rect 8312 1770 8380 1826
rect 8436 1770 8504 1826
rect 8560 1770 8628 1826
rect 8684 1770 8752 1826
rect 8808 1770 8876 1826
rect 8932 1770 9000 1826
rect 9056 1770 9124 1826
rect 9180 1770 9248 1826
rect 9304 1770 9372 1826
rect 9428 1770 9496 1826
rect 9552 1770 9620 1826
rect 9676 1770 9744 1826
rect 9800 1770 9810 1826
rect 7874 1702 9810 1770
rect 7874 1646 7884 1702
rect 7940 1646 8008 1702
rect 8064 1646 8132 1702
rect 8188 1646 8256 1702
rect 8312 1646 8380 1702
rect 8436 1646 8504 1702
rect 8560 1646 8628 1702
rect 8684 1646 8752 1702
rect 8808 1646 8876 1702
rect 8932 1646 9000 1702
rect 9056 1646 9124 1702
rect 9180 1646 9248 1702
rect 9304 1646 9372 1702
rect 9428 1646 9496 1702
rect 9552 1646 9620 1702
rect 9676 1646 9744 1702
rect 9800 1646 9810 1702
rect 7874 1636 9810 1646
rect 10244 4554 12180 4564
rect 10244 4498 10254 4554
rect 10310 4498 10378 4554
rect 10434 4498 10502 4554
rect 10558 4498 10626 4554
rect 10682 4498 10750 4554
rect 10806 4498 10874 4554
rect 10930 4498 10998 4554
rect 11054 4498 11122 4554
rect 11178 4498 11246 4554
rect 11302 4498 11370 4554
rect 11426 4498 11494 4554
rect 11550 4498 11618 4554
rect 11674 4498 11742 4554
rect 11798 4498 11866 4554
rect 11922 4498 11990 4554
rect 12046 4498 12114 4554
rect 12170 4498 12180 4554
rect 10244 4430 12180 4498
rect 10244 4374 10254 4430
rect 10310 4374 10378 4430
rect 10434 4374 10502 4430
rect 10558 4374 10626 4430
rect 10682 4374 10750 4430
rect 10806 4374 10874 4430
rect 10930 4374 10998 4430
rect 11054 4374 11122 4430
rect 11178 4374 11246 4430
rect 11302 4374 11370 4430
rect 11426 4374 11494 4430
rect 11550 4374 11618 4430
rect 11674 4374 11742 4430
rect 11798 4374 11866 4430
rect 11922 4374 11990 4430
rect 12046 4374 12114 4430
rect 12170 4374 12180 4430
rect 10244 4306 12180 4374
rect 10244 4250 10254 4306
rect 10310 4250 10378 4306
rect 10434 4250 10502 4306
rect 10558 4250 10626 4306
rect 10682 4250 10750 4306
rect 10806 4250 10874 4306
rect 10930 4250 10998 4306
rect 11054 4250 11122 4306
rect 11178 4250 11246 4306
rect 11302 4250 11370 4306
rect 11426 4250 11494 4306
rect 11550 4250 11618 4306
rect 11674 4250 11742 4306
rect 11798 4250 11866 4306
rect 11922 4250 11990 4306
rect 12046 4250 12114 4306
rect 12170 4250 12180 4306
rect 10244 4182 12180 4250
rect 10244 4126 10254 4182
rect 10310 4126 10378 4182
rect 10434 4126 10502 4182
rect 10558 4126 10626 4182
rect 10682 4126 10750 4182
rect 10806 4126 10874 4182
rect 10930 4126 10998 4182
rect 11054 4126 11122 4182
rect 11178 4126 11246 4182
rect 11302 4126 11370 4182
rect 11426 4126 11494 4182
rect 11550 4126 11618 4182
rect 11674 4126 11742 4182
rect 11798 4126 11866 4182
rect 11922 4126 11990 4182
rect 12046 4126 12114 4182
rect 12170 4126 12180 4182
rect 10244 4058 12180 4126
rect 10244 4002 10254 4058
rect 10310 4002 10378 4058
rect 10434 4002 10502 4058
rect 10558 4002 10626 4058
rect 10682 4002 10750 4058
rect 10806 4002 10874 4058
rect 10930 4002 10998 4058
rect 11054 4002 11122 4058
rect 11178 4002 11246 4058
rect 11302 4002 11370 4058
rect 11426 4002 11494 4058
rect 11550 4002 11618 4058
rect 11674 4002 11742 4058
rect 11798 4002 11866 4058
rect 11922 4002 11990 4058
rect 12046 4002 12114 4058
rect 12170 4002 12180 4058
rect 10244 3934 12180 4002
rect 10244 3878 10254 3934
rect 10310 3878 10378 3934
rect 10434 3878 10502 3934
rect 10558 3878 10626 3934
rect 10682 3878 10750 3934
rect 10806 3878 10874 3934
rect 10930 3878 10998 3934
rect 11054 3878 11122 3934
rect 11178 3878 11246 3934
rect 11302 3878 11370 3934
rect 11426 3878 11494 3934
rect 11550 3878 11618 3934
rect 11674 3878 11742 3934
rect 11798 3878 11866 3934
rect 11922 3878 11990 3934
rect 12046 3878 12114 3934
rect 12170 3878 12180 3934
rect 10244 3810 12180 3878
rect 10244 3754 10254 3810
rect 10310 3754 10378 3810
rect 10434 3754 10502 3810
rect 10558 3754 10626 3810
rect 10682 3754 10750 3810
rect 10806 3754 10874 3810
rect 10930 3754 10998 3810
rect 11054 3754 11122 3810
rect 11178 3754 11246 3810
rect 11302 3754 11370 3810
rect 11426 3754 11494 3810
rect 11550 3754 11618 3810
rect 11674 3754 11742 3810
rect 11798 3754 11866 3810
rect 11922 3754 11990 3810
rect 12046 3754 12114 3810
rect 12170 3754 12180 3810
rect 10244 3686 12180 3754
rect 10244 3630 10254 3686
rect 10310 3630 10378 3686
rect 10434 3630 10502 3686
rect 10558 3630 10626 3686
rect 10682 3630 10750 3686
rect 10806 3630 10874 3686
rect 10930 3630 10998 3686
rect 11054 3630 11122 3686
rect 11178 3630 11246 3686
rect 11302 3630 11370 3686
rect 11426 3630 11494 3686
rect 11550 3630 11618 3686
rect 11674 3630 11742 3686
rect 11798 3630 11866 3686
rect 11922 3630 11990 3686
rect 12046 3630 12114 3686
rect 12170 3630 12180 3686
rect 10244 3562 12180 3630
rect 10244 3506 10254 3562
rect 10310 3506 10378 3562
rect 10434 3506 10502 3562
rect 10558 3506 10626 3562
rect 10682 3506 10750 3562
rect 10806 3506 10874 3562
rect 10930 3506 10998 3562
rect 11054 3506 11122 3562
rect 11178 3506 11246 3562
rect 11302 3506 11370 3562
rect 11426 3506 11494 3562
rect 11550 3506 11618 3562
rect 11674 3506 11742 3562
rect 11798 3506 11866 3562
rect 11922 3506 11990 3562
rect 12046 3506 12114 3562
rect 12170 3506 12180 3562
rect 10244 3438 12180 3506
rect 10244 3382 10254 3438
rect 10310 3382 10378 3438
rect 10434 3382 10502 3438
rect 10558 3382 10626 3438
rect 10682 3382 10750 3438
rect 10806 3382 10874 3438
rect 10930 3382 10998 3438
rect 11054 3382 11122 3438
rect 11178 3382 11246 3438
rect 11302 3382 11370 3438
rect 11426 3382 11494 3438
rect 11550 3382 11618 3438
rect 11674 3382 11742 3438
rect 11798 3382 11866 3438
rect 11922 3382 11990 3438
rect 12046 3382 12114 3438
rect 12170 3382 12180 3438
rect 10244 3314 12180 3382
rect 10244 3258 10254 3314
rect 10310 3258 10378 3314
rect 10434 3258 10502 3314
rect 10558 3258 10626 3314
rect 10682 3258 10750 3314
rect 10806 3258 10874 3314
rect 10930 3258 10998 3314
rect 11054 3258 11122 3314
rect 11178 3258 11246 3314
rect 11302 3258 11370 3314
rect 11426 3258 11494 3314
rect 11550 3258 11618 3314
rect 11674 3258 11742 3314
rect 11798 3258 11866 3314
rect 11922 3258 11990 3314
rect 12046 3258 12114 3314
rect 12170 3258 12180 3314
rect 10244 3190 12180 3258
rect 10244 3134 10254 3190
rect 10310 3134 10378 3190
rect 10434 3134 10502 3190
rect 10558 3134 10626 3190
rect 10682 3134 10750 3190
rect 10806 3134 10874 3190
rect 10930 3134 10998 3190
rect 11054 3134 11122 3190
rect 11178 3134 11246 3190
rect 11302 3134 11370 3190
rect 11426 3134 11494 3190
rect 11550 3134 11618 3190
rect 11674 3134 11742 3190
rect 11798 3134 11866 3190
rect 11922 3134 11990 3190
rect 12046 3134 12114 3190
rect 12170 3134 12180 3190
rect 10244 3066 12180 3134
rect 10244 3010 10254 3066
rect 10310 3010 10378 3066
rect 10434 3010 10502 3066
rect 10558 3010 10626 3066
rect 10682 3010 10750 3066
rect 10806 3010 10874 3066
rect 10930 3010 10998 3066
rect 11054 3010 11122 3066
rect 11178 3010 11246 3066
rect 11302 3010 11370 3066
rect 11426 3010 11494 3066
rect 11550 3010 11618 3066
rect 11674 3010 11742 3066
rect 11798 3010 11866 3066
rect 11922 3010 11990 3066
rect 12046 3010 12114 3066
rect 12170 3010 12180 3066
rect 10244 2942 12180 3010
rect 10244 2886 10254 2942
rect 10310 2886 10378 2942
rect 10434 2886 10502 2942
rect 10558 2886 10626 2942
rect 10682 2886 10750 2942
rect 10806 2886 10874 2942
rect 10930 2886 10998 2942
rect 11054 2886 11122 2942
rect 11178 2886 11246 2942
rect 11302 2886 11370 2942
rect 11426 2886 11494 2942
rect 11550 2886 11618 2942
rect 11674 2886 11742 2942
rect 11798 2886 11866 2942
rect 11922 2886 11990 2942
rect 12046 2886 12114 2942
rect 12170 2886 12180 2942
rect 10244 2818 12180 2886
rect 10244 2762 10254 2818
rect 10310 2762 10378 2818
rect 10434 2762 10502 2818
rect 10558 2762 10626 2818
rect 10682 2762 10750 2818
rect 10806 2762 10874 2818
rect 10930 2762 10998 2818
rect 11054 2762 11122 2818
rect 11178 2762 11246 2818
rect 11302 2762 11370 2818
rect 11426 2762 11494 2818
rect 11550 2762 11618 2818
rect 11674 2762 11742 2818
rect 11798 2762 11866 2818
rect 11922 2762 11990 2818
rect 12046 2762 12114 2818
rect 12170 2762 12180 2818
rect 10244 2694 12180 2762
rect 10244 2638 10254 2694
rect 10310 2638 10378 2694
rect 10434 2638 10502 2694
rect 10558 2638 10626 2694
rect 10682 2638 10750 2694
rect 10806 2638 10874 2694
rect 10930 2638 10998 2694
rect 11054 2638 11122 2694
rect 11178 2638 11246 2694
rect 11302 2638 11370 2694
rect 11426 2638 11494 2694
rect 11550 2638 11618 2694
rect 11674 2638 11742 2694
rect 11798 2638 11866 2694
rect 11922 2638 11990 2694
rect 12046 2638 12114 2694
rect 12170 2638 12180 2694
rect 10244 2570 12180 2638
rect 10244 2514 10254 2570
rect 10310 2514 10378 2570
rect 10434 2514 10502 2570
rect 10558 2514 10626 2570
rect 10682 2514 10750 2570
rect 10806 2514 10874 2570
rect 10930 2514 10998 2570
rect 11054 2514 11122 2570
rect 11178 2514 11246 2570
rect 11302 2514 11370 2570
rect 11426 2514 11494 2570
rect 11550 2514 11618 2570
rect 11674 2514 11742 2570
rect 11798 2514 11866 2570
rect 11922 2514 11990 2570
rect 12046 2514 12114 2570
rect 12170 2514 12180 2570
rect 10244 2446 12180 2514
rect 10244 2390 10254 2446
rect 10310 2390 10378 2446
rect 10434 2390 10502 2446
rect 10558 2390 10626 2446
rect 10682 2390 10750 2446
rect 10806 2390 10874 2446
rect 10930 2390 10998 2446
rect 11054 2390 11122 2446
rect 11178 2390 11246 2446
rect 11302 2390 11370 2446
rect 11426 2390 11494 2446
rect 11550 2390 11618 2446
rect 11674 2390 11742 2446
rect 11798 2390 11866 2446
rect 11922 2390 11990 2446
rect 12046 2390 12114 2446
rect 12170 2390 12180 2446
rect 10244 2322 12180 2390
rect 10244 2266 10254 2322
rect 10310 2266 10378 2322
rect 10434 2266 10502 2322
rect 10558 2266 10626 2322
rect 10682 2266 10750 2322
rect 10806 2266 10874 2322
rect 10930 2266 10998 2322
rect 11054 2266 11122 2322
rect 11178 2266 11246 2322
rect 11302 2266 11370 2322
rect 11426 2266 11494 2322
rect 11550 2266 11618 2322
rect 11674 2266 11742 2322
rect 11798 2266 11866 2322
rect 11922 2266 11990 2322
rect 12046 2266 12114 2322
rect 12170 2266 12180 2322
rect 10244 2198 12180 2266
rect 10244 2142 10254 2198
rect 10310 2142 10378 2198
rect 10434 2142 10502 2198
rect 10558 2142 10626 2198
rect 10682 2142 10750 2198
rect 10806 2142 10874 2198
rect 10930 2142 10998 2198
rect 11054 2142 11122 2198
rect 11178 2142 11246 2198
rect 11302 2142 11370 2198
rect 11426 2142 11494 2198
rect 11550 2142 11618 2198
rect 11674 2142 11742 2198
rect 11798 2142 11866 2198
rect 11922 2142 11990 2198
rect 12046 2142 12114 2198
rect 12170 2142 12180 2198
rect 10244 2074 12180 2142
rect 10244 2018 10254 2074
rect 10310 2018 10378 2074
rect 10434 2018 10502 2074
rect 10558 2018 10626 2074
rect 10682 2018 10750 2074
rect 10806 2018 10874 2074
rect 10930 2018 10998 2074
rect 11054 2018 11122 2074
rect 11178 2018 11246 2074
rect 11302 2018 11370 2074
rect 11426 2018 11494 2074
rect 11550 2018 11618 2074
rect 11674 2018 11742 2074
rect 11798 2018 11866 2074
rect 11922 2018 11990 2074
rect 12046 2018 12114 2074
rect 12170 2018 12180 2074
rect 10244 1950 12180 2018
rect 10244 1894 10254 1950
rect 10310 1894 10378 1950
rect 10434 1894 10502 1950
rect 10558 1894 10626 1950
rect 10682 1894 10750 1950
rect 10806 1894 10874 1950
rect 10930 1894 10998 1950
rect 11054 1894 11122 1950
rect 11178 1894 11246 1950
rect 11302 1894 11370 1950
rect 11426 1894 11494 1950
rect 11550 1894 11618 1950
rect 11674 1894 11742 1950
rect 11798 1894 11866 1950
rect 11922 1894 11990 1950
rect 12046 1894 12114 1950
rect 12170 1894 12180 1950
rect 10244 1826 12180 1894
rect 10244 1770 10254 1826
rect 10310 1770 10378 1826
rect 10434 1770 10502 1826
rect 10558 1770 10626 1826
rect 10682 1770 10750 1826
rect 10806 1770 10874 1826
rect 10930 1770 10998 1826
rect 11054 1770 11122 1826
rect 11178 1770 11246 1826
rect 11302 1770 11370 1826
rect 11426 1770 11494 1826
rect 11550 1770 11618 1826
rect 11674 1770 11742 1826
rect 11798 1770 11866 1826
rect 11922 1770 11990 1826
rect 12046 1770 12114 1826
rect 12170 1770 12180 1826
rect 10244 1702 12180 1770
rect 10244 1646 10254 1702
rect 10310 1646 10378 1702
rect 10434 1646 10502 1702
rect 10558 1646 10626 1702
rect 10682 1646 10750 1702
rect 10806 1646 10874 1702
rect 10930 1646 10998 1702
rect 11054 1646 11122 1702
rect 11178 1646 11246 1702
rect 11302 1646 11370 1702
rect 11426 1646 11494 1702
rect 11550 1646 11618 1702
rect 11674 1646 11742 1702
rect 11798 1646 11866 1702
rect 11922 1646 11990 1702
rect 12046 1646 12114 1702
rect 12170 1646 12180 1702
rect 10244 1636 12180 1646
rect 12861 4554 14673 4564
rect 12861 4498 12871 4554
rect 12927 4498 12995 4554
rect 13051 4498 13119 4554
rect 13175 4498 13243 4554
rect 13299 4498 13367 4554
rect 13423 4498 13491 4554
rect 13547 4498 13615 4554
rect 13671 4498 13739 4554
rect 13795 4498 13863 4554
rect 13919 4498 13987 4554
rect 14043 4498 14111 4554
rect 14167 4498 14235 4554
rect 14291 4498 14359 4554
rect 14415 4498 14483 4554
rect 14539 4498 14607 4554
rect 14663 4498 14673 4554
rect 12861 4430 14673 4498
rect 12861 4374 12871 4430
rect 12927 4374 12995 4430
rect 13051 4374 13119 4430
rect 13175 4374 13243 4430
rect 13299 4374 13367 4430
rect 13423 4374 13491 4430
rect 13547 4374 13615 4430
rect 13671 4374 13739 4430
rect 13795 4374 13863 4430
rect 13919 4374 13987 4430
rect 14043 4374 14111 4430
rect 14167 4374 14235 4430
rect 14291 4374 14359 4430
rect 14415 4374 14483 4430
rect 14539 4374 14607 4430
rect 14663 4374 14673 4430
rect 12861 4306 14673 4374
rect 12861 4250 12871 4306
rect 12927 4250 12995 4306
rect 13051 4250 13119 4306
rect 13175 4250 13243 4306
rect 13299 4250 13367 4306
rect 13423 4250 13491 4306
rect 13547 4250 13615 4306
rect 13671 4250 13739 4306
rect 13795 4250 13863 4306
rect 13919 4250 13987 4306
rect 14043 4250 14111 4306
rect 14167 4250 14235 4306
rect 14291 4250 14359 4306
rect 14415 4250 14483 4306
rect 14539 4250 14607 4306
rect 14663 4250 14673 4306
rect 12861 4182 14673 4250
rect 12861 4126 12871 4182
rect 12927 4126 12995 4182
rect 13051 4126 13119 4182
rect 13175 4126 13243 4182
rect 13299 4126 13367 4182
rect 13423 4126 13491 4182
rect 13547 4126 13615 4182
rect 13671 4126 13739 4182
rect 13795 4126 13863 4182
rect 13919 4126 13987 4182
rect 14043 4126 14111 4182
rect 14167 4126 14235 4182
rect 14291 4126 14359 4182
rect 14415 4126 14483 4182
rect 14539 4126 14607 4182
rect 14663 4126 14673 4182
rect 12861 4058 14673 4126
rect 12861 4002 12871 4058
rect 12927 4002 12995 4058
rect 13051 4002 13119 4058
rect 13175 4002 13243 4058
rect 13299 4002 13367 4058
rect 13423 4002 13491 4058
rect 13547 4002 13615 4058
rect 13671 4002 13739 4058
rect 13795 4002 13863 4058
rect 13919 4002 13987 4058
rect 14043 4002 14111 4058
rect 14167 4002 14235 4058
rect 14291 4002 14359 4058
rect 14415 4002 14483 4058
rect 14539 4002 14607 4058
rect 14663 4002 14673 4058
rect 12861 3934 14673 4002
rect 12861 3878 12871 3934
rect 12927 3878 12995 3934
rect 13051 3878 13119 3934
rect 13175 3878 13243 3934
rect 13299 3878 13367 3934
rect 13423 3878 13491 3934
rect 13547 3878 13615 3934
rect 13671 3878 13739 3934
rect 13795 3878 13863 3934
rect 13919 3878 13987 3934
rect 14043 3878 14111 3934
rect 14167 3878 14235 3934
rect 14291 3878 14359 3934
rect 14415 3878 14483 3934
rect 14539 3878 14607 3934
rect 14663 3878 14673 3934
rect 12861 3810 14673 3878
rect 12861 3754 12871 3810
rect 12927 3754 12995 3810
rect 13051 3754 13119 3810
rect 13175 3754 13243 3810
rect 13299 3754 13367 3810
rect 13423 3754 13491 3810
rect 13547 3754 13615 3810
rect 13671 3754 13739 3810
rect 13795 3754 13863 3810
rect 13919 3754 13987 3810
rect 14043 3754 14111 3810
rect 14167 3754 14235 3810
rect 14291 3754 14359 3810
rect 14415 3754 14483 3810
rect 14539 3754 14607 3810
rect 14663 3754 14673 3810
rect 12861 3686 14673 3754
rect 12861 3630 12871 3686
rect 12927 3630 12995 3686
rect 13051 3630 13119 3686
rect 13175 3630 13243 3686
rect 13299 3630 13367 3686
rect 13423 3630 13491 3686
rect 13547 3630 13615 3686
rect 13671 3630 13739 3686
rect 13795 3630 13863 3686
rect 13919 3630 13987 3686
rect 14043 3630 14111 3686
rect 14167 3630 14235 3686
rect 14291 3630 14359 3686
rect 14415 3630 14483 3686
rect 14539 3630 14607 3686
rect 14663 3630 14673 3686
rect 12861 3562 14673 3630
rect 12861 3506 12871 3562
rect 12927 3506 12995 3562
rect 13051 3506 13119 3562
rect 13175 3506 13243 3562
rect 13299 3506 13367 3562
rect 13423 3506 13491 3562
rect 13547 3506 13615 3562
rect 13671 3506 13739 3562
rect 13795 3506 13863 3562
rect 13919 3506 13987 3562
rect 14043 3506 14111 3562
rect 14167 3506 14235 3562
rect 14291 3506 14359 3562
rect 14415 3506 14483 3562
rect 14539 3506 14607 3562
rect 14663 3506 14673 3562
rect 12861 3438 14673 3506
rect 12861 3382 12871 3438
rect 12927 3382 12995 3438
rect 13051 3382 13119 3438
rect 13175 3382 13243 3438
rect 13299 3382 13367 3438
rect 13423 3382 13491 3438
rect 13547 3382 13615 3438
rect 13671 3382 13739 3438
rect 13795 3382 13863 3438
rect 13919 3382 13987 3438
rect 14043 3382 14111 3438
rect 14167 3382 14235 3438
rect 14291 3382 14359 3438
rect 14415 3382 14483 3438
rect 14539 3382 14607 3438
rect 14663 3382 14673 3438
rect 12861 3314 14673 3382
rect 12861 3258 12871 3314
rect 12927 3258 12995 3314
rect 13051 3258 13119 3314
rect 13175 3258 13243 3314
rect 13299 3258 13367 3314
rect 13423 3258 13491 3314
rect 13547 3258 13615 3314
rect 13671 3258 13739 3314
rect 13795 3258 13863 3314
rect 13919 3258 13987 3314
rect 14043 3258 14111 3314
rect 14167 3258 14235 3314
rect 14291 3258 14359 3314
rect 14415 3258 14483 3314
rect 14539 3258 14607 3314
rect 14663 3258 14673 3314
rect 12861 3190 14673 3258
rect 12861 3134 12871 3190
rect 12927 3134 12995 3190
rect 13051 3134 13119 3190
rect 13175 3134 13243 3190
rect 13299 3134 13367 3190
rect 13423 3134 13491 3190
rect 13547 3134 13615 3190
rect 13671 3134 13739 3190
rect 13795 3134 13863 3190
rect 13919 3134 13987 3190
rect 14043 3134 14111 3190
rect 14167 3134 14235 3190
rect 14291 3134 14359 3190
rect 14415 3134 14483 3190
rect 14539 3134 14607 3190
rect 14663 3134 14673 3190
rect 12861 3066 14673 3134
rect 12861 3010 12871 3066
rect 12927 3010 12995 3066
rect 13051 3010 13119 3066
rect 13175 3010 13243 3066
rect 13299 3010 13367 3066
rect 13423 3010 13491 3066
rect 13547 3010 13615 3066
rect 13671 3010 13739 3066
rect 13795 3010 13863 3066
rect 13919 3010 13987 3066
rect 14043 3010 14111 3066
rect 14167 3010 14235 3066
rect 14291 3010 14359 3066
rect 14415 3010 14483 3066
rect 14539 3010 14607 3066
rect 14663 3010 14673 3066
rect 12861 2942 14673 3010
rect 12861 2886 12871 2942
rect 12927 2886 12995 2942
rect 13051 2886 13119 2942
rect 13175 2886 13243 2942
rect 13299 2886 13367 2942
rect 13423 2886 13491 2942
rect 13547 2886 13615 2942
rect 13671 2886 13739 2942
rect 13795 2886 13863 2942
rect 13919 2886 13987 2942
rect 14043 2886 14111 2942
rect 14167 2886 14235 2942
rect 14291 2886 14359 2942
rect 14415 2886 14483 2942
rect 14539 2886 14607 2942
rect 14663 2886 14673 2942
rect 12861 2818 14673 2886
rect 12861 2762 12871 2818
rect 12927 2762 12995 2818
rect 13051 2762 13119 2818
rect 13175 2762 13243 2818
rect 13299 2762 13367 2818
rect 13423 2762 13491 2818
rect 13547 2762 13615 2818
rect 13671 2762 13739 2818
rect 13795 2762 13863 2818
rect 13919 2762 13987 2818
rect 14043 2762 14111 2818
rect 14167 2762 14235 2818
rect 14291 2762 14359 2818
rect 14415 2762 14483 2818
rect 14539 2762 14607 2818
rect 14663 2762 14673 2818
rect 12861 2694 14673 2762
rect 12861 2638 12871 2694
rect 12927 2638 12995 2694
rect 13051 2638 13119 2694
rect 13175 2638 13243 2694
rect 13299 2638 13367 2694
rect 13423 2638 13491 2694
rect 13547 2638 13615 2694
rect 13671 2638 13739 2694
rect 13795 2638 13863 2694
rect 13919 2638 13987 2694
rect 14043 2638 14111 2694
rect 14167 2638 14235 2694
rect 14291 2638 14359 2694
rect 14415 2638 14483 2694
rect 14539 2638 14607 2694
rect 14663 2638 14673 2694
rect 12861 2570 14673 2638
rect 12861 2514 12871 2570
rect 12927 2514 12995 2570
rect 13051 2514 13119 2570
rect 13175 2514 13243 2570
rect 13299 2514 13367 2570
rect 13423 2514 13491 2570
rect 13547 2514 13615 2570
rect 13671 2514 13739 2570
rect 13795 2514 13863 2570
rect 13919 2514 13987 2570
rect 14043 2514 14111 2570
rect 14167 2514 14235 2570
rect 14291 2514 14359 2570
rect 14415 2514 14483 2570
rect 14539 2514 14607 2570
rect 14663 2514 14673 2570
rect 12861 2446 14673 2514
rect 12861 2390 12871 2446
rect 12927 2390 12995 2446
rect 13051 2390 13119 2446
rect 13175 2390 13243 2446
rect 13299 2390 13367 2446
rect 13423 2390 13491 2446
rect 13547 2390 13615 2446
rect 13671 2390 13739 2446
rect 13795 2390 13863 2446
rect 13919 2390 13987 2446
rect 14043 2390 14111 2446
rect 14167 2390 14235 2446
rect 14291 2390 14359 2446
rect 14415 2390 14483 2446
rect 14539 2390 14607 2446
rect 14663 2390 14673 2446
rect 12861 2322 14673 2390
rect 12861 2266 12871 2322
rect 12927 2266 12995 2322
rect 13051 2266 13119 2322
rect 13175 2266 13243 2322
rect 13299 2266 13367 2322
rect 13423 2266 13491 2322
rect 13547 2266 13615 2322
rect 13671 2266 13739 2322
rect 13795 2266 13863 2322
rect 13919 2266 13987 2322
rect 14043 2266 14111 2322
rect 14167 2266 14235 2322
rect 14291 2266 14359 2322
rect 14415 2266 14483 2322
rect 14539 2266 14607 2322
rect 14663 2266 14673 2322
rect 12861 2198 14673 2266
rect 12861 2142 12871 2198
rect 12927 2142 12995 2198
rect 13051 2142 13119 2198
rect 13175 2142 13243 2198
rect 13299 2142 13367 2198
rect 13423 2142 13491 2198
rect 13547 2142 13615 2198
rect 13671 2142 13739 2198
rect 13795 2142 13863 2198
rect 13919 2142 13987 2198
rect 14043 2142 14111 2198
rect 14167 2142 14235 2198
rect 14291 2142 14359 2198
rect 14415 2142 14483 2198
rect 14539 2142 14607 2198
rect 14663 2142 14673 2198
rect 12861 2074 14673 2142
rect 12861 2018 12871 2074
rect 12927 2018 12995 2074
rect 13051 2018 13119 2074
rect 13175 2018 13243 2074
rect 13299 2018 13367 2074
rect 13423 2018 13491 2074
rect 13547 2018 13615 2074
rect 13671 2018 13739 2074
rect 13795 2018 13863 2074
rect 13919 2018 13987 2074
rect 14043 2018 14111 2074
rect 14167 2018 14235 2074
rect 14291 2018 14359 2074
rect 14415 2018 14483 2074
rect 14539 2018 14607 2074
rect 14663 2018 14673 2074
rect 12861 1950 14673 2018
rect 12861 1894 12871 1950
rect 12927 1894 12995 1950
rect 13051 1894 13119 1950
rect 13175 1894 13243 1950
rect 13299 1894 13367 1950
rect 13423 1894 13491 1950
rect 13547 1894 13615 1950
rect 13671 1894 13739 1950
rect 13795 1894 13863 1950
rect 13919 1894 13987 1950
rect 14043 1894 14111 1950
rect 14167 1894 14235 1950
rect 14291 1894 14359 1950
rect 14415 1894 14483 1950
rect 14539 1894 14607 1950
rect 14663 1894 14673 1950
rect 12861 1826 14673 1894
rect 12861 1770 12871 1826
rect 12927 1770 12995 1826
rect 13051 1770 13119 1826
rect 13175 1770 13243 1826
rect 13299 1770 13367 1826
rect 13423 1770 13491 1826
rect 13547 1770 13615 1826
rect 13671 1770 13739 1826
rect 13795 1770 13863 1826
rect 13919 1770 13987 1826
rect 14043 1770 14111 1826
rect 14167 1770 14235 1826
rect 14291 1770 14359 1826
rect 14415 1770 14483 1826
rect 14539 1770 14607 1826
rect 14663 1770 14673 1826
rect 12861 1702 14673 1770
rect 12861 1646 12871 1702
rect 12927 1646 12995 1702
rect 13051 1646 13119 1702
rect 13175 1646 13243 1702
rect 13299 1646 13367 1702
rect 13423 1646 13491 1702
rect 13547 1646 13615 1702
rect 13671 1646 13739 1702
rect 13795 1646 13863 1702
rect 13919 1646 13987 1702
rect 14043 1646 14111 1702
rect 14167 1646 14235 1702
rect 14291 1646 14359 1702
rect 14415 1646 14483 1702
rect 14539 1646 14607 1702
rect 14663 1646 14673 1702
rect 12861 1636 14673 1646
rect -11 1604 86 1614
rect 14892 1614 14902 4586
rect 14958 1614 14989 4586
rect 14892 1604 14989 1614
rect 261 818 2161 1190
rect 261 766 321 818
rect 373 766 429 818
rect 481 766 537 818
rect 589 766 645 818
rect 697 766 753 818
rect 805 766 861 818
rect 913 766 969 818
rect 1021 766 1077 818
rect 1129 766 1185 818
rect 1237 766 1293 818
rect 1345 766 1401 818
rect 1453 766 1509 818
rect 1561 766 1617 818
rect 1669 766 1725 818
rect 1777 766 1833 818
rect 1885 766 1941 818
rect 1993 766 2049 818
rect 2101 766 2161 818
rect 261 0 2161 766
rect 2741 818 4791 1190
rect 2741 766 2876 818
rect 2928 766 2984 818
rect 3036 766 3092 818
rect 3144 766 3200 818
rect 3252 766 3308 818
rect 3360 766 3416 818
rect 3468 766 3524 818
rect 3576 766 3632 818
rect 3684 766 3740 818
rect 3792 766 3848 818
rect 3900 766 3956 818
rect 4008 766 4064 818
rect 4116 766 4172 818
rect 4224 766 4280 818
rect 4332 766 4388 818
rect 4440 766 4496 818
rect 4548 766 4604 818
rect 4656 766 4791 818
rect 2741 0 4791 766
rect 5111 818 7161 1190
rect 5111 766 5246 818
rect 5298 766 5354 818
rect 5406 766 5462 818
rect 5514 766 5570 818
rect 5622 766 5678 818
rect 5730 766 5786 818
rect 5838 766 5894 818
rect 5946 766 6002 818
rect 6054 766 6110 818
rect 6162 766 6218 818
rect 6270 766 6326 818
rect 6378 766 6434 818
rect 6486 766 6542 818
rect 6594 766 6650 818
rect 6702 766 6758 818
rect 6810 766 6866 818
rect 6918 766 6974 818
rect 7026 766 7161 818
rect 5111 0 7161 766
rect 7817 818 9867 1190
rect 7817 766 7952 818
rect 8004 766 8060 818
rect 8112 766 8168 818
rect 8220 766 8276 818
rect 8328 766 8384 818
rect 8436 766 8492 818
rect 8544 766 8600 818
rect 8652 766 8708 818
rect 8760 766 8816 818
rect 8868 766 8924 818
rect 8976 766 9032 818
rect 9084 766 9140 818
rect 9192 766 9248 818
rect 9300 766 9356 818
rect 9408 766 9464 818
rect 9516 766 9572 818
rect 9624 766 9680 818
rect 9732 766 9867 818
rect 7817 0 9867 766
rect 10187 818 12237 1190
rect 10187 766 10322 818
rect 10374 766 10430 818
rect 10482 766 10538 818
rect 10590 766 10646 818
rect 10698 766 10754 818
rect 10806 766 10862 818
rect 10914 766 10970 818
rect 11022 766 11078 818
rect 11130 766 11186 818
rect 11238 766 11294 818
rect 11346 766 11402 818
rect 11454 766 11510 818
rect 11562 766 11618 818
rect 11670 766 11726 818
rect 11778 766 11834 818
rect 11886 766 11942 818
rect 11994 766 12050 818
rect 12102 766 12237 818
rect 10187 0 12237 766
rect 12817 818 14717 1190
rect 12817 766 12877 818
rect 12929 766 12985 818
rect 13037 766 13093 818
rect 13145 766 13201 818
rect 13253 766 13309 818
rect 13361 766 13417 818
rect 13469 766 13525 818
rect 13577 766 13633 818
rect 13685 766 13741 818
rect 13793 766 13849 818
rect 13901 766 13957 818
rect 14009 766 14065 818
rect 14117 766 14173 818
rect 14225 766 14281 818
rect 14333 766 14389 818
rect 14441 766 14497 818
rect 14549 766 14605 818
rect 14657 766 14717 818
rect 12817 0 14717 766
<< via2 >>
rect 20 57259 76 57261
rect 20 57207 22 57259
rect 22 57207 74 57259
rect 74 57207 76 57259
rect 20 57151 76 57207
rect 20 57099 22 57151
rect 22 57099 74 57151
rect 74 57099 76 57151
rect 20 57043 76 57099
rect 20 56991 22 57043
rect 22 56991 74 57043
rect 74 56991 76 57043
rect 20 56935 76 56991
rect 20 56883 22 56935
rect 22 56883 74 56935
rect 74 56883 76 56935
rect 20 56827 76 56883
rect 20 56775 22 56827
rect 22 56775 74 56827
rect 74 56775 76 56827
rect 20 56719 76 56775
rect 20 56667 22 56719
rect 22 56667 74 56719
rect 74 56667 76 56719
rect 20 56611 76 56667
rect 20 56559 22 56611
rect 22 56559 74 56611
rect 74 56559 76 56611
rect 20 56503 76 56559
rect 20 56451 22 56503
rect 22 56451 74 56503
rect 74 56451 76 56503
rect 20 56395 76 56451
rect 20 56343 22 56395
rect 22 56343 74 56395
rect 74 56343 76 56395
rect 20 56287 76 56343
rect 20 56235 22 56287
rect 22 56235 74 56287
rect 74 56235 76 56287
rect 20 56179 76 56235
rect 20 56127 22 56179
rect 22 56127 74 56179
rect 74 56127 76 56179
rect 20 56071 76 56127
rect 20 56019 22 56071
rect 22 56019 74 56071
rect 74 56019 76 56071
rect 20 56017 76 56019
rect 315 57169 371 57225
rect 439 57169 495 57225
rect 563 57169 619 57225
rect 687 57169 743 57225
rect 811 57169 867 57225
rect 935 57169 991 57225
rect 1059 57169 1115 57225
rect 1183 57169 1239 57225
rect 1307 57169 1363 57225
rect 1431 57169 1487 57225
rect 1555 57169 1611 57225
rect 1679 57169 1735 57225
rect 1803 57169 1859 57225
rect 1927 57169 1983 57225
rect 2051 57169 2107 57225
rect 315 57045 371 57101
rect 439 57052 483 57101
rect 483 57052 495 57101
rect 563 57052 591 57101
rect 591 57052 619 57101
rect 687 57052 699 57101
rect 699 57052 743 57101
rect 811 57052 859 57101
rect 859 57052 867 57101
rect 935 57052 967 57101
rect 967 57052 991 57101
rect 1059 57052 1075 57101
rect 1075 57052 1115 57101
rect 439 57045 495 57052
rect 563 57045 619 57052
rect 687 57045 743 57052
rect 811 57045 867 57052
rect 935 57045 991 57052
rect 1059 57045 1115 57052
rect 1183 57045 1239 57101
rect 1307 57052 1347 57101
rect 1347 57052 1363 57101
rect 1431 57052 1455 57101
rect 1455 57052 1487 57101
rect 1555 57052 1563 57101
rect 1563 57052 1611 57101
rect 1679 57052 1723 57101
rect 1723 57052 1735 57101
rect 1803 57052 1831 57101
rect 1831 57052 1859 57101
rect 1927 57052 1939 57101
rect 1939 57052 1983 57101
rect 1307 57045 1363 57052
rect 1431 57045 1487 57052
rect 1555 57045 1611 57052
rect 1679 57045 1735 57052
rect 1803 57045 1859 57052
rect 1927 57045 1983 57052
rect 2051 57045 2107 57101
rect 315 56921 371 56977
rect 439 56921 495 56977
rect 563 56921 619 56977
rect 687 56921 743 56977
rect 811 56921 867 56977
rect 935 56921 991 56977
rect 1059 56921 1115 56977
rect 1183 56921 1239 56977
rect 1307 56921 1363 56977
rect 1431 56921 1487 56977
rect 1555 56921 1611 56977
rect 1679 56921 1735 56977
rect 1803 56921 1859 56977
rect 1927 56921 1983 56977
rect 2051 56921 2107 56977
rect 315 56797 371 56853
rect 439 56797 495 56853
rect 563 56797 619 56853
rect 687 56797 743 56853
rect 811 56797 867 56853
rect 935 56797 991 56853
rect 1059 56797 1115 56853
rect 1183 56797 1239 56853
rect 1307 56797 1363 56853
rect 1431 56797 1487 56853
rect 1555 56797 1611 56853
rect 1679 56797 1735 56853
rect 1803 56797 1859 56853
rect 1927 56797 1983 56853
rect 2051 56797 2107 56853
rect 315 56673 371 56729
rect 439 56673 495 56729
rect 563 56673 619 56729
rect 687 56673 743 56729
rect 811 56673 867 56729
rect 935 56673 991 56729
rect 1059 56673 1115 56729
rect 1183 56673 1239 56729
rect 1307 56673 1363 56729
rect 1431 56673 1487 56729
rect 1555 56673 1611 56729
rect 1679 56673 1735 56729
rect 1803 56673 1859 56729
rect 1927 56673 1983 56729
rect 2051 56673 2107 56729
rect 315 56591 369 56605
rect 369 56591 371 56605
rect 439 56591 493 56605
rect 493 56591 495 56605
rect 563 56591 617 56605
rect 617 56591 619 56605
rect 687 56591 741 56605
rect 741 56591 743 56605
rect 315 56549 371 56591
rect 439 56549 495 56591
rect 563 56549 619 56591
rect 687 56549 743 56591
rect 811 56549 867 56605
rect 935 56549 991 56605
rect 1059 56549 1115 56605
rect 1183 56549 1239 56605
rect 1307 56549 1363 56605
rect 1431 56549 1487 56605
rect 1555 56549 1611 56605
rect 1679 56549 1735 56605
rect 1803 56549 1859 56605
rect 1927 56549 1983 56605
rect 2051 56549 2107 56605
rect 315 56467 369 56481
rect 369 56467 371 56481
rect 439 56467 493 56481
rect 493 56467 495 56481
rect 563 56467 617 56481
rect 617 56467 619 56481
rect 687 56467 741 56481
rect 741 56467 743 56481
rect 315 56425 371 56467
rect 439 56425 495 56467
rect 563 56425 619 56467
rect 687 56425 743 56467
rect 811 56425 867 56481
rect 935 56425 991 56481
rect 1059 56425 1115 56481
rect 1183 56425 1239 56481
rect 1307 56425 1363 56481
rect 1431 56425 1487 56481
rect 1555 56425 1611 56481
rect 1679 56425 1735 56481
rect 1803 56425 1859 56481
rect 1927 56425 1983 56481
rect 2051 56425 2107 56481
rect 315 56343 369 56357
rect 369 56343 371 56357
rect 439 56343 493 56357
rect 493 56343 495 56357
rect 563 56343 617 56357
rect 617 56343 619 56357
rect 687 56343 741 56357
rect 741 56343 743 56357
rect 315 56301 371 56343
rect 439 56301 495 56343
rect 563 56301 619 56343
rect 687 56301 743 56343
rect 811 56301 867 56357
rect 935 56301 991 56357
rect 1059 56301 1115 56357
rect 1183 56301 1239 56357
rect 1307 56301 1363 56357
rect 1431 56301 1487 56357
rect 1555 56301 1611 56357
rect 1679 56301 1735 56357
rect 1803 56301 1859 56357
rect 1927 56301 1983 56357
rect 2051 56301 2107 56357
rect 315 56219 369 56233
rect 369 56219 371 56233
rect 439 56219 493 56233
rect 493 56219 495 56233
rect 563 56219 617 56233
rect 617 56219 619 56233
rect 687 56219 741 56233
rect 741 56219 743 56233
rect 315 56177 371 56219
rect 439 56177 495 56219
rect 563 56177 619 56219
rect 687 56177 743 56219
rect 811 56177 867 56233
rect 935 56177 991 56233
rect 1059 56177 1115 56233
rect 1183 56177 1239 56233
rect 1307 56177 1363 56233
rect 1431 56177 1487 56233
rect 1555 56177 1611 56233
rect 1679 56177 1735 56233
rect 1803 56177 1859 56233
rect 1927 56177 1983 56233
rect 2051 56177 2107 56233
rect 315 56095 369 56109
rect 369 56095 371 56109
rect 439 56095 493 56109
rect 493 56095 495 56109
rect 563 56095 617 56109
rect 617 56095 619 56109
rect 687 56095 741 56109
rect 741 56095 743 56109
rect 315 56053 371 56095
rect 439 56053 495 56095
rect 563 56053 619 56095
rect 687 56053 743 56095
rect 811 56053 867 56109
rect 935 56053 991 56109
rect 1059 56053 1115 56109
rect 1183 56053 1239 56109
rect 1307 56053 1363 56109
rect 1431 56053 1487 56109
rect 1555 56053 1611 56109
rect 1679 56053 1735 56109
rect 1803 56053 1859 56109
rect 1927 56053 1983 56109
rect 2051 56053 2107 56109
rect 20 54174 76 54176
rect 20 54122 22 54174
rect 22 54122 74 54174
rect 74 54122 76 54174
rect 20 54066 76 54122
rect 20 54014 22 54066
rect 22 54014 74 54066
rect 74 54014 76 54066
rect 20 53958 76 54014
rect 20 53906 22 53958
rect 22 53906 74 53958
rect 74 53906 76 53958
rect 20 53850 76 53906
rect 20 53798 22 53850
rect 22 53798 74 53850
rect 74 53798 76 53850
rect 20 53742 76 53798
rect 20 53690 22 53742
rect 22 53690 74 53742
rect 74 53690 76 53742
rect 20 53634 76 53690
rect 20 53582 22 53634
rect 22 53582 74 53634
rect 74 53582 76 53634
rect 20 53526 76 53582
rect 20 53474 22 53526
rect 22 53474 74 53526
rect 74 53474 76 53526
rect 20 53418 76 53474
rect 20 53366 22 53418
rect 22 53366 74 53418
rect 74 53366 76 53418
rect 20 53310 76 53366
rect 20 53258 22 53310
rect 22 53258 74 53310
rect 74 53258 76 53310
rect 20 53202 76 53258
rect 20 53150 22 53202
rect 22 53150 74 53202
rect 74 53150 76 53202
rect 20 53094 76 53150
rect 20 53042 22 53094
rect 22 53042 74 53094
rect 74 53042 76 53094
rect 20 52986 76 53042
rect 20 52934 22 52986
rect 22 52934 74 52986
rect 74 52934 76 52986
rect 20 52878 76 52934
rect 20 52826 22 52878
rect 22 52826 74 52878
rect 74 52826 76 52878
rect 20 52824 76 52826
rect 315 54111 369 54148
rect 369 54111 371 54148
rect 439 54111 493 54148
rect 493 54111 495 54148
rect 563 54111 617 54148
rect 617 54111 619 54148
rect 687 54111 741 54148
rect 741 54111 743 54148
rect 315 54092 371 54111
rect 439 54092 495 54111
rect 563 54092 619 54111
rect 687 54092 743 54111
rect 811 54092 867 54148
rect 935 54092 991 54148
rect 1059 54092 1115 54148
rect 1183 54092 1239 54148
rect 1307 54092 1363 54148
rect 1431 54092 1487 54148
rect 1555 54092 1611 54148
rect 1679 54092 1735 54148
rect 1803 54092 1859 54148
rect 1927 54092 1983 54148
rect 2051 54092 2107 54148
rect 315 53987 369 54024
rect 369 53987 371 54024
rect 439 53987 493 54024
rect 493 53987 495 54024
rect 563 53987 617 54024
rect 617 53987 619 54024
rect 687 53987 741 54024
rect 741 53987 743 54024
rect 315 53968 371 53987
rect 439 53968 495 53987
rect 563 53968 619 53987
rect 687 53968 743 53987
rect 811 53968 867 54024
rect 935 53968 991 54024
rect 1059 53968 1115 54024
rect 1183 53968 1239 54024
rect 1307 53968 1363 54024
rect 1431 53968 1487 54024
rect 1555 53968 1611 54024
rect 1679 53968 1735 54024
rect 1803 53968 1859 54024
rect 1927 53968 1983 54024
rect 2051 53968 2107 54024
rect 315 53863 369 53900
rect 369 53863 371 53900
rect 439 53863 493 53900
rect 493 53863 495 53900
rect 563 53863 617 53900
rect 617 53863 619 53900
rect 687 53863 741 53900
rect 741 53863 743 53900
rect 315 53844 371 53863
rect 439 53844 495 53863
rect 563 53844 619 53863
rect 687 53844 743 53863
rect 811 53844 867 53900
rect 935 53844 991 53900
rect 1059 53844 1115 53900
rect 1183 53844 1239 53900
rect 1307 53844 1363 53900
rect 1431 53844 1487 53900
rect 1555 53844 1611 53900
rect 1679 53844 1735 53900
rect 1803 53844 1859 53900
rect 1927 53844 1983 53900
rect 2051 53844 2107 53900
rect 315 53739 369 53776
rect 369 53739 371 53776
rect 439 53739 493 53776
rect 493 53739 495 53776
rect 563 53739 617 53776
rect 617 53739 619 53776
rect 687 53739 741 53776
rect 741 53739 743 53776
rect 315 53720 371 53739
rect 439 53720 495 53739
rect 563 53720 619 53739
rect 687 53720 743 53739
rect 811 53720 867 53776
rect 935 53720 991 53776
rect 1059 53720 1115 53776
rect 1183 53720 1239 53776
rect 1307 53720 1363 53776
rect 1431 53720 1487 53776
rect 1555 53720 1611 53776
rect 1679 53720 1735 53776
rect 1803 53720 1859 53776
rect 1927 53720 1983 53776
rect 2051 53720 2107 53776
rect 315 53615 369 53652
rect 369 53615 371 53652
rect 439 53615 493 53652
rect 493 53615 495 53652
rect 563 53615 617 53652
rect 617 53615 619 53652
rect 687 53615 741 53652
rect 741 53615 743 53652
rect 315 53596 371 53615
rect 439 53596 495 53615
rect 563 53596 619 53615
rect 687 53596 743 53615
rect 811 53596 867 53652
rect 935 53596 991 53652
rect 1059 53596 1115 53652
rect 1183 53596 1239 53652
rect 1307 53596 1363 53652
rect 1431 53596 1487 53652
rect 1555 53596 1611 53652
rect 1679 53596 1735 53652
rect 1803 53596 1859 53652
rect 1927 53596 1983 53652
rect 2051 53596 2107 53652
rect 315 53491 369 53528
rect 369 53491 371 53528
rect 439 53491 493 53528
rect 493 53491 495 53528
rect 563 53491 617 53528
rect 617 53491 619 53528
rect 687 53491 741 53528
rect 741 53491 743 53528
rect 315 53472 371 53491
rect 439 53472 495 53491
rect 563 53472 619 53491
rect 687 53472 743 53491
rect 811 53472 867 53528
rect 935 53483 991 53528
rect 1059 53483 1115 53528
rect 1183 53483 1239 53528
rect 1307 53483 1363 53528
rect 1431 53483 1487 53528
rect 1555 53483 1611 53528
rect 1679 53483 1735 53528
rect 1803 53483 1859 53528
rect 1927 53483 1983 53528
rect 2051 53483 2107 53528
rect 935 53472 977 53483
rect 977 53472 991 53483
rect 1059 53472 1085 53483
rect 1085 53472 1115 53483
rect 1183 53472 1193 53483
rect 1193 53472 1239 53483
rect 1307 53472 1353 53483
rect 1353 53472 1363 53483
rect 1431 53472 1461 53483
rect 1461 53472 1487 53483
rect 1555 53472 1569 53483
rect 1569 53472 1611 53483
rect 1679 53472 1733 53483
rect 1733 53472 1735 53483
rect 1803 53472 1841 53483
rect 1841 53472 1859 53483
rect 1927 53472 1949 53483
rect 1949 53472 1983 53483
rect 2051 53472 2057 53483
rect 2057 53472 2107 53483
rect 315 53367 369 53404
rect 369 53367 371 53404
rect 439 53367 493 53404
rect 493 53367 495 53404
rect 563 53367 617 53404
rect 617 53367 619 53404
rect 687 53367 741 53404
rect 741 53367 743 53404
rect 315 53348 371 53367
rect 439 53348 495 53367
rect 563 53348 619 53367
rect 687 53348 743 53367
rect 811 53348 867 53404
rect 935 53375 991 53404
rect 1059 53375 1115 53404
rect 1183 53375 1239 53404
rect 1307 53375 1363 53404
rect 1431 53375 1487 53404
rect 1555 53375 1611 53404
rect 1679 53375 1735 53404
rect 1803 53375 1859 53404
rect 1927 53375 1983 53404
rect 2051 53375 2107 53404
rect 935 53348 977 53375
rect 977 53348 991 53375
rect 1059 53348 1085 53375
rect 1085 53348 1115 53375
rect 1183 53348 1193 53375
rect 1193 53348 1239 53375
rect 1307 53348 1353 53375
rect 1353 53348 1363 53375
rect 1431 53348 1461 53375
rect 1461 53348 1487 53375
rect 1555 53348 1569 53375
rect 1569 53348 1611 53375
rect 1679 53348 1733 53375
rect 1733 53348 1735 53375
rect 1803 53348 1841 53375
rect 1841 53348 1859 53375
rect 1927 53348 1949 53375
rect 1949 53348 1983 53375
rect 2051 53348 2057 53375
rect 2057 53348 2107 53375
rect 315 53243 369 53280
rect 369 53243 371 53280
rect 439 53243 493 53280
rect 493 53243 495 53280
rect 563 53243 617 53280
rect 617 53243 619 53280
rect 687 53243 741 53280
rect 741 53243 743 53280
rect 315 53224 371 53243
rect 439 53224 495 53243
rect 563 53224 619 53243
rect 687 53224 743 53243
rect 811 53224 867 53280
rect 935 53267 991 53280
rect 1059 53267 1115 53280
rect 1183 53267 1239 53280
rect 1307 53267 1363 53280
rect 1431 53267 1487 53280
rect 1555 53267 1611 53280
rect 1679 53267 1735 53280
rect 1803 53267 1859 53280
rect 1927 53267 1983 53280
rect 2051 53267 2107 53280
rect 935 53224 977 53267
rect 977 53224 991 53267
rect 1059 53224 1085 53267
rect 1085 53224 1115 53267
rect 1183 53224 1193 53267
rect 1193 53224 1239 53267
rect 1307 53224 1353 53267
rect 1353 53224 1363 53267
rect 1431 53224 1461 53267
rect 1461 53224 1487 53267
rect 1555 53224 1569 53267
rect 1569 53224 1611 53267
rect 1679 53224 1733 53267
rect 1733 53224 1735 53267
rect 1803 53224 1841 53267
rect 1841 53224 1859 53267
rect 1927 53224 1949 53267
rect 1949 53224 1983 53267
rect 2051 53224 2057 53267
rect 2057 53224 2107 53267
rect 315 53100 371 53156
rect 439 53100 495 53156
rect 563 53100 619 53156
rect 687 53100 743 53156
rect 811 53100 867 53156
rect 935 53100 991 53156
rect 1059 53100 1115 53156
rect 1183 53100 1239 53156
rect 1307 53100 1363 53156
rect 1431 53100 1487 53156
rect 1555 53100 1611 53156
rect 1679 53100 1735 53156
rect 1803 53100 1859 53156
rect 1927 53100 1983 53156
rect 2051 53100 2107 53156
rect 315 52976 371 53032
rect 439 52976 495 53032
rect 563 52976 619 53032
rect 687 52976 743 53032
rect 811 52976 867 53032
rect 935 52976 991 53032
rect 1059 52976 1115 53032
rect 1183 52976 1239 53032
rect 1307 52976 1363 53032
rect 1431 52976 1487 53032
rect 1555 52976 1611 53032
rect 1679 52976 1735 53032
rect 1803 52976 1859 53032
rect 1927 52976 1983 53032
rect 2051 52976 2107 53032
rect 315 52852 371 52908
rect 439 52852 495 52908
rect 563 52852 619 52908
rect 687 52852 743 52908
rect 811 52852 867 52908
rect 935 52852 991 52908
rect 1059 52852 1115 52908
rect 1183 52852 1239 52908
rect 1307 52852 1363 52908
rect 1431 52852 1487 52908
rect 1555 52852 1611 52908
rect 1679 52852 1735 52908
rect 1803 52852 1859 52908
rect 1927 52852 1983 52908
rect 2051 52852 2107 52908
rect 20 52574 76 52576
rect 20 52522 22 52574
rect 22 52522 74 52574
rect 74 52522 76 52574
rect 20 52466 76 52522
rect 20 52414 22 52466
rect 22 52414 74 52466
rect 74 52414 76 52466
rect 20 52358 76 52414
rect 20 52306 22 52358
rect 22 52306 74 52358
rect 74 52306 76 52358
rect 20 52250 76 52306
rect 20 52198 22 52250
rect 22 52198 74 52250
rect 74 52198 76 52250
rect 20 52142 76 52198
rect 20 52090 22 52142
rect 22 52090 74 52142
rect 74 52090 76 52142
rect 20 52034 76 52090
rect 20 51982 22 52034
rect 22 51982 74 52034
rect 74 51982 76 52034
rect 20 51926 76 51982
rect 20 51874 22 51926
rect 22 51874 74 51926
rect 74 51874 76 51926
rect 20 51818 76 51874
rect 20 51766 22 51818
rect 22 51766 74 51818
rect 74 51766 76 51818
rect 20 51710 76 51766
rect 20 51658 22 51710
rect 22 51658 74 51710
rect 74 51658 76 51710
rect 20 51602 76 51658
rect 20 51550 22 51602
rect 22 51550 74 51602
rect 74 51550 76 51602
rect 20 51494 76 51550
rect 20 51442 22 51494
rect 22 51442 74 51494
rect 74 51442 76 51494
rect 20 51386 76 51442
rect 20 51334 22 51386
rect 22 51334 74 51386
rect 74 51334 76 51386
rect 20 51278 76 51334
rect 20 51226 22 51278
rect 22 51226 74 51278
rect 74 51226 76 51278
rect 20 51224 76 51226
rect 315 52492 371 52548
rect 439 52492 495 52548
rect 563 52492 619 52548
rect 687 52492 743 52548
rect 811 52492 867 52548
rect 935 52492 991 52548
rect 1059 52492 1115 52548
rect 1183 52492 1239 52548
rect 1307 52492 1363 52548
rect 1431 52492 1487 52548
rect 1555 52492 1611 52548
rect 1679 52492 1735 52548
rect 1803 52492 1859 52548
rect 1927 52492 1983 52548
rect 2051 52492 2107 52548
rect 315 52368 371 52424
rect 439 52368 495 52424
rect 563 52368 619 52424
rect 687 52368 743 52424
rect 811 52368 867 52424
rect 935 52368 991 52424
rect 1059 52368 1115 52424
rect 1183 52368 1239 52424
rect 1307 52368 1363 52424
rect 1431 52368 1487 52424
rect 1555 52368 1611 52424
rect 1679 52368 1735 52424
rect 1803 52368 1859 52424
rect 1927 52368 1983 52424
rect 2051 52368 2107 52424
rect 315 52244 371 52300
rect 439 52244 495 52300
rect 563 52244 619 52300
rect 687 52244 743 52300
rect 811 52244 867 52300
rect 935 52244 991 52300
rect 1059 52244 1115 52300
rect 1183 52244 1239 52300
rect 1307 52244 1363 52300
rect 1431 52244 1487 52300
rect 1555 52244 1611 52300
rect 1679 52244 1735 52300
rect 1803 52244 1859 52300
rect 1927 52244 1983 52300
rect 2051 52244 2107 52300
rect 315 52120 371 52176
rect 439 52120 495 52176
rect 563 52120 619 52176
rect 687 52120 743 52176
rect 811 52120 867 52176
rect 935 52120 991 52176
rect 1059 52120 1115 52176
rect 1183 52120 1239 52176
rect 1307 52120 1363 52176
rect 1431 52120 1487 52176
rect 1555 52120 1611 52176
rect 1679 52120 1735 52176
rect 1803 52120 1859 52176
rect 1927 52120 1983 52176
rect 2051 52120 2107 52176
rect 315 51996 371 52052
rect 439 51996 495 52052
rect 563 51996 619 52052
rect 687 51996 743 52052
rect 811 51996 867 52052
rect 935 51996 991 52052
rect 1059 51996 1115 52052
rect 1183 51996 1239 52052
rect 1307 51996 1363 52052
rect 1431 51996 1487 52052
rect 1555 51996 1611 52052
rect 1679 51996 1735 52052
rect 1803 51996 1859 52052
rect 1927 51996 1983 52052
rect 2051 51996 2107 52052
rect 315 51872 371 51928
rect 439 51872 495 51928
rect 563 51872 619 51928
rect 687 51872 743 51928
rect 811 51872 867 51928
rect 935 51872 991 51928
rect 1059 51872 1115 51928
rect 1183 51872 1239 51928
rect 1307 51872 1363 51928
rect 1431 51872 1487 51928
rect 1555 51872 1611 51928
rect 1679 51872 1735 51928
rect 1803 51872 1859 51928
rect 1927 51872 1983 51928
rect 2051 51872 2107 51928
rect 315 51748 371 51804
rect 439 51748 495 51804
rect 563 51748 619 51804
rect 687 51748 743 51804
rect 811 51748 867 51804
rect 935 51748 991 51804
rect 1059 51748 1115 51804
rect 1183 51748 1239 51804
rect 1307 51748 1363 51804
rect 1431 51748 1487 51804
rect 1555 51748 1611 51804
rect 1679 51748 1735 51804
rect 1803 51748 1859 51804
rect 1927 51748 1983 51804
rect 2051 51748 2107 51804
rect 315 51624 371 51680
rect 439 51624 495 51680
rect 563 51624 619 51680
rect 687 51624 743 51680
rect 811 51624 867 51680
rect 935 51624 991 51680
rect 1059 51624 1115 51680
rect 1183 51624 1239 51680
rect 1307 51624 1363 51680
rect 1431 51624 1487 51680
rect 1555 51624 1611 51680
rect 1679 51624 1735 51680
rect 1803 51624 1859 51680
rect 1927 51624 1983 51680
rect 2051 51624 2107 51680
rect 315 51500 371 51556
rect 439 51500 495 51556
rect 563 51500 619 51556
rect 687 51500 743 51556
rect 811 51500 867 51556
rect 935 51500 991 51556
rect 1059 51500 1115 51556
rect 1183 51500 1239 51556
rect 1307 51500 1363 51556
rect 1431 51500 1487 51556
rect 1555 51500 1611 51556
rect 1679 51500 1735 51556
rect 1803 51500 1859 51556
rect 1927 51500 1983 51556
rect 2051 51500 2107 51556
rect 315 51376 371 51432
rect 439 51376 495 51432
rect 563 51376 619 51432
rect 687 51376 743 51432
rect 811 51376 867 51432
rect 935 51376 991 51432
rect 1059 51376 1115 51432
rect 1183 51376 1239 51432
rect 1307 51376 1363 51432
rect 1431 51376 1487 51432
rect 1555 51376 1611 51432
rect 1679 51376 1735 51432
rect 1803 51376 1859 51432
rect 1927 51376 1983 51432
rect 2051 51376 2107 51432
rect 315 51252 371 51308
rect 439 51252 495 51308
rect 563 51252 619 51308
rect 687 51252 743 51308
rect 811 51252 867 51308
rect 935 51252 991 51308
rect 1059 51252 1115 51308
rect 1183 51252 1239 51308
rect 1307 51252 1363 51308
rect 1431 51252 1487 51308
rect 1555 51252 1611 51308
rect 1679 51252 1735 51308
rect 1803 51252 1859 51308
rect 1927 51252 1983 51308
rect 2051 51252 2107 51308
rect 20 49374 76 49376
rect 20 49322 22 49374
rect 22 49322 74 49374
rect 74 49322 76 49374
rect 20 49266 76 49322
rect 20 49214 22 49266
rect 22 49214 74 49266
rect 74 49214 76 49266
rect 20 49158 76 49214
rect 20 49106 22 49158
rect 22 49106 74 49158
rect 74 49106 76 49158
rect 20 49050 76 49106
rect 20 48998 22 49050
rect 22 48998 74 49050
rect 74 48998 76 49050
rect 20 48942 76 48998
rect 20 48890 22 48942
rect 22 48890 74 48942
rect 74 48890 76 48942
rect 20 48834 76 48890
rect 20 48782 22 48834
rect 22 48782 74 48834
rect 74 48782 76 48834
rect 20 48726 76 48782
rect 20 48674 22 48726
rect 22 48674 74 48726
rect 74 48674 76 48726
rect 20 48618 76 48674
rect 20 48566 22 48618
rect 22 48566 74 48618
rect 74 48566 76 48618
rect 20 48510 76 48566
rect 20 48458 22 48510
rect 22 48458 74 48510
rect 74 48458 76 48510
rect 20 48402 76 48458
rect 20 48350 22 48402
rect 22 48350 74 48402
rect 74 48350 76 48402
rect 20 48294 76 48350
rect 20 48242 22 48294
rect 22 48242 74 48294
rect 74 48242 76 48294
rect 20 48186 76 48242
rect 20 48134 22 48186
rect 22 48134 74 48186
rect 74 48134 76 48186
rect 20 48078 76 48134
rect 20 48026 22 48078
rect 22 48026 74 48078
rect 74 48026 76 48078
rect 20 48024 76 48026
rect 2491 55692 2547 55748
rect 2615 55692 2671 55748
rect 2491 55568 2547 55624
rect 2615 55568 2671 55624
rect 2491 55444 2547 55500
rect 2615 55444 2671 55500
rect 2491 55320 2547 55376
rect 2615 55320 2671 55376
rect 2491 55196 2547 55252
rect 2615 55196 2671 55252
rect 2491 55072 2547 55128
rect 2615 55072 2671 55128
rect 2491 54948 2547 55004
rect 2615 54948 2671 55004
rect 2491 54824 2547 54880
rect 2615 54824 2671 54880
rect 2491 54700 2547 54756
rect 2615 54700 2671 54756
rect 2491 54576 2547 54632
rect 2615 54576 2671 54632
rect 2491 54452 2547 54508
rect 2615 54452 2671 54508
rect 315 49292 371 49348
rect 439 49292 495 49348
rect 563 49292 619 49348
rect 687 49292 743 49348
rect 811 49292 867 49348
rect 935 49292 991 49348
rect 1059 49292 1115 49348
rect 1183 49292 1239 49348
rect 1307 49292 1363 49348
rect 1431 49292 1487 49348
rect 1555 49292 1611 49348
rect 1679 49292 1735 49348
rect 1803 49292 1859 49348
rect 1927 49292 1983 49348
rect 2051 49292 2107 49348
rect 315 49168 371 49224
rect 439 49168 495 49224
rect 563 49168 619 49224
rect 687 49168 743 49224
rect 811 49168 867 49224
rect 935 49168 991 49224
rect 1059 49168 1115 49224
rect 1183 49168 1239 49224
rect 1307 49168 1363 49224
rect 1431 49168 1487 49224
rect 1555 49168 1611 49224
rect 1679 49168 1735 49224
rect 1803 49168 1859 49224
rect 1927 49168 1983 49224
rect 2051 49168 2107 49224
rect 315 49044 371 49100
rect 439 49044 495 49100
rect 563 49044 619 49100
rect 687 49044 743 49100
rect 811 49044 867 49100
rect 935 49044 991 49100
rect 1059 49044 1115 49100
rect 1183 49044 1239 49100
rect 1307 49044 1363 49100
rect 1431 49044 1487 49100
rect 1555 49044 1611 49100
rect 1679 49044 1735 49100
rect 1803 49044 1859 49100
rect 1927 49044 1983 49100
rect 2051 49044 2107 49100
rect 315 48920 371 48976
rect 439 48920 495 48976
rect 563 48920 619 48976
rect 687 48920 743 48976
rect 811 48920 867 48976
rect 935 48920 991 48976
rect 1059 48920 1115 48976
rect 1183 48920 1239 48976
rect 1307 48920 1363 48976
rect 1431 48920 1487 48976
rect 1555 48920 1611 48976
rect 1679 48920 1735 48976
rect 1803 48920 1859 48976
rect 1927 48920 1983 48976
rect 2051 48920 2107 48976
rect 315 48796 371 48852
rect 439 48796 495 48852
rect 563 48796 619 48852
rect 687 48796 743 48852
rect 811 48796 867 48852
rect 935 48796 991 48852
rect 1059 48796 1115 48852
rect 1183 48796 1239 48852
rect 1307 48796 1363 48852
rect 1431 48796 1487 48852
rect 1555 48796 1611 48852
rect 1679 48796 1735 48852
rect 1803 48796 1859 48852
rect 1927 48796 1983 48852
rect 2051 48796 2107 48852
rect 315 48672 371 48728
rect 439 48672 495 48728
rect 563 48672 619 48728
rect 687 48672 743 48728
rect 811 48672 867 48728
rect 935 48672 991 48728
rect 1059 48672 1115 48728
rect 1183 48672 1239 48728
rect 1307 48672 1363 48728
rect 1431 48672 1487 48728
rect 1555 48672 1611 48728
rect 1679 48672 1735 48728
rect 1803 48672 1859 48728
rect 1927 48672 1983 48728
rect 2051 48672 2107 48728
rect 315 48548 371 48604
rect 439 48548 495 48604
rect 563 48548 619 48604
rect 687 48548 743 48604
rect 811 48548 867 48604
rect 935 48548 991 48604
rect 1059 48548 1115 48604
rect 1183 48548 1239 48604
rect 1307 48548 1363 48604
rect 1431 48548 1487 48604
rect 1555 48548 1611 48604
rect 1679 48548 1735 48604
rect 1803 48548 1859 48604
rect 1927 48548 1983 48604
rect 2051 48548 2107 48604
rect 315 48424 371 48480
rect 439 48424 495 48480
rect 563 48424 619 48480
rect 687 48424 743 48480
rect 811 48424 867 48480
rect 935 48424 991 48480
rect 1059 48424 1115 48480
rect 1183 48424 1239 48480
rect 1307 48424 1363 48480
rect 1431 48424 1487 48480
rect 1555 48424 1611 48480
rect 1679 48424 1735 48480
rect 1803 48424 1859 48480
rect 1927 48424 1983 48480
rect 2051 48424 2107 48480
rect 315 48300 371 48356
rect 439 48300 495 48356
rect 563 48300 619 48356
rect 687 48300 743 48356
rect 811 48300 867 48356
rect 935 48300 991 48356
rect 1059 48300 1115 48356
rect 1183 48300 1239 48356
rect 1307 48300 1363 48356
rect 1431 48300 1487 48356
rect 1555 48300 1611 48356
rect 1679 48300 1735 48356
rect 1803 48300 1859 48356
rect 1927 48300 1983 48356
rect 2051 48300 2107 48356
rect 315 48176 371 48232
rect 439 48176 495 48232
rect 563 48176 619 48232
rect 687 48176 743 48232
rect 811 48176 867 48232
rect 935 48176 991 48232
rect 1059 48176 1115 48232
rect 1183 48176 1239 48232
rect 1307 48176 1363 48232
rect 1431 48176 1487 48232
rect 1555 48176 1611 48232
rect 1679 48176 1735 48232
rect 1803 48176 1859 48232
rect 1927 48176 1983 48232
rect 2051 48176 2107 48232
rect 315 48052 371 48108
rect 439 48052 495 48108
rect 563 48052 619 48108
rect 687 48052 743 48108
rect 811 48052 867 48108
rect 935 48052 991 48108
rect 1059 48052 1115 48108
rect 1183 48052 1239 48108
rect 1307 48052 1363 48108
rect 1431 48052 1487 48108
rect 1555 48052 1611 48108
rect 1679 48052 1735 48108
rect 1803 48052 1859 48108
rect 1927 48052 1983 48108
rect 2051 48052 2107 48108
rect 2302 50870 2358 50926
rect 2302 50738 2358 50794
rect 2302 50606 2358 50662
rect 2302 50474 2358 50530
rect 2302 50342 2358 50398
rect 2302 50210 2358 50266
rect 2302 50078 2358 50134
rect 2302 49946 2358 50002
rect 2302 49814 2358 49870
rect 2302 49682 2358 49738
rect 20 46174 76 46176
rect 20 46122 22 46174
rect 22 46122 74 46174
rect 74 46122 76 46174
rect 20 46066 76 46122
rect 20 46014 22 46066
rect 22 46014 74 46066
rect 74 46014 76 46066
rect 20 45958 76 46014
rect 20 45906 22 45958
rect 22 45906 74 45958
rect 74 45906 76 45958
rect 20 45850 76 45906
rect 20 45798 22 45850
rect 22 45798 74 45850
rect 74 45798 76 45850
rect 20 45742 76 45798
rect 20 45690 22 45742
rect 22 45690 74 45742
rect 74 45690 76 45742
rect 20 45634 76 45690
rect 20 45582 22 45634
rect 22 45582 74 45634
rect 74 45582 76 45634
rect 20 45526 76 45582
rect 20 45474 22 45526
rect 22 45474 74 45526
rect 74 45474 76 45526
rect 20 45418 76 45474
rect 20 45366 22 45418
rect 22 45366 74 45418
rect 74 45366 76 45418
rect 20 45310 76 45366
rect 20 45258 22 45310
rect 22 45258 74 45310
rect 74 45258 76 45310
rect 20 45202 76 45258
rect 20 45150 22 45202
rect 22 45150 74 45202
rect 74 45150 76 45202
rect 20 45094 76 45150
rect 20 45042 22 45094
rect 22 45042 74 45094
rect 74 45042 76 45094
rect 20 44986 76 45042
rect 20 44934 22 44986
rect 22 44934 74 44986
rect 74 44934 76 44986
rect 20 44878 76 44934
rect 20 44826 22 44878
rect 22 44826 74 44878
rect 74 44826 76 44878
rect 20 44824 76 44826
rect 315 46092 371 46148
rect 439 46092 495 46148
rect 563 46092 619 46148
rect 687 46092 743 46148
rect 811 46092 867 46148
rect 935 46092 991 46148
rect 1059 46092 1115 46148
rect 1183 46092 1239 46148
rect 1307 46092 1363 46148
rect 1431 46092 1487 46148
rect 1555 46092 1611 46148
rect 1679 46092 1735 46148
rect 1803 46092 1859 46148
rect 1927 46092 1983 46148
rect 2051 46092 2107 46148
rect 315 45968 371 46024
rect 439 45968 495 46024
rect 563 45968 619 46024
rect 687 45968 743 46024
rect 811 45968 867 46024
rect 935 45968 991 46024
rect 1059 45968 1115 46024
rect 1183 45968 1239 46024
rect 1307 45968 1363 46024
rect 1431 45968 1487 46024
rect 1555 45968 1611 46024
rect 1679 45968 1735 46024
rect 1803 45968 1859 46024
rect 1927 45968 1983 46024
rect 2051 45968 2107 46024
rect 315 45844 371 45900
rect 439 45844 495 45900
rect 563 45844 619 45900
rect 687 45844 743 45900
rect 811 45844 867 45900
rect 935 45844 991 45900
rect 1059 45844 1115 45900
rect 1183 45844 1239 45900
rect 1307 45844 1363 45900
rect 1431 45844 1487 45900
rect 1555 45844 1611 45900
rect 1679 45844 1735 45900
rect 1803 45844 1859 45900
rect 1927 45844 1983 45900
rect 2051 45844 2107 45900
rect 315 45720 371 45776
rect 439 45720 495 45776
rect 563 45720 619 45776
rect 687 45720 743 45776
rect 811 45720 867 45776
rect 935 45720 991 45776
rect 1059 45720 1115 45776
rect 1183 45720 1239 45776
rect 1307 45720 1363 45776
rect 1431 45720 1487 45776
rect 1555 45720 1611 45776
rect 1679 45720 1735 45776
rect 1803 45720 1859 45776
rect 1927 45720 1983 45776
rect 2051 45720 2107 45776
rect 315 45596 371 45652
rect 439 45596 495 45652
rect 563 45596 619 45652
rect 687 45596 743 45652
rect 811 45596 867 45652
rect 935 45596 991 45652
rect 1059 45596 1115 45652
rect 1183 45596 1239 45652
rect 1307 45596 1363 45652
rect 1431 45596 1487 45652
rect 1555 45596 1611 45652
rect 1679 45596 1735 45652
rect 1803 45596 1859 45652
rect 1927 45596 1983 45652
rect 2051 45596 2107 45652
rect 315 45472 371 45528
rect 439 45472 495 45528
rect 563 45472 619 45528
rect 687 45472 743 45528
rect 811 45472 867 45528
rect 935 45472 991 45528
rect 1059 45472 1115 45528
rect 1183 45472 1239 45528
rect 1307 45472 1363 45528
rect 1431 45472 1487 45528
rect 1555 45472 1611 45528
rect 1679 45472 1735 45528
rect 1803 45472 1859 45528
rect 1927 45472 1983 45528
rect 2051 45472 2107 45528
rect 315 45348 371 45404
rect 439 45348 495 45404
rect 563 45348 619 45404
rect 687 45348 743 45404
rect 811 45348 867 45404
rect 935 45348 991 45404
rect 1059 45348 1115 45404
rect 1183 45348 1239 45404
rect 1307 45348 1363 45404
rect 1431 45348 1487 45404
rect 1555 45348 1611 45404
rect 1679 45348 1735 45404
rect 1803 45348 1859 45404
rect 1927 45348 1983 45404
rect 2051 45348 2107 45404
rect 315 45224 371 45280
rect 439 45224 495 45280
rect 563 45224 619 45280
rect 687 45224 743 45280
rect 811 45224 867 45280
rect 935 45224 991 45280
rect 1059 45224 1115 45280
rect 1183 45224 1239 45280
rect 1307 45224 1363 45280
rect 1431 45224 1487 45280
rect 1555 45224 1611 45280
rect 1679 45224 1735 45280
rect 1803 45224 1859 45280
rect 1927 45224 1983 45280
rect 2051 45224 2107 45280
rect 315 45100 371 45156
rect 439 45100 495 45156
rect 563 45100 619 45156
rect 687 45100 743 45156
rect 811 45100 867 45156
rect 935 45100 991 45156
rect 1059 45100 1115 45156
rect 1183 45100 1239 45156
rect 1307 45100 1363 45156
rect 1431 45100 1487 45156
rect 1555 45100 1611 45156
rect 1679 45100 1735 45156
rect 1803 45100 1859 45156
rect 1927 45100 1983 45156
rect 2051 45100 2107 45156
rect 315 44976 371 45032
rect 439 44976 495 45032
rect 563 44976 619 45032
rect 687 44976 743 45032
rect 811 44976 867 45032
rect 935 44976 991 45032
rect 1059 44976 1115 45032
rect 1183 44976 1239 45032
rect 1307 44976 1363 45032
rect 1431 44976 1487 45032
rect 1555 44976 1611 45032
rect 1679 44976 1735 45032
rect 1803 44976 1859 45032
rect 1927 44976 1983 45032
rect 2051 44976 2107 45032
rect 315 44852 371 44908
rect 439 44852 495 44908
rect 563 44852 619 44908
rect 687 44852 743 44908
rect 811 44852 867 44908
rect 935 44852 991 44908
rect 1059 44852 1115 44908
rect 1183 44852 1239 44908
rect 1307 44852 1363 44908
rect 1431 44852 1487 44908
rect 1555 44852 1611 44908
rect 1679 44852 1735 44908
rect 1803 44852 1859 44908
rect 1927 44852 1983 44908
rect 2051 44852 2107 44908
rect 2491 47692 2547 47748
rect 2615 47734 2671 47748
rect 2615 47692 2642 47734
rect 2642 47692 2671 47734
rect 2491 47568 2547 47624
rect 2615 47568 2671 47624
rect 2491 47444 2547 47500
rect 2615 47444 2671 47500
rect 2491 47320 2547 47376
rect 2615 47320 2671 47376
rect 2491 47196 2547 47252
rect 2615 47196 2671 47252
rect 2808 57169 2864 57225
rect 2932 57169 2988 57225
rect 3056 57169 3112 57225
rect 3180 57169 3236 57225
rect 3304 57169 3360 57225
rect 3428 57169 3484 57225
rect 3552 57169 3608 57225
rect 3676 57169 3732 57225
rect 3800 57169 3856 57225
rect 3924 57169 3980 57225
rect 4048 57169 4104 57225
rect 4172 57169 4228 57225
rect 4296 57169 4352 57225
rect 4420 57169 4476 57225
rect 4544 57169 4600 57225
rect 4668 57169 4724 57225
rect 2808 57052 2820 57101
rect 2820 57052 2864 57101
rect 2932 57052 2984 57101
rect 2984 57052 2988 57101
rect 3056 57052 3092 57101
rect 3092 57052 3112 57101
rect 3180 57052 3200 57101
rect 3200 57052 3236 57101
rect 3304 57052 3308 57101
rect 3308 57052 3360 57101
rect 3428 57052 3468 57101
rect 3468 57052 3484 57101
rect 3552 57052 3576 57101
rect 3576 57052 3608 57101
rect 3676 57052 3684 57101
rect 3684 57052 3732 57101
rect 3800 57052 3848 57101
rect 3848 57052 3856 57101
rect 3924 57052 3956 57101
rect 3956 57052 3980 57101
rect 4048 57052 4064 57101
rect 4064 57052 4104 57101
rect 4172 57052 4224 57101
rect 4224 57052 4228 57101
rect 4296 57052 4332 57101
rect 4332 57052 4352 57101
rect 4420 57052 4440 57101
rect 4440 57052 4476 57101
rect 4544 57052 4548 57101
rect 4548 57052 4600 57101
rect 4668 57052 4712 57101
rect 4712 57052 4724 57101
rect 2808 57045 2864 57052
rect 2932 57045 2988 57052
rect 3056 57045 3112 57052
rect 3180 57045 3236 57052
rect 3304 57045 3360 57052
rect 3428 57045 3484 57052
rect 3552 57045 3608 57052
rect 3676 57045 3732 57052
rect 3800 57045 3856 57052
rect 3924 57045 3980 57052
rect 4048 57045 4104 57052
rect 4172 57045 4228 57052
rect 4296 57045 4352 57052
rect 4420 57045 4476 57052
rect 4544 57045 4600 57052
rect 4668 57045 4724 57052
rect 2808 56921 2864 56977
rect 2932 56921 2988 56977
rect 3056 56921 3112 56977
rect 3180 56921 3236 56977
rect 3304 56921 3360 56977
rect 3428 56921 3484 56977
rect 3552 56921 3608 56977
rect 3676 56921 3732 56977
rect 3800 56921 3856 56977
rect 3924 56921 3980 56977
rect 4048 56921 4104 56977
rect 4172 56921 4228 56977
rect 4296 56921 4352 56977
rect 4420 56921 4476 56977
rect 4544 56921 4600 56977
rect 4668 56921 4724 56977
rect 2808 56797 2864 56853
rect 2932 56797 2988 56853
rect 3056 56797 3112 56853
rect 3180 56797 3236 56853
rect 3304 56797 3360 56853
rect 3428 56797 3484 56853
rect 3552 56797 3608 56853
rect 3676 56797 3732 56853
rect 3800 56797 3856 56853
rect 3924 56797 3980 56853
rect 4048 56797 4104 56853
rect 4172 56797 4228 56853
rect 4296 56797 4352 56853
rect 4420 56797 4476 56853
rect 4544 56797 4600 56853
rect 4668 56797 4724 56853
rect 2808 56673 2864 56729
rect 2932 56673 2988 56729
rect 3056 56673 3112 56729
rect 3180 56673 3236 56729
rect 3304 56673 3360 56729
rect 3428 56673 3484 56729
rect 3552 56673 3608 56729
rect 3676 56673 3732 56729
rect 3800 56673 3856 56729
rect 3924 56673 3980 56729
rect 4048 56673 4104 56729
rect 4172 56673 4228 56729
rect 4296 56673 4352 56729
rect 4420 56673 4476 56729
rect 4544 56673 4600 56729
rect 4668 56673 4724 56729
rect 2808 56549 2864 56605
rect 2932 56549 2988 56605
rect 3056 56549 3112 56605
rect 3180 56549 3236 56605
rect 3304 56549 3360 56605
rect 3428 56549 3484 56605
rect 3552 56549 3608 56605
rect 3676 56549 3732 56605
rect 3800 56549 3856 56605
rect 3924 56591 3955 56605
rect 3955 56591 3980 56605
rect 4048 56591 4079 56605
rect 4079 56591 4104 56605
rect 4172 56591 4203 56605
rect 4203 56591 4228 56605
rect 3924 56549 3980 56591
rect 4048 56549 4104 56591
rect 4172 56549 4228 56591
rect 4296 56549 4352 56605
rect 4420 56549 4476 56605
rect 4544 56549 4600 56605
rect 4668 56549 4724 56605
rect 2808 56425 2864 56481
rect 2932 56425 2988 56481
rect 3056 56425 3112 56481
rect 3180 56425 3236 56481
rect 3304 56425 3360 56481
rect 3428 56425 3484 56481
rect 3552 56425 3608 56481
rect 3676 56425 3732 56481
rect 3800 56425 3856 56481
rect 3924 56467 3955 56481
rect 3955 56467 3980 56481
rect 4048 56467 4079 56481
rect 4079 56467 4104 56481
rect 4172 56467 4203 56481
rect 4203 56467 4228 56481
rect 3924 56425 3980 56467
rect 4048 56425 4104 56467
rect 4172 56425 4228 56467
rect 4296 56425 4352 56481
rect 4420 56425 4476 56481
rect 4544 56425 4600 56481
rect 4668 56425 4724 56481
rect 2808 56301 2864 56357
rect 2932 56301 2988 56357
rect 3056 56301 3112 56357
rect 3180 56301 3236 56357
rect 3304 56301 3360 56357
rect 3428 56301 3484 56357
rect 3552 56301 3608 56357
rect 3676 56301 3732 56357
rect 3800 56301 3856 56357
rect 3924 56343 3955 56357
rect 3955 56343 3980 56357
rect 4048 56343 4079 56357
rect 4079 56343 4104 56357
rect 4172 56343 4203 56357
rect 4203 56343 4228 56357
rect 3924 56301 3980 56343
rect 4048 56301 4104 56343
rect 4172 56301 4228 56343
rect 4296 56301 4352 56357
rect 4420 56301 4476 56357
rect 4544 56301 4600 56357
rect 4668 56301 4724 56357
rect 2808 56177 2864 56233
rect 2932 56177 2988 56233
rect 3056 56177 3112 56233
rect 3180 56177 3236 56233
rect 3304 56177 3360 56233
rect 3428 56177 3484 56233
rect 3552 56177 3608 56233
rect 3676 56177 3732 56233
rect 3800 56177 3856 56233
rect 3924 56219 3955 56233
rect 3955 56219 3980 56233
rect 4048 56219 4079 56233
rect 4079 56219 4104 56233
rect 4172 56219 4203 56233
rect 4203 56219 4228 56233
rect 3924 56177 3980 56219
rect 4048 56177 4104 56219
rect 4172 56177 4228 56219
rect 4296 56177 4352 56233
rect 4420 56177 4476 56233
rect 4544 56177 4600 56233
rect 4668 56177 4724 56233
rect 2808 56053 2864 56109
rect 2932 56053 2988 56109
rect 3056 56053 3112 56109
rect 3180 56053 3236 56109
rect 3304 56053 3360 56109
rect 3428 56053 3484 56109
rect 3552 56053 3608 56109
rect 3676 56053 3732 56109
rect 3800 56053 3856 56109
rect 3924 56095 3955 56109
rect 3955 56095 3980 56109
rect 4048 56095 4079 56109
rect 4079 56095 4104 56109
rect 4172 56095 4203 56109
rect 4203 56095 4228 56109
rect 3924 56053 3980 56095
rect 4048 56053 4104 56095
rect 4172 56053 4228 56095
rect 4296 56053 4352 56109
rect 4420 56053 4476 56109
rect 4544 56053 4600 56109
rect 4668 56053 4724 56109
rect 2808 54092 2864 54148
rect 2932 54092 2988 54148
rect 3056 54092 3112 54148
rect 3180 54092 3236 54148
rect 3304 54092 3360 54148
rect 3428 54092 3484 54148
rect 3552 54092 3608 54148
rect 3676 54092 3732 54148
rect 3800 54092 3856 54148
rect 3924 54111 3955 54148
rect 3955 54111 3980 54148
rect 4048 54111 4079 54148
rect 4079 54111 4104 54148
rect 4172 54111 4203 54148
rect 4203 54111 4228 54148
rect 3924 54092 3980 54111
rect 4048 54092 4104 54111
rect 4172 54092 4228 54111
rect 4296 54092 4352 54148
rect 4420 54092 4476 54148
rect 4544 54092 4600 54148
rect 4668 54092 4724 54148
rect 2808 53968 2864 54024
rect 2932 53968 2988 54024
rect 3056 53968 3112 54024
rect 3180 53968 3236 54024
rect 3304 53968 3360 54024
rect 3428 53968 3484 54024
rect 3552 53968 3608 54024
rect 3676 53968 3732 54024
rect 3800 53968 3856 54024
rect 3924 53987 3955 54024
rect 3955 53987 3980 54024
rect 4048 53987 4079 54024
rect 4079 53987 4104 54024
rect 4172 53987 4203 54024
rect 4203 53987 4228 54024
rect 3924 53968 3980 53987
rect 4048 53968 4104 53987
rect 4172 53968 4228 53987
rect 4296 53968 4352 54024
rect 4420 53968 4476 54024
rect 4544 53968 4600 54024
rect 4668 53968 4724 54024
rect 2808 53844 2864 53900
rect 2932 53844 2988 53900
rect 3056 53844 3112 53900
rect 3180 53844 3236 53900
rect 3304 53844 3360 53900
rect 3428 53844 3484 53900
rect 3552 53844 3608 53900
rect 3676 53844 3732 53900
rect 3800 53844 3856 53900
rect 3924 53863 3955 53900
rect 3955 53863 3980 53900
rect 4048 53863 4079 53900
rect 4079 53863 4104 53900
rect 4172 53863 4203 53900
rect 4203 53863 4228 53900
rect 3924 53844 3980 53863
rect 4048 53844 4104 53863
rect 4172 53844 4228 53863
rect 4296 53844 4352 53900
rect 4420 53844 4476 53900
rect 4544 53844 4600 53900
rect 4668 53844 4724 53900
rect 2808 53720 2864 53776
rect 2932 53720 2988 53776
rect 3056 53720 3112 53776
rect 3180 53720 3236 53776
rect 3304 53720 3360 53776
rect 3428 53720 3484 53776
rect 3552 53720 3608 53776
rect 3676 53720 3732 53776
rect 3800 53720 3856 53776
rect 3924 53739 3955 53776
rect 3955 53739 3980 53776
rect 4048 53739 4079 53776
rect 4079 53739 4104 53776
rect 4172 53739 4203 53776
rect 4203 53739 4228 53776
rect 3924 53720 3980 53739
rect 4048 53720 4104 53739
rect 4172 53720 4228 53739
rect 4296 53720 4352 53776
rect 4420 53720 4476 53776
rect 4544 53720 4600 53776
rect 4668 53720 4724 53776
rect 2808 53596 2864 53652
rect 2932 53596 2988 53652
rect 3056 53596 3112 53652
rect 3180 53596 3236 53652
rect 3304 53596 3360 53652
rect 3428 53596 3484 53652
rect 3552 53596 3608 53652
rect 3676 53596 3732 53652
rect 3800 53596 3856 53652
rect 3924 53615 3955 53652
rect 3955 53615 3980 53652
rect 4048 53615 4079 53652
rect 4079 53615 4104 53652
rect 4172 53615 4203 53652
rect 4203 53615 4228 53652
rect 3924 53596 3980 53615
rect 4048 53596 4104 53615
rect 4172 53596 4228 53615
rect 4296 53596 4352 53652
rect 4420 53596 4476 53652
rect 4544 53596 4600 53652
rect 4668 53596 4724 53652
rect 2808 53483 2864 53528
rect 2932 53483 2988 53528
rect 3056 53483 3112 53528
rect 3180 53483 3236 53528
rect 3304 53483 3360 53528
rect 3428 53483 3484 53528
rect 3552 53483 3608 53528
rect 3676 53483 3732 53528
rect 2808 53472 2815 53483
rect 2815 53472 2864 53483
rect 2932 53472 2979 53483
rect 2979 53472 2988 53483
rect 3056 53472 3087 53483
rect 3087 53472 3112 53483
rect 3180 53472 3195 53483
rect 3195 53472 3236 53483
rect 3304 53472 3355 53483
rect 3355 53472 3360 53483
rect 3428 53472 3463 53483
rect 3463 53472 3484 53483
rect 3552 53472 3571 53483
rect 3571 53472 3608 53483
rect 3676 53472 3679 53483
rect 3679 53472 3732 53483
rect 3800 53472 3856 53528
rect 3924 53491 3955 53528
rect 3955 53491 3980 53528
rect 4048 53491 4079 53528
rect 4079 53491 4104 53528
rect 4172 53491 4203 53528
rect 4203 53491 4228 53528
rect 3924 53472 3980 53491
rect 4048 53472 4104 53491
rect 4172 53472 4228 53491
rect 4296 53472 4352 53528
rect 4420 53472 4476 53528
rect 4544 53472 4600 53528
rect 4668 53472 4724 53528
rect 2808 53375 2864 53404
rect 2932 53375 2988 53404
rect 3056 53375 3112 53404
rect 3180 53375 3236 53404
rect 3304 53375 3360 53404
rect 3428 53375 3484 53404
rect 3552 53375 3608 53404
rect 3676 53375 3732 53404
rect 2808 53348 2815 53375
rect 2815 53348 2864 53375
rect 2932 53348 2979 53375
rect 2979 53348 2988 53375
rect 3056 53348 3087 53375
rect 3087 53348 3112 53375
rect 3180 53348 3195 53375
rect 3195 53348 3236 53375
rect 3304 53348 3355 53375
rect 3355 53348 3360 53375
rect 3428 53348 3463 53375
rect 3463 53348 3484 53375
rect 3552 53348 3571 53375
rect 3571 53348 3608 53375
rect 3676 53348 3679 53375
rect 3679 53348 3732 53375
rect 3800 53348 3856 53404
rect 3924 53367 3955 53404
rect 3955 53367 3980 53404
rect 4048 53367 4079 53404
rect 4079 53367 4104 53404
rect 4172 53367 4203 53404
rect 4203 53367 4228 53404
rect 3924 53348 3980 53367
rect 4048 53348 4104 53367
rect 4172 53348 4228 53367
rect 4296 53348 4352 53404
rect 4420 53348 4476 53404
rect 4544 53348 4600 53404
rect 4668 53348 4724 53404
rect 2808 53267 2864 53280
rect 2932 53267 2988 53280
rect 3056 53267 3112 53280
rect 3180 53267 3236 53280
rect 3304 53267 3360 53280
rect 3428 53267 3484 53280
rect 3552 53267 3608 53280
rect 3676 53267 3732 53280
rect 2808 53224 2815 53267
rect 2815 53224 2864 53267
rect 2932 53224 2979 53267
rect 2979 53224 2988 53267
rect 3056 53224 3087 53267
rect 3087 53224 3112 53267
rect 3180 53224 3195 53267
rect 3195 53224 3236 53267
rect 3304 53224 3355 53267
rect 3355 53224 3360 53267
rect 3428 53224 3463 53267
rect 3463 53224 3484 53267
rect 3552 53224 3571 53267
rect 3571 53224 3608 53267
rect 3676 53224 3679 53267
rect 3679 53224 3732 53267
rect 3800 53224 3856 53280
rect 3924 53243 3955 53280
rect 3955 53243 3980 53280
rect 4048 53243 4079 53280
rect 4079 53243 4104 53280
rect 4172 53243 4203 53280
rect 4203 53243 4228 53280
rect 3924 53224 3980 53243
rect 4048 53224 4104 53243
rect 4172 53224 4228 53243
rect 4296 53224 4352 53280
rect 4420 53224 4476 53280
rect 4544 53224 4600 53280
rect 4668 53224 4724 53280
rect 2808 53100 2864 53156
rect 2932 53100 2988 53156
rect 3056 53100 3112 53156
rect 3180 53100 3236 53156
rect 3304 53100 3360 53156
rect 3428 53100 3484 53156
rect 3552 53100 3608 53156
rect 3676 53100 3732 53156
rect 3800 53100 3856 53156
rect 3924 53100 3980 53156
rect 4048 53100 4104 53156
rect 4172 53100 4228 53156
rect 4296 53100 4352 53156
rect 4420 53100 4476 53156
rect 4544 53100 4600 53156
rect 4668 53100 4724 53156
rect 2808 52976 2864 53032
rect 2932 52976 2988 53032
rect 3056 52976 3112 53032
rect 3180 52976 3236 53032
rect 3304 52976 3360 53032
rect 3428 52976 3484 53032
rect 3552 52976 3608 53032
rect 3676 52976 3732 53032
rect 3800 52976 3856 53032
rect 3924 52976 3980 53032
rect 4048 52976 4104 53032
rect 4172 52976 4228 53032
rect 4296 52976 4352 53032
rect 4420 52976 4476 53032
rect 4544 52976 4600 53032
rect 4668 52976 4724 53032
rect 2808 52852 2864 52908
rect 2932 52852 2988 52908
rect 3056 52852 3112 52908
rect 3180 52852 3236 52908
rect 3304 52852 3360 52908
rect 3428 52852 3484 52908
rect 3552 52852 3608 52908
rect 3676 52852 3732 52908
rect 3800 52852 3856 52908
rect 3924 52852 3980 52908
rect 4048 52852 4104 52908
rect 4172 52852 4228 52908
rect 4296 52852 4352 52908
rect 4420 52852 4476 52908
rect 4544 52852 4600 52908
rect 4668 52852 4724 52908
rect 2808 52492 2864 52548
rect 2932 52492 2988 52548
rect 3056 52492 3112 52548
rect 3180 52492 3236 52548
rect 3304 52492 3360 52548
rect 3428 52492 3484 52548
rect 3552 52492 3608 52548
rect 3676 52492 3732 52548
rect 3800 52492 3856 52548
rect 3924 52492 3980 52548
rect 4048 52492 4104 52548
rect 4172 52492 4228 52548
rect 4296 52492 4352 52548
rect 4420 52492 4476 52548
rect 4544 52492 4600 52548
rect 4668 52492 4724 52548
rect 2808 52368 2864 52424
rect 2932 52368 2988 52424
rect 3056 52368 3112 52424
rect 3180 52368 3236 52424
rect 3304 52368 3360 52424
rect 3428 52368 3484 52424
rect 3552 52368 3608 52424
rect 3676 52368 3732 52424
rect 3800 52368 3856 52424
rect 3924 52368 3980 52424
rect 4048 52368 4104 52424
rect 4172 52368 4228 52424
rect 4296 52368 4352 52424
rect 4420 52368 4476 52424
rect 4544 52368 4600 52424
rect 4668 52368 4724 52424
rect 2808 52244 2864 52300
rect 2932 52244 2988 52300
rect 3056 52244 3112 52300
rect 3180 52244 3236 52300
rect 3304 52244 3360 52300
rect 3428 52244 3484 52300
rect 3552 52244 3608 52300
rect 3676 52244 3732 52300
rect 3800 52244 3856 52300
rect 3924 52244 3980 52300
rect 4048 52244 4104 52300
rect 4172 52244 4228 52300
rect 4296 52244 4352 52300
rect 4420 52244 4476 52300
rect 4544 52244 4600 52300
rect 4668 52244 4724 52300
rect 2808 52120 2864 52176
rect 2932 52120 2988 52176
rect 3056 52120 3112 52176
rect 3180 52120 3236 52176
rect 3304 52120 3360 52176
rect 3428 52120 3484 52176
rect 3552 52120 3608 52176
rect 3676 52120 3732 52176
rect 3800 52120 3856 52176
rect 3924 52120 3980 52176
rect 4048 52120 4104 52176
rect 4172 52120 4228 52176
rect 4296 52120 4352 52176
rect 4420 52120 4476 52176
rect 4544 52120 4600 52176
rect 4668 52120 4724 52176
rect 2808 51996 2864 52052
rect 2932 51996 2988 52052
rect 3056 51996 3112 52052
rect 3180 52009 3236 52052
rect 3304 52009 3360 52052
rect 3428 52009 3484 52052
rect 3552 52009 3608 52052
rect 3676 52009 3732 52052
rect 3800 52009 3856 52052
rect 3924 52009 3980 52052
rect 4048 52009 4104 52052
rect 4172 52009 4228 52052
rect 4296 52009 4352 52052
rect 4420 52009 4476 52052
rect 4544 52009 4600 52052
rect 4668 52009 4724 52052
rect 3180 51996 3213 52009
rect 3213 51996 3236 52009
rect 3304 51996 3321 52009
rect 3321 51996 3360 52009
rect 3428 51996 3429 52009
rect 3429 51996 3484 52009
rect 3552 51996 3593 52009
rect 3593 51996 3608 52009
rect 3676 51996 3701 52009
rect 3701 51996 3732 52009
rect 3800 51996 3809 52009
rect 3809 51996 3856 52009
rect 3924 51996 3969 52009
rect 3969 51996 3980 52009
rect 4048 51996 4077 52009
rect 4077 51996 4104 52009
rect 4172 51996 4185 52009
rect 4185 51996 4228 52009
rect 4296 51996 4349 52009
rect 4349 51996 4352 52009
rect 4420 51996 4457 52009
rect 4457 51996 4476 52009
rect 4544 51996 4565 52009
rect 4565 51996 4600 52009
rect 4668 51996 4673 52009
rect 4673 51996 4724 52009
rect 2808 51872 2864 51928
rect 2932 51872 2988 51928
rect 3056 51872 3112 51928
rect 3180 51901 3236 51928
rect 3304 51901 3360 51928
rect 3428 51901 3484 51928
rect 3552 51901 3608 51928
rect 3676 51901 3732 51928
rect 3800 51901 3856 51928
rect 3924 51901 3980 51928
rect 4048 51901 4104 51928
rect 4172 51901 4228 51928
rect 4296 51901 4352 51928
rect 4420 51901 4476 51928
rect 4544 51901 4600 51928
rect 4668 51901 4724 51928
rect 3180 51872 3213 51901
rect 3213 51872 3236 51901
rect 3304 51872 3321 51901
rect 3321 51872 3360 51901
rect 3428 51872 3429 51901
rect 3429 51872 3484 51901
rect 3552 51872 3593 51901
rect 3593 51872 3608 51901
rect 3676 51872 3701 51901
rect 3701 51872 3732 51901
rect 3800 51872 3809 51901
rect 3809 51872 3856 51901
rect 3924 51872 3969 51901
rect 3969 51872 3980 51901
rect 4048 51872 4077 51901
rect 4077 51872 4104 51901
rect 4172 51872 4185 51901
rect 4185 51872 4228 51901
rect 4296 51872 4349 51901
rect 4349 51872 4352 51901
rect 4420 51872 4457 51901
rect 4457 51872 4476 51901
rect 4544 51872 4565 51901
rect 4565 51872 4600 51901
rect 4668 51872 4673 51901
rect 4673 51872 4724 51901
rect 2808 51748 2864 51804
rect 2932 51748 2988 51804
rect 3056 51748 3112 51804
rect 3180 51748 3236 51804
rect 3304 51748 3360 51804
rect 3428 51748 3484 51804
rect 3552 51748 3608 51804
rect 3676 51748 3732 51804
rect 3800 51748 3856 51804
rect 3924 51748 3980 51804
rect 4048 51748 4104 51804
rect 4172 51748 4228 51804
rect 4296 51748 4352 51804
rect 4420 51748 4476 51804
rect 4544 51748 4600 51804
rect 4668 51748 4724 51804
rect 2808 51624 2864 51680
rect 2932 51624 2988 51680
rect 3056 51624 3112 51680
rect 3180 51624 3236 51680
rect 3304 51624 3360 51680
rect 3428 51624 3484 51680
rect 3552 51624 3608 51680
rect 3676 51624 3732 51680
rect 3800 51624 3856 51680
rect 3924 51624 3980 51680
rect 4048 51624 4104 51680
rect 4172 51624 4228 51680
rect 4296 51624 4352 51680
rect 4420 51624 4476 51680
rect 4544 51624 4600 51680
rect 4668 51624 4724 51680
rect 2808 51500 2864 51556
rect 2932 51500 2988 51556
rect 3056 51500 3112 51556
rect 3180 51500 3236 51556
rect 3304 51500 3360 51556
rect 3428 51500 3484 51556
rect 3552 51500 3608 51556
rect 3676 51500 3732 51556
rect 3800 51500 3856 51556
rect 3924 51500 3980 51556
rect 4048 51500 4104 51556
rect 4172 51500 4228 51556
rect 4296 51500 4352 51556
rect 4420 51500 4476 51556
rect 4544 51500 4600 51556
rect 4668 51500 4724 51556
rect 2808 51376 2864 51432
rect 2932 51376 2988 51432
rect 3056 51376 3112 51432
rect 3180 51376 3236 51432
rect 3304 51376 3360 51432
rect 3428 51376 3484 51432
rect 3552 51376 3608 51432
rect 3676 51376 3732 51432
rect 3800 51376 3856 51432
rect 3924 51376 3980 51432
rect 4048 51376 4104 51432
rect 4172 51376 4228 51432
rect 4296 51376 4352 51432
rect 4420 51376 4476 51432
rect 4544 51376 4600 51432
rect 4668 51376 4724 51432
rect 2808 51252 2864 51308
rect 2932 51252 2988 51308
rect 3056 51252 3112 51308
rect 3180 51252 3236 51308
rect 3304 51252 3360 51308
rect 3428 51252 3484 51308
rect 3552 51252 3608 51308
rect 3676 51252 3732 51308
rect 3800 51252 3856 51308
rect 3924 51252 3980 51308
rect 4048 51252 4104 51308
rect 4172 51252 4228 51308
rect 4296 51252 4352 51308
rect 4420 51252 4476 51308
rect 4544 51252 4600 51308
rect 4668 51252 4724 51308
rect 2808 49292 2864 49348
rect 2932 49292 2988 49348
rect 3056 49292 3112 49348
rect 3180 49338 3236 49348
rect 3304 49338 3360 49348
rect 3428 49338 3484 49348
rect 3552 49338 3608 49348
rect 3676 49338 3732 49348
rect 3800 49338 3856 49348
rect 3924 49338 3980 49348
rect 4048 49338 4104 49348
rect 4172 49338 4228 49348
rect 4296 49338 4352 49348
rect 4420 49338 4476 49348
rect 4544 49338 4600 49348
rect 4668 49338 4724 49348
rect 3180 49292 3213 49338
rect 3213 49292 3236 49338
rect 3304 49292 3321 49338
rect 3321 49292 3360 49338
rect 3428 49292 3429 49338
rect 3429 49292 3484 49338
rect 3552 49292 3593 49338
rect 3593 49292 3608 49338
rect 3676 49292 3701 49338
rect 3701 49292 3732 49338
rect 3800 49292 3809 49338
rect 3809 49292 3856 49338
rect 3924 49292 3969 49338
rect 3969 49292 3980 49338
rect 4048 49292 4077 49338
rect 4077 49292 4104 49338
rect 4172 49292 4185 49338
rect 4185 49292 4228 49338
rect 4296 49292 4349 49338
rect 4349 49292 4352 49338
rect 4420 49292 4457 49338
rect 4457 49292 4476 49338
rect 4544 49292 4565 49338
rect 4565 49292 4600 49338
rect 4668 49292 4673 49338
rect 4673 49292 4724 49338
rect 2808 49168 2864 49224
rect 2932 49168 2988 49224
rect 3056 49168 3112 49224
rect 3180 49178 3213 49224
rect 3213 49178 3236 49224
rect 3304 49178 3321 49224
rect 3321 49178 3360 49224
rect 3428 49178 3429 49224
rect 3429 49178 3484 49224
rect 3552 49178 3593 49224
rect 3593 49178 3608 49224
rect 3676 49178 3701 49224
rect 3701 49178 3732 49224
rect 3800 49178 3809 49224
rect 3809 49178 3856 49224
rect 3924 49178 3969 49224
rect 3969 49178 3980 49224
rect 4048 49178 4077 49224
rect 4077 49178 4104 49224
rect 4172 49178 4185 49224
rect 4185 49178 4228 49224
rect 4296 49178 4349 49224
rect 4349 49178 4352 49224
rect 4420 49178 4457 49224
rect 4457 49178 4476 49224
rect 4544 49178 4565 49224
rect 4565 49178 4600 49224
rect 4668 49178 4673 49224
rect 4673 49178 4724 49224
rect 3180 49168 3236 49178
rect 3304 49168 3360 49178
rect 3428 49168 3484 49178
rect 3552 49168 3608 49178
rect 3676 49168 3732 49178
rect 3800 49168 3856 49178
rect 3924 49168 3980 49178
rect 4048 49168 4104 49178
rect 4172 49168 4228 49178
rect 4296 49168 4352 49178
rect 4420 49168 4476 49178
rect 4544 49168 4600 49178
rect 4668 49168 4724 49178
rect 2808 49044 2864 49100
rect 2932 49044 2988 49100
rect 3056 49044 3112 49100
rect 3180 49070 3213 49100
rect 3213 49070 3236 49100
rect 3304 49070 3321 49100
rect 3321 49070 3360 49100
rect 3428 49070 3429 49100
rect 3429 49070 3484 49100
rect 3552 49070 3593 49100
rect 3593 49070 3608 49100
rect 3676 49070 3701 49100
rect 3701 49070 3732 49100
rect 3800 49070 3809 49100
rect 3809 49070 3856 49100
rect 3924 49070 3969 49100
rect 3969 49070 3980 49100
rect 4048 49070 4077 49100
rect 4077 49070 4104 49100
rect 4172 49070 4185 49100
rect 4185 49070 4228 49100
rect 4296 49070 4349 49100
rect 4349 49070 4352 49100
rect 4420 49070 4457 49100
rect 4457 49070 4476 49100
rect 4544 49070 4565 49100
rect 4565 49070 4600 49100
rect 4668 49070 4673 49100
rect 4673 49070 4724 49100
rect 3180 49044 3236 49070
rect 3304 49044 3360 49070
rect 3428 49044 3484 49070
rect 3552 49044 3608 49070
rect 3676 49044 3732 49070
rect 3800 49044 3856 49070
rect 3924 49044 3980 49070
rect 4048 49044 4104 49070
rect 4172 49044 4228 49070
rect 4296 49044 4352 49070
rect 4420 49044 4476 49070
rect 4544 49044 4600 49070
rect 4668 49044 4724 49070
rect 2808 48920 2864 48976
rect 2932 48920 2988 48976
rect 3056 48920 3112 48976
rect 3180 48920 3236 48976
rect 3304 48920 3360 48976
rect 3428 48920 3484 48976
rect 3552 48920 3608 48976
rect 3676 48920 3732 48976
rect 3800 48920 3856 48976
rect 3924 48920 3980 48976
rect 4048 48920 4104 48976
rect 4172 48920 4228 48976
rect 4296 48920 4352 48976
rect 4420 48920 4476 48976
rect 4544 48920 4600 48976
rect 4668 48920 4724 48976
rect 2808 48796 2864 48852
rect 2932 48796 2988 48852
rect 3056 48796 3112 48852
rect 3180 48796 3236 48852
rect 3304 48796 3360 48852
rect 3428 48796 3484 48852
rect 3552 48796 3608 48852
rect 3676 48796 3732 48852
rect 3800 48796 3856 48852
rect 3924 48796 3980 48852
rect 4048 48796 4104 48852
rect 4172 48796 4228 48852
rect 4296 48796 4352 48852
rect 4420 48796 4476 48852
rect 4544 48796 4600 48852
rect 4668 48796 4724 48852
rect 2808 48672 2864 48728
rect 2932 48672 2988 48728
rect 3056 48672 3112 48728
rect 3180 48672 3236 48728
rect 3304 48672 3360 48728
rect 3428 48672 3484 48728
rect 3552 48672 3608 48728
rect 3676 48672 3732 48728
rect 3800 48672 3856 48728
rect 3924 48672 3980 48728
rect 4048 48672 4104 48728
rect 4172 48672 4228 48728
rect 4296 48672 4352 48728
rect 4420 48672 4476 48728
rect 4544 48672 4600 48728
rect 4668 48672 4724 48728
rect 2808 48548 2864 48604
rect 2932 48548 2988 48604
rect 3056 48548 3112 48604
rect 3180 48548 3236 48604
rect 3304 48548 3360 48604
rect 3428 48548 3484 48604
rect 3552 48548 3608 48604
rect 3676 48548 3732 48604
rect 3800 48548 3856 48604
rect 3924 48548 3980 48604
rect 4048 48548 4104 48604
rect 4172 48548 4228 48604
rect 4296 48548 4352 48604
rect 4420 48548 4476 48604
rect 4544 48548 4600 48604
rect 4668 48548 4724 48604
rect 2808 48424 2864 48480
rect 2932 48424 2988 48480
rect 3056 48424 3112 48480
rect 3180 48427 3236 48480
rect 3304 48427 3360 48480
rect 3428 48427 3484 48480
rect 3552 48427 3608 48480
rect 3676 48427 3732 48480
rect 3800 48427 3856 48480
rect 3924 48427 3980 48480
rect 4048 48427 4104 48480
rect 4172 48427 4228 48480
rect 4296 48427 4352 48480
rect 4420 48427 4476 48480
rect 4544 48427 4600 48480
rect 4668 48427 4724 48480
rect 3180 48424 3213 48427
rect 3213 48424 3236 48427
rect 3304 48424 3321 48427
rect 3321 48424 3360 48427
rect 3428 48424 3429 48427
rect 3429 48424 3484 48427
rect 3552 48424 3593 48427
rect 3593 48424 3608 48427
rect 3676 48424 3701 48427
rect 3701 48424 3732 48427
rect 3800 48424 3809 48427
rect 3809 48424 3856 48427
rect 3924 48424 3969 48427
rect 3969 48424 3980 48427
rect 4048 48424 4077 48427
rect 4077 48424 4104 48427
rect 4172 48424 4185 48427
rect 4185 48424 4228 48427
rect 4296 48424 4349 48427
rect 4349 48424 4352 48427
rect 4420 48424 4457 48427
rect 4457 48424 4476 48427
rect 4544 48424 4565 48427
rect 4565 48424 4600 48427
rect 4668 48424 4673 48427
rect 4673 48424 4724 48427
rect 2808 48300 2864 48356
rect 2932 48300 2988 48356
rect 3056 48300 3112 48356
rect 3180 48319 3236 48356
rect 3304 48319 3360 48356
rect 3428 48319 3484 48356
rect 3552 48319 3608 48356
rect 3676 48319 3732 48356
rect 3800 48319 3856 48356
rect 3924 48319 3980 48356
rect 4048 48319 4104 48356
rect 4172 48319 4228 48356
rect 4296 48319 4352 48356
rect 4420 48319 4476 48356
rect 4544 48319 4600 48356
rect 4668 48319 4724 48356
rect 3180 48300 3213 48319
rect 3213 48300 3236 48319
rect 3304 48300 3321 48319
rect 3321 48300 3360 48319
rect 3428 48300 3429 48319
rect 3429 48300 3484 48319
rect 3552 48300 3593 48319
rect 3593 48300 3608 48319
rect 3676 48300 3701 48319
rect 3701 48300 3732 48319
rect 3800 48300 3809 48319
rect 3809 48300 3856 48319
rect 3924 48300 3969 48319
rect 3969 48300 3980 48319
rect 4048 48300 4077 48319
rect 4077 48300 4104 48319
rect 4172 48300 4185 48319
rect 4185 48300 4228 48319
rect 4296 48300 4349 48319
rect 4349 48300 4352 48319
rect 4420 48300 4457 48319
rect 4457 48300 4476 48319
rect 4544 48300 4565 48319
rect 4565 48300 4600 48319
rect 4668 48300 4673 48319
rect 4673 48300 4724 48319
rect 2808 48176 2864 48232
rect 2932 48176 2988 48232
rect 3056 48176 3112 48232
rect 3180 48176 3236 48232
rect 3304 48176 3360 48232
rect 3428 48176 3484 48232
rect 3552 48176 3608 48232
rect 3676 48176 3732 48232
rect 3800 48176 3856 48232
rect 3924 48176 3980 48232
rect 4048 48176 4104 48232
rect 4172 48176 4228 48232
rect 4296 48176 4352 48232
rect 4420 48176 4476 48232
rect 4544 48176 4600 48232
rect 4668 48176 4724 48232
rect 2808 48052 2864 48108
rect 2932 48052 2988 48108
rect 3056 48052 3112 48108
rect 3180 48052 3236 48108
rect 3304 48052 3360 48108
rect 3428 48052 3484 48108
rect 3552 48052 3608 48108
rect 3676 48052 3732 48108
rect 3800 48052 3856 48108
rect 3924 48052 3980 48108
rect 4048 48052 4104 48108
rect 4172 48052 4228 48108
rect 4296 48052 4352 48108
rect 4420 48052 4476 48108
rect 4544 48052 4600 48108
rect 4668 48052 4724 48108
rect 4861 55721 4917 55748
rect 4985 55721 5041 55748
rect 4861 55692 4871 55721
rect 4871 55692 4917 55721
rect 4985 55692 5031 55721
rect 5031 55692 5041 55721
rect 4861 55613 4917 55624
rect 4985 55613 5041 55624
rect 4861 55568 4871 55613
rect 4871 55568 4917 55613
rect 4985 55568 5031 55613
rect 5031 55568 5041 55613
rect 4861 55453 4871 55500
rect 4871 55453 4917 55500
rect 4985 55453 5031 55500
rect 5031 55453 5041 55500
rect 4861 55444 4917 55453
rect 4985 55444 5041 55453
rect 4861 55345 4871 55376
rect 4871 55345 4917 55376
rect 4985 55345 5031 55376
rect 5031 55345 5041 55376
rect 4861 55320 4917 55345
rect 4985 55320 5041 55345
rect 4861 55237 4871 55252
rect 4871 55237 4917 55252
rect 4985 55237 5031 55252
rect 5031 55237 5041 55252
rect 4861 55196 4917 55237
rect 4985 55196 5041 55237
rect 4861 55073 4917 55128
rect 4985 55073 5041 55128
rect 4861 55072 4871 55073
rect 4871 55072 4917 55073
rect 4985 55072 5031 55073
rect 5031 55072 5041 55073
rect 4861 54965 4917 55004
rect 4985 54965 5041 55004
rect 4861 54948 4871 54965
rect 4871 54948 4917 54965
rect 4985 54948 5031 54965
rect 5031 54948 5041 54965
rect 4861 54857 4917 54880
rect 4985 54857 5041 54880
rect 4861 54824 4871 54857
rect 4871 54824 4917 54857
rect 4985 54824 5031 54857
rect 5031 54824 5041 54857
rect 4861 54749 4917 54756
rect 4985 54749 5041 54756
rect 4861 54700 4871 54749
rect 4871 54700 4917 54749
rect 4985 54700 5031 54749
rect 5031 54700 5041 54749
rect 4861 54589 4871 54632
rect 4871 54589 4917 54632
rect 4985 54589 5031 54632
rect 5031 54589 5041 54632
rect 4861 54576 4917 54589
rect 4985 54576 5041 54589
rect 4861 54481 4871 54508
rect 4871 54481 4917 54508
rect 4985 54481 5031 54508
rect 5031 54481 5041 54508
rect 4861 54452 4917 54481
rect 4985 54452 5041 54481
rect 4861 47704 4871 47748
rect 4871 47704 4917 47748
rect 4985 47704 5031 47748
rect 5031 47704 5041 47748
rect 4861 47692 4917 47704
rect 4985 47692 5041 47704
rect 4861 47568 4917 47624
rect 4985 47568 5041 47624
rect 4861 47444 4917 47500
rect 4985 47444 5041 47500
rect 4861 47320 4917 47376
rect 4985 47320 5041 47376
rect 4861 47196 4917 47252
rect 4985 47196 5041 47252
rect 2491 47072 2547 47128
rect 2615 47072 2671 47128
rect 2491 46948 2547 47004
rect 2615 46948 2671 47004
rect 2491 46824 2547 46880
rect 2615 46824 2671 46880
rect 2491 46700 2547 46756
rect 2615 46700 2671 46756
rect 2491 46576 2547 46632
rect 2615 46576 2671 46632
rect 2491 46452 2547 46508
rect 2615 46452 2671 46508
rect 5178 57169 5234 57225
rect 5302 57169 5358 57225
rect 5426 57169 5482 57225
rect 5550 57169 5606 57225
rect 5674 57169 5730 57225
rect 5798 57169 5854 57225
rect 5922 57169 5978 57225
rect 6046 57169 6102 57225
rect 6170 57169 6226 57225
rect 6294 57169 6350 57225
rect 6418 57169 6474 57225
rect 6542 57169 6598 57225
rect 6666 57169 6722 57225
rect 6790 57169 6846 57225
rect 6914 57169 6970 57225
rect 7038 57169 7094 57225
rect 5178 57052 5190 57101
rect 5190 57052 5234 57101
rect 5302 57052 5354 57101
rect 5354 57052 5358 57101
rect 5426 57052 5462 57101
rect 5462 57052 5482 57101
rect 5550 57052 5570 57101
rect 5570 57052 5606 57101
rect 5674 57052 5678 57101
rect 5678 57052 5730 57101
rect 5798 57052 5838 57101
rect 5838 57052 5854 57101
rect 5922 57052 5946 57101
rect 5946 57052 5978 57101
rect 6046 57052 6054 57101
rect 6054 57052 6102 57101
rect 6170 57052 6218 57101
rect 6218 57052 6226 57101
rect 6294 57052 6326 57101
rect 6326 57052 6350 57101
rect 6418 57052 6434 57101
rect 6434 57052 6474 57101
rect 6542 57052 6594 57101
rect 6594 57052 6598 57101
rect 6666 57052 6702 57101
rect 6702 57052 6722 57101
rect 6790 57052 6810 57101
rect 6810 57052 6846 57101
rect 6914 57052 6918 57101
rect 6918 57052 6970 57101
rect 7038 57052 7082 57101
rect 7082 57052 7094 57101
rect 5178 57045 5234 57052
rect 5302 57045 5358 57052
rect 5426 57045 5482 57052
rect 5550 57045 5606 57052
rect 5674 57045 5730 57052
rect 5798 57045 5854 57052
rect 5922 57045 5978 57052
rect 6046 57045 6102 57052
rect 6170 57045 6226 57052
rect 6294 57045 6350 57052
rect 6418 57045 6474 57052
rect 6542 57045 6598 57052
rect 6666 57045 6722 57052
rect 6790 57045 6846 57052
rect 6914 57045 6970 57052
rect 7038 57045 7094 57052
rect 5178 56921 5234 56977
rect 5302 56921 5358 56977
rect 5426 56921 5482 56977
rect 5550 56921 5606 56977
rect 5674 56921 5730 56977
rect 5798 56921 5854 56977
rect 5922 56921 5978 56977
rect 6046 56921 6102 56977
rect 6170 56921 6226 56977
rect 6294 56921 6350 56977
rect 6418 56921 6474 56977
rect 6542 56921 6598 56977
rect 6666 56921 6722 56977
rect 6790 56921 6846 56977
rect 6914 56921 6970 56977
rect 7038 56921 7094 56977
rect 5178 56797 5234 56853
rect 5302 56797 5358 56853
rect 5426 56797 5482 56853
rect 5550 56797 5606 56853
rect 5674 56797 5730 56853
rect 5798 56797 5854 56853
rect 5922 56797 5978 56853
rect 6046 56797 6102 56853
rect 6170 56797 6226 56853
rect 6294 56797 6350 56853
rect 6418 56797 6474 56853
rect 6542 56797 6598 56853
rect 6666 56797 6722 56853
rect 6790 56797 6846 56853
rect 6914 56797 6970 56853
rect 7038 56797 7094 56853
rect 5178 56673 5234 56729
rect 5302 56673 5358 56729
rect 5426 56673 5482 56729
rect 5550 56673 5606 56729
rect 5674 56673 5730 56729
rect 5798 56673 5854 56729
rect 5922 56673 5978 56729
rect 6046 56673 6102 56729
rect 6170 56673 6226 56729
rect 6294 56673 6350 56729
rect 6418 56673 6474 56729
rect 6542 56673 6598 56729
rect 6666 56673 6722 56729
rect 6790 56673 6846 56729
rect 6914 56673 6970 56729
rect 7038 56673 7094 56729
rect 5178 56549 5234 56605
rect 5302 56549 5358 56605
rect 5426 56549 5482 56605
rect 5550 56549 5606 56605
rect 5674 56549 5730 56605
rect 5798 56549 5854 56605
rect 5922 56549 5978 56605
rect 6046 56549 6102 56605
rect 6170 56549 6226 56605
rect 6294 56549 6350 56605
rect 6418 56549 6474 56605
rect 6542 56549 6598 56605
rect 6666 56549 6722 56605
rect 6790 56549 6846 56605
rect 6914 56549 6970 56605
rect 7038 56549 7094 56605
rect 5178 56425 5234 56481
rect 5302 56425 5358 56481
rect 5426 56425 5482 56481
rect 5550 56425 5606 56481
rect 5674 56425 5730 56481
rect 5798 56425 5854 56481
rect 5922 56425 5978 56481
rect 6046 56425 6102 56481
rect 6170 56425 6226 56481
rect 6294 56425 6350 56481
rect 6418 56425 6474 56481
rect 6542 56425 6598 56481
rect 6666 56425 6722 56481
rect 6790 56425 6846 56481
rect 6914 56425 6970 56481
rect 7038 56425 7094 56481
rect 5178 56301 5234 56357
rect 5302 56301 5358 56357
rect 5426 56301 5482 56357
rect 5550 56301 5606 56357
rect 5674 56301 5730 56357
rect 5798 56301 5854 56357
rect 5922 56301 5978 56357
rect 6046 56301 6102 56357
rect 6170 56301 6226 56357
rect 6294 56301 6350 56357
rect 6418 56301 6474 56357
rect 6542 56301 6598 56357
rect 6666 56301 6722 56357
rect 6790 56301 6846 56357
rect 6914 56301 6970 56357
rect 7038 56301 7094 56357
rect 5178 56177 5234 56233
rect 5302 56177 5358 56233
rect 5426 56177 5482 56233
rect 5550 56177 5606 56233
rect 5674 56177 5730 56233
rect 5798 56177 5854 56233
rect 5922 56177 5978 56233
rect 6046 56177 6102 56233
rect 6170 56177 6226 56233
rect 6294 56177 6350 56233
rect 6418 56177 6474 56233
rect 6542 56177 6598 56233
rect 6666 56177 6722 56233
rect 6790 56177 6846 56233
rect 6914 56177 6970 56233
rect 7038 56177 7094 56233
rect 5178 56053 5234 56109
rect 5302 56053 5358 56109
rect 5426 56053 5482 56109
rect 5550 56053 5606 56109
rect 5674 56053 5730 56109
rect 5798 56053 5854 56109
rect 5922 56053 5978 56109
rect 6046 56053 6102 56109
rect 6170 56053 6226 56109
rect 6294 56053 6350 56109
rect 6418 56053 6474 56109
rect 6542 56053 6598 56109
rect 6666 56053 6722 56109
rect 6790 56053 6846 56109
rect 6914 56053 6970 56109
rect 7038 56053 7094 56109
rect 5178 54092 5234 54148
rect 5302 54092 5358 54148
rect 5426 54092 5482 54148
rect 5550 54092 5606 54148
rect 5674 54092 5730 54148
rect 5798 54092 5854 54148
rect 5922 54092 5978 54148
rect 6046 54092 6102 54148
rect 6170 54092 6226 54148
rect 6294 54092 6350 54148
rect 6418 54092 6474 54148
rect 6542 54092 6598 54148
rect 6666 54092 6722 54148
rect 6790 54092 6846 54148
rect 6914 54092 6970 54148
rect 7038 54092 7094 54148
rect 5178 53968 5234 54024
rect 5302 53968 5358 54024
rect 5426 53968 5482 54024
rect 5550 53968 5606 54024
rect 5674 53968 5730 54024
rect 5798 53968 5854 54024
rect 5922 53968 5978 54024
rect 6046 53968 6102 54024
rect 6170 53968 6226 54024
rect 6294 53968 6350 54024
rect 6418 53968 6474 54024
rect 6542 53968 6598 54024
rect 6666 53968 6722 54024
rect 6790 53968 6846 54024
rect 6914 53968 6970 54024
rect 7038 53968 7094 54024
rect 5178 53844 5234 53900
rect 5302 53844 5358 53900
rect 5426 53844 5482 53900
rect 5550 53844 5606 53900
rect 5674 53844 5730 53900
rect 5798 53844 5854 53900
rect 5922 53844 5978 53900
rect 6046 53844 6102 53900
rect 6170 53844 6226 53900
rect 6294 53844 6350 53900
rect 6418 53844 6474 53900
rect 6542 53844 6598 53900
rect 6666 53844 6722 53900
rect 6790 53844 6846 53900
rect 6914 53844 6970 53900
rect 7038 53844 7094 53900
rect 5178 53720 5234 53776
rect 5302 53720 5358 53776
rect 5426 53720 5482 53776
rect 5550 53720 5606 53776
rect 5674 53720 5730 53776
rect 5798 53720 5854 53776
rect 5922 53720 5978 53776
rect 6046 53720 6102 53776
rect 6170 53720 6226 53776
rect 6294 53720 6350 53776
rect 6418 53720 6474 53776
rect 6542 53720 6598 53776
rect 6666 53720 6722 53776
rect 6790 53720 6846 53776
rect 6914 53720 6970 53776
rect 7038 53720 7094 53776
rect 5178 53596 5234 53652
rect 5302 53596 5358 53652
rect 5426 53596 5482 53652
rect 5550 53596 5606 53652
rect 5674 53596 5730 53652
rect 5798 53596 5854 53652
rect 5922 53596 5978 53652
rect 6046 53596 6102 53652
rect 6170 53596 6226 53652
rect 6294 53596 6350 53652
rect 6418 53596 6474 53652
rect 6542 53596 6598 53652
rect 6666 53596 6722 53652
rect 6790 53596 6846 53652
rect 6914 53596 6970 53652
rect 7038 53596 7094 53652
rect 5178 53483 5234 53528
rect 5302 53483 5358 53528
rect 5426 53483 5482 53528
rect 5550 53483 5606 53528
rect 5674 53483 5730 53528
rect 5798 53483 5854 53528
rect 5922 53483 5978 53528
rect 6046 53483 6102 53528
rect 6170 53483 6226 53528
rect 6294 53483 6350 53528
rect 6418 53483 6474 53528
rect 6542 53483 6598 53528
rect 6666 53483 6722 53528
rect 6790 53483 6846 53528
rect 6914 53483 6970 53528
rect 7038 53483 7094 53528
rect 5178 53472 5190 53483
rect 5190 53472 5234 53483
rect 5302 53472 5354 53483
rect 5354 53472 5358 53483
rect 5426 53472 5462 53483
rect 5462 53472 5482 53483
rect 5550 53472 5570 53483
rect 5570 53472 5606 53483
rect 5674 53472 5678 53483
rect 5678 53472 5730 53483
rect 5798 53472 5838 53483
rect 5838 53472 5854 53483
rect 5922 53472 5946 53483
rect 5946 53472 5978 53483
rect 6046 53472 6054 53483
rect 6054 53472 6102 53483
rect 6170 53472 6218 53483
rect 6218 53472 6226 53483
rect 6294 53472 6326 53483
rect 6326 53472 6350 53483
rect 6418 53472 6434 53483
rect 6434 53472 6474 53483
rect 6542 53472 6594 53483
rect 6594 53472 6598 53483
rect 6666 53472 6702 53483
rect 6702 53472 6722 53483
rect 6790 53472 6810 53483
rect 6810 53472 6846 53483
rect 6914 53472 6918 53483
rect 6918 53472 6970 53483
rect 7038 53472 7082 53483
rect 7082 53472 7094 53483
rect 5178 53375 5234 53404
rect 5302 53375 5358 53404
rect 5426 53375 5482 53404
rect 5550 53375 5606 53404
rect 5674 53375 5730 53404
rect 5798 53375 5854 53404
rect 5922 53375 5978 53404
rect 6046 53375 6102 53404
rect 6170 53375 6226 53404
rect 6294 53375 6350 53404
rect 6418 53375 6474 53404
rect 6542 53375 6598 53404
rect 6666 53375 6722 53404
rect 6790 53375 6846 53404
rect 6914 53375 6970 53404
rect 7038 53375 7094 53404
rect 5178 53348 5190 53375
rect 5190 53348 5234 53375
rect 5302 53348 5354 53375
rect 5354 53348 5358 53375
rect 5426 53348 5462 53375
rect 5462 53348 5482 53375
rect 5550 53348 5570 53375
rect 5570 53348 5606 53375
rect 5674 53348 5678 53375
rect 5678 53348 5730 53375
rect 5798 53348 5838 53375
rect 5838 53348 5854 53375
rect 5922 53348 5946 53375
rect 5946 53348 5978 53375
rect 6046 53348 6054 53375
rect 6054 53348 6102 53375
rect 6170 53348 6218 53375
rect 6218 53348 6226 53375
rect 6294 53348 6326 53375
rect 6326 53348 6350 53375
rect 6418 53348 6434 53375
rect 6434 53348 6474 53375
rect 6542 53348 6594 53375
rect 6594 53348 6598 53375
rect 6666 53348 6702 53375
rect 6702 53348 6722 53375
rect 6790 53348 6810 53375
rect 6810 53348 6846 53375
rect 6914 53348 6918 53375
rect 6918 53348 6970 53375
rect 7038 53348 7082 53375
rect 7082 53348 7094 53375
rect 5178 53267 5234 53280
rect 5302 53267 5358 53280
rect 5426 53267 5482 53280
rect 5550 53267 5606 53280
rect 5674 53267 5730 53280
rect 5798 53267 5854 53280
rect 5922 53267 5978 53280
rect 6046 53267 6102 53280
rect 6170 53267 6226 53280
rect 6294 53267 6350 53280
rect 6418 53267 6474 53280
rect 6542 53267 6598 53280
rect 6666 53267 6722 53280
rect 6790 53267 6846 53280
rect 6914 53267 6970 53280
rect 7038 53267 7094 53280
rect 5178 53224 5190 53267
rect 5190 53224 5234 53267
rect 5302 53224 5354 53267
rect 5354 53224 5358 53267
rect 5426 53224 5462 53267
rect 5462 53224 5482 53267
rect 5550 53224 5570 53267
rect 5570 53224 5606 53267
rect 5674 53224 5678 53267
rect 5678 53224 5730 53267
rect 5798 53224 5838 53267
rect 5838 53224 5854 53267
rect 5922 53224 5946 53267
rect 5946 53224 5978 53267
rect 6046 53224 6054 53267
rect 6054 53224 6102 53267
rect 6170 53224 6218 53267
rect 6218 53224 6226 53267
rect 6294 53224 6326 53267
rect 6326 53224 6350 53267
rect 6418 53224 6434 53267
rect 6434 53224 6474 53267
rect 6542 53224 6594 53267
rect 6594 53224 6598 53267
rect 6666 53224 6702 53267
rect 6702 53224 6722 53267
rect 6790 53224 6810 53267
rect 6810 53224 6846 53267
rect 6914 53224 6918 53267
rect 6918 53224 6970 53267
rect 7038 53224 7082 53267
rect 7082 53224 7094 53267
rect 5178 53100 5234 53156
rect 5302 53100 5358 53156
rect 5426 53100 5482 53156
rect 5550 53100 5606 53156
rect 5674 53100 5730 53156
rect 5798 53100 5854 53156
rect 5922 53100 5978 53156
rect 6046 53100 6102 53156
rect 6170 53100 6226 53156
rect 6294 53100 6350 53156
rect 6418 53100 6474 53156
rect 6542 53100 6598 53156
rect 6666 53100 6722 53156
rect 6790 53100 6846 53156
rect 6914 53100 6970 53156
rect 7038 53100 7094 53156
rect 5178 52976 5234 53032
rect 5302 52976 5358 53032
rect 5426 52976 5482 53032
rect 5550 52976 5606 53032
rect 5674 52976 5730 53032
rect 5798 52976 5854 53032
rect 5922 52976 5978 53032
rect 6046 52976 6102 53032
rect 6170 52976 6226 53032
rect 6294 52976 6350 53032
rect 6418 52976 6474 53032
rect 6542 52976 6598 53032
rect 6666 52976 6722 53032
rect 6790 52976 6846 53032
rect 6914 52976 6970 53032
rect 7038 52976 7094 53032
rect 5178 52852 5234 52908
rect 5302 52852 5358 52908
rect 5426 52852 5482 52908
rect 5550 52852 5606 52908
rect 5674 52852 5730 52908
rect 5798 52852 5854 52908
rect 5922 52852 5978 52908
rect 6046 52852 6102 52908
rect 6170 52852 6226 52908
rect 6294 52852 6350 52908
rect 6418 52852 6474 52908
rect 6542 52852 6598 52908
rect 6666 52852 6722 52908
rect 6790 52852 6846 52908
rect 6914 52852 6970 52908
rect 7038 52852 7094 52908
rect 5178 52492 5234 52548
rect 5302 52492 5358 52548
rect 5426 52492 5482 52548
rect 5550 52492 5606 52548
rect 5674 52492 5730 52548
rect 5798 52492 5854 52548
rect 5922 52492 5978 52548
rect 6046 52492 6102 52548
rect 6170 52492 6226 52548
rect 6294 52492 6350 52548
rect 6418 52492 6474 52548
rect 6542 52492 6598 52548
rect 6666 52492 6722 52548
rect 6790 52492 6846 52548
rect 6914 52492 6970 52548
rect 7038 52492 7094 52548
rect 5178 52368 5234 52424
rect 5302 52368 5358 52424
rect 5426 52368 5482 52424
rect 5550 52368 5606 52424
rect 5674 52368 5730 52424
rect 5798 52368 5854 52424
rect 5922 52368 5978 52424
rect 6046 52368 6102 52424
rect 6170 52368 6226 52424
rect 6294 52368 6350 52424
rect 6418 52368 6474 52424
rect 6542 52368 6598 52424
rect 6666 52368 6722 52424
rect 6790 52368 6846 52424
rect 6914 52368 6970 52424
rect 7038 52368 7094 52424
rect 5178 52244 5234 52300
rect 5302 52244 5358 52300
rect 5426 52244 5482 52300
rect 5550 52244 5606 52300
rect 5674 52244 5730 52300
rect 5798 52244 5854 52300
rect 5922 52244 5978 52300
rect 6046 52244 6102 52300
rect 6170 52244 6226 52300
rect 6294 52244 6350 52300
rect 6418 52244 6474 52300
rect 6542 52244 6598 52300
rect 6666 52244 6722 52300
rect 6790 52244 6846 52300
rect 6914 52244 6970 52300
rect 7038 52244 7094 52300
rect 5178 52120 5234 52176
rect 5302 52120 5358 52176
rect 5426 52120 5482 52176
rect 5550 52120 5606 52176
rect 5674 52120 5730 52176
rect 5798 52120 5854 52176
rect 5922 52120 5978 52176
rect 6046 52120 6102 52176
rect 6170 52120 6226 52176
rect 6294 52120 6350 52176
rect 6418 52120 6474 52176
rect 6542 52120 6598 52176
rect 6666 52120 6722 52176
rect 6790 52120 6846 52176
rect 6914 52120 6970 52176
rect 7038 52120 7094 52176
rect 5178 52009 5234 52052
rect 5302 52009 5358 52052
rect 5426 52009 5482 52052
rect 5550 52009 5606 52052
rect 5674 52009 5730 52052
rect 5798 52009 5854 52052
rect 5922 52009 5978 52052
rect 6046 52009 6102 52052
rect 6170 52009 6226 52052
rect 6294 52009 6350 52052
rect 6418 52009 6474 52052
rect 6542 52009 6598 52052
rect 6666 52009 6722 52052
rect 6790 52009 6846 52052
rect 6914 52009 6970 52052
rect 7038 52009 7094 52052
rect 5178 51996 5190 52009
rect 5190 51996 5234 52009
rect 5302 51996 5354 52009
rect 5354 51996 5358 52009
rect 5426 51996 5462 52009
rect 5462 51996 5482 52009
rect 5550 51996 5570 52009
rect 5570 51996 5606 52009
rect 5674 51996 5678 52009
rect 5678 51996 5730 52009
rect 5798 51996 5838 52009
rect 5838 51996 5854 52009
rect 5922 51996 5946 52009
rect 5946 51996 5978 52009
rect 6046 51996 6054 52009
rect 6054 51996 6102 52009
rect 6170 51996 6218 52009
rect 6218 51996 6226 52009
rect 6294 51996 6326 52009
rect 6326 51996 6350 52009
rect 6418 51996 6434 52009
rect 6434 51996 6474 52009
rect 6542 51996 6594 52009
rect 6594 51996 6598 52009
rect 6666 51996 6702 52009
rect 6702 51996 6722 52009
rect 6790 51996 6810 52009
rect 6810 51996 6846 52009
rect 6914 51996 6918 52009
rect 6918 51996 6970 52009
rect 7038 51996 7082 52009
rect 7082 51996 7094 52009
rect 5178 51901 5234 51928
rect 5302 51901 5358 51928
rect 5426 51901 5482 51928
rect 5550 51901 5606 51928
rect 5674 51901 5730 51928
rect 5798 51901 5854 51928
rect 5922 51901 5978 51928
rect 6046 51901 6102 51928
rect 6170 51901 6226 51928
rect 6294 51901 6350 51928
rect 6418 51901 6474 51928
rect 6542 51901 6598 51928
rect 6666 51901 6722 51928
rect 6790 51901 6846 51928
rect 6914 51901 6970 51928
rect 7038 51901 7094 51928
rect 5178 51872 5190 51901
rect 5190 51872 5234 51901
rect 5302 51872 5354 51901
rect 5354 51872 5358 51901
rect 5426 51872 5462 51901
rect 5462 51872 5482 51901
rect 5550 51872 5570 51901
rect 5570 51872 5606 51901
rect 5674 51872 5678 51901
rect 5678 51872 5730 51901
rect 5798 51872 5838 51901
rect 5838 51872 5854 51901
rect 5922 51872 5946 51901
rect 5946 51872 5978 51901
rect 6046 51872 6054 51901
rect 6054 51872 6102 51901
rect 6170 51872 6218 51901
rect 6218 51872 6226 51901
rect 6294 51872 6326 51901
rect 6326 51872 6350 51901
rect 6418 51872 6434 51901
rect 6434 51872 6474 51901
rect 6542 51872 6594 51901
rect 6594 51872 6598 51901
rect 6666 51872 6702 51901
rect 6702 51872 6722 51901
rect 6790 51872 6810 51901
rect 6810 51872 6846 51901
rect 6914 51872 6918 51901
rect 6918 51872 6970 51901
rect 7038 51872 7082 51901
rect 7082 51872 7094 51901
rect 5178 51748 5234 51804
rect 5302 51748 5358 51804
rect 5426 51748 5482 51804
rect 5550 51748 5606 51804
rect 5674 51748 5730 51804
rect 5798 51748 5854 51804
rect 5922 51748 5978 51804
rect 6046 51748 6102 51804
rect 6170 51748 6226 51804
rect 6294 51748 6350 51804
rect 6418 51748 6474 51804
rect 6542 51748 6598 51804
rect 6666 51748 6722 51804
rect 6790 51748 6846 51804
rect 6914 51748 6970 51804
rect 7038 51748 7094 51804
rect 5178 51624 5234 51680
rect 5302 51624 5358 51680
rect 5426 51624 5482 51680
rect 5550 51624 5606 51680
rect 5674 51624 5730 51680
rect 5798 51624 5854 51680
rect 5922 51624 5978 51680
rect 6046 51624 6102 51680
rect 6170 51624 6226 51680
rect 6294 51624 6350 51680
rect 6418 51624 6474 51680
rect 6542 51624 6598 51680
rect 6666 51624 6722 51680
rect 6790 51624 6846 51680
rect 6914 51624 6970 51680
rect 7038 51624 7094 51680
rect 5178 51500 5234 51556
rect 5302 51500 5358 51556
rect 5426 51500 5482 51556
rect 5550 51500 5606 51556
rect 5674 51500 5730 51556
rect 5798 51500 5854 51556
rect 5922 51500 5978 51556
rect 6046 51500 6102 51556
rect 6170 51500 6226 51556
rect 6294 51500 6350 51556
rect 6418 51500 6474 51556
rect 6542 51500 6598 51556
rect 6666 51500 6722 51556
rect 6790 51500 6846 51556
rect 6914 51500 6970 51556
rect 7038 51500 7094 51556
rect 5178 51376 5234 51432
rect 5302 51376 5358 51432
rect 5426 51376 5482 51432
rect 5550 51376 5606 51432
rect 5674 51376 5730 51432
rect 5798 51376 5854 51432
rect 5922 51376 5978 51432
rect 6046 51376 6102 51432
rect 6170 51376 6226 51432
rect 6294 51376 6350 51432
rect 6418 51376 6474 51432
rect 6542 51376 6598 51432
rect 6666 51376 6722 51432
rect 6790 51376 6846 51432
rect 6914 51376 6970 51432
rect 7038 51376 7094 51432
rect 5178 51252 5234 51308
rect 5302 51252 5358 51308
rect 5426 51252 5482 51308
rect 5550 51252 5606 51308
rect 5674 51252 5730 51308
rect 5798 51252 5854 51308
rect 5922 51252 5978 51308
rect 6046 51252 6102 51308
rect 6170 51252 6226 51308
rect 6294 51252 6350 51308
rect 6418 51252 6474 51308
rect 6542 51252 6598 51308
rect 6666 51252 6722 51308
rect 6790 51252 6846 51308
rect 6914 51252 6970 51308
rect 7038 51252 7094 51308
rect 5178 49338 5234 49348
rect 5302 49338 5358 49348
rect 5426 49338 5482 49348
rect 5550 49338 5606 49348
rect 5674 49338 5730 49348
rect 5798 49338 5854 49348
rect 5922 49338 5978 49348
rect 6046 49338 6102 49348
rect 6170 49338 6226 49348
rect 6294 49338 6350 49348
rect 6418 49338 6474 49348
rect 6542 49338 6598 49348
rect 6666 49338 6722 49348
rect 6790 49338 6846 49348
rect 6914 49338 6970 49348
rect 7038 49338 7094 49348
rect 5178 49292 5190 49338
rect 5190 49292 5234 49338
rect 5302 49292 5354 49338
rect 5354 49292 5358 49338
rect 5426 49292 5462 49338
rect 5462 49292 5482 49338
rect 5550 49292 5570 49338
rect 5570 49292 5606 49338
rect 5674 49292 5678 49338
rect 5678 49292 5730 49338
rect 5798 49292 5838 49338
rect 5838 49292 5854 49338
rect 5922 49292 5946 49338
rect 5946 49292 5978 49338
rect 6046 49292 6054 49338
rect 6054 49292 6102 49338
rect 6170 49292 6218 49338
rect 6218 49292 6226 49338
rect 6294 49292 6326 49338
rect 6326 49292 6350 49338
rect 6418 49292 6434 49338
rect 6434 49292 6474 49338
rect 6542 49292 6594 49338
rect 6594 49292 6598 49338
rect 6666 49292 6702 49338
rect 6702 49292 6722 49338
rect 6790 49292 6810 49338
rect 6810 49292 6846 49338
rect 6914 49292 6918 49338
rect 6918 49292 6970 49338
rect 7038 49292 7082 49338
rect 7082 49292 7094 49338
rect 5178 49178 5190 49224
rect 5190 49178 5234 49224
rect 5302 49178 5354 49224
rect 5354 49178 5358 49224
rect 5426 49178 5462 49224
rect 5462 49178 5482 49224
rect 5550 49178 5570 49224
rect 5570 49178 5606 49224
rect 5674 49178 5678 49224
rect 5678 49178 5730 49224
rect 5798 49178 5838 49224
rect 5838 49178 5854 49224
rect 5922 49178 5946 49224
rect 5946 49178 5978 49224
rect 6046 49178 6054 49224
rect 6054 49178 6102 49224
rect 6170 49178 6218 49224
rect 6218 49178 6226 49224
rect 6294 49178 6326 49224
rect 6326 49178 6350 49224
rect 6418 49178 6434 49224
rect 6434 49178 6474 49224
rect 6542 49178 6594 49224
rect 6594 49178 6598 49224
rect 6666 49178 6702 49224
rect 6702 49178 6722 49224
rect 6790 49178 6810 49224
rect 6810 49178 6846 49224
rect 6914 49178 6918 49224
rect 6918 49178 6970 49224
rect 7038 49178 7082 49224
rect 7082 49178 7094 49224
rect 5178 49168 5234 49178
rect 5302 49168 5358 49178
rect 5426 49168 5482 49178
rect 5550 49168 5606 49178
rect 5674 49168 5730 49178
rect 5798 49168 5854 49178
rect 5922 49168 5978 49178
rect 6046 49168 6102 49178
rect 6170 49168 6226 49178
rect 6294 49168 6350 49178
rect 6418 49168 6474 49178
rect 6542 49168 6598 49178
rect 6666 49168 6722 49178
rect 6790 49168 6846 49178
rect 6914 49168 6970 49178
rect 7038 49168 7094 49178
rect 5178 49070 5190 49100
rect 5190 49070 5234 49100
rect 5302 49070 5354 49100
rect 5354 49070 5358 49100
rect 5426 49070 5462 49100
rect 5462 49070 5482 49100
rect 5550 49070 5570 49100
rect 5570 49070 5606 49100
rect 5674 49070 5678 49100
rect 5678 49070 5730 49100
rect 5798 49070 5838 49100
rect 5838 49070 5854 49100
rect 5922 49070 5946 49100
rect 5946 49070 5978 49100
rect 6046 49070 6054 49100
rect 6054 49070 6102 49100
rect 6170 49070 6218 49100
rect 6218 49070 6226 49100
rect 6294 49070 6326 49100
rect 6326 49070 6350 49100
rect 6418 49070 6434 49100
rect 6434 49070 6474 49100
rect 6542 49070 6594 49100
rect 6594 49070 6598 49100
rect 6666 49070 6702 49100
rect 6702 49070 6722 49100
rect 6790 49070 6810 49100
rect 6810 49070 6846 49100
rect 6914 49070 6918 49100
rect 6918 49070 6970 49100
rect 7038 49070 7082 49100
rect 7082 49070 7094 49100
rect 5178 49044 5234 49070
rect 5302 49044 5358 49070
rect 5426 49044 5482 49070
rect 5550 49044 5606 49070
rect 5674 49044 5730 49070
rect 5798 49044 5854 49070
rect 5922 49044 5978 49070
rect 6046 49044 6102 49070
rect 6170 49044 6226 49070
rect 6294 49044 6350 49070
rect 6418 49044 6474 49070
rect 6542 49044 6598 49070
rect 6666 49044 6722 49070
rect 6790 49044 6846 49070
rect 6914 49044 6970 49070
rect 7038 49044 7094 49070
rect 5178 48920 5234 48976
rect 5302 48920 5358 48976
rect 5426 48920 5482 48976
rect 5550 48920 5606 48976
rect 5674 48920 5730 48976
rect 5798 48920 5854 48976
rect 5922 48920 5978 48976
rect 6046 48920 6102 48976
rect 6170 48920 6226 48976
rect 6294 48920 6350 48976
rect 6418 48920 6474 48976
rect 6542 48920 6598 48976
rect 6666 48920 6722 48976
rect 6790 48920 6846 48976
rect 6914 48920 6970 48976
rect 7038 48920 7094 48976
rect 5178 48796 5234 48852
rect 5302 48796 5358 48852
rect 5426 48796 5482 48852
rect 5550 48796 5606 48852
rect 5674 48796 5730 48852
rect 5798 48796 5854 48852
rect 5922 48796 5978 48852
rect 6046 48796 6102 48852
rect 6170 48796 6226 48852
rect 6294 48796 6350 48852
rect 6418 48796 6474 48852
rect 6542 48796 6598 48852
rect 6666 48796 6722 48852
rect 6790 48796 6846 48852
rect 6914 48796 6970 48852
rect 7038 48796 7094 48852
rect 5178 48672 5234 48728
rect 5302 48672 5358 48728
rect 5426 48672 5482 48728
rect 5550 48672 5606 48728
rect 5674 48672 5730 48728
rect 5798 48672 5854 48728
rect 5922 48672 5978 48728
rect 6046 48672 6102 48728
rect 6170 48672 6226 48728
rect 6294 48672 6350 48728
rect 6418 48672 6474 48728
rect 6542 48672 6598 48728
rect 6666 48672 6722 48728
rect 6790 48672 6846 48728
rect 6914 48672 6970 48728
rect 7038 48672 7094 48728
rect 5178 48548 5234 48604
rect 5302 48548 5358 48604
rect 5426 48548 5482 48604
rect 5550 48548 5606 48604
rect 5674 48548 5730 48604
rect 5798 48548 5854 48604
rect 5922 48548 5978 48604
rect 6046 48548 6102 48604
rect 6170 48548 6226 48604
rect 6294 48548 6350 48604
rect 6418 48548 6474 48604
rect 6542 48548 6598 48604
rect 6666 48548 6722 48604
rect 6790 48548 6846 48604
rect 6914 48548 6970 48604
rect 7038 48548 7094 48604
rect 5178 48427 5234 48480
rect 5302 48427 5358 48480
rect 5426 48427 5482 48480
rect 5550 48427 5606 48480
rect 5674 48427 5730 48480
rect 5798 48427 5854 48480
rect 5922 48427 5978 48480
rect 6046 48427 6102 48480
rect 6170 48427 6226 48480
rect 6294 48427 6350 48480
rect 6418 48427 6474 48480
rect 6542 48427 6598 48480
rect 6666 48427 6722 48480
rect 6790 48427 6846 48480
rect 6914 48427 6970 48480
rect 7038 48427 7094 48480
rect 5178 48424 5190 48427
rect 5190 48424 5234 48427
rect 5302 48424 5354 48427
rect 5354 48424 5358 48427
rect 5426 48424 5462 48427
rect 5462 48424 5482 48427
rect 5550 48424 5570 48427
rect 5570 48424 5606 48427
rect 5674 48424 5678 48427
rect 5678 48424 5730 48427
rect 5798 48424 5838 48427
rect 5838 48424 5854 48427
rect 5922 48424 5946 48427
rect 5946 48424 5978 48427
rect 6046 48424 6054 48427
rect 6054 48424 6102 48427
rect 6170 48424 6218 48427
rect 6218 48424 6226 48427
rect 6294 48424 6326 48427
rect 6326 48424 6350 48427
rect 6418 48424 6434 48427
rect 6434 48424 6474 48427
rect 6542 48424 6594 48427
rect 6594 48424 6598 48427
rect 6666 48424 6702 48427
rect 6702 48424 6722 48427
rect 6790 48424 6810 48427
rect 6810 48424 6846 48427
rect 6914 48424 6918 48427
rect 6918 48424 6970 48427
rect 7038 48424 7082 48427
rect 7082 48424 7094 48427
rect 5178 48319 5234 48356
rect 5302 48319 5358 48356
rect 5426 48319 5482 48356
rect 5550 48319 5606 48356
rect 5674 48319 5730 48356
rect 5798 48319 5854 48356
rect 5922 48319 5978 48356
rect 6046 48319 6102 48356
rect 6170 48319 6226 48356
rect 6294 48319 6350 48356
rect 6418 48319 6474 48356
rect 6542 48319 6598 48356
rect 6666 48319 6722 48356
rect 6790 48319 6846 48356
rect 6914 48319 6970 48356
rect 7038 48319 7094 48356
rect 5178 48300 5190 48319
rect 5190 48300 5234 48319
rect 5302 48300 5354 48319
rect 5354 48300 5358 48319
rect 5426 48300 5462 48319
rect 5462 48300 5482 48319
rect 5550 48300 5570 48319
rect 5570 48300 5606 48319
rect 5674 48300 5678 48319
rect 5678 48300 5730 48319
rect 5798 48300 5838 48319
rect 5838 48300 5854 48319
rect 5922 48300 5946 48319
rect 5946 48300 5978 48319
rect 6046 48300 6054 48319
rect 6054 48300 6102 48319
rect 6170 48300 6218 48319
rect 6218 48300 6226 48319
rect 6294 48300 6326 48319
rect 6326 48300 6350 48319
rect 6418 48300 6434 48319
rect 6434 48300 6474 48319
rect 6542 48300 6594 48319
rect 6594 48300 6598 48319
rect 6666 48300 6702 48319
rect 6702 48300 6722 48319
rect 6790 48300 6810 48319
rect 6810 48300 6846 48319
rect 6914 48300 6918 48319
rect 6918 48300 6970 48319
rect 7038 48300 7082 48319
rect 7082 48300 7094 48319
rect 5178 48176 5234 48232
rect 5302 48176 5358 48232
rect 5426 48176 5482 48232
rect 5550 48176 5606 48232
rect 5674 48176 5730 48232
rect 5798 48176 5854 48232
rect 5922 48176 5978 48232
rect 6046 48176 6102 48232
rect 6170 48176 6226 48232
rect 6294 48176 6350 48232
rect 6418 48176 6474 48232
rect 6542 48176 6598 48232
rect 6666 48176 6722 48232
rect 6790 48176 6846 48232
rect 6914 48176 6970 48232
rect 7038 48176 7094 48232
rect 5178 48052 5234 48108
rect 5302 48052 5358 48108
rect 5426 48052 5482 48108
rect 5550 48052 5606 48108
rect 5674 48052 5730 48108
rect 5798 48052 5854 48108
rect 5922 48052 5978 48108
rect 6046 48052 6102 48108
rect 6170 48052 6226 48108
rect 6294 48052 6350 48108
rect 6418 48052 6474 48108
rect 6542 48052 6598 48108
rect 6666 48052 6722 48108
rect 6790 48052 6846 48108
rect 6914 48052 6970 48108
rect 7038 48052 7094 48108
rect 7275 55692 7331 55748
rect 7399 55692 7455 55748
rect 7523 55692 7579 55748
rect 7647 55692 7703 55748
rect 7275 55568 7331 55624
rect 7399 55568 7455 55624
rect 7523 55568 7579 55624
rect 7647 55568 7703 55624
rect 7275 55444 7331 55500
rect 7399 55444 7455 55500
rect 7523 55444 7579 55500
rect 7647 55444 7703 55500
rect 7275 55320 7331 55376
rect 7399 55320 7455 55376
rect 7523 55320 7579 55376
rect 7647 55320 7703 55376
rect 7275 55196 7331 55252
rect 7399 55196 7455 55252
rect 7523 55196 7579 55252
rect 7647 55196 7703 55252
rect 7275 55072 7331 55128
rect 7399 55072 7455 55128
rect 7523 55072 7579 55128
rect 7647 55072 7703 55128
rect 7275 54948 7331 55004
rect 7399 54948 7455 55004
rect 7523 54948 7579 55004
rect 7647 54948 7703 55004
rect 7275 54824 7331 54880
rect 7399 54824 7455 54880
rect 7523 54824 7579 54880
rect 7647 54824 7703 54880
rect 7275 54700 7331 54756
rect 7399 54700 7455 54756
rect 7523 54700 7579 54756
rect 7647 54700 7703 54756
rect 7275 54576 7331 54632
rect 7399 54576 7455 54632
rect 7523 54576 7579 54632
rect 7647 54576 7703 54632
rect 7275 54452 7331 54508
rect 7399 54452 7455 54508
rect 7523 54452 7579 54508
rect 7647 54452 7703 54508
rect 7275 47704 7299 47748
rect 7299 47704 7331 47748
rect 7399 47704 7407 47748
rect 7407 47704 7455 47748
rect 7523 47704 7571 47748
rect 7571 47704 7579 47748
rect 7647 47704 7679 47748
rect 7679 47704 7703 47748
rect 7275 47692 7331 47704
rect 7399 47692 7455 47704
rect 7523 47692 7579 47704
rect 7647 47692 7703 47704
rect 7275 47568 7331 47624
rect 7399 47568 7455 47624
rect 7523 47568 7579 47624
rect 7647 47568 7703 47624
rect 7275 47444 7331 47500
rect 7399 47444 7455 47500
rect 7523 47444 7579 47500
rect 7647 47444 7703 47500
rect 7275 47320 7331 47376
rect 7399 47320 7455 47376
rect 7523 47320 7579 47376
rect 7647 47320 7703 47376
rect 7275 47196 7331 47252
rect 7399 47196 7455 47252
rect 7523 47196 7579 47252
rect 7647 47196 7703 47252
rect 7884 57169 7940 57225
rect 8008 57169 8064 57225
rect 8132 57169 8188 57225
rect 8256 57169 8312 57225
rect 8380 57169 8436 57225
rect 8504 57169 8560 57225
rect 8628 57169 8684 57225
rect 8752 57169 8808 57225
rect 8876 57169 8932 57225
rect 9000 57169 9056 57225
rect 9124 57169 9180 57225
rect 9248 57169 9304 57225
rect 9372 57169 9428 57225
rect 9496 57169 9552 57225
rect 9620 57169 9676 57225
rect 9744 57169 9800 57225
rect 7884 57052 7896 57101
rect 7896 57052 7940 57101
rect 8008 57052 8060 57101
rect 8060 57052 8064 57101
rect 8132 57052 8168 57101
rect 8168 57052 8188 57101
rect 8256 57052 8276 57101
rect 8276 57052 8312 57101
rect 8380 57052 8384 57101
rect 8384 57052 8436 57101
rect 8504 57052 8544 57101
rect 8544 57052 8560 57101
rect 8628 57052 8652 57101
rect 8652 57052 8684 57101
rect 8752 57052 8760 57101
rect 8760 57052 8808 57101
rect 8876 57052 8924 57101
rect 8924 57052 8932 57101
rect 9000 57052 9032 57101
rect 9032 57052 9056 57101
rect 9124 57052 9140 57101
rect 9140 57052 9180 57101
rect 9248 57052 9300 57101
rect 9300 57052 9304 57101
rect 9372 57052 9408 57101
rect 9408 57052 9428 57101
rect 9496 57052 9516 57101
rect 9516 57052 9552 57101
rect 9620 57052 9624 57101
rect 9624 57052 9676 57101
rect 9744 57052 9788 57101
rect 9788 57052 9800 57101
rect 7884 57045 7940 57052
rect 8008 57045 8064 57052
rect 8132 57045 8188 57052
rect 8256 57045 8312 57052
rect 8380 57045 8436 57052
rect 8504 57045 8560 57052
rect 8628 57045 8684 57052
rect 8752 57045 8808 57052
rect 8876 57045 8932 57052
rect 9000 57045 9056 57052
rect 9124 57045 9180 57052
rect 9248 57045 9304 57052
rect 9372 57045 9428 57052
rect 9496 57045 9552 57052
rect 9620 57045 9676 57052
rect 9744 57045 9800 57052
rect 7884 56921 7940 56977
rect 8008 56921 8064 56977
rect 8132 56921 8188 56977
rect 8256 56921 8312 56977
rect 8380 56921 8436 56977
rect 8504 56921 8560 56977
rect 8628 56921 8684 56977
rect 8752 56921 8808 56977
rect 8876 56921 8932 56977
rect 9000 56921 9056 56977
rect 9124 56921 9180 56977
rect 9248 56921 9304 56977
rect 9372 56921 9428 56977
rect 9496 56921 9552 56977
rect 9620 56921 9676 56977
rect 9744 56921 9800 56977
rect 7884 56797 7940 56853
rect 8008 56797 8064 56853
rect 8132 56797 8188 56853
rect 8256 56797 8312 56853
rect 8380 56797 8436 56853
rect 8504 56797 8560 56853
rect 8628 56797 8684 56853
rect 8752 56797 8808 56853
rect 8876 56797 8932 56853
rect 9000 56797 9056 56853
rect 9124 56797 9180 56853
rect 9248 56797 9304 56853
rect 9372 56797 9428 56853
rect 9496 56797 9552 56853
rect 9620 56797 9676 56853
rect 9744 56797 9800 56853
rect 7884 56673 7940 56729
rect 8008 56673 8064 56729
rect 8132 56673 8188 56729
rect 8256 56673 8312 56729
rect 8380 56673 8436 56729
rect 8504 56673 8560 56729
rect 8628 56673 8684 56729
rect 8752 56673 8808 56729
rect 8876 56673 8932 56729
rect 9000 56673 9056 56729
rect 9124 56673 9180 56729
rect 9248 56673 9304 56729
rect 9372 56673 9428 56729
rect 9496 56673 9552 56729
rect 9620 56673 9676 56729
rect 9744 56673 9800 56729
rect 7884 56549 7940 56605
rect 8008 56549 8064 56605
rect 8132 56549 8188 56605
rect 8256 56549 8312 56605
rect 8380 56549 8436 56605
rect 8504 56549 8560 56605
rect 8628 56549 8684 56605
rect 8752 56549 8808 56605
rect 8876 56549 8932 56605
rect 9000 56549 9056 56605
rect 9124 56549 9180 56605
rect 9248 56549 9304 56605
rect 9372 56549 9428 56605
rect 9496 56549 9552 56605
rect 9620 56549 9676 56605
rect 9744 56549 9800 56605
rect 7884 56425 7940 56481
rect 8008 56425 8064 56481
rect 8132 56425 8188 56481
rect 8256 56425 8312 56481
rect 8380 56425 8436 56481
rect 8504 56425 8560 56481
rect 8628 56425 8684 56481
rect 8752 56425 8808 56481
rect 8876 56425 8932 56481
rect 9000 56425 9056 56481
rect 9124 56425 9180 56481
rect 9248 56425 9304 56481
rect 9372 56425 9428 56481
rect 9496 56425 9552 56481
rect 9620 56425 9676 56481
rect 9744 56425 9800 56481
rect 7884 56301 7940 56357
rect 8008 56301 8064 56357
rect 8132 56301 8188 56357
rect 8256 56301 8312 56357
rect 8380 56301 8436 56357
rect 8504 56301 8560 56357
rect 8628 56301 8684 56357
rect 8752 56301 8808 56357
rect 8876 56301 8932 56357
rect 9000 56301 9056 56357
rect 9124 56301 9180 56357
rect 9248 56301 9304 56357
rect 9372 56301 9428 56357
rect 9496 56301 9552 56357
rect 9620 56301 9676 56357
rect 9744 56301 9800 56357
rect 7884 56177 7940 56233
rect 8008 56177 8064 56233
rect 8132 56177 8188 56233
rect 8256 56177 8312 56233
rect 8380 56177 8436 56233
rect 8504 56177 8560 56233
rect 8628 56177 8684 56233
rect 8752 56177 8808 56233
rect 8876 56177 8932 56233
rect 9000 56177 9056 56233
rect 9124 56177 9180 56233
rect 9248 56177 9304 56233
rect 9372 56177 9428 56233
rect 9496 56177 9552 56233
rect 9620 56177 9676 56233
rect 9744 56177 9800 56233
rect 7884 56053 7940 56109
rect 8008 56053 8064 56109
rect 8132 56053 8188 56109
rect 8256 56053 8312 56109
rect 8380 56053 8436 56109
rect 8504 56053 8560 56109
rect 8628 56053 8684 56109
rect 8752 56053 8808 56109
rect 8876 56053 8932 56109
rect 9000 56053 9056 56109
rect 9124 56053 9180 56109
rect 9248 56053 9304 56109
rect 9372 56053 9428 56109
rect 9496 56053 9552 56109
rect 9620 56053 9676 56109
rect 9744 56053 9800 56109
rect 7884 54092 7940 54148
rect 8008 54092 8064 54148
rect 8132 54092 8188 54148
rect 8256 54092 8312 54148
rect 8380 54092 8436 54148
rect 8504 54092 8560 54148
rect 8628 54092 8684 54148
rect 8752 54092 8808 54148
rect 8876 54092 8932 54148
rect 9000 54092 9056 54148
rect 9124 54092 9180 54148
rect 9248 54092 9304 54148
rect 9372 54092 9428 54148
rect 9496 54092 9552 54148
rect 9620 54092 9676 54148
rect 9744 54092 9800 54148
rect 7884 53968 7940 54024
rect 8008 53968 8064 54024
rect 8132 53968 8188 54024
rect 8256 53968 8312 54024
rect 8380 53968 8436 54024
rect 8504 53968 8560 54024
rect 8628 53968 8684 54024
rect 8752 53968 8808 54024
rect 8876 53968 8932 54024
rect 9000 53968 9056 54024
rect 9124 53968 9180 54024
rect 9248 53968 9304 54024
rect 9372 53968 9428 54024
rect 9496 53968 9552 54024
rect 9620 53968 9676 54024
rect 9744 53968 9800 54024
rect 7884 53844 7940 53900
rect 8008 53844 8064 53900
rect 8132 53844 8188 53900
rect 8256 53844 8312 53900
rect 8380 53844 8436 53900
rect 8504 53844 8560 53900
rect 8628 53844 8684 53900
rect 8752 53844 8808 53900
rect 8876 53844 8932 53900
rect 9000 53844 9056 53900
rect 9124 53844 9180 53900
rect 9248 53844 9304 53900
rect 9372 53844 9428 53900
rect 9496 53844 9552 53900
rect 9620 53844 9676 53900
rect 9744 53844 9800 53900
rect 7884 53720 7940 53776
rect 8008 53720 8064 53776
rect 8132 53720 8188 53776
rect 8256 53720 8312 53776
rect 8380 53720 8436 53776
rect 8504 53720 8560 53776
rect 8628 53720 8684 53776
rect 8752 53720 8808 53776
rect 8876 53720 8932 53776
rect 9000 53720 9056 53776
rect 9124 53720 9180 53776
rect 9248 53720 9304 53776
rect 9372 53720 9428 53776
rect 9496 53720 9552 53776
rect 9620 53720 9676 53776
rect 9744 53720 9800 53776
rect 7884 53596 7940 53652
rect 8008 53596 8064 53652
rect 8132 53596 8188 53652
rect 8256 53596 8312 53652
rect 8380 53596 8436 53652
rect 8504 53596 8560 53652
rect 8628 53596 8684 53652
rect 8752 53596 8808 53652
rect 8876 53596 8932 53652
rect 9000 53596 9056 53652
rect 9124 53596 9180 53652
rect 9248 53596 9304 53652
rect 9372 53596 9428 53652
rect 9496 53596 9552 53652
rect 9620 53596 9676 53652
rect 9744 53596 9800 53652
rect 7884 53483 7940 53528
rect 8008 53483 8064 53528
rect 8132 53483 8188 53528
rect 8256 53483 8312 53528
rect 8380 53483 8436 53528
rect 8504 53483 8560 53528
rect 8628 53483 8684 53528
rect 8752 53483 8808 53528
rect 8876 53483 8932 53528
rect 9000 53483 9056 53528
rect 9124 53483 9180 53528
rect 9248 53483 9304 53528
rect 9372 53483 9428 53528
rect 9496 53483 9552 53528
rect 9620 53483 9676 53528
rect 9744 53483 9800 53528
rect 7884 53472 7896 53483
rect 7896 53472 7940 53483
rect 8008 53472 8060 53483
rect 8060 53472 8064 53483
rect 8132 53472 8168 53483
rect 8168 53472 8188 53483
rect 8256 53472 8276 53483
rect 8276 53472 8312 53483
rect 8380 53472 8384 53483
rect 8384 53472 8436 53483
rect 8504 53472 8544 53483
rect 8544 53472 8560 53483
rect 8628 53472 8652 53483
rect 8652 53472 8684 53483
rect 8752 53472 8760 53483
rect 8760 53472 8808 53483
rect 8876 53472 8924 53483
rect 8924 53472 8932 53483
rect 9000 53472 9032 53483
rect 9032 53472 9056 53483
rect 9124 53472 9140 53483
rect 9140 53472 9180 53483
rect 9248 53472 9300 53483
rect 9300 53472 9304 53483
rect 9372 53472 9408 53483
rect 9408 53472 9428 53483
rect 9496 53472 9516 53483
rect 9516 53472 9552 53483
rect 9620 53472 9624 53483
rect 9624 53472 9676 53483
rect 9744 53472 9788 53483
rect 9788 53472 9800 53483
rect 7884 53375 7940 53404
rect 8008 53375 8064 53404
rect 8132 53375 8188 53404
rect 8256 53375 8312 53404
rect 8380 53375 8436 53404
rect 8504 53375 8560 53404
rect 8628 53375 8684 53404
rect 8752 53375 8808 53404
rect 8876 53375 8932 53404
rect 9000 53375 9056 53404
rect 9124 53375 9180 53404
rect 9248 53375 9304 53404
rect 9372 53375 9428 53404
rect 9496 53375 9552 53404
rect 9620 53375 9676 53404
rect 9744 53375 9800 53404
rect 7884 53348 7896 53375
rect 7896 53348 7940 53375
rect 8008 53348 8060 53375
rect 8060 53348 8064 53375
rect 8132 53348 8168 53375
rect 8168 53348 8188 53375
rect 8256 53348 8276 53375
rect 8276 53348 8312 53375
rect 8380 53348 8384 53375
rect 8384 53348 8436 53375
rect 8504 53348 8544 53375
rect 8544 53348 8560 53375
rect 8628 53348 8652 53375
rect 8652 53348 8684 53375
rect 8752 53348 8760 53375
rect 8760 53348 8808 53375
rect 8876 53348 8924 53375
rect 8924 53348 8932 53375
rect 9000 53348 9032 53375
rect 9032 53348 9056 53375
rect 9124 53348 9140 53375
rect 9140 53348 9180 53375
rect 9248 53348 9300 53375
rect 9300 53348 9304 53375
rect 9372 53348 9408 53375
rect 9408 53348 9428 53375
rect 9496 53348 9516 53375
rect 9516 53348 9552 53375
rect 9620 53348 9624 53375
rect 9624 53348 9676 53375
rect 9744 53348 9788 53375
rect 9788 53348 9800 53375
rect 7884 53267 7940 53280
rect 8008 53267 8064 53280
rect 8132 53267 8188 53280
rect 8256 53267 8312 53280
rect 8380 53267 8436 53280
rect 8504 53267 8560 53280
rect 8628 53267 8684 53280
rect 8752 53267 8808 53280
rect 8876 53267 8932 53280
rect 9000 53267 9056 53280
rect 9124 53267 9180 53280
rect 9248 53267 9304 53280
rect 9372 53267 9428 53280
rect 9496 53267 9552 53280
rect 9620 53267 9676 53280
rect 9744 53267 9800 53280
rect 7884 53224 7896 53267
rect 7896 53224 7940 53267
rect 8008 53224 8060 53267
rect 8060 53224 8064 53267
rect 8132 53224 8168 53267
rect 8168 53224 8188 53267
rect 8256 53224 8276 53267
rect 8276 53224 8312 53267
rect 8380 53224 8384 53267
rect 8384 53224 8436 53267
rect 8504 53224 8544 53267
rect 8544 53224 8560 53267
rect 8628 53224 8652 53267
rect 8652 53224 8684 53267
rect 8752 53224 8760 53267
rect 8760 53224 8808 53267
rect 8876 53224 8924 53267
rect 8924 53224 8932 53267
rect 9000 53224 9032 53267
rect 9032 53224 9056 53267
rect 9124 53224 9140 53267
rect 9140 53224 9180 53267
rect 9248 53224 9300 53267
rect 9300 53224 9304 53267
rect 9372 53224 9408 53267
rect 9408 53224 9428 53267
rect 9496 53224 9516 53267
rect 9516 53224 9552 53267
rect 9620 53224 9624 53267
rect 9624 53224 9676 53267
rect 9744 53224 9788 53267
rect 9788 53224 9800 53267
rect 7884 53100 7940 53156
rect 8008 53100 8064 53156
rect 8132 53100 8188 53156
rect 8256 53100 8312 53156
rect 8380 53100 8436 53156
rect 8504 53100 8560 53156
rect 8628 53100 8684 53156
rect 8752 53100 8808 53156
rect 8876 53100 8932 53156
rect 9000 53100 9056 53156
rect 9124 53100 9180 53156
rect 9248 53100 9304 53156
rect 9372 53100 9428 53156
rect 9496 53100 9552 53156
rect 9620 53100 9676 53156
rect 9744 53100 9800 53156
rect 7884 52976 7940 53032
rect 8008 52976 8064 53032
rect 8132 52976 8188 53032
rect 8256 52976 8312 53032
rect 8380 52976 8436 53032
rect 8504 52976 8560 53032
rect 8628 52976 8684 53032
rect 8752 52976 8808 53032
rect 8876 52976 8932 53032
rect 9000 52976 9056 53032
rect 9124 52976 9180 53032
rect 9248 52976 9304 53032
rect 9372 52976 9428 53032
rect 9496 52976 9552 53032
rect 9620 52976 9676 53032
rect 9744 52976 9800 53032
rect 7884 52852 7940 52908
rect 8008 52852 8064 52908
rect 8132 52852 8188 52908
rect 8256 52852 8312 52908
rect 8380 52852 8436 52908
rect 8504 52852 8560 52908
rect 8628 52852 8684 52908
rect 8752 52852 8808 52908
rect 8876 52852 8932 52908
rect 9000 52852 9056 52908
rect 9124 52852 9180 52908
rect 9248 52852 9304 52908
rect 9372 52852 9428 52908
rect 9496 52852 9552 52908
rect 9620 52852 9676 52908
rect 9744 52852 9800 52908
rect 7884 52492 7940 52548
rect 8008 52492 8064 52548
rect 8132 52492 8188 52548
rect 8256 52492 8312 52548
rect 8380 52492 8436 52548
rect 8504 52492 8560 52548
rect 8628 52492 8684 52548
rect 8752 52492 8808 52548
rect 8876 52492 8932 52548
rect 9000 52492 9056 52548
rect 9124 52492 9180 52548
rect 9248 52492 9304 52548
rect 9372 52492 9428 52548
rect 9496 52492 9552 52548
rect 9620 52492 9676 52548
rect 9744 52492 9800 52548
rect 7884 52368 7940 52424
rect 8008 52368 8064 52424
rect 8132 52368 8188 52424
rect 8256 52368 8312 52424
rect 8380 52368 8436 52424
rect 8504 52368 8560 52424
rect 8628 52368 8684 52424
rect 8752 52368 8808 52424
rect 8876 52368 8932 52424
rect 9000 52368 9056 52424
rect 9124 52368 9180 52424
rect 9248 52368 9304 52424
rect 9372 52368 9428 52424
rect 9496 52368 9552 52424
rect 9620 52368 9676 52424
rect 9744 52368 9800 52424
rect 7884 52244 7940 52300
rect 8008 52244 8064 52300
rect 8132 52244 8188 52300
rect 8256 52244 8312 52300
rect 8380 52244 8436 52300
rect 8504 52244 8560 52300
rect 8628 52244 8684 52300
rect 8752 52244 8808 52300
rect 8876 52244 8932 52300
rect 9000 52244 9056 52300
rect 9124 52244 9180 52300
rect 9248 52244 9304 52300
rect 9372 52244 9428 52300
rect 9496 52244 9552 52300
rect 9620 52244 9676 52300
rect 9744 52244 9800 52300
rect 7884 52120 7940 52176
rect 8008 52120 8064 52176
rect 8132 52120 8188 52176
rect 8256 52120 8312 52176
rect 8380 52120 8436 52176
rect 8504 52120 8560 52176
rect 8628 52120 8684 52176
rect 8752 52120 8808 52176
rect 8876 52120 8932 52176
rect 9000 52120 9056 52176
rect 9124 52120 9180 52176
rect 9248 52120 9304 52176
rect 9372 52120 9428 52176
rect 9496 52120 9552 52176
rect 9620 52120 9676 52176
rect 9744 52120 9800 52176
rect 7884 52009 7940 52052
rect 8008 52009 8064 52052
rect 8132 52009 8188 52052
rect 8256 52009 8312 52052
rect 8380 52009 8436 52052
rect 8504 52009 8560 52052
rect 8628 52009 8684 52052
rect 8752 52009 8808 52052
rect 8876 52009 8932 52052
rect 9000 52009 9056 52052
rect 9124 52009 9180 52052
rect 9248 52009 9304 52052
rect 9372 52009 9428 52052
rect 9496 52009 9552 52052
rect 9620 52009 9676 52052
rect 9744 52009 9800 52052
rect 7884 51996 7896 52009
rect 7896 51996 7940 52009
rect 8008 51996 8060 52009
rect 8060 51996 8064 52009
rect 8132 51996 8168 52009
rect 8168 51996 8188 52009
rect 8256 51996 8276 52009
rect 8276 51996 8312 52009
rect 8380 51996 8384 52009
rect 8384 51996 8436 52009
rect 8504 51996 8544 52009
rect 8544 51996 8560 52009
rect 8628 51996 8652 52009
rect 8652 51996 8684 52009
rect 8752 51996 8760 52009
rect 8760 51996 8808 52009
rect 8876 51996 8924 52009
rect 8924 51996 8932 52009
rect 9000 51996 9032 52009
rect 9032 51996 9056 52009
rect 9124 51996 9140 52009
rect 9140 51996 9180 52009
rect 9248 51996 9300 52009
rect 9300 51996 9304 52009
rect 9372 51996 9408 52009
rect 9408 51996 9428 52009
rect 9496 51996 9516 52009
rect 9516 51996 9552 52009
rect 9620 51996 9624 52009
rect 9624 51996 9676 52009
rect 9744 51996 9788 52009
rect 9788 51996 9800 52009
rect 7884 51901 7940 51928
rect 8008 51901 8064 51928
rect 8132 51901 8188 51928
rect 8256 51901 8312 51928
rect 8380 51901 8436 51928
rect 8504 51901 8560 51928
rect 8628 51901 8684 51928
rect 8752 51901 8808 51928
rect 8876 51901 8932 51928
rect 9000 51901 9056 51928
rect 9124 51901 9180 51928
rect 9248 51901 9304 51928
rect 9372 51901 9428 51928
rect 9496 51901 9552 51928
rect 9620 51901 9676 51928
rect 9744 51901 9800 51928
rect 7884 51872 7896 51901
rect 7896 51872 7940 51901
rect 8008 51872 8060 51901
rect 8060 51872 8064 51901
rect 8132 51872 8168 51901
rect 8168 51872 8188 51901
rect 8256 51872 8276 51901
rect 8276 51872 8312 51901
rect 8380 51872 8384 51901
rect 8384 51872 8436 51901
rect 8504 51872 8544 51901
rect 8544 51872 8560 51901
rect 8628 51872 8652 51901
rect 8652 51872 8684 51901
rect 8752 51872 8760 51901
rect 8760 51872 8808 51901
rect 8876 51872 8924 51901
rect 8924 51872 8932 51901
rect 9000 51872 9032 51901
rect 9032 51872 9056 51901
rect 9124 51872 9140 51901
rect 9140 51872 9180 51901
rect 9248 51872 9300 51901
rect 9300 51872 9304 51901
rect 9372 51872 9408 51901
rect 9408 51872 9428 51901
rect 9496 51872 9516 51901
rect 9516 51872 9552 51901
rect 9620 51872 9624 51901
rect 9624 51872 9676 51901
rect 9744 51872 9788 51901
rect 9788 51872 9800 51901
rect 7884 51748 7940 51804
rect 8008 51748 8064 51804
rect 8132 51748 8188 51804
rect 8256 51748 8312 51804
rect 8380 51748 8436 51804
rect 8504 51748 8560 51804
rect 8628 51748 8684 51804
rect 8752 51748 8808 51804
rect 8876 51748 8932 51804
rect 9000 51748 9056 51804
rect 9124 51748 9180 51804
rect 9248 51748 9304 51804
rect 9372 51748 9428 51804
rect 9496 51748 9552 51804
rect 9620 51748 9676 51804
rect 9744 51748 9800 51804
rect 7884 51624 7940 51680
rect 8008 51624 8064 51680
rect 8132 51624 8188 51680
rect 8256 51624 8312 51680
rect 8380 51624 8436 51680
rect 8504 51624 8560 51680
rect 8628 51624 8684 51680
rect 8752 51624 8808 51680
rect 8876 51624 8932 51680
rect 9000 51624 9056 51680
rect 9124 51624 9180 51680
rect 9248 51624 9304 51680
rect 9372 51624 9428 51680
rect 9496 51624 9552 51680
rect 9620 51624 9676 51680
rect 9744 51624 9800 51680
rect 7884 51500 7940 51556
rect 8008 51500 8064 51556
rect 8132 51500 8188 51556
rect 8256 51500 8312 51556
rect 8380 51500 8436 51556
rect 8504 51500 8560 51556
rect 8628 51500 8684 51556
rect 8752 51500 8808 51556
rect 8876 51500 8932 51556
rect 9000 51500 9056 51556
rect 9124 51500 9180 51556
rect 9248 51500 9304 51556
rect 9372 51500 9428 51556
rect 9496 51500 9552 51556
rect 9620 51500 9676 51556
rect 9744 51500 9800 51556
rect 7884 51376 7940 51432
rect 8008 51376 8064 51432
rect 8132 51376 8188 51432
rect 8256 51376 8312 51432
rect 8380 51376 8436 51432
rect 8504 51376 8560 51432
rect 8628 51376 8684 51432
rect 8752 51376 8808 51432
rect 8876 51376 8932 51432
rect 9000 51376 9056 51432
rect 9124 51376 9180 51432
rect 9248 51376 9304 51432
rect 9372 51376 9428 51432
rect 9496 51376 9552 51432
rect 9620 51376 9676 51432
rect 9744 51376 9800 51432
rect 7884 51252 7940 51308
rect 8008 51252 8064 51308
rect 8132 51252 8188 51308
rect 8256 51252 8312 51308
rect 8380 51252 8436 51308
rect 8504 51252 8560 51308
rect 8628 51252 8684 51308
rect 8752 51252 8808 51308
rect 8876 51252 8932 51308
rect 9000 51252 9056 51308
rect 9124 51252 9180 51308
rect 9248 51252 9304 51308
rect 9372 51252 9428 51308
rect 9496 51252 9552 51308
rect 9620 51252 9676 51308
rect 9744 51252 9800 51308
rect 7884 49338 7940 49348
rect 8008 49338 8064 49348
rect 8132 49338 8188 49348
rect 8256 49338 8312 49348
rect 8380 49338 8436 49348
rect 8504 49338 8560 49348
rect 8628 49338 8684 49348
rect 8752 49338 8808 49348
rect 8876 49338 8932 49348
rect 9000 49338 9056 49348
rect 9124 49338 9180 49348
rect 9248 49338 9304 49348
rect 9372 49338 9428 49348
rect 9496 49338 9552 49348
rect 9620 49338 9676 49348
rect 9744 49338 9800 49348
rect 7884 49292 7896 49338
rect 7896 49292 7940 49338
rect 8008 49292 8060 49338
rect 8060 49292 8064 49338
rect 8132 49292 8168 49338
rect 8168 49292 8188 49338
rect 8256 49292 8276 49338
rect 8276 49292 8312 49338
rect 8380 49292 8384 49338
rect 8384 49292 8436 49338
rect 8504 49292 8544 49338
rect 8544 49292 8560 49338
rect 8628 49292 8652 49338
rect 8652 49292 8684 49338
rect 8752 49292 8760 49338
rect 8760 49292 8808 49338
rect 8876 49292 8924 49338
rect 8924 49292 8932 49338
rect 9000 49292 9032 49338
rect 9032 49292 9056 49338
rect 9124 49292 9140 49338
rect 9140 49292 9180 49338
rect 9248 49292 9300 49338
rect 9300 49292 9304 49338
rect 9372 49292 9408 49338
rect 9408 49292 9428 49338
rect 9496 49292 9516 49338
rect 9516 49292 9552 49338
rect 9620 49292 9624 49338
rect 9624 49292 9676 49338
rect 9744 49292 9788 49338
rect 9788 49292 9800 49338
rect 7884 49178 7896 49224
rect 7896 49178 7940 49224
rect 8008 49178 8060 49224
rect 8060 49178 8064 49224
rect 8132 49178 8168 49224
rect 8168 49178 8188 49224
rect 8256 49178 8276 49224
rect 8276 49178 8312 49224
rect 8380 49178 8384 49224
rect 8384 49178 8436 49224
rect 8504 49178 8544 49224
rect 8544 49178 8560 49224
rect 8628 49178 8652 49224
rect 8652 49178 8684 49224
rect 8752 49178 8760 49224
rect 8760 49178 8808 49224
rect 8876 49178 8924 49224
rect 8924 49178 8932 49224
rect 9000 49178 9032 49224
rect 9032 49178 9056 49224
rect 9124 49178 9140 49224
rect 9140 49178 9180 49224
rect 9248 49178 9300 49224
rect 9300 49178 9304 49224
rect 9372 49178 9408 49224
rect 9408 49178 9428 49224
rect 9496 49178 9516 49224
rect 9516 49178 9552 49224
rect 9620 49178 9624 49224
rect 9624 49178 9676 49224
rect 9744 49178 9788 49224
rect 9788 49178 9800 49224
rect 7884 49168 7940 49178
rect 8008 49168 8064 49178
rect 8132 49168 8188 49178
rect 8256 49168 8312 49178
rect 8380 49168 8436 49178
rect 8504 49168 8560 49178
rect 8628 49168 8684 49178
rect 8752 49168 8808 49178
rect 8876 49168 8932 49178
rect 9000 49168 9056 49178
rect 9124 49168 9180 49178
rect 9248 49168 9304 49178
rect 9372 49168 9428 49178
rect 9496 49168 9552 49178
rect 9620 49168 9676 49178
rect 9744 49168 9800 49178
rect 7884 49070 7896 49100
rect 7896 49070 7940 49100
rect 8008 49070 8060 49100
rect 8060 49070 8064 49100
rect 8132 49070 8168 49100
rect 8168 49070 8188 49100
rect 8256 49070 8276 49100
rect 8276 49070 8312 49100
rect 8380 49070 8384 49100
rect 8384 49070 8436 49100
rect 8504 49070 8544 49100
rect 8544 49070 8560 49100
rect 8628 49070 8652 49100
rect 8652 49070 8684 49100
rect 8752 49070 8760 49100
rect 8760 49070 8808 49100
rect 8876 49070 8924 49100
rect 8924 49070 8932 49100
rect 9000 49070 9032 49100
rect 9032 49070 9056 49100
rect 9124 49070 9140 49100
rect 9140 49070 9180 49100
rect 9248 49070 9300 49100
rect 9300 49070 9304 49100
rect 9372 49070 9408 49100
rect 9408 49070 9428 49100
rect 9496 49070 9516 49100
rect 9516 49070 9552 49100
rect 9620 49070 9624 49100
rect 9624 49070 9676 49100
rect 9744 49070 9788 49100
rect 9788 49070 9800 49100
rect 7884 49044 7940 49070
rect 8008 49044 8064 49070
rect 8132 49044 8188 49070
rect 8256 49044 8312 49070
rect 8380 49044 8436 49070
rect 8504 49044 8560 49070
rect 8628 49044 8684 49070
rect 8752 49044 8808 49070
rect 8876 49044 8932 49070
rect 9000 49044 9056 49070
rect 9124 49044 9180 49070
rect 9248 49044 9304 49070
rect 9372 49044 9428 49070
rect 9496 49044 9552 49070
rect 9620 49044 9676 49070
rect 9744 49044 9800 49070
rect 7884 48920 7940 48976
rect 8008 48920 8064 48976
rect 8132 48920 8188 48976
rect 8256 48920 8312 48976
rect 8380 48920 8436 48976
rect 8504 48920 8560 48976
rect 8628 48920 8684 48976
rect 8752 48920 8808 48976
rect 8876 48920 8932 48976
rect 9000 48920 9056 48976
rect 9124 48920 9180 48976
rect 9248 48920 9304 48976
rect 9372 48920 9428 48976
rect 9496 48920 9552 48976
rect 9620 48920 9676 48976
rect 9744 48920 9800 48976
rect 7884 48796 7940 48852
rect 8008 48796 8064 48852
rect 8132 48796 8188 48852
rect 8256 48796 8312 48852
rect 8380 48796 8436 48852
rect 8504 48796 8560 48852
rect 8628 48796 8684 48852
rect 8752 48796 8808 48852
rect 8876 48796 8932 48852
rect 9000 48796 9056 48852
rect 9124 48796 9180 48852
rect 9248 48796 9304 48852
rect 9372 48796 9428 48852
rect 9496 48796 9552 48852
rect 9620 48796 9676 48852
rect 9744 48796 9800 48852
rect 7884 48672 7940 48728
rect 8008 48672 8064 48728
rect 8132 48672 8188 48728
rect 8256 48672 8312 48728
rect 8380 48672 8436 48728
rect 8504 48672 8560 48728
rect 8628 48672 8684 48728
rect 8752 48672 8808 48728
rect 8876 48672 8932 48728
rect 9000 48672 9056 48728
rect 9124 48672 9180 48728
rect 9248 48672 9304 48728
rect 9372 48672 9428 48728
rect 9496 48672 9552 48728
rect 9620 48672 9676 48728
rect 9744 48672 9800 48728
rect 7884 48548 7940 48604
rect 8008 48548 8064 48604
rect 8132 48548 8188 48604
rect 8256 48548 8312 48604
rect 8380 48548 8436 48604
rect 8504 48548 8560 48604
rect 8628 48548 8684 48604
rect 8752 48548 8808 48604
rect 8876 48548 8932 48604
rect 9000 48548 9056 48604
rect 9124 48548 9180 48604
rect 9248 48548 9304 48604
rect 9372 48548 9428 48604
rect 9496 48548 9552 48604
rect 9620 48548 9676 48604
rect 9744 48548 9800 48604
rect 7884 48427 7940 48480
rect 8008 48427 8064 48480
rect 8132 48427 8188 48480
rect 8256 48427 8312 48480
rect 8380 48427 8436 48480
rect 8504 48427 8560 48480
rect 8628 48427 8684 48480
rect 8752 48427 8808 48480
rect 8876 48427 8932 48480
rect 9000 48427 9056 48480
rect 9124 48427 9180 48480
rect 9248 48427 9304 48480
rect 9372 48427 9428 48480
rect 9496 48427 9552 48480
rect 9620 48427 9676 48480
rect 9744 48427 9800 48480
rect 7884 48424 7896 48427
rect 7896 48424 7940 48427
rect 8008 48424 8060 48427
rect 8060 48424 8064 48427
rect 8132 48424 8168 48427
rect 8168 48424 8188 48427
rect 8256 48424 8276 48427
rect 8276 48424 8312 48427
rect 8380 48424 8384 48427
rect 8384 48424 8436 48427
rect 8504 48424 8544 48427
rect 8544 48424 8560 48427
rect 8628 48424 8652 48427
rect 8652 48424 8684 48427
rect 8752 48424 8760 48427
rect 8760 48424 8808 48427
rect 8876 48424 8924 48427
rect 8924 48424 8932 48427
rect 9000 48424 9032 48427
rect 9032 48424 9056 48427
rect 9124 48424 9140 48427
rect 9140 48424 9180 48427
rect 9248 48424 9300 48427
rect 9300 48424 9304 48427
rect 9372 48424 9408 48427
rect 9408 48424 9428 48427
rect 9496 48424 9516 48427
rect 9516 48424 9552 48427
rect 9620 48424 9624 48427
rect 9624 48424 9676 48427
rect 9744 48424 9788 48427
rect 9788 48424 9800 48427
rect 7884 48319 7940 48356
rect 8008 48319 8064 48356
rect 8132 48319 8188 48356
rect 8256 48319 8312 48356
rect 8380 48319 8436 48356
rect 8504 48319 8560 48356
rect 8628 48319 8684 48356
rect 8752 48319 8808 48356
rect 8876 48319 8932 48356
rect 9000 48319 9056 48356
rect 9124 48319 9180 48356
rect 9248 48319 9304 48356
rect 9372 48319 9428 48356
rect 9496 48319 9552 48356
rect 9620 48319 9676 48356
rect 9744 48319 9800 48356
rect 7884 48300 7896 48319
rect 7896 48300 7940 48319
rect 8008 48300 8060 48319
rect 8060 48300 8064 48319
rect 8132 48300 8168 48319
rect 8168 48300 8188 48319
rect 8256 48300 8276 48319
rect 8276 48300 8312 48319
rect 8380 48300 8384 48319
rect 8384 48300 8436 48319
rect 8504 48300 8544 48319
rect 8544 48300 8560 48319
rect 8628 48300 8652 48319
rect 8652 48300 8684 48319
rect 8752 48300 8760 48319
rect 8760 48300 8808 48319
rect 8876 48300 8924 48319
rect 8924 48300 8932 48319
rect 9000 48300 9032 48319
rect 9032 48300 9056 48319
rect 9124 48300 9140 48319
rect 9140 48300 9180 48319
rect 9248 48300 9300 48319
rect 9300 48300 9304 48319
rect 9372 48300 9408 48319
rect 9408 48300 9428 48319
rect 9496 48300 9516 48319
rect 9516 48300 9552 48319
rect 9620 48300 9624 48319
rect 9624 48300 9676 48319
rect 9744 48300 9788 48319
rect 9788 48300 9800 48319
rect 7884 48176 7940 48232
rect 8008 48176 8064 48232
rect 8132 48176 8188 48232
rect 8256 48176 8312 48232
rect 8380 48176 8436 48232
rect 8504 48176 8560 48232
rect 8628 48176 8684 48232
rect 8752 48176 8808 48232
rect 8876 48176 8932 48232
rect 9000 48176 9056 48232
rect 9124 48176 9180 48232
rect 9248 48176 9304 48232
rect 9372 48176 9428 48232
rect 9496 48176 9552 48232
rect 9620 48176 9676 48232
rect 9744 48176 9800 48232
rect 7884 48052 7940 48108
rect 8008 48052 8064 48108
rect 8132 48052 8188 48108
rect 8256 48052 8312 48108
rect 8380 48052 8436 48108
rect 8504 48052 8560 48108
rect 8628 48052 8684 48108
rect 8752 48052 8808 48108
rect 8876 48052 8932 48108
rect 9000 48052 9056 48108
rect 9124 48052 9180 48108
rect 9248 48052 9304 48108
rect 9372 48052 9428 48108
rect 9496 48052 9552 48108
rect 9620 48052 9676 48108
rect 9744 48052 9800 48108
rect 9937 55721 9993 55748
rect 10061 55721 10117 55748
rect 9937 55692 9947 55721
rect 9947 55692 9993 55721
rect 10061 55692 10107 55721
rect 10107 55692 10117 55721
rect 9937 55613 9993 55624
rect 10061 55613 10117 55624
rect 9937 55568 9947 55613
rect 9947 55568 9993 55613
rect 10061 55568 10107 55613
rect 10107 55568 10117 55613
rect 9937 55453 9947 55500
rect 9947 55453 9993 55500
rect 10061 55453 10107 55500
rect 10107 55453 10117 55500
rect 9937 55444 9993 55453
rect 10061 55444 10117 55453
rect 9937 55345 9947 55376
rect 9947 55345 9993 55376
rect 10061 55345 10107 55376
rect 10107 55345 10117 55376
rect 9937 55320 9993 55345
rect 10061 55320 10117 55345
rect 9937 55237 9947 55252
rect 9947 55237 9993 55252
rect 10061 55237 10107 55252
rect 10107 55237 10117 55252
rect 9937 55196 9993 55237
rect 10061 55196 10117 55237
rect 9937 55073 9993 55128
rect 10061 55073 10117 55128
rect 9937 55072 9947 55073
rect 9947 55072 9993 55073
rect 10061 55072 10107 55073
rect 10107 55072 10117 55073
rect 9937 54965 9993 55004
rect 10061 54965 10117 55004
rect 9937 54948 9947 54965
rect 9947 54948 9993 54965
rect 10061 54948 10107 54965
rect 10107 54948 10117 54965
rect 9937 54857 9993 54880
rect 10061 54857 10117 54880
rect 9937 54824 9947 54857
rect 9947 54824 9993 54857
rect 10061 54824 10107 54857
rect 10107 54824 10117 54857
rect 9937 54749 9993 54756
rect 10061 54749 10117 54756
rect 9937 54700 9947 54749
rect 9947 54700 9993 54749
rect 10061 54700 10107 54749
rect 10107 54700 10117 54749
rect 9937 54589 9947 54632
rect 9947 54589 9993 54632
rect 10061 54589 10107 54632
rect 10107 54589 10117 54632
rect 9937 54576 9993 54589
rect 10061 54576 10117 54589
rect 9937 54481 9947 54508
rect 9947 54481 9993 54508
rect 10061 54481 10107 54508
rect 10107 54481 10117 54508
rect 9937 54452 9993 54481
rect 10061 54452 10117 54481
rect 9937 47704 9947 47748
rect 9947 47704 9993 47748
rect 10061 47704 10107 47748
rect 10107 47704 10117 47748
rect 9937 47692 9993 47704
rect 10061 47692 10117 47704
rect 9937 47568 9993 47624
rect 10061 47568 10117 47624
rect 9937 47444 9993 47500
rect 10061 47444 10117 47500
rect 9937 47320 9993 47376
rect 10061 47320 10117 47376
rect 9937 47196 9993 47252
rect 10061 47196 10117 47252
rect 4861 47072 4917 47128
rect 4985 47072 5041 47128
rect 4861 46948 4917 47004
rect 4985 46948 5041 47004
rect 4861 46824 4917 46880
rect 4985 46824 5041 46880
rect 4861 46700 4917 46756
rect 4985 46700 5041 46756
rect 4861 46576 4917 46632
rect 4985 46576 5041 46632
rect 4861 46452 4917 46508
rect 4985 46452 5041 46508
rect 7275 47072 7331 47128
rect 7399 47072 7455 47128
rect 7523 47072 7579 47128
rect 7647 47072 7703 47128
rect 7275 46948 7331 47004
rect 7399 46948 7455 47004
rect 7523 46948 7579 47004
rect 7647 46948 7703 47004
rect 7275 46824 7331 46880
rect 7399 46824 7455 46880
rect 7523 46824 7579 46880
rect 7647 46824 7703 46880
rect 7275 46700 7331 46756
rect 7399 46700 7455 46756
rect 7523 46700 7579 46756
rect 7647 46700 7703 46756
rect 7275 46576 7331 46632
rect 7399 46576 7455 46632
rect 7523 46576 7579 46632
rect 7647 46576 7703 46632
rect 7275 46452 7331 46508
rect 7399 46452 7455 46508
rect 7523 46452 7579 46508
rect 7647 46452 7703 46508
rect 10254 57169 10310 57225
rect 10378 57169 10434 57225
rect 10502 57169 10558 57225
rect 10626 57169 10682 57225
rect 10750 57169 10806 57225
rect 10874 57169 10930 57225
rect 10998 57169 11054 57225
rect 11122 57169 11178 57225
rect 11246 57169 11302 57225
rect 11370 57169 11426 57225
rect 11494 57169 11550 57225
rect 11618 57169 11674 57225
rect 11742 57169 11798 57225
rect 11866 57169 11922 57225
rect 11990 57169 12046 57225
rect 12114 57169 12170 57225
rect 10254 57052 10266 57101
rect 10266 57052 10310 57101
rect 10378 57052 10430 57101
rect 10430 57052 10434 57101
rect 10502 57052 10538 57101
rect 10538 57052 10558 57101
rect 10626 57052 10646 57101
rect 10646 57052 10682 57101
rect 10750 57052 10754 57101
rect 10754 57052 10806 57101
rect 10874 57052 10914 57101
rect 10914 57052 10930 57101
rect 10998 57052 11022 57101
rect 11022 57052 11054 57101
rect 11122 57052 11130 57101
rect 11130 57052 11178 57101
rect 11246 57052 11294 57101
rect 11294 57052 11302 57101
rect 11370 57052 11402 57101
rect 11402 57052 11426 57101
rect 11494 57052 11510 57101
rect 11510 57052 11550 57101
rect 11618 57052 11670 57101
rect 11670 57052 11674 57101
rect 11742 57052 11778 57101
rect 11778 57052 11798 57101
rect 11866 57052 11886 57101
rect 11886 57052 11922 57101
rect 11990 57052 11994 57101
rect 11994 57052 12046 57101
rect 12114 57052 12158 57101
rect 12158 57052 12170 57101
rect 10254 57045 10310 57052
rect 10378 57045 10434 57052
rect 10502 57045 10558 57052
rect 10626 57045 10682 57052
rect 10750 57045 10806 57052
rect 10874 57045 10930 57052
rect 10998 57045 11054 57052
rect 11122 57045 11178 57052
rect 11246 57045 11302 57052
rect 11370 57045 11426 57052
rect 11494 57045 11550 57052
rect 11618 57045 11674 57052
rect 11742 57045 11798 57052
rect 11866 57045 11922 57052
rect 11990 57045 12046 57052
rect 12114 57045 12170 57052
rect 10254 56921 10310 56977
rect 10378 56921 10434 56977
rect 10502 56921 10558 56977
rect 10626 56921 10682 56977
rect 10750 56921 10806 56977
rect 10874 56921 10930 56977
rect 10998 56921 11054 56977
rect 11122 56921 11178 56977
rect 11246 56921 11302 56977
rect 11370 56921 11426 56977
rect 11494 56921 11550 56977
rect 11618 56921 11674 56977
rect 11742 56921 11798 56977
rect 11866 56921 11922 56977
rect 11990 56921 12046 56977
rect 12114 56921 12170 56977
rect 10254 56797 10310 56853
rect 10378 56797 10434 56853
rect 10502 56797 10558 56853
rect 10626 56797 10682 56853
rect 10750 56797 10806 56853
rect 10874 56797 10930 56853
rect 10998 56797 11054 56853
rect 11122 56797 11178 56853
rect 11246 56797 11302 56853
rect 11370 56797 11426 56853
rect 11494 56797 11550 56853
rect 11618 56797 11674 56853
rect 11742 56797 11798 56853
rect 11866 56797 11922 56853
rect 11990 56797 12046 56853
rect 12114 56797 12170 56853
rect 10254 56673 10310 56729
rect 10378 56673 10434 56729
rect 10502 56673 10558 56729
rect 10626 56673 10682 56729
rect 10750 56673 10806 56729
rect 10874 56673 10930 56729
rect 10998 56673 11054 56729
rect 11122 56673 11178 56729
rect 11246 56673 11302 56729
rect 11370 56673 11426 56729
rect 11494 56673 11550 56729
rect 11618 56673 11674 56729
rect 11742 56673 11798 56729
rect 11866 56673 11922 56729
rect 11990 56673 12046 56729
rect 12114 56673 12170 56729
rect 10254 56549 10310 56605
rect 10378 56549 10434 56605
rect 10502 56549 10558 56605
rect 10626 56549 10682 56605
rect 10750 56591 10775 56605
rect 10775 56591 10806 56605
rect 10874 56591 10899 56605
rect 10899 56591 10930 56605
rect 10998 56591 11023 56605
rect 11023 56591 11054 56605
rect 10750 56549 10806 56591
rect 10874 56549 10930 56591
rect 10998 56549 11054 56591
rect 11122 56549 11178 56605
rect 11246 56549 11302 56605
rect 11370 56549 11426 56605
rect 11494 56549 11550 56605
rect 11618 56549 11674 56605
rect 11742 56549 11798 56605
rect 11866 56549 11922 56605
rect 11990 56549 12046 56605
rect 12114 56549 12170 56605
rect 10254 56425 10310 56481
rect 10378 56425 10434 56481
rect 10502 56425 10558 56481
rect 10626 56425 10682 56481
rect 10750 56467 10775 56481
rect 10775 56467 10806 56481
rect 10874 56467 10899 56481
rect 10899 56467 10930 56481
rect 10998 56467 11023 56481
rect 11023 56467 11054 56481
rect 10750 56425 10806 56467
rect 10874 56425 10930 56467
rect 10998 56425 11054 56467
rect 11122 56425 11178 56481
rect 11246 56425 11302 56481
rect 11370 56425 11426 56481
rect 11494 56425 11550 56481
rect 11618 56425 11674 56481
rect 11742 56425 11798 56481
rect 11866 56425 11922 56481
rect 11990 56425 12046 56481
rect 12114 56425 12170 56481
rect 10254 56301 10310 56357
rect 10378 56301 10434 56357
rect 10502 56301 10558 56357
rect 10626 56301 10682 56357
rect 10750 56343 10775 56357
rect 10775 56343 10806 56357
rect 10874 56343 10899 56357
rect 10899 56343 10930 56357
rect 10998 56343 11023 56357
rect 11023 56343 11054 56357
rect 10750 56301 10806 56343
rect 10874 56301 10930 56343
rect 10998 56301 11054 56343
rect 11122 56301 11178 56357
rect 11246 56301 11302 56357
rect 11370 56301 11426 56357
rect 11494 56301 11550 56357
rect 11618 56301 11674 56357
rect 11742 56301 11798 56357
rect 11866 56301 11922 56357
rect 11990 56301 12046 56357
rect 12114 56301 12170 56357
rect 10254 56177 10310 56233
rect 10378 56177 10434 56233
rect 10502 56177 10558 56233
rect 10626 56177 10682 56233
rect 10750 56219 10775 56233
rect 10775 56219 10806 56233
rect 10874 56219 10899 56233
rect 10899 56219 10930 56233
rect 10998 56219 11023 56233
rect 11023 56219 11054 56233
rect 10750 56177 10806 56219
rect 10874 56177 10930 56219
rect 10998 56177 11054 56219
rect 11122 56177 11178 56233
rect 11246 56177 11302 56233
rect 11370 56177 11426 56233
rect 11494 56177 11550 56233
rect 11618 56177 11674 56233
rect 11742 56177 11798 56233
rect 11866 56177 11922 56233
rect 11990 56177 12046 56233
rect 12114 56177 12170 56233
rect 10254 56053 10310 56109
rect 10378 56053 10434 56109
rect 10502 56053 10558 56109
rect 10626 56053 10682 56109
rect 10750 56095 10775 56109
rect 10775 56095 10806 56109
rect 10874 56095 10899 56109
rect 10899 56095 10930 56109
rect 10998 56095 11023 56109
rect 11023 56095 11054 56109
rect 10750 56053 10806 56095
rect 10874 56053 10930 56095
rect 10998 56053 11054 56095
rect 11122 56053 11178 56109
rect 11246 56053 11302 56109
rect 11370 56053 11426 56109
rect 11494 56053 11550 56109
rect 11618 56053 11674 56109
rect 11742 56053 11798 56109
rect 11866 56053 11922 56109
rect 11990 56053 12046 56109
rect 12114 56053 12170 56109
rect 10254 54092 10310 54148
rect 10378 54092 10434 54148
rect 10502 54092 10558 54148
rect 10626 54092 10682 54148
rect 10750 54111 10775 54148
rect 10775 54111 10806 54148
rect 10874 54111 10899 54148
rect 10899 54111 10930 54148
rect 10998 54111 11023 54148
rect 11023 54111 11054 54148
rect 10750 54092 10806 54111
rect 10874 54092 10930 54111
rect 10998 54092 11054 54111
rect 11122 54092 11178 54148
rect 11246 54092 11302 54148
rect 11370 54092 11426 54148
rect 11494 54092 11550 54148
rect 11618 54092 11674 54148
rect 11742 54092 11798 54148
rect 11866 54092 11922 54148
rect 11990 54092 12046 54148
rect 12114 54092 12170 54148
rect 10254 53968 10310 54024
rect 10378 53968 10434 54024
rect 10502 53968 10558 54024
rect 10626 53968 10682 54024
rect 10750 53987 10775 54024
rect 10775 53987 10806 54024
rect 10874 53987 10899 54024
rect 10899 53987 10930 54024
rect 10998 53987 11023 54024
rect 11023 53987 11054 54024
rect 10750 53968 10806 53987
rect 10874 53968 10930 53987
rect 10998 53968 11054 53987
rect 11122 53968 11178 54024
rect 11246 53968 11302 54024
rect 11370 53968 11426 54024
rect 11494 53968 11550 54024
rect 11618 53968 11674 54024
rect 11742 53968 11798 54024
rect 11866 53968 11922 54024
rect 11990 53968 12046 54024
rect 12114 53968 12170 54024
rect 10254 53844 10310 53900
rect 10378 53844 10434 53900
rect 10502 53844 10558 53900
rect 10626 53844 10682 53900
rect 10750 53863 10775 53900
rect 10775 53863 10806 53900
rect 10874 53863 10899 53900
rect 10899 53863 10930 53900
rect 10998 53863 11023 53900
rect 11023 53863 11054 53900
rect 10750 53844 10806 53863
rect 10874 53844 10930 53863
rect 10998 53844 11054 53863
rect 11122 53844 11178 53900
rect 11246 53844 11302 53900
rect 11370 53844 11426 53900
rect 11494 53844 11550 53900
rect 11618 53844 11674 53900
rect 11742 53844 11798 53900
rect 11866 53844 11922 53900
rect 11990 53844 12046 53900
rect 12114 53844 12170 53900
rect 10254 53720 10310 53776
rect 10378 53720 10434 53776
rect 10502 53720 10558 53776
rect 10626 53720 10682 53776
rect 10750 53739 10775 53776
rect 10775 53739 10806 53776
rect 10874 53739 10899 53776
rect 10899 53739 10930 53776
rect 10998 53739 11023 53776
rect 11023 53739 11054 53776
rect 10750 53720 10806 53739
rect 10874 53720 10930 53739
rect 10998 53720 11054 53739
rect 11122 53720 11178 53776
rect 11246 53720 11302 53776
rect 11370 53720 11426 53776
rect 11494 53720 11550 53776
rect 11618 53720 11674 53776
rect 11742 53720 11798 53776
rect 11866 53720 11922 53776
rect 11990 53720 12046 53776
rect 12114 53720 12170 53776
rect 10254 53596 10310 53652
rect 10378 53596 10434 53652
rect 10502 53596 10558 53652
rect 10626 53596 10682 53652
rect 10750 53615 10775 53652
rect 10775 53615 10806 53652
rect 10874 53615 10899 53652
rect 10899 53615 10930 53652
rect 10998 53615 11023 53652
rect 11023 53615 11054 53652
rect 10750 53596 10806 53615
rect 10874 53596 10930 53615
rect 10998 53596 11054 53615
rect 11122 53596 11178 53652
rect 11246 53596 11302 53652
rect 11370 53596 11426 53652
rect 11494 53596 11550 53652
rect 11618 53596 11674 53652
rect 11742 53596 11798 53652
rect 11866 53596 11922 53652
rect 11990 53596 12046 53652
rect 12114 53596 12170 53652
rect 10254 53472 10310 53528
rect 10378 53472 10434 53528
rect 10502 53472 10558 53528
rect 10626 53472 10682 53528
rect 10750 53491 10775 53528
rect 10775 53491 10806 53528
rect 10874 53491 10899 53528
rect 10899 53491 10930 53528
rect 10998 53491 11023 53528
rect 11023 53491 11054 53528
rect 10750 53472 10806 53491
rect 10874 53472 10930 53491
rect 10998 53472 11054 53491
rect 11122 53472 11178 53528
rect 11246 53483 11302 53528
rect 11370 53483 11426 53528
rect 11494 53483 11550 53528
rect 11618 53483 11674 53528
rect 11742 53483 11798 53528
rect 11866 53483 11922 53528
rect 11990 53483 12046 53528
rect 12114 53483 12170 53528
rect 11246 53472 11299 53483
rect 11299 53472 11302 53483
rect 11370 53472 11407 53483
rect 11407 53472 11426 53483
rect 11494 53472 11515 53483
rect 11515 53472 11550 53483
rect 11618 53472 11623 53483
rect 11623 53472 11674 53483
rect 11742 53472 11783 53483
rect 11783 53472 11798 53483
rect 11866 53472 11891 53483
rect 11891 53472 11922 53483
rect 11990 53472 11999 53483
rect 11999 53472 12046 53483
rect 12114 53472 12163 53483
rect 12163 53472 12170 53483
rect 10254 53348 10310 53404
rect 10378 53348 10434 53404
rect 10502 53348 10558 53404
rect 10626 53348 10682 53404
rect 10750 53367 10775 53404
rect 10775 53367 10806 53404
rect 10874 53367 10899 53404
rect 10899 53367 10930 53404
rect 10998 53367 11023 53404
rect 11023 53367 11054 53404
rect 10750 53348 10806 53367
rect 10874 53348 10930 53367
rect 10998 53348 11054 53367
rect 11122 53348 11178 53404
rect 11246 53375 11302 53404
rect 11370 53375 11426 53404
rect 11494 53375 11550 53404
rect 11618 53375 11674 53404
rect 11742 53375 11798 53404
rect 11866 53375 11922 53404
rect 11990 53375 12046 53404
rect 12114 53375 12170 53404
rect 11246 53348 11299 53375
rect 11299 53348 11302 53375
rect 11370 53348 11407 53375
rect 11407 53348 11426 53375
rect 11494 53348 11515 53375
rect 11515 53348 11550 53375
rect 11618 53348 11623 53375
rect 11623 53348 11674 53375
rect 11742 53348 11783 53375
rect 11783 53348 11798 53375
rect 11866 53348 11891 53375
rect 11891 53348 11922 53375
rect 11990 53348 11999 53375
rect 11999 53348 12046 53375
rect 12114 53348 12163 53375
rect 12163 53348 12170 53375
rect 10254 53224 10310 53280
rect 10378 53224 10434 53280
rect 10502 53224 10558 53280
rect 10626 53224 10682 53280
rect 10750 53243 10775 53280
rect 10775 53243 10806 53280
rect 10874 53243 10899 53280
rect 10899 53243 10930 53280
rect 10998 53243 11023 53280
rect 11023 53243 11054 53280
rect 10750 53224 10806 53243
rect 10874 53224 10930 53243
rect 10998 53224 11054 53243
rect 11122 53224 11178 53280
rect 11246 53267 11302 53280
rect 11370 53267 11426 53280
rect 11494 53267 11550 53280
rect 11618 53267 11674 53280
rect 11742 53267 11798 53280
rect 11866 53267 11922 53280
rect 11990 53267 12046 53280
rect 12114 53267 12170 53280
rect 11246 53224 11299 53267
rect 11299 53224 11302 53267
rect 11370 53224 11407 53267
rect 11407 53224 11426 53267
rect 11494 53224 11515 53267
rect 11515 53224 11550 53267
rect 11618 53224 11623 53267
rect 11623 53224 11674 53267
rect 11742 53224 11783 53267
rect 11783 53224 11798 53267
rect 11866 53224 11891 53267
rect 11891 53224 11922 53267
rect 11990 53224 11999 53267
rect 11999 53224 12046 53267
rect 12114 53224 12163 53267
rect 12163 53224 12170 53267
rect 10254 53100 10310 53156
rect 10378 53100 10434 53156
rect 10502 53100 10558 53156
rect 10626 53100 10682 53156
rect 10750 53100 10806 53156
rect 10874 53100 10930 53156
rect 10998 53100 11054 53156
rect 11122 53100 11178 53156
rect 11246 53100 11302 53156
rect 11370 53100 11426 53156
rect 11494 53100 11550 53156
rect 11618 53100 11674 53156
rect 11742 53100 11798 53156
rect 11866 53100 11922 53156
rect 11990 53100 12046 53156
rect 12114 53100 12170 53156
rect 10254 52976 10310 53032
rect 10378 52976 10434 53032
rect 10502 52976 10558 53032
rect 10626 52976 10682 53032
rect 10750 52976 10806 53032
rect 10874 52976 10930 53032
rect 10998 52976 11054 53032
rect 11122 52976 11178 53032
rect 11246 52976 11302 53032
rect 11370 52976 11426 53032
rect 11494 52976 11550 53032
rect 11618 52976 11674 53032
rect 11742 52976 11798 53032
rect 11866 52976 11922 53032
rect 11990 52976 12046 53032
rect 12114 52976 12170 53032
rect 10254 52852 10310 52908
rect 10378 52852 10434 52908
rect 10502 52852 10558 52908
rect 10626 52852 10682 52908
rect 10750 52852 10806 52908
rect 10874 52852 10930 52908
rect 10998 52852 11054 52908
rect 11122 52852 11178 52908
rect 11246 52852 11302 52908
rect 11370 52852 11426 52908
rect 11494 52852 11550 52908
rect 11618 52852 11674 52908
rect 11742 52852 11798 52908
rect 11866 52852 11922 52908
rect 11990 52852 12046 52908
rect 12114 52852 12170 52908
rect 10254 52492 10310 52548
rect 10378 52492 10434 52548
rect 10502 52492 10558 52548
rect 10626 52492 10682 52548
rect 10750 52492 10806 52548
rect 10874 52492 10930 52548
rect 10998 52492 11054 52548
rect 11122 52492 11178 52548
rect 11246 52492 11302 52548
rect 11370 52492 11426 52548
rect 11494 52492 11550 52548
rect 11618 52492 11674 52548
rect 11742 52492 11798 52548
rect 11866 52492 11922 52548
rect 11990 52492 12046 52548
rect 12114 52492 12170 52548
rect 10254 52368 10310 52424
rect 10378 52368 10434 52424
rect 10502 52368 10558 52424
rect 10626 52368 10682 52424
rect 10750 52368 10806 52424
rect 10874 52368 10930 52424
rect 10998 52368 11054 52424
rect 11122 52368 11178 52424
rect 11246 52368 11302 52424
rect 11370 52368 11426 52424
rect 11494 52368 11550 52424
rect 11618 52368 11674 52424
rect 11742 52368 11798 52424
rect 11866 52368 11922 52424
rect 11990 52368 12046 52424
rect 12114 52368 12170 52424
rect 10254 52244 10310 52300
rect 10378 52244 10434 52300
rect 10502 52244 10558 52300
rect 10626 52244 10682 52300
rect 10750 52244 10806 52300
rect 10874 52244 10930 52300
rect 10998 52244 11054 52300
rect 11122 52244 11178 52300
rect 11246 52244 11302 52300
rect 11370 52244 11426 52300
rect 11494 52244 11550 52300
rect 11618 52244 11674 52300
rect 11742 52244 11798 52300
rect 11866 52244 11922 52300
rect 11990 52244 12046 52300
rect 12114 52244 12170 52300
rect 10254 52120 10310 52176
rect 10378 52120 10434 52176
rect 10502 52120 10558 52176
rect 10626 52120 10682 52176
rect 10750 52120 10806 52176
rect 10874 52120 10930 52176
rect 10998 52120 11054 52176
rect 11122 52120 11178 52176
rect 11246 52120 11302 52176
rect 11370 52120 11426 52176
rect 11494 52120 11550 52176
rect 11618 52120 11674 52176
rect 11742 52120 11798 52176
rect 11866 52120 11922 52176
rect 11990 52120 12046 52176
rect 12114 52120 12170 52176
rect 10254 52009 10310 52052
rect 10378 52009 10434 52052
rect 10502 52009 10558 52052
rect 10626 52009 10682 52052
rect 10750 52009 10806 52052
rect 10874 52009 10930 52052
rect 10998 52009 11054 52052
rect 11122 52009 11178 52052
rect 11246 52009 11302 52052
rect 11370 52009 11426 52052
rect 11494 52009 11550 52052
rect 11618 52009 11674 52052
rect 11742 52009 11798 52052
rect 10254 51996 10305 52009
rect 10305 51996 10310 52009
rect 10378 51996 10413 52009
rect 10413 51996 10434 52009
rect 10502 51996 10521 52009
rect 10521 51996 10558 52009
rect 10626 51996 10629 52009
rect 10629 51996 10682 52009
rect 10750 51996 10793 52009
rect 10793 51996 10806 52009
rect 10874 51996 10901 52009
rect 10901 51996 10930 52009
rect 10998 51996 11009 52009
rect 11009 51996 11054 52009
rect 11122 51996 11169 52009
rect 11169 51996 11178 52009
rect 11246 51996 11277 52009
rect 11277 51996 11302 52009
rect 11370 51996 11385 52009
rect 11385 51996 11426 52009
rect 11494 51996 11549 52009
rect 11549 51996 11550 52009
rect 11618 51996 11657 52009
rect 11657 51996 11674 52009
rect 11742 51996 11765 52009
rect 11765 51996 11798 52009
rect 11866 51996 11922 52052
rect 11990 51996 12046 52052
rect 12114 51996 12170 52052
rect 10254 51901 10310 51928
rect 10378 51901 10434 51928
rect 10502 51901 10558 51928
rect 10626 51901 10682 51928
rect 10750 51901 10806 51928
rect 10874 51901 10930 51928
rect 10998 51901 11054 51928
rect 11122 51901 11178 51928
rect 11246 51901 11302 51928
rect 11370 51901 11426 51928
rect 11494 51901 11550 51928
rect 11618 51901 11674 51928
rect 11742 51901 11798 51928
rect 10254 51872 10305 51901
rect 10305 51872 10310 51901
rect 10378 51872 10413 51901
rect 10413 51872 10434 51901
rect 10502 51872 10521 51901
rect 10521 51872 10558 51901
rect 10626 51872 10629 51901
rect 10629 51872 10682 51901
rect 10750 51872 10793 51901
rect 10793 51872 10806 51901
rect 10874 51872 10901 51901
rect 10901 51872 10930 51901
rect 10998 51872 11009 51901
rect 11009 51872 11054 51901
rect 11122 51872 11169 51901
rect 11169 51872 11178 51901
rect 11246 51872 11277 51901
rect 11277 51872 11302 51901
rect 11370 51872 11385 51901
rect 11385 51872 11426 51901
rect 11494 51872 11549 51901
rect 11549 51872 11550 51901
rect 11618 51872 11657 51901
rect 11657 51872 11674 51901
rect 11742 51872 11765 51901
rect 11765 51872 11798 51901
rect 11866 51872 11922 51928
rect 11990 51872 12046 51928
rect 12114 51872 12170 51928
rect 10254 51748 10310 51804
rect 10378 51748 10434 51804
rect 10502 51748 10558 51804
rect 10626 51748 10682 51804
rect 10750 51748 10806 51804
rect 10874 51748 10930 51804
rect 10998 51748 11054 51804
rect 11122 51748 11178 51804
rect 11246 51748 11302 51804
rect 11370 51748 11426 51804
rect 11494 51748 11550 51804
rect 11618 51748 11674 51804
rect 11742 51748 11798 51804
rect 11866 51748 11922 51804
rect 11990 51748 12046 51804
rect 12114 51748 12170 51804
rect 10254 51624 10310 51680
rect 10378 51624 10434 51680
rect 10502 51624 10558 51680
rect 10626 51624 10682 51680
rect 10750 51624 10806 51680
rect 10874 51624 10930 51680
rect 10998 51624 11054 51680
rect 11122 51624 11178 51680
rect 11246 51624 11302 51680
rect 11370 51624 11426 51680
rect 11494 51624 11550 51680
rect 11618 51624 11674 51680
rect 11742 51624 11798 51680
rect 11866 51624 11922 51680
rect 11990 51624 12046 51680
rect 12114 51624 12170 51680
rect 10254 51500 10310 51556
rect 10378 51500 10434 51556
rect 10502 51500 10558 51556
rect 10626 51500 10682 51556
rect 10750 51500 10806 51556
rect 10874 51500 10930 51556
rect 10998 51500 11054 51556
rect 11122 51500 11178 51556
rect 11246 51500 11302 51556
rect 11370 51500 11426 51556
rect 11494 51500 11550 51556
rect 11618 51500 11674 51556
rect 11742 51500 11798 51556
rect 11866 51500 11922 51556
rect 11990 51500 12046 51556
rect 12114 51500 12170 51556
rect 10254 51376 10310 51432
rect 10378 51376 10434 51432
rect 10502 51376 10558 51432
rect 10626 51376 10682 51432
rect 10750 51376 10806 51432
rect 10874 51376 10930 51432
rect 10998 51376 11054 51432
rect 11122 51376 11178 51432
rect 11246 51376 11302 51432
rect 11370 51376 11426 51432
rect 11494 51376 11550 51432
rect 11618 51376 11674 51432
rect 11742 51376 11798 51432
rect 11866 51376 11922 51432
rect 11990 51376 12046 51432
rect 12114 51376 12170 51432
rect 10254 51252 10310 51308
rect 10378 51252 10434 51308
rect 10502 51252 10558 51308
rect 10626 51252 10682 51308
rect 10750 51252 10806 51308
rect 10874 51252 10930 51308
rect 10998 51252 11054 51308
rect 11122 51252 11178 51308
rect 11246 51252 11302 51308
rect 11370 51252 11426 51308
rect 11494 51252 11550 51308
rect 11618 51252 11674 51308
rect 11742 51252 11798 51308
rect 11866 51252 11922 51308
rect 11990 51252 12046 51308
rect 12114 51252 12170 51308
rect 10254 49338 10310 49348
rect 10378 49338 10434 49348
rect 10502 49338 10558 49348
rect 10626 49338 10682 49348
rect 10750 49338 10806 49348
rect 10874 49338 10930 49348
rect 10998 49338 11054 49348
rect 11122 49338 11178 49348
rect 11246 49338 11302 49348
rect 11370 49338 11426 49348
rect 11494 49338 11550 49348
rect 11618 49338 11674 49348
rect 11742 49338 11798 49348
rect 10254 49292 10305 49338
rect 10305 49292 10310 49338
rect 10378 49292 10413 49338
rect 10413 49292 10434 49338
rect 10502 49292 10521 49338
rect 10521 49292 10558 49338
rect 10626 49292 10629 49338
rect 10629 49292 10682 49338
rect 10750 49292 10793 49338
rect 10793 49292 10806 49338
rect 10874 49292 10901 49338
rect 10901 49292 10930 49338
rect 10998 49292 11009 49338
rect 11009 49292 11054 49338
rect 11122 49292 11169 49338
rect 11169 49292 11178 49338
rect 11246 49292 11277 49338
rect 11277 49292 11302 49338
rect 11370 49292 11385 49338
rect 11385 49292 11426 49338
rect 11494 49292 11549 49338
rect 11549 49292 11550 49338
rect 11618 49292 11657 49338
rect 11657 49292 11674 49338
rect 11742 49292 11765 49338
rect 11765 49292 11798 49338
rect 11866 49292 11922 49348
rect 11990 49292 12046 49348
rect 12114 49292 12170 49348
rect 10254 49178 10305 49224
rect 10305 49178 10310 49224
rect 10378 49178 10413 49224
rect 10413 49178 10434 49224
rect 10502 49178 10521 49224
rect 10521 49178 10558 49224
rect 10626 49178 10629 49224
rect 10629 49178 10682 49224
rect 10750 49178 10793 49224
rect 10793 49178 10806 49224
rect 10874 49178 10901 49224
rect 10901 49178 10930 49224
rect 10998 49178 11009 49224
rect 11009 49178 11054 49224
rect 11122 49178 11169 49224
rect 11169 49178 11178 49224
rect 11246 49178 11277 49224
rect 11277 49178 11302 49224
rect 11370 49178 11385 49224
rect 11385 49178 11426 49224
rect 11494 49178 11549 49224
rect 11549 49178 11550 49224
rect 11618 49178 11657 49224
rect 11657 49178 11674 49224
rect 11742 49178 11765 49224
rect 11765 49178 11798 49224
rect 10254 49168 10310 49178
rect 10378 49168 10434 49178
rect 10502 49168 10558 49178
rect 10626 49168 10682 49178
rect 10750 49168 10806 49178
rect 10874 49168 10930 49178
rect 10998 49168 11054 49178
rect 11122 49168 11178 49178
rect 11246 49168 11302 49178
rect 11370 49168 11426 49178
rect 11494 49168 11550 49178
rect 11618 49168 11674 49178
rect 11742 49168 11798 49178
rect 11866 49168 11922 49224
rect 11990 49168 12046 49224
rect 12114 49168 12170 49224
rect 10254 49070 10305 49100
rect 10305 49070 10310 49100
rect 10378 49070 10413 49100
rect 10413 49070 10434 49100
rect 10502 49070 10521 49100
rect 10521 49070 10558 49100
rect 10626 49070 10629 49100
rect 10629 49070 10682 49100
rect 10750 49070 10793 49100
rect 10793 49070 10806 49100
rect 10874 49070 10901 49100
rect 10901 49070 10930 49100
rect 10998 49070 11009 49100
rect 11009 49070 11054 49100
rect 11122 49070 11169 49100
rect 11169 49070 11178 49100
rect 11246 49070 11277 49100
rect 11277 49070 11302 49100
rect 11370 49070 11385 49100
rect 11385 49070 11426 49100
rect 11494 49070 11549 49100
rect 11549 49070 11550 49100
rect 11618 49070 11657 49100
rect 11657 49070 11674 49100
rect 11742 49070 11765 49100
rect 11765 49070 11798 49100
rect 10254 49044 10310 49070
rect 10378 49044 10434 49070
rect 10502 49044 10558 49070
rect 10626 49044 10682 49070
rect 10750 49044 10806 49070
rect 10874 49044 10930 49070
rect 10998 49044 11054 49070
rect 11122 49044 11178 49070
rect 11246 49044 11302 49070
rect 11370 49044 11426 49070
rect 11494 49044 11550 49070
rect 11618 49044 11674 49070
rect 11742 49044 11798 49070
rect 11866 49044 11922 49100
rect 11990 49044 12046 49100
rect 12114 49044 12170 49100
rect 10254 48920 10310 48976
rect 10378 48920 10434 48976
rect 10502 48920 10558 48976
rect 10626 48920 10682 48976
rect 10750 48920 10806 48976
rect 10874 48920 10930 48976
rect 10998 48920 11054 48976
rect 11122 48920 11178 48976
rect 11246 48920 11302 48976
rect 11370 48920 11426 48976
rect 11494 48920 11550 48976
rect 11618 48920 11674 48976
rect 11742 48920 11798 48976
rect 11866 48920 11922 48976
rect 11990 48920 12046 48976
rect 12114 48920 12170 48976
rect 10254 48796 10310 48852
rect 10378 48796 10434 48852
rect 10502 48796 10558 48852
rect 10626 48796 10682 48852
rect 10750 48796 10806 48852
rect 10874 48796 10930 48852
rect 10998 48796 11054 48852
rect 11122 48796 11178 48852
rect 11246 48796 11302 48852
rect 11370 48796 11426 48852
rect 11494 48796 11550 48852
rect 11618 48796 11674 48852
rect 11742 48796 11798 48852
rect 11866 48796 11922 48852
rect 11990 48796 12046 48852
rect 12114 48796 12170 48852
rect 10254 48672 10310 48728
rect 10378 48672 10434 48728
rect 10502 48672 10558 48728
rect 10626 48672 10682 48728
rect 10750 48672 10806 48728
rect 10874 48672 10930 48728
rect 10998 48672 11054 48728
rect 11122 48672 11178 48728
rect 11246 48672 11302 48728
rect 11370 48672 11426 48728
rect 11494 48672 11550 48728
rect 11618 48672 11674 48728
rect 11742 48672 11798 48728
rect 11866 48672 11922 48728
rect 11990 48672 12046 48728
rect 12114 48672 12170 48728
rect 10254 48548 10310 48604
rect 10378 48548 10434 48604
rect 10502 48548 10558 48604
rect 10626 48548 10682 48604
rect 10750 48548 10806 48604
rect 10874 48548 10930 48604
rect 10998 48548 11054 48604
rect 11122 48548 11178 48604
rect 11246 48548 11302 48604
rect 11370 48548 11426 48604
rect 11494 48548 11550 48604
rect 11618 48548 11674 48604
rect 11742 48548 11798 48604
rect 11866 48548 11922 48604
rect 11990 48548 12046 48604
rect 12114 48548 12170 48604
rect 10254 48427 10310 48480
rect 10378 48427 10434 48480
rect 10502 48427 10558 48480
rect 10626 48427 10682 48480
rect 10750 48427 10806 48480
rect 10874 48427 10930 48480
rect 10998 48427 11054 48480
rect 11122 48427 11178 48480
rect 11246 48427 11302 48480
rect 11370 48427 11426 48480
rect 11494 48427 11550 48480
rect 11618 48427 11674 48480
rect 11742 48427 11798 48480
rect 10254 48424 10305 48427
rect 10305 48424 10310 48427
rect 10378 48424 10413 48427
rect 10413 48424 10434 48427
rect 10502 48424 10521 48427
rect 10521 48424 10558 48427
rect 10626 48424 10629 48427
rect 10629 48424 10682 48427
rect 10750 48424 10793 48427
rect 10793 48424 10806 48427
rect 10874 48424 10901 48427
rect 10901 48424 10930 48427
rect 10998 48424 11009 48427
rect 11009 48424 11054 48427
rect 11122 48424 11169 48427
rect 11169 48424 11178 48427
rect 11246 48424 11277 48427
rect 11277 48424 11302 48427
rect 11370 48424 11385 48427
rect 11385 48424 11426 48427
rect 11494 48424 11549 48427
rect 11549 48424 11550 48427
rect 11618 48424 11657 48427
rect 11657 48424 11674 48427
rect 11742 48424 11765 48427
rect 11765 48424 11798 48427
rect 11866 48424 11922 48480
rect 11990 48424 12046 48480
rect 12114 48424 12170 48480
rect 10254 48319 10310 48356
rect 10378 48319 10434 48356
rect 10502 48319 10558 48356
rect 10626 48319 10682 48356
rect 10750 48319 10806 48356
rect 10874 48319 10930 48356
rect 10998 48319 11054 48356
rect 11122 48319 11178 48356
rect 11246 48319 11302 48356
rect 11370 48319 11426 48356
rect 11494 48319 11550 48356
rect 11618 48319 11674 48356
rect 11742 48319 11798 48356
rect 10254 48300 10305 48319
rect 10305 48300 10310 48319
rect 10378 48300 10413 48319
rect 10413 48300 10434 48319
rect 10502 48300 10521 48319
rect 10521 48300 10558 48319
rect 10626 48300 10629 48319
rect 10629 48300 10682 48319
rect 10750 48300 10793 48319
rect 10793 48300 10806 48319
rect 10874 48300 10901 48319
rect 10901 48300 10930 48319
rect 10998 48300 11009 48319
rect 11009 48300 11054 48319
rect 11122 48300 11169 48319
rect 11169 48300 11178 48319
rect 11246 48300 11277 48319
rect 11277 48300 11302 48319
rect 11370 48300 11385 48319
rect 11385 48300 11426 48319
rect 11494 48300 11549 48319
rect 11549 48300 11550 48319
rect 11618 48300 11657 48319
rect 11657 48300 11674 48319
rect 11742 48300 11765 48319
rect 11765 48300 11798 48319
rect 11866 48300 11922 48356
rect 11990 48300 12046 48356
rect 12114 48300 12170 48356
rect 10254 48176 10310 48232
rect 10378 48176 10434 48232
rect 10502 48176 10558 48232
rect 10626 48176 10682 48232
rect 10750 48176 10806 48232
rect 10874 48176 10930 48232
rect 10998 48176 11054 48232
rect 11122 48176 11178 48232
rect 11246 48176 11302 48232
rect 11370 48176 11426 48232
rect 11494 48176 11550 48232
rect 11618 48176 11674 48232
rect 11742 48176 11798 48232
rect 11866 48176 11922 48232
rect 11990 48176 12046 48232
rect 12114 48176 12170 48232
rect 10254 48052 10310 48108
rect 10378 48052 10434 48108
rect 10502 48052 10558 48108
rect 10626 48052 10682 48108
rect 10750 48052 10806 48108
rect 10874 48052 10930 48108
rect 10998 48052 11054 48108
rect 11122 48052 11178 48108
rect 11246 48052 11302 48108
rect 11370 48052 11426 48108
rect 11494 48052 11550 48108
rect 11618 48052 11674 48108
rect 11742 48052 11798 48108
rect 11866 48052 11922 48108
rect 11990 48052 12046 48108
rect 12114 48052 12170 48108
rect 12307 55692 12363 55748
rect 12431 55692 12487 55748
rect 12307 55568 12363 55624
rect 12431 55568 12487 55624
rect 12307 55444 12363 55500
rect 12431 55444 12487 55500
rect 12307 55320 12363 55376
rect 12431 55320 12487 55376
rect 12307 55196 12363 55252
rect 12431 55196 12487 55252
rect 12307 55072 12363 55128
rect 12431 55072 12487 55128
rect 12307 54948 12363 55004
rect 12431 54948 12487 55004
rect 12307 54824 12363 54880
rect 12431 54824 12487 54880
rect 12307 54700 12363 54756
rect 12431 54700 12487 54756
rect 12307 54576 12363 54632
rect 12431 54576 12487 54632
rect 12307 54452 12363 54508
rect 12431 54452 12487 54508
rect 12307 47734 12363 47748
rect 12307 47692 12336 47734
rect 12336 47692 12363 47734
rect 12431 47692 12487 47748
rect 12307 47568 12363 47624
rect 12431 47568 12487 47624
rect 12307 47444 12363 47500
rect 12431 47444 12487 47500
rect 12307 47320 12363 47376
rect 12431 47320 12487 47376
rect 12307 47196 12363 47252
rect 12431 47196 12487 47252
rect 9937 47072 9993 47128
rect 10061 47072 10117 47128
rect 9937 46948 9993 47004
rect 10061 46948 10117 47004
rect 9937 46824 9993 46880
rect 10061 46824 10117 46880
rect 9937 46700 9993 46756
rect 10061 46700 10117 46756
rect 9937 46576 9993 46632
rect 10061 46576 10117 46632
rect 9937 46452 9993 46508
rect 10061 46452 10117 46508
rect 12871 57169 12927 57225
rect 12995 57169 13051 57225
rect 13119 57169 13175 57225
rect 13243 57169 13299 57225
rect 13367 57169 13423 57225
rect 13491 57169 13547 57225
rect 13615 57169 13671 57225
rect 13739 57169 13795 57225
rect 13863 57169 13919 57225
rect 13987 57169 14043 57225
rect 14111 57169 14167 57225
rect 14235 57169 14291 57225
rect 14359 57169 14415 57225
rect 14483 57169 14539 57225
rect 14607 57169 14663 57225
rect 12871 57045 12927 57101
rect 12995 57052 13039 57101
rect 13039 57052 13051 57101
rect 13119 57052 13147 57101
rect 13147 57052 13175 57101
rect 13243 57052 13255 57101
rect 13255 57052 13299 57101
rect 13367 57052 13415 57101
rect 13415 57052 13423 57101
rect 13491 57052 13523 57101
rect 13523 57052 13547 57101
rect 13615 57052 13631 57101
rect 13631 57052 13671 57101
rect 12995 57045 13051 57052
rect 13119 57045 13175 57052
rect 13243 57045 13299 57052
rect 13367 57045 13423 57052
rect 13491 57045 13547 57052
rect 13615 57045 13671 57052
rect 13739 57045 13795 57101
rect 13863 57052 13903 57101
rect 13903 57052 13919 57101
rect 13987 57052 14011 57101
rect 14011 57052 14043 57101
rect 14111 57052 14119 57101
rect 14119 57052 14167 57101
rect 14235 57052 14279 57101
rect 14279 57052 14291 57101
rect 14359 57052 14387 57101
rect 14387 57052 14415 57101
rect 14483 57052 14495 57101
rect 14495 57052 14539 57101
rect 13863 57045 13919 57052
rect 13987 57045 14043 57052
rect 14111 57045 14167 57052
rect 14235 57045 14291 57052
rect 14359 57045 14415 57052
rect 14483 57045 14539 57052
rect 14607 57045 14663 57101
rect 12871 56921 12927 56977
rect 12995 56921 13051 56977
rect 13119 56921 13175 56977
rect 13243 56921 13299 56977
rect 13367 56921 13423 56977
rect 13491 56921 13547 56977
rect 13615 56921 13671 56977
rect 13739 56921 13795 56977
rect 13863 56921 13919 56977
rect 13987 56921 14043 56977
rect 14111 56921 14167 56977
rect 14235 56921 14291 56977
rect 14359 56921 14415 56977
rect 14483 56921 14539 56977
rect 14607 56921 14663 56977
rect 12871 56797 12927 56853
rect 12995 56797 13051 56853
rect 13119 56797 13175 56853
rect 13243 56797 13299 56853
rect 13367 56797 13423 56853
rect 13491 56797 13547 56853
rect 13615 56797 13671 56853
rect 13739 56797 13795 56853
rect 13863 56797 13919 56853
rect 13987 56797 14043 56853
rect 14111 56797 14167 56853
rect 14235 56797 14291 56853
rect 14359 56797 14415 56853
rect 14483 56797 14539 56853
rect 14607 56797 14663 56853
rect 12871 56673 12927 56729
rect 12995 56673 13051 56729
rect 13119 56673 13175 56729
rect 13243 56673 13299 56729
rect 13367 56673 13423 56729
rect 13491 56673 13547 56729
rect 13615 56673 13671 56729
rect 13739 56673 13795 56729
rect 13863 56673 13919 56729
rect 13987 56673 14043 56729
rect 14111 56673 14167 56729
rect 14235 56673 14291 56729
rect 14359 56673 14415 56729
rect 14483 56673 14539 56729
rect 14607 56673 14663 56729
rect 12871 56549 12927 56605
rect 12995 56549 13051 56605
rect 13119 56549 13175 56605
rect 13243 56549 13299 56605
rect 13367 56549 13423 56605
rect 13491 56549 13547 56605
rect 13615 56549 13671 56605
rect 13739 56549 13795 56605
rect 13863 56549 13919 56605
rect 13987 56549 14043 56605
rect 14111 56549 14167 56605
rect 14235 56591 14237 56605
rect 14237 56591 14291 56605
rect 14359 56591 14361 56605
rect 14361 56591 14415 56605
rect 14483 56591 14485 56605
rect 14485 56591 14539 56605
rect 14607 56591 14609 56605
rect 14609 56591 14663 56605
rect 14235 56549 14291 56591
rect 14359 56549 14415 56591
rect 14483 56549 14539 56591
rect 14607 56549 14663 56591
rect 12871 56425 12927 56481
rect 12995 56425 13051 56481
rect 13119 56425 13175 56481
rect 13243 56425 13299 56481
rect 13367 56425 13423 56481
rect 13491 56425 13547 56481
rect 13615 56425 13671 56481
rect 13739 56425 13795 56481
rect 13863 56425 13919 56481
rect 13987 56425 14043 56481
rect 14111 56425 14167 56481
rect 14235 56467 14237 56481
rect 14237 56467 14291 56481
rect 14359 56467 14361 56481
rect 14361 56467 14415 56481
rect 14483 56467 14485 56481
rect 14485 56467 14539 56481
rect 14607 56467 14609 56481
rect 14609 56467 14663 56481
rect 14235 56425 14291 56467
rect 14359 56425 14415 56467
rect 14483 56425 14539 56467
rect 14607 56425 14663 56467
rect 12871 56301 12927 56357
rect 12995 56301 13051 56357
rect 13119 56301 13175 56357
rect 13243 56301 13299 56357
rect 13367 56301 13423 56357
rect 13491 56301 13547 56357
rect 13615 56301 13671 56357
rect 13739 56301 13795 56357
rect 13863 56301 13919 56357
rect 13987 56301 14043 56357
rect 14111 56301 14167 56357
rect 14235 56343 14237 56357
rect 14237 56343 14291 56357
rect 14359 56343 14361 56357
rect 14361 56343 14415 56357
rect 14483 56343 14485 56357
rect 14485 56343 14539 56357
rect 14607 56343 14609 56357
rect 14609 56343 14663 56357
rect 14235 56301 14291 56343
rect 14359 56301 14415 56343
rect 14483 56301 14539 56343
rect 14607 56301 14663 56343
rect 12871 56177 12927 56233
rect 12995 56177 13051 56233
rect 13119 56177 13175 56233
rect 13243 56177 13299 56233
rect 13367 56177 13423 56233
rect 13491 56177 13547 56233
rect 13615 56177 13671 56233
rect 13739 56177 13795 56233
rect 13863 56177 13919 56233
rect 13987 56177 14043 56233
rect 14111 56177 14167 56233
rect 14235 56219 14237 56233
rect 14237 56219 14291 56233
rect 14359 56219 14361 56233
rect 14361 56219 14415 56233
rect 14483 56219 14485 56233
rect 14485 56219 14539 56233
rect 14607 56219 14609 56233
rect 14609 56219 14663 56233
rect 14235 56177 14291 56219
rect 14359 56177 14415 56219
rect 14483 56177 14539 56219
rect 14607 56177 14663 56219
rect 12871 56053 12927 56109
rect 12995 56053 13051 56109
rect 13119 56053 13175 56109
rect 13243 56053 13299 56109
rect 13367 56053 13423 56109
rect 13491 56053 13547 56109
rect 13615 56053 13671 56109
rect 13739 56053 13795 56109
rect 13863 56053 13919 56109
rect 13987 56053 14043 56109
rect 14111 56053 14167 56109
rect 14235 56095 14237 56109
rect 14237 56095 14291 56109
rect 14359 56095 14361 56109
rect 14361 56095 14415 56109
rect 14483 56095 14485 56109
rect 14485 56095 14539 56109
rect 14607 56095 14609 56109
rect 14609 56095 14663 56109
rect 14235 56053 14291 56095
rect 14359 56053 14415 56095
rect 14483 56053 14539 56095
rect 14607 56053 14663 56095
rect 14902 57259 14958 57261
rect 14902 57207 14904 57259
rect 14904 57207 14956 57259
rect 14956 57207 14958 57259
rect 14902 57151 14958 57207
rect 14902 57099 14904 57151
rect 14904 57099 14956 57151
rect 14956 57099 14958 57151
rect 14902 57043 14958 57099
rect 14902 56991 14904 57043
rect 14904 56991 14956 57043
rect 14956 56991 14958 57043
rect 14902 56935 14958 56991
rect 14902 56883 14904 56935
rect 14904 56883 14956 56935
rect 14956 56883 14958 56935
rect 14902 56827 14958 56883
rect 14902 56775 14904 56827
rect 14904 56775 14956 56827
rect 14956 56775 14958 56827
rect 14902 56719 14958 56775
rect 14902 56667 14904 56719
rect 14904 56667 14956 56719
rect 14956 56667 14958 56719
rect 14902 56611 14958 56667
rect 14902 56559 14904 56611
rect 14904 56559 14956 56611
rect 14956 56559 14958 56611
rect 14902 56503 14958 56559
rect 14902 56451 14904 56503
rect 14904 56451 14956 56503
rect 14956 56451 14958 56503
rect 14902 56395 14958 56451
rect 14902 56343 14904 56395
rect 14904 56343 14956 56395
rect 14956 56343 14958 56395
rect 14902 56287 14958 56343
rect 14902 56235 14904 56287
rect 14904 56235 14956 56287
rect 14956 56235 14958 56287
rect 14902 56179 14958 56235
rect 14902 56127 14904 56179
rect 14904 56127 14956 56179
rect 14956 56127 14958 56179
rect 14902 56071 14958 56127
rect 14902 56019 14904 56071
rect 14904 56019 14956 56071
rect 14956 56019 14958 56071
rect 14902 56017 14958 56019
rect 12871 54092 12927 54148
rect 12995 54092 13051 54148
rect 13119 54092 13175 54148
rect 13243 54092 13299 54148
rect 13367 54092 13423 54148
rect 13491 54092 13547 54148
rect 13615 54092 13671 54148
rect 13739 54092 13795 54148
rect 13863 54092 13919 54148
rect 13987 54092 14043 54148
rect 14111 54092 14167 54148
rect 14235 54111 14237 54148
rect 14237 54111 14291 54148
rect 14359 54111 14361 54148
rect 14361 54111 14415 54148
rect 14483 54111 14485 54148
rect 14485 54111 14539 54148
rect 14607 54111 14609 54148
rect 14609 54111 14663 54148
rect 14235 54092 14291 54111
rect 14359 54092 14415 54111
rect 14483 54092 14539 54111
rect 14607 54092 14663 54111
rect 12871 53968 12927 54024
rect 12995 53968 13051 54024
rect 13119 53968 13175 54024
rect 13243 53968 13299 54024
rect 13367 53968 13423 54024
rect 13491 53968 13547 54024
rect 13615 53968 13671 54024
rect 13739 53968 13795 54024
rect 13863 53968 13919 54024
rect 13987 53968 14043 54024
rect 14111 53968 14167 54024
rect 14235 53987 14237 54024
rect 14237 53987 14291 54024
rect 14359 53987 14361 54024
rect 14361 53987 14415 54024
rect 14483 53987 14485 54024
rect 14485 53987 14539 54024
rect 14607 53987 14609 54024
rect 14609 53987 14663 54024
rect 14235 53968 14291 53987
rect 14359 53968 14415 53987
rect 14483 53968 14539 53987
rect 14607 53968 14663 53987
rect 12871 53844 12927 53900
rect 12995 53844 13051 53900
rect 13119 53844 13175 53900
rect 13243 53844 13299 53900
rect 13367 53844 13423 53900
rect 13491 53844 13547 53900
rect 13615 53844 13671 53900
rect 13739 53844 13795 53900
rect 13863 53844 13919 53900
rect 13987 53844 14043 53900
rect 14111 53844 14167 53900
rect 14235 53863 14237 53900
rect 14237 53863 14291 53900
rect 14359 53863 14361 53900
rect 14361 53863 14415 53900
rect 14483 53863 14485 53900
rect 14485 53863 14539 53900
rect 14607 53863 14609 53900
rect 14609 53863 14663 53900
rect 14235 53844 14291 53863
rect 14359 53844 14415 53863
rect 14483 53844 14539 53863
rect 14607 53844 14663 53863
rect 12871 53720 12927 53776
rect 12995 53720 13051 53776
rect 13119 53720 13175 53776
rect 13243 53720 13299 53776
rect 13367 53720 13423 53776
rect 13491 53720 13547 53776
rect 13615 53720 13671 53776
rect 13739 53720 13795 53776
rect 13863 53720 13919 53776
rect 13987 53720 14043 53776
rect 14111 53720 14167 53776
rect 14235 53739 14237 53776
rect 14237 53739 14291 53776
rect 14359 53739 14361 53776
rect 14361 53739 14415 53776
rect 14483 53739 14485 53776
rect 14485 53739 14539 53776
rect 14607 53739 14609 53776
rect 14609 53739 14663 53776
rect 14235 53720 14291 53739
rect 14359 53720 14415 53739
rect 14483 53720 14539 53739
rect 14607 53720 14663 53739
rect 12871 53596 12927 53652
rect 12995 53596 13051 53652
rect 13119 53596 13175 53652
rect 13243 53596 13299 53652
rect 13367 53596 13423 53652
rect 13491 53596 13547 53652
rect 13615 53596 13671 53652
rect 13739 53596 13795 53652
rect 13863 53596 13919 53652
rect 13987 53596 14043 53652
rect 14111 53596 14167 53652
rect 14235 53615 14237 53652
rect 14237 53615 14291 53652
rect 14359 53615 14361 53652
rect 14361 53615 14415 53652
rect 14483 53615 14485 53652
rect 14485 53615 14539 53652
rect 14607 53615 14609 53652
rect 14609 53615 14663 53652
rect 14235 53596 14291 53615
rect 14359 53596 14415 53615
rect 14483 53596 14539 53615
rect 14607 53596 14663 53615
rect 12871 53483 12927 53528
rect 12995 53483 13051 53528
rect 13119 53483 13175 53528
rect 13243 53483 13299 53528
rect 13367 53483 13423 53528
rect 13491 53483 13547 53528
rect 13615 53483 13671 53528
rect 13739 53483 13795 53528
rect 13863 53483 13919 53528
rect 13987 53483 14043 53528
rect 12871 53472 12921 53483
rect 12921 53472 12927 53483
rect 12995 53472 13029 53483
rect 13029 53472 13051 53483
rect 13119 53472 13137 53483
rect 13137 53472 13175 53483
rect 13243 53472 13245 53483
rect 13245 53472 13299 53483
rect 13367 53472 13409 53483
rect 13409 53472 13423 53483
rect 13491 53472 13517 53483
rect 13517 53472 13547 53483
rect 13615 53472 13625 53483
rect 13625 53472 13671 53483
rect 13739 53472 13785 53483
rect 13785 53472 13795 53483
rect 13863 53472 13893 53483
rect 13893 53472 13919 53483
rect 13987 53472 14001 53483
rect 14001 53472 14043 53483
rect 14111 53472 14167 53528
rect 14235 53491 14237 53528
rect 14237 53491 14291 53528
rect 14359 53491 14361 53528
rect 14361 53491 14415 53528
rect 14483 53491 14485 53528
rect 14485 53491 14539 53528
rect 14607 53491 14609 53528
rect 14609 53491 14663 53528
rect 14235 53472 14291 53491
rect 14359 53472 14415 53491
rect 14483 53472 14539 53491
rect 14607 53472 14663 53491
rect 12871 53375 12927 53404
rect 12995 53375 13051 53404
rect 13119 53375 13175 53404
rect 13243 53375 13299 53404
rect 13367 53375 13423 53404
rect 13491 53375 13547 53404
rect 13615 53375 13671 53404
rect 13739 53375 13795 53404
rect 13863 53375 13919 53404
rect 13987 53375 14043 53404
rect 12871 53348 12921 53375
rect 12921 53348 12927 53375
rect 12995 53348 13029 53375
rect 13029 53348 13051 53375
rect 13119 53348 13137 53375
rect 13137 53348 13175 53375
rect 13243 53348 13245 53375
rect 13245 53348 13299 53375
rect 13367 53348 13409 53375
rect 13409 53348 13423 53375
rect 13491 53348 13517 53375
rect 13517 53348 13547 53375
rect 13615 53348 13625 53375
rect 13625 53348 13671 53375
rect 13739 53348 13785 53375
rect 13785 53348 13795 53375
rect 13863 53348 13893 53375
rect 13893 53348 13919 53375
rect 13987 53348 14001 53375
rect 14001 53348 14043 53375
rect 14111 53348 14167 53404
rect 14235 53367 14237 53404
rect 14237 53367 14291 53404
rect 14359 53367 14361 53404
rect 14361 53367 14415 53404
rect 14483 53367 14485 53404
rect 14485 53367 14539 53404
rect 14607 53367 14609 53404
rect 14609 53367 14663 53404
rect 14235 53348 14291 53367
rect 14359 53348 14415 53367
rect 14483 53348 14539 53367
rect 14607 53348 14663 53367
rect 12871 53267 12927 53280
rect 12995 53267 13051 53280
rect 13119 53267 13175 53280
rect 13243 53267 13299 53280
rect 13367 53267 13423 53280
rect 13491 53267 13547 53280
rect 13615 53267 13671 53280
rect 13739 53267 13795 53280
rect 13863 53267 13919 53280
rect 13987 53267 14043 53280
rect 12871 53224 12921 53267
rect 12921 53224 12927 53267
rect 12995 53224 13029 53267
rect 13029 53224 13051 53267
rect 13119 53224 13137 53267
rect 13137 53224 13175 53267
rect 13243 53224 13245 53267
rect 13245 53224 13299 53267
rect 13367 53224 13409 53267
rect 13409 53224 13423 53267
rect 13491 53224 13517 53267
rect 13517 53224 13547 53267
rect 13615 53224 13625 53267
rect 13625 53224 13671 53267
rect 13739 53224 13785 53267
rect 13785 53224 13795 53267
rect 13863 53224 13893 53267
rect 13893 53224 13919 53267
rect 13987 53224 14001 53267
rect 14001 53224 14043 53267
rect 14111 53224 14167 53280
rect 14235 53243 14237 53280
rect 14237 53243 14291 53280
rect 14359 53243 14361 53280
rect 14361 53243 14415 53280
rect 14483 53243 14485 53280
rect 14485 53243 14539 53280
rect 14607 53243 14609 53280
rect 14609 53243 14663 53280
rect 14235 53224 14291 53243
rect 14359 53224 14415 53243
rect 14483 53224 14539 53243
rect 14607 53224 14663 53243
rect 12871 53100 12927 53156
rect 12995 53100 13051 53156
rect 13119 53100 13175 53156
rect 13243 53100 13299 53156
rect 13367 53100 13423 53156
rect 13491 53100 13547 53156
rect 13615 53100 13671 53156
rect 13739 53100 13795 53156
rect 13863 53100 13919 53156
rect 13987 53100 14043 53156
rect 14111 53100 14167 53156
rect 14235 53100 14291 53156
rect 14359 53100 14415 53156
rect 14483 53100 14539 53156
rect 14607 53100 14663 53156
rect 12871 52976 12927 53032
rect 12995 52976 13051 53032
rect 13119 52976 13175 53032
rect 13243 52976 13299 53032
rect 13367 52976 13423 53032
rect 13491 52976 13547 53032
rect 13615 52976 13671 53032
rect 13739 52976 13795 53032
rect 13863 52976 13919 53032
rect 13987 52976 14043 53032
rect 14111 52976 14167 53032
rect 14235 52976 14291 53032
rect 14359 52976 14415 53032
rect 14483 52976 14539 53032
rect 14607 52976 14663 53032
rect 12871 52852 12927 52908
rect 12995 52852 13051 52908
rect 13119 52852 13175 52908
rect 13243 52852 13299 52908
rect 13367 52852 13423 52908
rect 13491 52852 13547 52908
rect 13615 52852 13671 52908
rect 13739 52852 13795 52908
rect 13863 52852 13919 52908
rect 13987 52852 14043 52908
rect 14111 52852 14167 52908
rect 14235 52852 14291 52908
rect 14359 52852 14415 52908
rect 14483 52852 14539 52908
rect 14607 52852 14663 52908
rect 14902 54174 14958 54176
rect 14902 54122 14904 54174
rect 14904 54122 14956 54174
rect 14956 54122 14958 54174
rect 14902 54066 14958 54122
rect 14902 54014 14904 54066
rect 14904 54014 14956 54066
rect 14956 54014 14958 54066
rect 14902 53958 14958 54014
rect 14902 53906 14904 53958
rect 14904 53906 14956 53958
rect 14956 53906 14958 53958
rect 14902 53850 14958 53906
rect 14902 53798 14904 53850
rect 14904 53798 14956 53850
rect 14956 53798 14958 53850
rect 14902 53742 14958 53798
rect 14902 53690 14904 53742
rect 14904 53690 14956 53742
rect 14956 53690 14958 53742
rect 14902 53634 14958 53690
rect 14902 53582 14904 53634
rect 14904 53582 14956 53634
rect 14956 53582 14958 53634
rect 14902 53526 14958 53582
rect 14902 53474 14904 53526
rect 14904 53474 14956 53526
rect 14956 53474 14958 53526
rect 14902 53418 14958 53474
rect 14902 53366 14904 53418
rect 14904 53366 14956 53418
rect 14956 53366 14958 53418
rect 14902 53310 14958 53366
rect 14902 53258 14904 53310
rect 14904 53258 14956 53310
rect 14956 53258 14958 53310
rect 14902 53202 14958 53258
rect 14902 53150 14904 53202
rect 14904 53150 14956 53202
rect 14956 53150 14958 53202
rect 14902 53094 14958 53150
rect 14902 53042 14904 53094
rect 14904 53042 14956 53094
rect 14956 53042 14958 53094
rect 14902 52986 14958 53042
rect 14902 52934 14904 52986
rect 14904 52934 14956 52986
rect 14956 52934 14958 52986
rect 14902 52878 14958 52934
rect 14902 52826 14904 52878
rect 14904 52826 14956 52878
rect 14956 52826 14958 52878
rect 14902 52824 14958 52826
rect 12871 52492 12927 52548
rect 12995 52492 13051 52548
rect 13119 52492 13175 52548
rect 13243 52492 13299 52548
rect 13367 52492 13423 52548
rect 13491 52492 13547 52548
rect 13615 52492 13671 52548
rect 13739 52492 13795 52548
rect 13863 52492 13919 52548
rect 13987 52492 14043 52548
rect 14111 52492 14167 52548
rect 14235 52492 14291 52548
rect 14359 52492 14415 52548
rect 14483 52492 14539 52548
rect 14607 52492 14663 52548
rect 12871 52368 12927 52424
rect 12995 52368 13051 52424
rect 13119 52368 13175 52424
rect 13243 52368 13299 52424
rect 13367 52368 13423 52424
rect 13491 52368 13547 52424
rect 13615 52368 13671 52424
rect 13739 52368 13795 52424
rect 13863 52368 13919 52424
rect 13987 52368 14043 52424
rect 14111 52368 14167 52424
rect 14235 52368 14291 52424
rect 14359 52368 14415 52424
rect 14483 52368 14539 52424
rect 14607 52368 14663 52424
rect 12871 52244 12927 52300
rect 12995 52244 13051 52300
rect 13119 52244 13175 52300
rect 13243 52244 13299 52300
rect 13367 52244 13423 52300
rect 13491 52244 13547 52300
rect 13615 52244 13671 52300
rect 13739 52244 13795 52300
rect 13863 52244 13919 52300
rect 13987 52244 14043 52300
rect 14111 52244 14167 52300
rect 14235 52244 14291 52300
rect 14359 52244 14415 52300
rect 14483 52244 14539 52300
rect 14607 52244 14663 52300
rect 12871 52120 12927 52176
rect 12995 52120 13051 52176
rect 13119 52120 13175 52176
rect 13243 52120 13299 52176
rect 13367 52120 13423 52176
rect 13491 52120 13547 52176
rect 13615 52120 13671 52176
rect 13739 52120 13795 52176
rect 13863 52120 13919 52176
rect 13987 52120 14043 52176
rect 14111 52120 14167 52176
rect 14235 52120 14291 52176
rect 14359 52120 14415 52176
rect 14483 52120 14539 52176
rect 14607 52120 14663 52176
rect 12871 51996 12927 52052
rect 12995 51996 13051 52052
rect 13119 51996 13175 52052
rect 13243 51996 13299 52052
rect 13367 51996 13423 52052
rect 13491 51996 13547 52052
rect 13615 51996 13671 52052
rect 13739 51996 13795 52052
rect 13863 51996 13919 52052
rect 13987 51996 14043 52052
rect 14111 51996 14167 52052
rect 14235 51996 14291 52052
rect 14359 51996 14415 52052
rect 14483 51996 14539 52052
rect 14607 51996 14663 52052
rect 12871 51872 12927 51928
rect 12995 51872 13051 51928
rect 13119 51872 13175 51928
rect 13243 51872 13299 51928
rect 13367 51872 13423 51928
rect 13491 51872 13547 51928
rect 13615 51872 13671 51928
rect 13739 51872 13795 51928
rect 13863 51872 13919 51928
rect 13987 51872 14043 51928
rect 14111 51872 14167 51928
rect 14235 51872 14291 51928
rect 14359 51872 14415 51928
rect 14483 51872 14539 51928
rect 14607 51872 14663 51928
rect 12871 51748 12927 51804
rect 12995 51748 13051 51804
rect 13119 51748 13175 51804
rect 13243 51748 13299 51804
rect 13367 51748 13423 51804
rect 13491 51748 13547 51804
rect 13615 51748 13671 51804
rect 13739 51748 13795 51804
rect 13863 51748 13919 51804
rect 13987 51748 14043 51804
rect 14111 51748 14167 51804
rect 14235 51748 14291 51804
rect 14359 51748 14415 51804
rect 14483 51748 14539 51804
rect 14607 51748 14663 51804
rect 12871 51624 12927 51680
rect 12995 51624 13051 51680
rect 13119 51624 13175 51680
rect 13243 51624 13299 51680
rect 13367 51624 13423 51680
rect 13491 51624 13547 51680
rect 13615 51624 13671 51680
rect 13739 51624 13795 51680
rect 13863 51624 13919 51680
rect 13987 51624 14043 51680
rect 14111 51624 14167 51680
rect 14235 51624 14291 51680
rect 14359 51624 14415 51680
rect 14483 51624 14539 51680
rect 14607 51624 14663 51680
rect 12871 51500 12927 51556
rect 12995 51500 13051 51556
rect 13119 51500 13175 51556
rect 13243 51500 13299 51556
rect 13367 51500 13423 51556
rect 13491 51500 13547 51556
rect 13615 51500 13671 51556
rect 13739 51500 13795 51556
rect 13863 51500 13919 51556
rect 13987 51500 14043 51556
rect 14111 51500 14167 51556
rect 14235 51500 14291 51556
rect 14359 51500 14415 51556
rect 14483 51500 14539 51556
rect 14607 51500 14663 51556
rect 12871 51376 12927 51432
rect 12995 51376 13051 51432
rect 13119 51376 13175 51432
rect 13243 51376 13299 51432
rect 13367 51376 13423 51432
rect 13491 51376 13547 51432
rect 13615 51376 13671 51432
rect 13739 51376 13795 51432
rect 13863 51376 13919 51432
rect 13987 51376 14043 51432
rect 14111 51376 14167 51432
rect 14235 51376 14291 51432
rect 14359 51376 14415 51432
rect 14483 51376 14539 51432
rect 14607 51376 14663 51432
rect 12871 51252 12927 51308
rect 12995 51252 13051 51308
rect 13119 51252 13175 51308
rect 13243 51252 13299 51308
rect 13367 51252 13423 51308
rect 13491 51252 13547 51308
rect 13615 51252 13671 51308
rect 13739 51252 13795 51308
rect 13863 51252 13919 51308
rect 13987 51252 14043 51308
rect 14111 51252 14167 51308
rect 14235 51252 14291 51308
rect 14359 51252 14415 51308
rect 14483 51252 14539 51308
rect 14607 51252 14663 51308
rect 14902 52574 14958 52576
rect 14902 52522 14904 52574
rect 14904 52522 14956 52574
rect 14956 52522 14958 52574
rect 14902 52466 14958 52522
rect 14902 52414 14904 52466
rect 14904 52414 14956 52466
rect 14956 52414 14958 52466
rect 14902 52358 14958 52414
rect 14902 52306 14904 52358
rect 14904 52306 14956 52358
rect 14956 52306 14958 52358
rect 14902 52250 14958 52306
rect 14902 52198 14904 52250
rect 14904 52198 14956 52250
rect 14956 52198 14958 52250
rect 14902 52142 14958 52198
rect 14902 52090 14904 52142
rect 14904 52090 14956 52142
rect 14956 52090 14958 52142
rect 14902 52034 14958 52090
rect 14902 51982 14904 52034
rect 14904 51982 14956 52034
rect 14956 51982 14958 52034
rect 14902 51926 14958 51982
rect 14902 51874 14904 51926
rect 14904 51874 14956 51926
rect 14956 51874 14958 51926
rect 14902 51818 14958 51874
rect 14902 51766 14904 51818
rect 14904 51766 14956 51818
rect 14956 51766 14958 51818
rect 14902 51710 14958 51766
rect 14902 51658 14904 51710
rect 14904 51658 14956 51710
rect 14956 51658 14958 51710
rect 14902 51602 14958 51658
rect 14902 51550 14904 51602
rect 14904 51550 14956 51602
rect 14956 51550 14958 51602
rect 14902 51494 14958 51550
rect 14902 51442 14904 51494
rect 14904 51442 14956 51494
rect 14956 51442 14958 51494
rect 14902 51386 14958 51442
rect 14902 51334 14904 51386
rect 14904 51334 14956 51386
rect 14956 51334 14958 51386
rect 14902 51278 14958 51334
rect 14902 51226 14904 51278
rect 14904 51226 14956 51278
rect 14956 51226 14958 51278
rect 14902 51224 14958 51226
rect 12871 49292 12927 49348
rect 12995 49292 13051 49348
rect 13119 49292 13175 49348
rect 13243 49292 13299 49348
rect 13367 49292 13423 49348
rect 13491 49292 13547 49348
rect 13615 49292 13671 49348
rect 13739 49292 13795 49348
rect 13863 49292 13919 49348
rect 13987 49292 14043 49348
rect 14111 49292 14167 49348
rect 14235 49292 14291 49348
rect 14359 49292 14415 49348
rect 14483 49292 14539 49348
rect 14607 49292 14663 49348
rect 12871 49168 12927 49224
rect 12995 49168 13051 49224
rect 13119 49168 13175 49224
rect 13243 49168 13299 49224
rect 13367 49168 13423 49224
rect 13491 49168 13547 49224
rect 13615 49168 13671 49224
rect 13739 49168 13795 49224
rect 13863 49168 13919 49224
rect 13987 49168 14043 49224
rect 14111 49168 14167 49224
rect 14235 49168 14291 49224
rect 14359 49168 14415 49224
rect 14483 49168 14539 49224
rect 14607 49168 14663 49224
rect 12871 49044 12927 49100
rect 12995 49044 13051 49100
rect 13119 49044 13175 49100
rect 13243 49044 13299 49100
rect 13367 49044 13423 49100
rect 13491 49044 13547 49100
rect 13615 49044 13671 49100
rect 13739 49044 13795 49100
rect 13863 49044 13919 49100
rect 13987 49044 14043 49100
rect 14111 49044 14167 49100
rect 14235 49044 14291 49100
rect 14359 49044 14415 49100
rect 14483 49044 14539 49100
rect 14607 49044 14663 49100
rect 12871 48920 12927 48976
rect 12995 48920 13051 48976
rect 13119 48920 13175 48976
rect 13243 48920 13299 48976
rect 13367 48920 13423 48976
rect 13491 48920 13547 48976
rect 13615 48920 13671 48976
rect 13739 48920 13795 48976
rect 13863 48920 13919 48976
rect 13987 48920 14043 48976
rect 14111 48920 14167 48976
rect 14235 48920 14291 48976
rect 14359 48920 14415 48976
rect 14483 48920 14539 48976
rect 14607 48920 14663 48976
rect 12871 48796 12927 48852
rect 12995 48796 13051 48852
rect 13119 48796 13175 48852
rect 13243 48796 13299 48852
rect 13367 48796 13423 48852
rect 13491 48796 13547 48852
rect 13615 48796 13671 48852
rect 13739 48796 13795 48852
rect 13863 48796 13919 48852
rect 13987 48796 14043 48852
rect 14111 48796 14167 48852
rect 14235 48796 14291 48852
rect 14359 48796 14415 48852
rect 14483 48796 14539 48852
rect 14607 48796 14663 48852
rect 12871 48672 12927 48728
rect 12995 48672 13051 48728
rect 13119 48672 13175 48728
rect 13243 48672 13299 48728
rect 13367 48672 13423 48728
rect 13491 48672 13547 48728
rect 13615 48672 13671 48728
rect 13739 48672 13795 48728
rect 13863 48672 13919 48728
rect 13987 48672 14043 48728
rect 14111 48672 14167 48728
rect 14235 48672 14291 48728
rect 14359 48672 14415 48728
rect 14483 48672 14539 48728
rect 14607 48672 14663 48728
rect 12871 48548 12927 48604
rect 12995 48548 13051 48604
rect 13119 48548 13175 48604
rect 13243 48548 13299 48604
rect 13367 48548 13423 48604
rect 13491 48548 13547 48604
rect 13615 48548 13671 48604
rect 13739 48548 13795 48604
rect 13863 48548 13919 48604
rect 13987 48548 14043 48604
rect 14111 48548 14167 48604
rect 14235 48548 14291 48604
rect 14359 48548 14415 48604
rect 14483 48548 14539 48604
rect 14607 48548 14663 48604
rect 12871 48424 12927 48480
rect 12995 48424 13051 48480
rect 13119 48424 13175 48480
rect 13243 48424 13299 48480
rect 13367 48424 13423 48480
rect 13491 48424 13547 48480
rect 13615 48424 13671 48480
rect 13739 48424 13795 48480
rect 13863 48424 13919 48480
rect 13987 48424 14043 48480
rect 14111 48424 14167 48480
rect 14235 48424 14291 48480
rect 14359 48424 14415 48480
rect 14483 48424 14539 48480
rect 14607 48424 14663 48480
rect 12871 48300 12927 48356
rect 12995 48300 13051 48356
rect 13119 48300 13175 48356
rect 13243 48300 13299 48356
rect 13367 48300 13423 48356
rect 13491 48300 13547 48356
rect 13615 48300 13671 48356
rect 13739 48300 13795 48356
rect 13863 48300 13919 48356
rect 13987 48300 14043 48356
rect 14111 48300 14167 48356
rect 14235 48300 14291 48356
rect 14359 48300 14415 48356
rect 14483 48300 14539 48356
rect 14607 48300 14663 48356
rect 12871 48176 12927 48232
rect 12995 48176 13051 48232
rect 13119 48176 13175 48232
rect 13243 48176 13299 48232
rect 13367 48176 13423 48232
rect 13491 48176 13547 48232
rect 13615 48176 13671 48232
rect 13739 48176 13795 48232
rect 13863 48176 13919 48232
rect 13987 48176 14043 48232
rect 14111 48176 14167 48232
rect 14235 48176 14291 48232
rect 14359 48176 14415 48232
rect 14483 48176 14539 48232
rect 14607 48176 14663 48232
rect 12871 48052 12927 48108
rect 12995 48052 13051 48108
rect 13119 48052 13175 48108
rect 13243 48052 13299 48108
rect 13367 48052 13423 48108
rect 13491 48052 13547 48108
rect 13615 48052 13671 48108
rect 13739 48052 13795 48108
rect 13863 48052 13919 48108
rect 13987 48052 14043 48108
rect 14111 48052 14167 48108
rect 14235 48052 14291 48108
rect 14359 48052 14415 48108
rect 14483 48052 14539 48108
rect 14607 48052 14663 48108
rect 14902 49374 14958 49376
rect 14902 49322 14904 49374
rect 14904 49322 14956 49374
rect 14956 49322 14958 49374
rect 14902 49266 14958 49322
rect 14902 49214 14904 49266
rect 14904 49214 14956 49266
rect 14956 49214 14958 49266
rect 14902 49158 14958 49214
rect 14902 49106 14904 49158
rect 14904 49106 14956 49158
rect 14956 49106 14958 49158
rect 14902 49050 14958 49106
rect 14902 48998 14904 49050
rect 14904 48998 14956 49050
rect 14956 48998 14958 49050
rect 14902 48942 14958 48998
rect 14902 48890 14904 48942
rect 14904 48890 14956 48942
rect 14956 48890 14958 48942
rect 14902 48834 14958 48890
rect 14902 48782 14904 48834
rect 14904 48782 14956 48834
rect 14956 48782 14958 48834
rect 14902 48726 14958 48782
rect 14902 48674 14904 48726
rect 14904 48674 14956 48726
rect 14956 48674 14958 48726
rect 14902 48618 14958 48674
rect 14902 48566 14904 48618
rect 14904 48566 14956 48618
rect 14956 48566 14958 48618
rect 14902 48510 14958 48566
rect 14902 48458 14904 48510
rect 14904 48458 14956 48510
rect 14956 48458 14958 48510
rect 14902 48402 14958 48458
rect 14902 48350 14904 48402
rect 14904 48350 14956 48402
rect 14956 48350 14958 48402
rect 14902 48294 14958 48350
rect 14902 48242 14904 48294
rect 14904 48242 14956 48294
rect 14956 48242 14958 48294
rect 14902 48186 14958 48242
rect 14902 48134 14904 48186
rect 14904 48134 14956 48186
rect 14956 48134 14958 48186
rect 14902 48078 14958 48134
rect 14902 48026 14904 48078
rect 14904 48026 14956 48078
rect 14956 48026 14958 48078
rect 14902 48024 14958 48026
rect 12307 47072 12363 47128
rect 12431 47072 12487 47128
rect 12307 46948 12363 47004
rect 12431 46948 12487 47004
rect 12307 46824 12363 46880
rect 12431 46824 12487 46880
rect 12307 46700 12363 46756
rect 12431 46700 12487 46756
rect 12307 46576 12363 46632
rect 12431 46576 12487 46632
rect 12307 46452 12363 46508
rect 12431 46452 12487 46508
rect 2808 46092 2864 46148
rect 2932 46092 2988 46148
rect 3056 46092 3112 46148
rect 3180 46092 3236 46148
rect 3304 46092 3360 46148
rect 3428 46092 3484 46148
rect 3552 46092 3608 46148
rect 3676 46092 3732 46148
rect 3800 46092 3856 46148
rect 3924 46092 3980 46148
rect 4048 46092 4104 46148
rect 4172 46092 4228 46148
rect 4296 46092 4352 46148
rect 4420 46092 4476 46148
rect 4544 46092 4600 46148
rect 4668 46092 4724 46148
rect 2808 45968 2864 46024
rect 2932 45968 2988 46024
rect 3056 45968 3112 46024
rect 3180 45968 3236 46024
rect 3304 45968 3360 46024
rect 3428 45968 3484 46024
rect 3552 45968 3608 46024
rect 3676 45968 3732 46024
rect 3800 45968 3856 46024
rect 3924 45968 3980 46024
rect 4048 45968 4104 46024
rect 4172 45968 4228 46024
rect 4296 45968 4352 46024
rect 4420 45968 4476 46024
rect 4544 45968 4600 46024
rect 4668 45968 4724 46024
rect 2808 45844 2864 45900
rect 2932 45844 2988 45900
rect 3056 45844 3112 45900
rect 3180 45844 3236 45900
rect 3304 45844 3360 45900
rect 3428 45844 3484 45900
rect 3552 45844 3608 45900
rect 3676 45844 3732 45900
rect 3800 45844 3856 45900
rect 3924 45844 3980 45900
rect 4048 45844 4104 45900
rect 4172 45844 4228 45900
rect 4296 45844 4352 45900
rect 4420 45844 4476 45900
rect 4544 45844 4600 45900
rect 4668 45844 4724 45900
rect 2808 45720 2864 45776
rect 2932 45720 2988 45776
rect 3056 45720 3112 45776
rect 3180 45720 3236 45776
rect 3304 45720 3360 45776
rect 3428 45720 3484 45776
rect 3552 45720 3608 45776
rect 3676 45720 3732 45776
rect 3800 45720 3856 45776
rect 3924 45720 3980 45776
rect 4048 45720 4104 45776
rect 4172 45720 4228 45776
rect 4296 45720 4352 45776
rect 4420 45720 4476 45776
rect 4544 45720 4600 45776
rect 4668 45720 4724 45776
rect 2808 45596 2864 45652
rect 2932 45596 2988 45652
rect 3056 45596 3112 45652
rect 3180 45596 3236 45652
rect 3304 45596 3360 45652
rect 3428 45596 3484 45652
rect 3552 45596 3608 45652
rect 3676 45596 3732 45652
rect 3800 45596 3856 45652
rect 3924 45596 3980 45652
rect 4048 45596 4104 45652
rect 4172 45596 4228 45652
rect 4296 45596 4352 45652
rect 4420 45596 4476 45652
rect 4544 45596 4600 45652
rect 4668 45596 4724 45652
rect 2808 45472 2864 45528
rect 2932 45472 2988 45528
rect 3056 45472 3112 45528
rect 3180 45472 3236 45528
rect 3304 45472 3360 45528
rect 3428 45472 3484 45528
rect 3552 45472 3608 45528
rect 3676 45472 3732 45528
rect 3800 45472 3856 45528
rect 3924 45472 3980 45528
rect 4048 45472 4104 45528
rect 4172 45472 4228 45528
rect 4296 45472 4352 45528
rect 4420 45472 4476 45528
rect 4544 45472 4600 45528
rect 4668 45472 4724 45528
rect 2808 45348 2864 45404
rect 2932 45348 2988 45404
rect 3056 45348 3112 45404
rect 3180 45348 3236 45404
rect 3304 45348 3360 45404
rect 3428 45348 3484 45404
rect 3552 45348 3608 45404
rect 3676 45348 3732 45404
rect 3800 45348 3856 45404
rect 3924 45348 3980 45404
rect 4048 45348 4104 45404
rect 4172 45348 4228 45404
rect 4296 45348 4352 45404
rect 4420 45348 4476 45404
rect 4544 45348 4600 45404
rect 4668 45348 4724 45404
rect 2808 45224 2864 45280
rect 2932 45224 2988 45280
rect 3056 45224 3112 45280
rect 3180 45224 3236 45280
rect 3304 45224 3360 45280
rect 3428 45224 3484 45280
rect 3552 45224 3608 45280
rect 3676 45224 3732 45280
rect 3800 45224 3856 45280
rect 3924 45224 3980 45280
rect 4048 45224 4104 45280
rect 4172 45224 4228 45280
rect 4296 45224 4352 45280
rect 4420 45224 4476 45280
rect 4544 45224 4600 45280
rect 4668 45224 4724 45280
rect 2808 45100 2864 45156
rect 2932 45100 2988 45156
rect 3056 45100 3112 45156
rect 3180 45100 3236 45156
rect 3304 45100 3360 45156
rect 3428 45100 3484 45156
rect 3552 45100 3608 45156
rect 3676 45100 3732 45156
rect 3800 45100 3856 45156
rect 3924 45100 3980 45156
rect 4048 45100 4104 45156
rect 4172 45100 4228 45156
rect 4296 45100 4352 45156
rect 4420 45100 4476 45156
rect 4544 45100 4600 45156
rect 4668 45100 4724 45156
rect 2808 44976 2864 45032
rect 2932 44976 2988 45032
rect 3056 44976 3112 45032
rect 3180 44976 3236 45032
rect 3304 44976 3360 45032
rect 3428 44976 3484 45032
rect 3552 44976 3608 45032
rect 3676 44976 3732 45032
rect 3800 44976 3856 45032
rect 3924 44976 3980 45032
rect 4048 44976 4104 45032
rect 4172 44976 4228 45032
rect 4296 44976 4352 45032
rect 4420 44976 4476 45032
rect 4544 44976 4600 45032
rect 4668 44976 4724 45032
rect 2808 44852 2864 44908
rect 2932 44852 2988 44908
rect 3056 44852 3112 44908
rect 3180 44852 3236 44908
rect 3304 44852 3360 44908
rect 3428 44852 3484 44908
rect 3552 44852 3608 44908
rect 3676 44852 3732 44908
rect 3800 44852 3856 44908
rect 3924 44852 3980 44908
rect 4048 44852 4104 44908
rect 4172 44852 4228 44908
rect 4296 44852 4352 44908
rect 4420 44852 4476 44908
rect 4544 44852 4600 44908
rect 4668 44852 4724 44908
rect 5178 46092 5234 46148
rect 5302 46092 5358 46148
rect 5426 46092 5482 46148
rect 5550 46092 5606 46148
rect 5674 46092 5730 46148
rect 5798 46092 5854 46148
rect 5922 46092 5978 46148
rect 6046 46092 6102 46148
rect 6170 46092 6226 46148
rect 6294 46092 6350 46148
rect 6418 46092 6474 46148
rect 6542 46092 6598 46148
rect 6666 46092 6722 46148
rect 6790 46092 6846 46148
rect 6914 46092 6970 46148
rect 7038 46092 7094 46148
rect 5178 45968 5234 46024
rect 5302 45968 5358 46024
rect 5426 45968 5482 46024
rect 5550 45968 5606 46024
rect 5674 45968 5730 46024
rect 5798 45968 5854 46024
rect 5922 45968 5978 46024
rect 6046 45968 6102 46024
rect 6170 45968 6226 46024
rect 6294 45968 6350 46024
rect 6418 45968 6474 46024
rect 6542 45968 6598 46024
rect 6666 45968 6722 46024
rect 6790 45968 6846 46024
rect 6914 45968 6970 46024
rect 7038 45968 7094 46024
rect 5178 45844 5234 45900
rect 5302 45844 5358 45900
rect 5426 45844 5482 45900
rect 5550 45844 5606 45900
rect 5674 45844 5730 45900
rect 5798 45844 5854 45900
rect 5922 45844 5978 45900
rect 6046 45844 6102 45900
rect 6170 45844 6226 45900
rect 6294 45844 6350 45900
rect 6418 45844 6474 45900
rect 6542 45844 6598 45900
rect 6666 45844 6722 45900
rect 6790 45844 6846 45900
rect 6914 45844 6970 45900
rect 7038 45844 7094 45900
rect 5178 45720 5234 45776
rect 5302 45720 5358 45776
rect 5426 45720 5482 45776
rect 5550 45720 5606 45776
rect 5674 45720 5730 45776
rect 5798 45720 5854 45776
rect 5922 45720 5978 45776
rect 6046 45720 6102 45776
rect 6170 45720 6226 45776
rect 6294 45720 6350 45776
rect 6418 45720 6474 45776
rect 6542 45720 6598 45776
rect 6666 45720 6722 45776
rect 6790 45720 6846 45776
rect 6914 45720 6970 45776
rect 7038 45720 7094 45776
rect 5178 45596 5234 45652
rect 5302 45596 5358 45652
rect 5426 45596 5482 45652
rect 5550 45596 5606 45652
rect 5674 45596 5730 45652
rect 5798 45596 5854 45652
rect 5922 45596 5978 45652
rect 6046 45596 6102 45652
rect 6170 45596 6226 45652
rect 6294 45596 6350 45652
rect 6418 45596 6474 45652
rect 6542 45596 6598 45652
rect 6666 45596 6722 45652
rect 6790 45596 6846 45652
rect 6914 45596 6970 45652
rect 7038 45596 7094 45652
rect 5178 45472 5234 45528
rect 5302 45472 5358 45528
rect 5426 45472 5482 45528
rect 5550 45472 5606 45528
rect 5674 45472 5730 45528
rect 5798 45472 5854 45528
rect 5922 45472 5978 45528
rect 6046 45472 6102 45528
rect 6170 45472 6226 45528
rect 6294 45472 6350 45528
rect 6418 45472 6474 45528
rect 6542 45472 6598 45528
rect 6666 45472 6722 45528
rect 6790 45472 6846 45528
rect 6914 45472 6970 45528
rect 7038 45472 7094 45528
rect 5178 45348 5234 45404
rect 5302 45348 5358 45404
rect 5426 45348 5482 45404
rect 5550 45348 5606 45404
rect 5674 45348 5730 45404
rect 5798 45348 5854 45404
rect 5922 45348 5978 45404
rect 6046 45348 6102 45404
rect 6170 45348 6226 45404
rect 6294 45348 6350 45404
rect 6418 45348 6474 45404
rect 6542 45348 6598 45404
rect 6666 45348 6722 45404
rect 6790 45348 6846 45404
rect 6914 45348 6970 45404
rect 7038 45348 7094 45404
rect 5178 45224 5234 45280
rect 5302 45224 5358 45280
rect 5426 45224 5482 45280
rect 5550 45224 5606 45280
rect 5674 45224 5730 45280
rect 5798 45224 5854 45280
rect 5922 45224 5978 45280
rect 6046 45224 6102 45280
rect 6170 45224 6226 45280
rect 6294 45224 6350 45280
rect 6418 45224 6474 45280
rect 6542 45224 6598 45280
rect 6666 45224 6722 45280
rect 6790 45224 6846 45280
rect 6914 45224 6970 45280
rect 7038 45224 7094 45280
rect 5178 45100 5234 45156
rect 5302 45100 5358 45156
rect 5426 45100 5482 45156
rect 5550 45100 5606 45156
rect 5674 45100 5730 45156
rect 5798 45100 5854 45156
rect 5922 45100 5978 45156
rect 6046 45100 6102 45156
rect 6170 45100 6226 45156
rect 6294 45100 6350 45156
rect 6418 45100 6474 45156
rect 6542 45100 6598 45156
rect 6666 45100 6722 45156
rect 6790 45100 6846 45156
rect 6914 45100 6970 45156
rect 7038 45100 7094 45156
rect 5178 44976 5234 45032
rect 5302 44976 5358 45032
rect 5426 44976 5482 45032
rect 5550 44976 5606 45032
rect 5674 44976 5730 45032
rect 5798 44976 5854 45032
rect 5922 44976 5978 45032
rect 6046 44976 6102 45032
rect 6170 44976 6226 45032
rect 6294 44976 6350 45032
rect 6418 44976 6474 45032
rect 6542 44976 6598 45032
rect 6666 44976 6722 45032
rect 6790 44976 6846 45032
rect 6914 44976 6970 45032
rect 7038 44976 7094 45032
rect 5178 44852 5234 44908
rect 5302 44852 5358 44908
rect 5426 44852 5482 44908
rect 5550 44852 5606 44908
rect 5674 44852 5730 44908
rect 5798 44852 5854 44908
rect 5922 44852 5978 44908
rect 6046 44852 6102 44908
rect 6170 44852 6226 44908
rect 6294 44852 6350 44908
rect 6418 44852 6474 44908
rect 6542 44852 6598 44908
rect 6666 44852 6722 44908
rect 6790 44852 6846 44908
rect 6914 44852 6970 44908
rect 7038 44852 7094 44908
rect 7884 46092 7940 46148
rect 8008 46092 8064 46148
rect 8132 46092 8188 46148
rect 8256 46092 8312 46148
rect 8380 46092 8436 46148
rect 8504 46092 8560 46148
rect 8628 46092 8684 46148
rect 8752 46092 8808 46148
rect 8876 46092 8932 46148
rect 9000 46092 9056 46148
rect 9124 46092 9180 46148
rect 9248 46092 9304 46148
rect 9372 46092 9428 46148
rect 9496 46092 9552 46148
rect 9620 46092 9676 46148
rect 9744 46092 9800 46148
rect 7884 45968 7940 46024
rect 8008 45968 8064 46024
rect 8132 45968 8188 46024
rect 8256 45968 8312 46024
rect 8380 45968 8436 46024
rect 8504 45968 8560 46024
rect 8628 45968 8684 46024
rect 8752 45968 8808 46024
rect 8876 45968 8932 46024
rect 9000 45968 9056 46024
rect 9124 45968 9180 46024
rect 9248 45968 9304 46024
rect 9372 45968 9428 46024
rect 9496 45968 9552 46024
rect 9620 45968 9676 46024
rect 9744 45968 9800 46024
rect 7884 45844 7940 45900
rect 8008 45844 8064 45900
rect 8132 45844 8188 45900
rect 8256 45844 8312 45900
rect 8380 45844 8436 45900
rect 8504 45844 8560 45900
rect 8628 45844 8684 45900
rect 8752 45844 8808 45900
rect 8876 45844 8932 45900
rect 9000 45844 9056 45900
rect 9124 45844 9180 45900
rect 9248 45844 9304 45900
rect 9372 45844 9428 45900
rect 9496 45844 9552 45900
rect 9620 45844 9676 45900
rect 9744 45844 9800 45900
rect 7884 45720 7940 45776
rect 8008 45720 8064 45776
rect 8132 45720 8188 45776
rect 8256 45720 8312 45776
rect 8380 45720 8436 45776
rect 8504 45720 8560 45776
rect 8628 45720 8684 45776
rect 8752 45720 8808 45776
rect 8876 45720 8932 45776
rect 9000 45720 9056 45776
rect 9124 45720 9180 45776
rect 9248 45720 9304 45776
rect 9372 45720 9428 45776
rect 9496 45720 9552 45776
rect 9620 45720 9676 45776
rect 9744 45720 9800 45776
rect 7884 45596 7940 45652
rect 8008 45596 8064 45652
rect 8132 45596 8188 45652
rect 8256 45596 8312 45652
rect 8380 45596 8436 45652
rect 8504 45596 8560 45652
rect 8628 45596 8684 45652
rect 8752 45596 8808 45652
rect 8876 45596 8932 45652
rect 9000 45596 9056 45652
rect 9124 45596 9180 45652
rect 9248 45596 9304 45652
rect 9372 45596 9428 45652
rect 9496 45596 9552 45652
rect 9620 45596 9676 45652
rect 9744 45596 9800 45652
rect 7884 45472 7940 45528
rect 8008 45472 8064 45528
rect 8132 45472 8188 45528
rect 8256 45472 8312 45528
rect 8380 45472 8436 45528
rect 8504 45472 8560 45528
rect 8628 45472 8684 45528
rect 8752 45472 8808 45528
rect 8876 45472 8932 45528
rect 9000 45472 9056 45528
rect 9124 45472 9180 45528
rect 9248 45472 9304 45528
rect 9372 45472 9428 45528
rect 9496 45472 9552 45528
rect 9620 45472 9676 45528
rect 9744 45472 9800 45528
rect 7884 45348 7940 45404
rect 8008 45348 8064 45404
rect 8132 45348 8188 45404
rect 8256 45348 8312 45404
rect 8380 45348 8436 45404
rect 8504 45348 8560 45404
rect 8628 45348 8684 45404
rect 8752 45348 8808 45404
rect 8876 45348 8932 45404
rect 9000 45348 9056 45404
rect 9124 45348 9180 45404
rect 9248 45348 9304 45404
rect 9372 45348 9428 45404
rect 9496 45348 9552 45404
rect 9620 45348 9676 45404
rect 9744 45348 9800 45404
rect 7884 45224 7940 45280
rect 8008 45224 8064 45280
rect 8132 45224 8188 45280
rect 8256 45224 8312 45280
rect 8380 45224 8436 45280
rect 8504 45224 8560 45280
rect 8628 45224 8684 45280
rect 8752 45224 8808 45280
rect 8876 45224 8932 45280
rect 9000 45224 9056 45280
rect 9124 45224 9180 45280
rect 9248 45224 9304 45280
rect 9372 45224 9428 45280
rect 9496 45224 9552 45280
rect 9620 45224 9676 45280
rect 9744 45224 9800 45280
rect 7884 45100 7940 45156
rect 8008 45100 8064 45156
rect 8132 45100 8188 45156
rect 8256 45100 8312 45156
rect 8380 45100 8436 45156
rect 8504 45100 8560 45156
rect 8628 45100 8684 45156
rect 8752 45100 8808 45156
rect 8876 45100 8932 45156
rect 9000 45100 9056 45156
rect 9124 45100 9180 45156
rect 9248 45100 9304 45156
rect 9372 45100 9428 45156
rect 9496 45100 9552 45156
rect 9620 45100 9676 45156
rect 9744 45100 9800 45156
rect 7884 44976 7940 45032
rect 8008 44976 8064 45032
rect 8132 44976 8188 45032
rect 8256 44976 8312 45032
rect 8380 44976 8436 45032
rect 8504 44976 8560 45032
rect 8628 44976 8684 45032
rect 8752 44976 8808 45032
rect 8876 44976 8932 45032
rect 9000 44976 9056 45032
rect 9124 44976 9180 45032
rect 9248 44976 9304 45032
rect 9372 44976 9428 45032
rect 9496 44976 9552 45032
rect 9620 44976 9676 45032
rect 9744 44976 9800 45032
rect 7884 44852 7940 44908
rect 8008 44852 8064 44908
rect 8132 44852 8188 44908
rect 8256 44852 8312 44908
rect 8380 44852 8436 44908
rect 8504 44852 8560 44908
rect 8628 44852 8684 44908
rect 8752 44852 8808 44908
rect 8876 44852 8932 44908
rect 9000 44852 9056 44908
rect 9124 44852 9180 44908
rect 9248 44852 9304 44908
rect 9372 44852 9428 44908
rect 9496 44852 9552 44908
rect 9620 44852 9676 44908
rect 9744 44852 9800 44908
rect 10254 46092 10310 46148
rect 10378 46092 10434 46148
rect 10502 46092 10558 46148
rect 10626 46092 10682 46148
rect 10750 46092 10806 46148
rect 10874 46092 10930 46148
rect 10998 46092 11054 46148
rect 11122 46092 11178 46148
rect 11246 46092 11302 46148
rect 11370 46092 11426 46148
rect 11494 46092 11550 46148
rect 11618 46092 11674 46148
rect 11742 46092 11798 46148
rect 11866 46092 11922 46148
rect 11990 46092 12046 46148
rect 12114 46092 12170 46148
rect 10254 45968 10310 46024
rect 10378 45968 10434 46024
rect 10502 45968 10558 46024
rect 10626 45968 10682 46024
rect 10750 45968 10806 46024
rect 10874 45968 10930 46024
rect 10998 45968 11054 46024
rect 11122 45968 11178 46024
rect 11246 45968 11302 46024
rect 11370 45968 11426 46024
rect 11494 45968 11550 46024
rect 11618 45968 11674 46024
rect 11742 45968 11798 46024
rect 11866 45968 11922 46024
rect 11990 45968 12046 46024
rect 12114 45968 12170 46024
rect 10254 45844 10310 45900
rect 10378 45844 10434 45900
rect 10502 45844 10558 45900
rect 10626 45844 10682 45900
rect 10750 45844 10806 45900
rect 10874 45844 10930 45900
rect 10998 45844 11054 45900
rect 11122 45844 11178 45900
rect 11246 45844 11302 45900
rect 11370 45844 11426 45900
rect 11494 45844 11550 45900
rect 11618 45844 11674 45900
rect 11742 45844 11798 45900
rect 11866 45844 11922 45900
rect 11990 45844 12046 45900
rect 12114 45844 12170 45900
rect 10254 45720 10310 45776
rect 10378 45720 10434 45776
rect 10502 45720 10558 45776
rect 10626 45720 10682 45776
rect 10750 45720 10806 45776
rect 10874 45720 10930 45776
rect 10998 45720 11054 45776
rect 11122 45720 11178 45776
rect 11246 45720 11302 45776
rect 11370 45720 11426 45776
rect 11494 45720 11550 45776
rect 11618 45720 11674 45776
rect 11742 45720 11798 45776
rect 11866 45720 11922 45776
rect 11990 45720 12046 45776
rect 12114 45720 12170 45776
rect 10254 45596 10310 45652
rect 10378 45596 10434 45652
rect 10502 45596 10558 45652
rect 10626 45596 10682 45652
rect 10750 45596 10806 45652
rect 10874 45596 10930 45652
rect 10998 45596 11054 45652
rect 11122 45596 11178 45652
rect 11246 45596 11302 45652
rect 11370 45596 11426 45652
rect 11494 45596 11550 45652
rect 11618 45596 11674 45652
rect 11742 45596 11798 45652
rect 11866 45596 11922 45652
rect 11990 45596 12046 45652
rect 12114 45596 12170 45652
rect 10254 45472 10310 45528
rect 10378 45472 10434 45528
rect 10502 45472 10558 45528
rect 10626 45472 10682 45528
rect 10750 45472 10806 45528
rect 10874 45472 10930 45528
rect 10998 45472 11054 45528
rect 11122 45472 11178 45528
rect 11246 45472 11302 45528
rect 11370 45472 11426 45528
rect 11494 45472 11550 45528
rect 11618 45472 11674 45528
rect 11742 45472 11798 45528
rect 11866 45472 11922 45528
rect 11990 45472 12046 45528
rect 12114 45472 12170 45528
rect 10254 45348 10310 45404
rect 10378 45348 10434 45404
rect 10502 45348 10558 45404
rect 10626 45348 10682 45404
rect 10750 45348 10806 45404
rect 10874 45348 10930 45404
rect 10998 45348 11054 45404
rect 11122 45348 11178 45404
rect 11246 45348 11302 45404
rect 11370 45348 11426 45404
rect 11494 45348 11550 45404
rect 11618 45348 11674 45404
rect 11742 45348 11798 45404
rect 11866 45348 11922 45404
rect 11990 45348 12046 45404
rect 12114 45348 12170 45404
rect 10254 45224 10310 45280
rect 10378 45224 10434 45280
rect 10502 45224 10558 45280
rect 10626 45224 10682 45280
rect 10750 45224 10806 45280
rect 10874 45224 10930 45280
rect 10998 45224 11054 45280
rect 11122 45224 11178 45280
rect 11246 45224 11302 45280
rect 11370 45224 11426 45280
rect 11494 45224 11550 45280
rect 11618 45224 11674 45280
rect 11742 45224 11798 45280
rect 11866 45224 11922 45280
rect 11990 45224 12046 45280
rect 12114 45224 12170 45280
rect 10254 45100 10310 45156
rect 10378 45100 10434 45156
rect 10502 45100 10558 45156
rect 10626 45100 10682 45156
rect 10750 45100 10806 45156
rect 10874 45100 10930 45156
rect 10998 45100 11054 45156
rect 11122 45100 11178 45156
rect 11246 45100 11302 45156
rect 11370 45100 11426 45156
rect 11494 45100 11550 45156
rect 11618 45100 11674 45156
rect 11742 45100 11798 45156
rect 11866 45100 11922 45156
rect 11990 45100 12046 45156
rect 12114 45100 12170 45156
rect 10254 44976 10310 45032
rect 10378 44976 10434 45032
rect 10502 44976 10558 45032
rect 10626 44976 10682 45032
rect 10750 44976 10806 45032
rect 10874 44976 10930 45032
rect 10998 44976 11054 45032
rect 11122 44976 11178 45032
rect 11246 44976 11302 45032
rect 11370 44976 11426 45032
rect 11494 44976 11550 45032
rect 11618 44976 11674 45032
rect 11742 44976 11798 45032
rect 11866 44976 11922 45032
rect 11990 44976 12046 45032
rect 12114 44976 12170 45032
rect 10254 44852 10310 44908
rect 10378 44852 10434 44908
rect 10502 44852 10558 44908
rect 10626 44852 10682 44908
rect 10750 44852 10806 44908
rect 10874 44852 10930 44908
rect 10998 44852 11054 44908
rect 11122 44852 11178 44908
rect 11246 44852 11302 44908
rect 11370 44852 11426 44908
rect 11494 44852 11550 44908
rect 11618 44852 11674 44908
rect 11742 44852 11798 44908
rect 11866 44852 11922 44908
rect 11990 44852 12046 44908
rect 12114 44852 12170 44908
rect 12871 46092 12927 46148
rect 12995 46092 13051 46148
rect 13119 46092 13175 46148
rect 13243 46092 13299 46148
rect 13367 46092 13423 46148
rect 13491 46092 13547 46148
rect 13615 46092 13671 46148
rect 13739 46092 13795 46148
rect 13863 46092 13919 46148
rect 13987 46092 14043 46148
rect 14111 46092 14167 46148
rect 14235 46092 14291 46148
rect 14359 46092 14415 46148
rect 14483 46092 14539 46148
rect 14607 46092 14663 46148
rect 12871 45968 12927 46024
rect 12995 45968 13051 46024
rect 13119 45968 13175 46024
rect 13243 45968 13299 46024
rect 13367 45968 13423 46024
rect 13491 45968 13547 46024
rect 13615 45968 13671 46024
rect 13739 45968 13795 46024
rect 13863 45968 13919 46024
rect 13987 45968 14043 46024
rect 14111 45968 14167 46024
rect 14235 45968 14291 46024
rect 14359 45968 14415 46024
rect 14483 45968 14539 46024
rect 14607 45968 14663 46024
rect 12871 45844 12927 45900
rect 12995 45844 13051 45900
rect 13119 45844 13175 45900
rect 13243 45844 13299 45900
rect 13367 45844 13423 45900
rect 13491 45844 13547 45900
rect 13615 45844 13671 45900
rect 13739 45844 13795 45900
rect 13863 45844 13919 45900
rect 13987 45844 14043 45900
rect 14111 45844 14167 45900
rect 14235 45844 14291 45900
rect 14359 45844 14415 45900
rect 14483 45844 14539 45900
rect 14607 45844 14663 45900
rect 12871 45720 12927 45776
rect 12995 45720 13051 45776
rect 13119 45720 13175 45776
rect 13243 45720 13299 45776
rect 13367 45720 13423 45776
rect 13491 45720 13547 45776
rect 13615 45720 13671 45776
rect 13739 45720 13795 45776
rect 13863 45720 13919 45776
rect 13987 45720 14043 45776
rect 14111 45720 14167 45776
rect 14235 45720 14291 45776
rect 14359 45720 14415 45776
rect 14483 45720 14539 45776
rect 14607 45720 14663 45776
rect 12871 45596 12927 45652
rect 12995 45596 13051 45652
rect 13119 45596 13175 45652
rect 13243 45596 13299 45652
rect 13367 45596 13423 45652
rect 13491 45596 13547 45652
rect 13615 45596 13671 45652
rect 13739 45596 13795 45652
rect 13863 45596 13919 45652
rect 13987 45596 14043 45652
rect 14111 45596 14167 45652
rect 14235 45596 14291 45652
rect 14359 45596 14415 45652
rect 14483 45596 14539 45652
rect 14607 45596 14663 45652
rect 12871 45472 12927 45528
rect 12995 45472 13051 45528
rect 13119 45472 13175 45528
rect 13243 45472 13299 45528
rect 13367 45472 13423 45528
rect 13491 45472 13547 45528
rect 13615 45472 13671 45528
rect 13739 45472 13795 45528
rect 13863 45472 13919 45528
rect 13987 45472 14043 45528
rect 14111 45472 14167 45528
rect 14235 45472 14291 45528
rect 14359 45472 14415 45528
rect 14483 45472 14539 45528
rect 14607 45472 14663 45528
rect 12871 45348 12927 45404
rect 12995 45348 13051 45404
rect 13119 45348 13175 45404
rect 13243 45348 13299 45404
rect 13367 45348 13423 45404
rect 13491 45348 13547 45404
rect 13615 45348 13671 45404
rect 13739 45348 13795 45404
rect 13863 45348 13919 45404
rect 13987 45348 14043 45404
rect 14111 45348 14167 45404
rect 14235 45348 14291 45404
rect 14359 45348 14415 45404
rect 14483 45348 14539 45404
rect 14607 45348 14663 45404
rect 12871 45224 12927 45280
rect 12995 45224 13051 45280
rect 13119 45224 13175 45280
rect 13243 45224 13299 45280
rect 13367 45224 13423 45280
rect 13491 45224 13547 45280
rect 13615 45224 13671 45280
rect 13739 45224 13795 45280
rect 13863 45224 13919 45280
rect 13987 45224 14043 45280
rect 14111 45224 14167 45280
rect 14235 45224 14291 45280
rect 14359 45224 14415 45280
rect 14483 45224 14539 45280
rect 14607 45224 14663 45280
rect 12871 45100 12927 45156
rect 12995 45100 13051 45156
rect 13119 45100 13175 45156
rect 13243 45100 13299 45156
rect 13367 45100 13423 45156
rect 13491 45100 13547 45156
rect 13615 45100 13671 45156
rect 13739 45100 13795 45156
rect 13863 45100 13919 45156
rect 13987 45100 14043 45156
rect 14111 45100 14167 45156
rect 14235 45100 14291 45156
rect 14359 45100 14415 45156
rect 14483 45100 14539 45156
rect 14607 45100 14663 45156
rect 12871 44976 12927 45032
rect 12995 44976 13051 45032
rect 13119 44976 13175 45032
rect 13243 44976 13299 45032
rect 13367 44976 13423 45032
rect 13491 44976 13547 45032
rect 13615 44976 13671 45032
rect 13739 44976 13795 45032
rect 13863 44976 13919 45032
rect 13987 44976 14043 45032
rect 14111 44976 14167 45032
rect 14235 44976 14291 45032
rect 14359 44976 14415 45032
rect 14483 44976 14539 45032
rect 14607 44976 14663 45032
rect 12871 44852 12927 44908
rect 12995 44852 13051 44908
rect 13119 44852 13175 44908
rect 13243 44852 13299 44908
rect 13367 44852 13423 44908
rect 13491 44852 13547 44908
rect 13615 44852 13671 44908
rect 13739 44852 13795 44908
rect 13863 44852 13919 44908
rect 13987 44852 14043 44908
rect 14111 44852 14167 44908
rect 14235 44852 14291 44908
rect 14359 44852 14415 44908
rect 14483 44852 14539 44908
rect 14607 44852 14663 44908
rect 14902 46174 14958 46176
rect 14902 46122 14904 46174
rect 14904 46122 14956 46174
rect 14956 46122 14958 46174
rect 14902 46066 14958 46122
rect 14902 46014 14904 46066
rect 14904 46014 14956 46066
rect 14956 46014 14958 46066
rect 14902 45958 14958 46014
rect 14902 45906 14904 45958
rect 14904 45906 14956 45958
rect 14956 45906 14958 45958
rect 14902 45850 14958 45906
rect 14902 45798 14904 45850
rect 14904 45798 14956 45850
rect 14956 45798 14958 45850
rect 14902 45742 14958 45798
rect 14902 45690 14904 45742
rect 14904 45690 14956 45742
rect 14956 45690 14958 45742
rect 14902 45634 14958 45690
rect 14902 45582 14904 45634
rect 14904 45582 14956 45634
rect 14956 45582 14958 45634
rect 14902 45526 14958 45582
rect 14902 45474 14904 45526
rect 14904 45474 14956 45526
rect 14956 45474 14958 45526
rect 14902 45418 14958 45474
rect 14902 45366 14904 45418
rect 14904 45366 14956 45418
rect 14956 45366 14958 45418
rect 14902 45310 14958 45366
rect 14902 45258 14904 45310
rect 14904 45258 14956 45310
rect 14956 45258 14958 45310
rect 14902 45202 14958 45258
rect 14902 45150 14904 45202
rect 14904 45150 14956 45202
rect 14956 45150 14958 45202
rect 14902 45094 14958 45150
rect 14902 45042 14904 45094
rect 14904 45042 14956 45094
rect 14956 45042 14958 45094
rect 14902 44986 14958 45042
rect 14902 44934 14904 44986
rect 14904 44934 14956 44986
rect 14956 44934 14958 44986
rect 14902 44878 14958 44934
rect 14902 44826 14904 44878
rect 14904 44826 14956 44878
rect 14956 44826 14958 44878
rect 14902 44824 14958 44826
rect 2491 44492 2547 44548
rect 2615 44492 2671 44548
rect 2491 44368 2547 44424
rect 2615 44368 2671 44424
rect 2491 44244 2547 44300
rect 2615 44244 2671 44300
rect 2491 44120 2547 44176
rect 2615 44120 2671 44176
rect 2491 43996 2547 44052
rect 2615 43996 2671 44052
rect 2491 43872 2547 43928
rect 2615 43872 2671 43928
rect 2491 43748 2547 43804
rect 2615 43748 2671 43804
rect 2491 43624 2547 43680
rect 2615 43624 2671 43680
rect 2491 43500 2547 43556
rect 2615 43500 2671 43556
rect 2491 43376 2547 43432
rect 2615 43376 2671 43432
rect 2491 43252 2547 43308
rect 2615 43252 2671 43308
rect 4861 44492 4917 44548
rect 4985 44492 5041 44548
rect 4861 44368 4917 44424
rect 4985 44368 5041 44424
rect 4861 44244 4917 44300
rect 4985 44244 5041 44300
rect 4861 44120 4917 44176
rect 4985 44120 5041 44176
rect 4861 43996 4917 44052
rect 4985 43996 5041 44052
rect 4861 43872 4917 43928
rect 4985 43872 5041 43928
rect 4861 43748 4917 43804
rect 4985 43748 5041 43804
rect 4861 43624 4917 43680
rect 4985 43624 5041 43680
rect 4861 43500 4917 43556
rect 4985 43500 5041 43556
rect 4861 43376 4917 43432
rect 4985 43376 5041 43432
rect 4861 43252 4917 43308
rect 4985 43252 5041 43308
rect 7275 44492 7331 44548
rect 7399 44492 7455 44548
rect 7523 44492 7579 44548
rect 7647 44492 7703 44548
rect 7275 44368 7331 44424
rect 7399 44368 7455 44424
rect 7523 44368 7579 44424
rect 7647 44368 7703 44424
rect 7275 44244 7331 44300
rect 7399 44244 7455 44300
rect 7523 44244 7579 44300
rect 7647 44244 7703 44300
rect 7275 44120 7331 44176
rect 7399 44120 7455 44176
rect 7523 44120 7579 44176
rect 7647 44120 7703 44176
rect 7275 43996 7331 44052
rect 7399 43996 7455 44052
rect 7523 43996 7579 44052
rect 7647 43996 7703 44052
rect 7275 43872 7331 43928
rect 7399 43872 7455 43928
rect 7523 43872 7579 43928
rect 7647 43872 7703 43928
rect 7275 43748 7331 43804
rect 7399 43748 7455 43804
rect 7523 43748 7579 43804
rect 7647 43748 7703 43804
rect 7275 43624 7331 43680
rect 7399 43624 7455 43680
rect 7523 43624 7579 43680
rect 7647 43624 7703 43680
rect 7275 43500 7331 43556
rect 7399 43500 7455 43556
rect 7523 43500 7579 43556
rect 7647 43500 7703 43556
rect 7275 43376 7331 43432
rect 7399 43376 7455 43432
rect 7523 43376 7579 43432
rect 7647 43376 7703 43432
rect 7275 43252 7331 43308
rect 7399 43252 7455 43308
rect 7523 43252 7579 43308
rect 7647 43252 7703 43308
rect 9937 44492 9993 44548
rect 10061 44492 10117 44548
rect 9937 44368 9993 44424
rect 10061 44368 10117 44424
rect 9937 44244 9993 44300
rect 10061 44244 10117 44300
rect 9937 44120 9993 44176
rect 10061 44120 10117 44176
rect 9937 43996 9993 44052
rect 10061 43996 10117 44052
rect 9937 43872 9993 43928
rect 10061 43872 10117 43928
rect 9937 43748 9993 43804
rect 10061 43748 10117 43804
rect 9937 43624 9993 43680
rect 10061 43624 10117 43680
rect 9937 43500 9993 43556
rect 10061 43500 10117 43556
rect 9937 43376 9993 43432
rect 10061 43376 10117 43432
rect 9937 43252 9993 43308
rect 10061 43252 10117 43308
rect 12307 44492 12363 44548
rect 12431 44492 12487 44548
rect 12307 44368 12363 44424
rect 12431 44368 12487 44424
rect 12307 44244 12363 44300
rect 12431 44244 12487 44300
rect 12307 44120 12363 44176
rect 12431 44120 12487 44176
rect 12307 43996 12363 44052
rect 12431 43996 12487 44052
rect 12307 43872 12363 43928
rect 12431 43872 12487 43928
rect 12307 43748 12363 43804
rect 12431 43748 12487 43804
rect 12307 43624 12363 43680
rect 12431 43624 12487 43680
rect 12307 43500 12363 43556
rect 12431 43500 12487 43556
rect 12307 43376 12363 43432
rect 12431 43376 12487 43432
rect 12307 43252 12363 43308
rect 12431 43252 12487 43308
rect 2491 42892 2547 42948
rect 2615 42892 2671 42948
rect 2491 42768 2547 42824
rect 2615 42768 2671 42824
rect 2491 42644 2547 42700
rect 2615 42644 2671 42700
rect 2491 42520 2547 42576
rect 2615 42520 2671 42576
rect 2491 42396 2547 42452
rect 2615 42396 2671 42452
rect 2491 42272 2547 42328
rect 2615 42272 2671 42328
rect 2491 42148 2547 42204
rect 2615 42148 2671 42204
rect 2491 42024 2547 42080
rect 2615 42024 2671 42080
rect 2491 41900 2547 41956
rect 2615 41900 2671 41956
rect 2491 41776 2547 41832
rect 2615 41776 2671 41832
rect 2491 41652 2547 41708
rect 2615 41652 2671 41708
rect 4861 42892 4917 42948
rect 4985 42892 5041 42948
rect 4861 42768 4917 42824
rect 4985 42768 5041 42824
rect 4861 42644 4917 42700
rect 4985 42644 5041 42700
rect 4861 42520 4917 42576
rect 4985 42520 5041 42576
rect 4861 42396 4917 42452
rect 4985 42396 5041 42452
rect 4861 42272 4917 42328
rect 4985 42272 5041 42328
rect 4861 42148 4917 42204
rect 4985 42148 5041 42204
rect 4861 42024 4917 42080
rect 4985 42024 5041 42080
rect 4861 41900 4917 41956
rect 4985 41900 5041 41956
rect 4861 41776 4917 41832
rect 4985 41776 5041 41832
rect 4861 41652 4917 41708
rect 4985 41652 5041 41708
rect 7275 42892 7331 42948
rect 7399 42892 7455 42948
rect 7523 42892 7579 42948
rect 7647 42892 7703 42948
rect 7275 42768 7331 42824
rect 7399 42768 7455 42824
rect 7523 42768 7579 42824
rect 7647 42768 7703 42824
rect 7275 42644 7331 42700
rect 7399 42644 7455 42700
rect 7523 42644 7579 42700
rect 7647 42644 7703 42700
rect 7275 42520 7331 42576
rect 7399 42520 7455 42576
rect 7523 42520 7579 42576
rect 7647 42520 7703 42576
rect 7275 42396 7331 42452
rect 7399 42396 7455 42452
rect 7523 42396 7579 42452
rect 7647 42396 7703 42452
rect 7275 42272 7331 42328
rect 7399 42272 7455 42328
rect 7523 42272 7579 42328
rect 7647 42272 7703 42328
rect 7275 42148 7331 42204
rect 7399 42148 7455 42204
rect 7523 42148 7579 42204
rect 7647 42148 7703 42204
rect 7275 42024 7331 42080
rect 7399 42024 7455 42080
rect 7523 42024 7579 42080
rect 7647 42024 7703 42080
rect 7275 41900 7331 41956
rect 7399 41900 7455 41956
rect 7523 41900 7579 41956
rect 7647 41900 7703 41956
rect 7275 41776 7331 41832
rect 7399 41776 7455 41832
rect 7523 41776 7579 41832
rect 7647 41776 7703 41832
rect 7275 41652 7331 41708
rect 7399 41652 7455 41708
rect 7523 41652 7579 41708
rect 7647 41652 7703 41708
rect 9937 42892 9993 42948
rect 10061 42892 10117 42948
rect 9937 42768 9993 42824
rect 10061 42768 10117 42824
rect 9937 42644 9993 42700
rect 10061 42644 10117 42700
rect 9937 42520 9993 42576
rect 10061 42520 10117 42576
rect 9937 42396 9993 42452
rect 10061 42396 10117 42452
rect 9937 42272 9993 42328
rect 10061 42272 10117 42328
rect 9937 42148 9993 42204
rect 10061 42148 10117 42204
rect 9937 42024 9993 42080
rect 10061 42024 10117 42080
rect 9937 41900 9993 41956
rect 10061 41900 10117 41956
rect 9937 41776 9993 41832
rect 10061 41776 10117 41832
rect 9937 41652 9993 41708
rect 10061 41652 10117 41708
rect 12307 42892 12363 42948
rect 12431 42892 12487 42948
rect 12307 42768 12363 42824
rect 12431 42768 12487 42824
rect 12307 42644 12363 42700
rect 12431 42644 12487 42700
rect 12307 42520 12363 42576
rect 12431 42520 12487 42576
rect 12307 42396 12363 42452
rect 12431 42396 12487 42452
rect 12307 42272 12363 42328
rect 12431 42272 12487 42328
rect 12307 42148 12363 42204
rect 12431 42148 12487 42204
rect 12307 42024 12363 42080
rect 12431 42024 12487 42080
rect 12307 41900 12363 41956
rect 12431 41900 12487 41956
rect 12307 41776 12363 41832
rect 12431 41776 12487 41832
rect 12307 41652 12363 41708
rect 12431 41652 12487 41708
rect 2491 41292 2547 41348
rect 2615 41292 2671 41348
rect 2491 41168 2547 41224
rect 2615 41168 2671 41224
rect 2491 41044 2547 41100
rect 2615 41044 2671 41100
rect 2491 40920 2547 40976
rect 2615 40920 2671 40976
rect 2491 40796 2547 40852
rect 2615 40796 2671 40852
rect 2491 40672 2547 40728
rect 2615 40672 2671 40728
rect 2491 40548 2547 40604
rect 2615 40548 2671 40604
rect 2491 40424 2547 40480
rect 2615 40424 2671 40480
rect 2491 40300 2547 40356
rect 2615 40300 2671 40356
rect 2491 40176 2547 40232
rect 2615 40176 2671 40232
rect 2491 40052 2547 40108
rect 2615 40052 2671 40108
rect 4861 41292 4917 41348
rect 4985 41292 5041 41348
rect 4861 41168 4917 41224
rect 4985 41168 5041 41224
rect 4861 41044 4917 41100
rect 4985 41044 5041 41100
rect 4861 40920 4917 40976
rect 4985 40920 5041 40976
rect 4861 40796 4917 40852
rect 4985 40796 5041 40852
rect 4861 40672 4917 40728
rect 4985 40672 5041 40728
rect 4861 40548 4917 40604
rect 4985 40548 5041 40604
rect 4861 40424 4917 40480
rect 4985 40424 5041 40480
rect 4861 40300 4917 40356
rect 4985 40300 5041 40356
rect 4861 40176 4917 40232
rect 4985 40176 5041 40232
rect 4861 40052 4917 40108
rect 4985 40052 5041 40108
rect 7275 41292 7331 41348
rect 7399 41292 7455 41348
rect 7523 41292 7579 41348
rect 7647 41292 7703 41348
rect 7275 41168 7331 41224
rect 7399 41168 7455 41224
rect 7523 41168 7579 41224
rect 7647 41168 7703 41224
rect 7275 41044 7331 41100
rect 7399 41044 7455 41100
rect 7523 41044 7579 41100
rect 7647 41044 7703 41100
rect 7275 40920 7331 40976
rect 7399 40920 7455 40976
rect 7523 40920 7579 40976
rect 7647 40920 7703 40976
rect 7275 40796 7331 40852
rect 7399 40796 7455 40852
rect 7523 40796 7579 40852
rect 7647 40796 7703 40852
rect 7275 40672 7331 40728
rect 7399 40672 7455 40728
rect 7523 40672 7579 40728
rect 7647 40672 7703 40728
rect 7275 40548 7331 40604
rect 7399 40548 7455 40604
rect 7523 40548 7579 40604
rect 7647 40548 7703 40604
rect 7275 40424 7331 40480
rect 7399 40424 7455 40480
rect 7523 40424 7579 40480
rect 7647 40424 7703 40480
rect 7275 40300 7331 40356
rect 7399 40300 7455 40356
rect 7523 40300 7579 40356
rect 7647 40300 7703 40356
rect 7275 40176 7331 40232
rect 7399 40176 7455 40232
rect 7523 40176 7579 40232
rect 7647 40176 7703 40232
rect 7275 40052 7331 40108
rect 7399 40052 7455 40108
rect 7523 40052 7579 40108
rect 7647 40052 7703 40108
rect 9937 41292 9993 41348
rect 10061 41292 10117 41348
rect 9937 41168 9993 41224
rect 10061 41168 10117 41224
rect 9937 41044 9993 41100
rect 10061 41044 10117 41100
rect 9937 40920 9993 40976
rect 10061 40920 10117 40976
rect 9937 40796 9993 40852
rect 10061 40796 10117 40852
rect 9937 40672 9993 40728
rect 10061 40672 10117 40728
rect 9937 40548 9993 40604
rect 10061 40548 10117 40604
rect 9937 40424 9993 40480
rect 10061 40424 10117 40480
rect 9937 40300 9993 40356
rect 10061 40300 10117 40356
rect 9937 40176 9993 40232
rect 10061 40176 10117 40232
rect 9937 40052 9993 40108
rect 10061 40052 10117 40108
rect 12307 41292 12363 41348
rect 12431 41292 12487 41348
rect 12307 41168 12363 41224
rect 12431 41168 12487 41224
rect 12307 41044 12363 41100
rect 12431 41044 12487 41100
rect 12307 40920 12363 40976
rect 12431 40920 12487 40976
rect 12307 40796 12363 40852
rect 12431 40796 12487 40852
rect 12307 40672 12363 40728
rect 12431 40672 12487 40728
rect 12307 40548 12363 40604
rect 12431 40548 12487 40604
rect 12307 40424 12363 40480
rect 12431 40424 12487 40480
rect 12307 40300 12363 40356
rect 12431 40300 12487 40356
rect 12307 40176 12363 40232
rect 12431 40176 12487 40232
rect 12307 40052 12363 40108
rect 12431 40052 12487 40108
rect 2302 39671 2358 39727
rect 2302 39539 2358 39595
rect 2302 39407 2358 39463
rect 2302 39275 2358 39331
rect 2302 39143 2358 39199
rect 2302 39011 2358 39067
rect 2302 38879 2358 38935
rect 2302 38747 2358 38803
rect 2302 38615 2358 38671
rect 2302 38483 2358 38539
rect 20 38174 76 38176
rect 20 38122 22 38174
rect 22 38122 74 38174
rect 74 38122 76 38174
rect 20 38066 76 38122
rect 20 38014 22 38066
rect 22 38014 74 38066
rect 74 38014 76 38066
rect 20 37958 76 38014
rect 20 37906 22 37958
rect 22 37906 74 37958
rect 74 37906 76 37958
rect 20 37850 76 37906
rect 20 37798 22 37850
rect 22 37798 74 37850
rect 74 37798 76 37850
rect 20 37742 76 37798
rect 20 37690 22 37742
rect 22 37690 74 37742
rect 74 37690 76 37742
rect 20 37634 76 37690
rect 20 37582 22 37634
rect 22 37582 74 37634
rect 74 37582 76 37634
rect 20 37526 76 37582
rect 20 37474 22 37526
rect 22 37474 74 37526
rect 74 37474 76 37526
rect 20 37418 76 37474
rect 20 37366 22 37418
rect 22 37366 74 37418
rect 74 37366 76 37418
rect 20 37310 76 37366
rect 20 37258 22 37310
rect 22 37258 74 37310
rect 74 37258 76 37310
rect 20 37202 76 37258
rect 20 37150 22 37202
rect 22 37150 74 37202
rect 74 37150 76 37202
rect 20 37094 76 37150
rect 20 37042 22 37094
rect 22 37042 74 37094
rect 74 37042 76 37094
rect 20 36986 76 37042
rect 20 36934 22 36986
rect 22 36934 74 36986
rect 74 36934 76 36986
rect 20 36878 76 36934
rect 20 36826 22 36878
rect 22 36826 74 36878
rect 74 36826 76 36878
rect 20 36824 76 36826
rect 315 38092 371 38148
rect 439 38092 495 38148
rect 563 38092 619 38148
rect 687 38092 743 38148
rect 811 38092 867 38148
rect 935 38092 991 38148
rect 1059 38092 1115 38148
rect 1183 38092 1239 38148
rect 1307 38092 1363 38148
rect 1431 38092 1487 38148
rect 1555 38092 1611 38148
rect 1679 38092 1735 38148
rect 1803 38092 1859 38148
rect 1927 38092 1983 38148
rect 2051 38092 2107 38148
rect 315 37968 371 38024
rect 439 37968 495 38024
rect 563 37968 619 38024
rect 687 37968 743 38024
rect 811 37968 867 38024
rect 935 37968 991 38024
rect 1059 37968 1115 38024
rect 1183 37968 1239 38024
rect 1307 37968 1363 38024
rect 1431 37968 1487 38024
rect 1555 37968 1611 38024
rect 1679 37968 1735 38024
rect 1803 37968 1859 38024
rect 1927 37968 1983 38024
rect 2051 37968 2107 38024
rect 315 37844 371 37900
rect 439 37844 495 37900
rect 563 37844 619 37900
rect 687 37844 743 37900
rect 811 37844 867 37900
rect 935 37844 991 37900
rect 1059 37844 1115 37900
rect 1183 37844 1239 37900
rect 1307 37844 1363 37900
rect 1431 37844 1487 37900
rect 1555 37844 1611 37900
rect 1679 37844 1735 37900
rect 1803 37844 1859 37900
rect 1927 37844 1983 37900
rect 2051 37844 2107 37900
rect 315 37720 371 37776
rect 439 37720 495 37776
rect 563 37720 619 37776
rect 687 37720 743 37776
rect 811 37720 867 37776
rect 935 37720 991 37776
rect 1059 37720 1115 37776
rect 1183 37720 1239 37776
rect 1307 37720 1363 37776
rect 1431 37720 1487 37776
rect 1555 37720 1611 37776
rect 1679 37720 1735 37776
rect 1803 37720 1859 37776
rect 1927 37720 1983 37776
rect 2051 37720 2107 37776
rect 315 37596 371 37652
rect 439 37596 495 37652
rect 563 37596 619 37652
rect 687 37596 743 37652
rect 811 37596 867 37652
rect 935 37596 991 37652
rect 1059 37596 1115 37652
rect 1183 37596 1239 37652
rect 1307 37596 1363 37652
rect 1431 37596 1487 37652
rect 1555 37596 1611 37652
rect 1679 37596 1735 37652
rect 1803 37596 1859 37652
rect 1927 37596 1983 37652
rect 2051 37596 2107 37652
rect 315 37472 371 37528
rect 439 37472 495 37528
rect 563 37472 619 37528
rect 687 37472 743 37528
rect 811 37472 867 37528
rect 935 37472 991 37528
rect 1059 37472 1115 37528
rect 1183 37472 1239 37528
rect 1307 37472 1363 37528
rect 1431 37472 1487 37528
rect 1555 37472 1611 37528
rect 1679 37472 1735 37528
rect 1803 37472 1859 37528
rect 1927 37472 1983 37528
rect 2051 37472 2107 37528
rect 315 37348 371 37404
rect 439 37348 495 37404
rect 563 37348 619 37404
rect 687 37348 743 37404
rect 811 37348 867 37404
rect 935 37348 991 37404
rect 1059 37348 1115 37404
rect 1183 37348 1239 37404
rect 1307 37348 1363 37404
rect 1431 37348 1487 37404
rect 1555 37348 1611 37404
rect 1679 37348 1735 37404
rect 1803 37348 1859 37404
rect 1927 37348 1983 37404
rect 2051 37348 2107 37404
rect 315 37224 371 37280
rect 439 37224 495 37280
rect 563 37224 619 37280
rect 687 37224 743 37280
rect 811 37224 867 37280
rect 935 37224 991 37280
rect 1059 37224 1115 37280
rect 1183 37224 1239 37280
rect 1307 37224 1363 37280
rect 1431 37224 1487 37280
rect 1555 37224 1611 37280
rect 1679 37224 1735 37280
rect 1803 37224 1859 37280
rect 1927 37224 1983 37280
rect 2051 37224 2107 37280
rect 315 37100 371 37156
rect 439 37100 495 37156
rect 563 37100 619 37156
rect 687 37100 743 37156
rect 811 37100 867 37156
rect 935 37100 991 37156
rect 1059 37100 1115 37156
rect 1183 37100 1239 37156
rect 1307 37100 1363 37156
rect 1431 37100 1487 37156
rect 1555 37100 1611 37156
rect 1679 37100 1735 37156
rect 1803 37100 1859 37156
rect 1927 37100 1983 37156
rect 2051 37100 2107 37156
rect 315 36976 371 37032
rect 439 36976 495 37032
rect 563 36976 619 37032
rect 687 36976 743 37032
rect 811 36976 867 37032
rect 935 36976 991 37032
rect 1059 36976 1115 37032
rect 1183 36976 1239 37032
rect 1307 36976 1363 37032
rect 1431 36976 1487 37032
rect 1555 36976 1611 37032
rect 1679 36976 1735 37032
rect 1803 36976 1859 37032
rect 1927 36976 1983 37032
rect 2051 36976 2107 37032
rect 315 36852 371 36908
rect 439 36852 495 36908
rect 563 36852 619 36908
rect 687 36852 743 36908
rect 811 36852 867 36908
rect 935 36852 991 36908
rect 1059 36852 1115 36908
rect 1183 36852 1239 36908
rect 1307 36852 1363 36908
rect 1431 36852 1487 36908
rect 1555 36852 1611 36908
rect 1679 36852 1735 36908
rect 1803 36852 1859 36908
rect 1927 36852 1983 36908
rect 2051 36852 2107 36908
rect 2808 38092 2864 38148
rect 2932 38092 2988 38148
rect 3056 38092 3112 38148
rect 3180 38092 3236 38148
rect 3304 38092 3360 38148
rect 3428 38092 3484 38148
rect 3552 38092 3608 38148
rect 3676 38092 3732 38148
rect 3800 38092 3856 38148
rect 3924 38092 3980 38148
rect 4048 38092 4104 38148
rect 4172 38092 4228 38148
rect 4296 38092 4352 38148
rect 4420 38092 4476 38148
rect 4544 38092 4600 38148
rect 4668 38092 4724 38148
rect 2808 37968 2864 38024
rect 2932 37968 2988 38024
rect 3056 37968 3112 38024
rect 3180 37968 3236 38024
rect 3304 37968 3360 38024
rect 3428 37968 3484 38024
rect 3552 37968 3608 38024
rect 3676 37968 3732 38024
rect 3800 37968 3856 38024
rect 3924 37968 3980 38024
rect 4048 37968 4104 38024
rect 4172 37968 4228 38024
rect 4296 37968 4352 38024
rect 4420 37968 4476 38024
rect 4544 37968 4600 38024
rect 4668 37968 4724 38024
rect 2808 37844 2864 37900
rect 2932 37844 2988 37900
rect 3056 37844 3112 37900
rect 3180 37844 3236 37900
rect 3304 37844 3360 37900
rect 3428 37844 3484 37900
rect 3552 37844 3608 37900
rect 3676 37844 3732 37900
rect 3800 37844 3856 37900
rect 3924 37844 3980 37900
rect 4048 37844 4104 37900
rect 4172 37844 4228 37900
rect 4296 37844 4352 37900
rect 4420 37844 4476 37900
rect 4544 37844 4600 37900
rect 4668 37844 4724 37900
rect 2808 37720 2864 37776
rect 2932 37720 2988 37776
rect 3056 37720 3112 37776
rect 3180 37720 3236 37776
rect 3304 37720 3360 37776
rect 3428 37720 3484 37776
rect 3552 37720 3608 37776
rect 3676 37720 3732 37776
rect 3800 37720 3856 37776
rect 3924 37720 3980 37776
rect 4048 37720 4104 37776
rect 4172 37720 4228 37776
rect 4296 37720 4352 37776
rect 4420 37720 4476 37776
rect 4544 37720 4600 37776
rect 4668 37720 4724 37776
rect 2808 37596 2864 37652
rect 2932 37596 2988 37652
rect 3056 37596 3112 37652
rect 3180 37596 3236 37652
rect 3304 37596 3360 37652
rect 3428 37596 3484 37652
rect 3552 37596 3608 37652
rect 3676 37596 3732 37652
rect 3800 37596 3856 37652
rect 3924 37596 3980 37652
rect 4048 37596 4104 37652
rect 4172 37596 4228 37652
rect 4296 37596 4352 37652
rect 4420 37596 4476 37652
rect 4544 37596 4600 37652
rect 4668 37596 4724 37652
rect 2808 37472 2864 37528
rect 2932 37472 2988 37528
rect 3056 37472 3112 37528
rect 3180 37472 3236 37528
rect 3304 37472 3360 37528
rect 3428 37472 3484 37528
rect 3552 37472 3608 37528
rect 3676 37472 3732 37528
rect 3800 37472 3856 37528
rect 3924 37472 3980 37528
rect 4048 37472 4104 37528
rect 4172 37472 4228 37528
rect 4296 37472 4352 37528
rect 4420 37472 4476 37528
rect 4544 37472 4600 37528
rect 4668 37472 4724 37528
rect 2808 37348 2864 37404
rect 2932 37348 2988 37404
rect 3056 37348 3112 37404
rect 3180 37348 3236 37404
rect 3304 37348 3360 37404
rect 3428 37348 3484 37404
rect 3552 37348 3608 37404
rect 3676 37348 3732 37404
rect 3800 37348 3856 37404
rect 3924 37348 3980 37404
rect 4048 37348 4104 37404
rect 4172 37348 4228 37404
rect 4296 37348 4352 37404
rect 4420 37348 4476 37404
rect 4544 37348 4600 37404
rect 4668 37348 4724 37404
rect 2808 37224 2864 37280
rect 2932 37224 2988 37280
rect 3056 37224 3112 37280
rect 3180 37224 3236 37280
rect 3304 37224 3360 37280
rect 3428 37224 3484 37280
rect 3552 37224 3608 37280
rect 3676 37224 3732 37280
rect 3800 37224 3856 37280
rect 3924 37224 3980 37280
rect 4048 37224 4104 37280
rect 4172 37224 4228 37280
rect 4296 37224 4352 37280
rect 4420 37224 4476 37280
rect 4544 37224 4600 37280
rect 4668 37224 4724 37280
rect 2808 37100 2864 37156
rect 2932 37100 2988 37156
rect 3056 37100 3112 37156
rect 3180 37100 3236 37156
rect 3304 37100 3360 37156
rect 3428 37100 3484 37156
rect 3552 37100 3608 37156
rect 3676 37100 3732 37156
rect 3800 37100 3856 37156
rect 3924 37100 3980 37156
rect 4048 37100 4104 37156
rect 4172 37100 4228 37156
rect 4296 37100 4352 37156
rect 4420 37100 4476 37156
rect 4544 37100 4600 37156
rect 4668 37100 4724 37156
rect 2808 36976 2864 37032
rect 2932 36976 2988 37032
rect 3056 36976 3112 37032
rect 3180 36976 3236 37032
rect 3304 36976 3360 37032
rect 3428 36976 3484 37032
rect 3552 36976 3608 37032
rect 3676 36976 3732 37032
rect 3800 36976 3856 37032
rect 3924 36976 3980 37032
rect 4048 36976 4104 37032
rect 4172 36976 4228 37032
rect 4296 36976 4352 37032
rect 4420 36976 4476 37032
rect 4544 36976 4600 37032
rect 4668 36976 4724 37032
rect 2808 36852 2864 36908
rect 2932 36852 2988 36908
rect 3056 36852 3112 36908
rect 3180 36852 3236 36908
rect 3304 36852 3360 36908
rect 3428 36852 3484 36908
rect 3552 36852 3608 36908
rect 3676 36852 3732 36908
rect 3800 36852 3856 36908
rect 3924 36852 3980 36908
rect 4048 36852 4104 36908
rect 4172 36852 4228 36908
rect 4296 36852 4352 36908
rect 4420 36852 4476 36908
rect 4544 36852 4600 36908
rect 4668 36852 4724 36908
rect 5178 38092 5234 38148
rect 5302 38092 5358 38148
rect 5426 38092 5482 38148
rect 5550 38092 5606 38148
rect 5674 38092 5730 38148
rect 5798 38092 5854 38148
rect 5922 38092 5978 38148
rect 6046 38092 6102 38148
rect 6170 38092 6226 38148
rect 6294 38092 6350 38148
rect 6418 38092 6474 38148
rect 6542 38092 6598 38148
rect 6666 38092 6722 38148
rect 6790 38092 6846 38148
rect 6914 38092 6970 38148
rect 7038 38092 7094 38148
rect 5178 37968 5234 38024
rect 5302 37968 5358 38024
rect 5426 37968 5482 38024
rect 5550 37968 5606 38024
rect 5674 37968 5730 38024
rect 5798 37968 5854 38024
rect 5922 37968 5978 38024
rect 6046 37968 6102 38024
rect 6170 37968 6226 38024
rect 6294 37968 6350 38024
rect 6418 37968 6474 38024
rect 6542 37968 6598 38024
rect 6666 37968 6722 38024
rect 6790 37968 6846 38024
rect 6914 37968 6970 38024
rect 7038 37968 7094 38024
rect 5178 37844 5234 37900
rect 5302 37844 5358 37900
rect 5426 37844 5482 37900
rect 5550 37844 5606 37900
rect 5674 37844 5730 37900
rect 5798 37844 5854 37900
rect 5922 37844 5978 37900
rect 6046 37844 6102 37900
rect 6170 37844 6226 37900
rect 6294 37844 6350 37900
rect 6418 37844 6474 37900
rect 6542 37844 6598 37900
rect 6666 37844 6722 37900
rect 6790 37844 6846 37900
rect 6914 37844 6970 37900
rect 7038 37844 7094 37900
rect 5178 37720 5234 37776
rect 5302 37720 5358 37776
rect 5426 37720 5482 37776
rect 5550 37720 5606 37776
rect 5674 37720 5730 37776
rect 5798 37720 5854 37776
rect 5922 37720 5978 37776
rect 6046 37720 6102 37776
rect 6170 37720 6226 37776
rect 6294 37720 6350 37776
rect 6418 37720 6474 37776
rect 6542 37720 6598 37776
rect 6666 37720 6722 37776
rect 6790 37720 6846 37776
rect 6914 37720 6970 37776
rect 7038 37720 7094 37776
rect 5178 37596 5234 37652
rect 5302 37596 5358 37652
rect 5426 37596 5482 37652
rect 5550 37596 5606 37652
rect 5674 37596 5730 37652
rect 5798 37596 5854 37652
rect 5922 37596 5978 37652
rect 6046 37596 6102 37652
rect 6170 37596 6226 37652
rect 6294 37596 6350 37652
rect 6418 37596 6474 37652
rect 6542 37596 6598 37652
rect 6666 37596 6722 37652
rect 6790 37596 6846 37652
rect 6914 37596 6970 37652
rect 7038 37596 7094 37652
rect 5178 37472 5234 37528
rect 5302 37472 5358 37528
rect 5426 37472 5482 37528
rect 5550 37472 5606 37528
rect 5674 37472 5730 37528
rect 5798 37472 5854 37528
rect 5922 37472 5978 37528
rect 6046 37472 6102 37528
rect 6170 37472 6226 37528
rect 6294 37472 6350 37528
rect 6418 37472 6474 37528
rect 6542 37472 6598 37528
rect 6666 37472 6722 37528
rect 6790 37472 6846 37528
rect 6914 37472 6970 37528
rect 7038 37472 7094 37528
rect 5178 37348 5234 37404
rect 5302 37348 5358 37404
rect 5426 37348 5482 37404
rect 5550 37348 5606 37404
rect 5674 37348 5730 37404
rect 5798 37348 5854 37404
rect 5922 37348 5978 37404
rect 6046 37348 6102 37404
rect 6170 37348 6226 37404
rect 6294 37348 6350 37404
rect 6418 37348 6474 37404
rect 6542 37348 6598 37404
rect 6666 37348 6722 37404
rect 6790 37348 6846 37404
rect 6914 37348 6970 37404
rect 7038 37348 7094 37404
rect 5178 37224 5234 37280
rect 5302 37224 5358 37280
rect 5426 37224 5482 37280
rect 5550 37224 5606 37280
rect 5674 37224 5730 37280
rect 5798 37224 5854 37280
rect 5922 37224 5978 37280
rect 6046 37224 6102 37280
rect 6170 37224 6226 37280
rect 6294 37224 6350 37280
rect 6418 37224 6474 37280
rect 6542 37224 6598 37280
rect 6666 37224 6722 37280
rect 6790 37224 6846 37280
rect 6914 37224 6970 37280
rect 7038 37224 7094 37280
rect 5178 37100 5234 37156
rect 5302 37100 5358 37156
rect 5426 37100 5482 37156
rect 5550 37100 5606 37156
rect 5674 37100 5730 37156
rect 5798 37100 5854 37156
rect 5922 37100 5978 37156
rect 6046 37100 6102 37156
rect 6170 37100 6226 37156
rect 6294 37100 6350 37156
rect 6418 37100 6474 37156
rect 6542 37100 6598 37156
rect 6666 37100 6722 37156
rect 6790 37100 6846 37156
rect 6914 37100 6970 37156
rect 7038 37100 7094 37156
rect 5178 36976 5234 37032
rect 5302 36976 5358 37032
rect 5426 36976 5482 37032
rect 5550 36976 5606 37032
rect 5674 36976 5730 37032
rect 5798 36976 5854 37032
rect 5922 36976 5978 37032
rect 6046 36976 6102 37032
rect 6170 36976 6226 37032
rect 6294 36976 6350 37032
rect 6418 36976 6474 37032
rect 6542 36976 6598 37032
rect 6666 36976 6722 37032
rect 6790 36976 6846 37032
rect 6914 36976 6970 37032
rect 7038 36976 7094 37032
rect 5178 36852 5234 36908
rect 5302 36852 5358 36908
rect 5426 36852 5482 36908
rect 5550 36852 5606 36908
rect 5674 36852 5730 36908
rect 5798 36852 5854 36908
rect 5922 36852 5978 36908
rect 6046 36852 6102 36908
rect 6170 36852 6226 36908
rect 6294 36852 6350 36908
rect 6418 36852 6474 36908
rect 6542 36852 6598 36908
rect 6666 36852 6722 36908
rect 6790 36852 6846 36908
rect 6914 36852 6970 36908
rect 7038 36852 7094 36908
rect 7884 38092 7940 38148
rect 8008 38092 8064 38148
rect 8132 38092 8188 38148
rect 8256 38092 8312 38148
rect 8380 38092 8436 38148
rect 8504 38092 8560 38148
rect 8628 38092 8684 38148
rect 8752 38092 8808 38148
rect 8876 38092 8932 38148
rect 9000 38092 9056 38148
rect 9124 38092 9180 38148
rect 9248 38092 9304 38148
rect 9372 38092 9428 38148
rect 9496 38092 9552 38148
rect 9620 38092 9676 38148
rect 9744 38092 9800 38148
rect 7884 37968 7940 38024
rect 8008 37968 8064 38024
rect 8132 37968 8188 38024
rect 8256 37968 8312 38024
rect 8380 37968 8436 38024
rect 8504 37968 8560 38024
rect 8628 37968 8684 38024
rect 8752 37968 8808 38024
rect 8876 37968 8932 38024
rect 9000 37968 9056 38024
rect 9124 37968 9180 38024
rect 9248 37968 9304 38024
rect 9372 37968 9428 38024
rect 9496 37968 9552 38024
rect 9620 37968 9676 38024
rect 9744 37968 9800 38024
rect 7884 37844 7940 37900
rect 8008 37844 8064 37900
rect 8132 37844 8188 37900
rect 8256 37844 8312 37900
rect 8380 37844 8436 37900
rect 8504 37844 8560 37900
rect 8628 37844 8684 37900
rect 8752 37844 8808 37900
rect 8876 37844 8932 37900
rect 9000 37844 9056 37900
rect 9124 37844 9180 37900
rect 9248 37844 9304 37900
rect 9372 37844 9428 37900
rect 9496 37844 9552 37900
rect 9620 37844 9676 37900
rect 9744 37844 9800 37900
rect 7884 37720 7940 37776
rect 8008 37720 8064 37776
rect 8132 37720 8188 37776
rect 8256 37720 8312 37776
rect 8380 37720 8436 37776
rect 8504 37720 8560 37776
rect 8628 37720 8684 37776
rect 8752 37720 8808 37776
rect 8876 37720 8932 37776
rect 9000 37720 9056 37776
rect 9124 37720 9180 37776
rect 9248 37720 9304 37776
rect 9372 37720 9428 37776
rect 9496 37720 9552 37776
rect 9620 37720 9676 37776
rect 9744 37720 9800 37776
rect 7884 37596 7940 37652
rect 8008 37596 8064 37652
rect 8132 37596 8188 37652
rect 8256 37596 8312 37652
rect 8380 37596 8436 37652
rect 8504 37596 8560 37652
rect 8628 37596 8684 37652
rect 8752 37596 8808 37652
rect 8876 37596 8932 37652
rect 9000 37596 9056 37652
rect 9124 37596 9180 37652
rect 9248 37596 9304 37652
rect 9372 37596 9428 37652
rect 9496 37596 9552 37652
rect 9620 37596 9676 37652
rect 9744 37596 9800 37652
rect 7884 37472 7940 37528
rect 8008 37472 8064 37528
rect 8132 37472 8188 37528
rect 8256 37472 8312 37528
rect 8380 37472 8436 37528
rect 8504 37472 8560 37528
rect 8628 37472 8684 37528
rect 8752 37472 8808 37528
rect 8876 37472 8932 37528
rect 9000 37472 9056 37528
rect 9124 37472 9180 37528
rect 9248 37472 9304 37528
rect 9372 37472 9428 37528
rect 9496 37472 9552 37528
rect 9620 37472 9676 37528
rect 9744 37472 9800 37528
rect 7884 37348 7940 37404
rect 8008 37348 8064 37404
rect 8132 37348 8188 37404
rect 8256 37348 8312 37404
rect 8380 37348 8436 37404
rect 8504 37348 8560 37404
rect 8628 37348 8684 37404
rect 8752 37348 8808 37404
rect 8876 37348 8932 37404
rect 9000 37348 9056 37404
rect 9124 37348 9180 37404
rect 9248 37348 9304 37404
rect 9372 37348 9428 37404
rect 9496 37348 9552 37404
rect 9620 37348 9676 37404
rect 9744 37348 9800 37404
rect 7884 37224 7940 37280
rect 8008 37224 8064 37280
rect 8132 37224 8188 37280
rect 8256 37224 8312 37280
rect 8380 37224 8436 37280
rect 8504 37224 8560 37280
rect 8628 37224 8684 37280
rect 8752 37224 8808 37280
rect 8876 37224 8932 37280
rect 9000 37224 9056 37280
rect 9124 37224 9180 37280
rect 9248 37224 9304 37280
rect 9372 37224 9428 37280
rect 9496 37224 9552 37280
rect 9620 37224 9676 37280
rect 9744 37224 9800 37280
rect 7884 37100 7940 37156
rect 8008 37100 8064 37156
rect 8132 37100 8188 37156
rect 8256 37100 8312 37156
rect 8380 37100 8436 37156
rect 8504 37100 8560 37156
rect 8628 37100 8684 37156
rect 8752 37100 8808 37156
rect 8876 37100 8932 37156
rect 9000 37100 9056 37156
rect 9124 37100 9180 37156
rect 9248 37100 9304 37156
rect 9372 37100 9428 37156
rect 9496 37100 9552 37156
rect 9620 37100 9676 37156
rect 9744 37100 9800 37156
rect 7884 36976 7940 37032
rect 8008 36976 8064 37032
rect 8132 36976 8188 37032
rect 8256 36976 8312 37032
rect 8380 36976 8436 37032
rect 8504 36976 8560 37032
rect 8628 36976 8684 37032
rect 8752 36976 8808 37032
rect 8876 36976 8932 37032
rect 9000 36976 9056 37032
rect 9124 36976 9180 37032
rect 9248 36976 9304 37032
rect 9372 36976 9428 37032
rect 9496 36976 9552 37032
rect 9620 36976 9676 37032
rect 9744 36976 9800 37032
rect 7884 36852 7940 36908
rect 8008 36852 8064 36908
rect 8132 36852 8188 36908
rect 8256 36852 8312 36908
rect 8380 36852 8436 36908
rect 8504 36852 8560 36908
rect 8628 36852 8684 36908
rect 8752 36852 8808 36908
rect 8876 36852 8932 36908
rect 9000 36852 9056 36908
rect 9124 36852 9180 36908
rect 9248 36852 9304 36908
rect 9372 36852 9428 36908
rect 9496 36852 9552 36908
rect 9620 36852 9676 36908
rect 9744 36852 9800 36908
rect 10254 38092 10310 38148
rect 10378 38092 10434 38148
rect 10502 38092 10558 38148
rect 10626 38092 10682 38148
rect 10750 38092 10806 38148
rect 10874 38092 10930 38148
rect 10998 38092 11054 38148
rect 11122 38092 11178 38148
rect 11246 38092 11302 38148
rect 11370 38092 11426 38148
rect 11494 38092 11550 38148
rect 11618 38092 11674 38148
rect 11742 38092 11798 38148
rect 11866 38092 11922 38148
rect 11990 38092 12046 38148
rect 12114 38092 12170 38148
rect 10254 37968 10310 38024
rect 10378 37968 10434 38024
rect 10502 37968 10558 38024
rect 10626 37968 10682 38024
rect 10750 37968 10806 38024
rect 10874 37968 10930 38024
rect 10998 37968 11054 38024
rect 11122 37968 11178 38024
rect 11246 37968 11302 38024
rect 11370 37968 11426 38024
rect 11494 37968 11550 38024
rect 11618 37968 11674 38024
rect 11742 37968 11798 38024
rect 11866 37968 11922 38024
rect 11990 37968 12046 38024
rect 12114 37968 12170 38024
rect 10254 37844 10310 37900
rect 10378 37844 10434 37900
rect 10502 37844 10558 37900
rect 10626 37844 10682 37900
rect 10750 37844 10806 37900
rect 10874 37844 10930 37900
rect 10998 37844 11054 37900
rect 11122 37844 11178 37900
rect 11246 37844 11302 37900
rect 11370 37844 11426 37900
rect 11494 37844 11550 37900
rect 11618 37844 11674 37900
rect 11742 37844 11798 37900
rect 11866 37844 11922 37900
rect 11990 37844 12046 37900
rect 12114 37844 12170 37900
rect 10254 37720 10310 37776
rect 10378 37720 10434 37776
rect 10502 37720 10558 37776
rect 10626 37720 10682 37776
rect 10750 37720 10806 37776
rect 10874 37720 10930 37776
rect 10998 37720 11054 37776
rect 11122 37720 11178 37776
rect 11246 37720 11302 37776
rect 11370 37720 11426 37776
rect 11494 37720 11550 37776
rect 11618 37720 11674 37776
rect 11742 37720 11798 37776
rect 11866 37720 11922 37776
rect 11990 37720 12046 37776
rect 12114 37720 12170 37776
rect 10254 37596 10310 37652
rect 10378 37596 10434 37652
rect 10502 37596 10558 37652
rect 10626 37596 10682 37652
rect 10750 37596 10806 37652
rect 10874 37596 10930 37652
rect 10998 37596 11054 37652
rect 11122 37596 11178 37652
rect 11246 37596 11302 37652
rect 11370 37596 11426 37652
rect 11494 37596 11550 37652
rect 11618 37596 11674 37652
rect 11742 37596 11798 37652
rect 11866 37596 11922 37652
rect 11990 37596 12046 37652
rect 12114 37596 12170 37652
rect 10254 37472 10310 37528
rect 10378 37472 10434 37528
rect 10502 37472 10558 37528
rect 10626 37472 10682 37528
rect 10750 37472 10806 37528
rect 10874 37472 10930 37528
rect 10998 37472 11054 37528
rect 11122 37472 11178 37528
rect 11246 37472 11302 37528
rect 11370 37472 11426 37528
rect 11494 37472 11550 37528
rect 11618 37472 11674 37528
rect 11742 37472 11798 37528
rect 11866 37472 11922 37528
rect 11990 37472 12046 37528
rect 12114 37472 12170 37528
rect 10254 37348 10310 37404
rect 10378 37348 10434 37404
rect 10502 37348 10558 37404
rect 10626 37348 10682 37404
rect 10750 37348 10806 37404
rect 10874 37348 10930 37404
rect 10998 37348 11054 37404
rect 11122 37348 11178 37404
rect 11246 37348 11302 37404
rect 11370 37348 11426 37404
rect 11494 37348 11550 37404
rect 11618 37348 11674 37404
rect 11742 37348 11798 37404
rect 11866 37348 11922 37404
rect 11990 37348 12046 37404
rect 12114 37348 12170 37404
rect 10254 37224 10310 37280
rect 10378 37224 10434 37280
rect 10502 37224 10558 37280
rect 10626 37224 10682 37280
rect 10750 37224 10806 37280
rect 10874 37224 10930 37280
rect 10998 37224 11054 37280
rect 11122 37224 11178 37280
rect 11246 37224 11302 37280
rect 11370 37224 11426 37280
rect 11494 37224 11550 37280
rect 11618 37224 11674 37280
rect 11742 37224 11798 37280
rect 11866 37224 11922 37280
rect 11990 37224 12046 37280
rect 12114 37224 12170 37280
rect 10254 37100 10310 37156
rect 10378 37100 10434 37156
rect 10502 37100 10558 37156
rect 10626 37100 10682 37156
rect 10750 37100 10806 37156
rect 10874 37100 10930 37156
rect 10998 37100 11054 37156
rect 11122 37100 11178 37156
rect 11246 37100 11302 37156
rect 11370 37100 11426 37156
rect 11494 37100 11550 37156
rect 11618 37100 11674 37156
rect 11742 37100 11798 37156
rect 11866 37100 11922 37156
rect 11990 37100 12046 37156
rect 12114 37100 12170 37156
rect 10254 36976 10310 37032
rect 10378 36976 10434 37032
rect 10502 36976 10558 37032
rect 10626 36976 10682 37032
rect 10750 36976 10806 37032
rect 10874 36976 10930 37032
rect 10998 36976 11054 37032
rect 11122 36976 11178 37032
rect 11246 36976 11302 37032
rect 11370 36976 11426 37032
rect 11494 36976 11550 37032
rect 11618 36976 11674 37032
rect 11742 36976 11798 37032
rect 11866 36976 11922 37032
rect 11990 36976 12046 37032
rect 12114 36976 12170 37032
rect 10254 36852 10310 36908
rect 10378 36852 10434 36908
rect 10502 36852 10558 36908
rect 10626 36852 10682 36908
rect 10750 36852 10806 36908
rect 10874 36852 10930 36908
rect 10998 36852 11054 36908
rect 11122 36852 11178 36908
rect 11246 36852 11302 36908
rect 11370 36852 11426 36908
rect 11494 36852 11550 36908
rect 11618 36852 11674 36908
rect 11742 36852 11798 36908
rect 11866 36852 11922 36908
rect 11990 36852 12046 36908
rect 12114 36852 12170 36908
rect 12871 38092 12927 38148
rect 12995 38092 13051 38148
rect 13119 38092 13175 38148
rect 13243 38092 13299 38148
rect 13367 38092 13423 38148
rect 13491 38092 13547 38148
rect 13615 38092 13671 38148
rect 13739 38092 13795 38148
rect 13863 38092 13919 38148
rect 13987 38092 14043 38148
rect 14111 38092 14167 38148
rect 14235 38092 14291 38148
rect 14359 38092 14415 38148
rect 14483 38092 14539 38148
rect 14607 38092 14663 38148
rect 12871 37968 12927 38024
rect 12995 37968 13051 38024
rect 13119 37968 13175 38024
rect 13243 37968 13299 38024
rect 13367 37968 13423 38024
rect 13491 37968 13547 38024
rect 13615 37968 13671 38024
rect 13739 37968 13795 38024
rect 13863 37968 13919 38024
rect 13987 37968 14043 38024
rect 14111 37968 14167 38024
rect 14235 37968 14291 38024
rect 14359 37968 14415 38024
rect 14483 37968 14539 38024
rect 14607 37968 14663 38024
rect 12871 37844 12927 37900
rect 12995 37844 13051 37900
rect 13119 37844 13175 37900
rect 13243 37844 13299 37900
rect 13367 37844 13423 37900
rect 13491 37844 13547 37900
rect 13615 37844 13671 37900
rect 13739 37844 13795 37900
rect 13863 37844 13919 37900
rect 13987 37844 14043 37900
rect 14111 37844 14167 37900
rect 14235 37844 14291 37900
rect 14359 37844 14415 37900
rect 14483 37844 14539 37900
rect 14607 37844 14663 37900
rect 12871 37720 12927 37776
rect 12995 37720 13051 37776
rect 13119 37720 13175 37776
rect 13243 37720 13299 37776
rect 13367 37720 13423 37776
rect 13491 37720 13547 37776
rect 13615 37720 13671 37776
rect 13739 37720 13795 37776
rect 13863 37720 13919 37776
rect 13987 37720 14043 37776
rect 14111 37720 14167 37776
rect 14235 37720 14291 37776
rect 14359 37720 14415 37776
rect 14483 37720 14539 37776
rect 14607 37720 14663 37776
rect 12871 37596 12927 37652
rect 12995 37596 13051 37652
rect 13119 37596 13175 37652
rect 13243 37596 13299 37652
rect 13367 37596 13423 37652
rect 13491 37596 13547 37652
rect 13615 37596 13671 37652
rect 13739 37596 13795 37652
rect 13863 37596 13919 37652
rect 13987 37596 14043 37652
rect 14111 37596 14167 37652
rect 14235 37596 14291 37652
rect 14359 37596 14415 37652
rect 14483 37596 14539 37652
rect 14607 37596 14663 37652
rect 12871 37472 12927 37528
rect 12995 37472 13051 37528
rect 13119 37472 13175 37528
rect 13243 37472 13299 37528
rect 13367 37472 13423 37528
rect 13491 37472 13547 37528
rect 13615 37472 13671 37528
rect 13739 37472 13795 37528
rect 13863 37472 13919 37528
rect 13987 37472 14043 37528
rect 14111 37472 14167 37528
rect 14235 37472 14291 37528
rect 14359 37472 14415 37528
rect 14483 37472 14539 37528
rect 14607 37472 14663 37528
rect 12871 37348 12927 37404
rect 12995 37348 13051 37404
rect 13119 37348 13175 37404
rect 13243 37348 13299 37404
rect 13367 37348 13423 37404
rect 13491 37348 13547 37404
rect 13615 37348 13671 37404
rect 13739 37348 13795 37404
rect 13863 37348 13919 37404
rect 13987 37348 14043 37404
rect 14111 37348 14167 37404
rect 14235 37348 14291 37404
rect 14359 37348 14415 37404
rect 14483 37348 14539 37404
rect 14607 37348 14663 37404
rect 12871 37224 12927 37280
rect 12995 37224 13051 37280
rect 13119 37224 13175 37280
rect 13243 37224 13299 37280
rect 13367 37224 13423 37280
rect 13491 37224 13547 37280
rect 13615 37224 13671 37280
rect 13739 37224 13795 37280
rect 13863 37224 13919 37280
rect 13987 37224 14043 37280
rect 14111 37224 14167 37280
rect 14235 37224 14291 37280
rect 14359 37224 14415 37280
rect 14483 37224 14539 37280
rect 14607 37224 14663 37280
rect 12871 37100 12927 37156
rect 12995 37100 13051 37156
rect 13119 37100 13175 37156
rect 13243 37100 13299 37156
rect 13367 37100 13423 37156
rect 13491 37100 13547 37156
rect 13615 37100 13671 37156
rect 13739 37100 13795 37156
rect 13863 37100 13919 37156
rect 13987 37100 14043 37156
rect 14111 37100 14167 37156
rect 14235 37100 14291 37156
rect 14359 37100 14415 37156
rect 14483 37100 14539 37156
rect 14607 37100 14663 37156
rect 12871 36976 12927 37032
rect 12995 36976 13051 37032
rect 13119 36976 13175 37032
rect 13243 36976 13299 37032
rect 13367 36976 13423 37032
rect 13491 36976 13547 37032
rect 13615 36976 13671 37032
rect 13739 36976 13795 37032
rect 13863 36976 13919 37032
rect 13987 36976 14043 37032
rect 14111 36976 14167 37032
rect 14235 36976 14291 37032
rect 14359 36976 14415 37032
rect 14483 36976 14539 37032
rect 14607 36976 14663 37032
rect 12871 36852 12927 36908
rect 12995 36852 13051 36908
rect 13119 36852 13175 36908
rect 13243 36852 13299 36908
rect 13367 36852 13423 36908
rect 13491 36852 13547 36908
rect 13615 36852 13671 36908
rect 13739 36852 13795 36908
rect 13863 36852 13919 36908
rect 13987 36852 14043 36908
rect 14111 36852 14167 36908
rect 14235 36852 14291 36908
rect 14359 36852 14415 36908
rect 14483 36852 14539 36908
rect 14607 36852 14663 36908
rect 14902 38174 14958 38176
rect 14902 38122 14904 38174
rect 14904 38122 14956 38174
rect 14956 38122 14958 38174
rect 14902 38066 14958 38122
rect 14902 38014 14904 38066
rect 14904 38014 14956 38066
rect 14956 38014 14958 38066
rect 14902 37958 14958 38014
rect 14902 37906 14904 37958
rect 14904 37906 14956 37958
rect 14956 37906 14958 37958
rect 14902 37850 14958 37906
rect 14902 37798 14904 37850
rect 14904 37798 14956 37850
rect 14956 37798 14958 37850
rect 14902 37742 14958 37798
rect 14902 37690 14904 37742
rect 14904 37690 14956 37742
rect 14956 37690 14958 37742
rect 14902 37634 14958 37690
rect 14902 37582 14904 37634
rect 14904 37582 14956 37634
rect 14956 37582 14958 37634
rect 14902 37526 14958 37582
rect 14902 37474 14904 37526
rect 14904 37474 14956 37526
rect 14956 37474 14958 37526
rect 14902 37418 14958 37474
rect 14902 37366 14904 37418
rect 14904 37366 14956 37418
rect 14956 37366 14958 37418
rect 14902 37310 14958 37366
rect 14902 37258 14904 37310
rect 14904 37258 14956 37310
rect 14956 37258 14958 37310
rect 14902 37202 14958 37258
rect 14902 37150 14904 37202
rect 14904 37150 14956 37202
rect 14956 37150 14958 37202
rect 14902 37094 14958 37150
rect 14902 37042 14904 37094
rect 14904 37042 14956 37094
rect 14956 37042 14958 37094
rect 14902 36986 14958 37042
rect 14902 36934 14904 36986
rect 14904 36934 14956 36986
rect 14956 36934 14958 36986
rect 14902 36878 14958 36934
rect 14902 36826 14904 36878
rect 14904 36826 14956 36878
rect 14956 36826 14958 36878
rect 14902 36824 14958 36826
rect 20 36584 76 36586
rect 20 36532 22 36584
rect 22 36532 74 36584
rect 74 36532 76 36584
rect 20 36476 76 36532
rect 20 36424 22 36476
rect 22 36424 74 36476
rect 74 36424 76 36476
rect 20 36368 76 36424
rect 20 36316 22 36368
rect 22 36316 74 36368
rect 74 36316 76 36368
rect 20 36260 76 36316
rect 20 36208 22 36260
rect 22 36208 74 36260
rect 74 36208 76 36260
rect 20 36152 76 36208
rect 20 36100 22 36152
rect 22 36100 74 36152
rect 74 36100 76 36152
rect 20 36044 76 36100
rect 20 35992 22 36044
rect 22 35992 74 36044
rect 74 35992 76 36044
rect 20 35936 76 35992
rect 20 35884 22 35936
rect 22 35884 74 35936
rect 74 35884 76 35936
rect 20 35828 76 35884
rect 20 35776 22 35828
rect 22 35776 74 35828
rect 74 35776 76 35828
rect 20 35720 76 35776
rect 20 35668 22 35720
rect 22 35668 74 35720
rect 74 35668 76 35720
rect 20 35612 76 35668
rect 20 35560 22 35612
rect 22 35560 74 35612
rect 74 35560 76 35612
rect 20 35504 76 35560
rect 20 35452 22 35504
rect 22 35452 74 35504
rect 74 35452 76 35504
rect 20 35396 76 35452
rect 20 35344 22 35396
rect 22 35344 74 35396
rect 74 35344 76 35396
rect 20 35288 76 35344
rect 20 35236 22 35288
rect 22 35236 74 35288
rect 74 35236 76 35288
rect 20 35180 76 35236
rect 20 35128 22 35180
rect 22 35128 74 35180
rect 74 35128 76 35180
rect 20 35072 76 35128
rect 20 35020 22 35072
rect 22 35020 74 35072
rect 74 35020 76 35072
rect 20 34964 76 35020
rect 20 34912 22 34964
rect 22 34912 74 34964
rect 74 34912 76 34964
rect 20 34856 76 34912
rect 20 34804 22 34856
rect 22 34804 74 34856
rect 74 34804 76 34856
rect 20 34748 76 34804
rect 20 34696 22 34748
rect 22 34696 74 34748
rect 74 34696 76 34748
rect 20 34640 76 34696
rect 20 34588 22 34640
rect 22 34588 74 34640
rect 74 34588 76 34640
rect 20 34532 76 34588
rect 20 34480 22 34532
rect 22 34480 74 34532
rect 74 34480 76 34532
rect 20 34424 76 34480
rect 20 34372 22 34424
rect 22 34372 74 34424
rect 74 34372 76 34424
rect 20 34316 76 34372
rect 20 34264 22 34316
rect 22 34264 74 34316
rect 74 34264 76 34316
rect 20 34208 76 34264
rect 20 34156 22 34208
rect 22 34156 74 34208
rect 74 34156 76 34208
rect 20 34100 76 34156
rect 20 34048 22 34100
rect 22 34048 74 34100
rect 74 34048 76 34100
rect 20 33992 76 34048
rect 20 33940 22 33992
rect 22 33940 74 33992
rect 74 33940 76 33992
rect 20 33884 76 33940
rect 20 33832 22 33884
rect 22 33832 74 33884
rect 74 33832 76 33884
rect 20 33776 76 33832
rect 20 33724 22 33776
rect 22 33724 74 33776
rect 74 33724 76 33776
rect 20 33668 76 33724
rect 20 33616 22 33668
rect 22 33616 74 33668
rect 74 33616 76 33668
rect 20 33614 76 33616
rect 315 36498 371 36554
rect 439 36498 495 36554
rect 563 36498 619 36554
rect 687 36498 743 36554
rect 811 36498 867 36554
rect 935 36498 991 36554
rect 1059 36498 1115 36554
rect 1183 36498 1239 36554
rect 1307 36498 1363 36554
rect 1431 36498 1487 36554
rect 1555 36498 1611 36554
rect 1679 36498 1735 36554
rect 1803 36498 1859 36554
rect 1927 36498 1983 36554
rect 2051 36498 2107 36554
rect 315 36374 371 36430
rect 439 36374 495 36430
rect 563 36374 619 36430
rect 687 36374 743 36430
rect 811 36374 867 36430
rect 935 36374 991 36430
rect 1059 36374 1115 36430
rect 1183 36374 1239 36430
rect 1307 36374 1363 36430
rect 1431 36374 1487 36430
rect 1555 36374 1611 36430
rect 1679 36374 1735 36430
rect 1803 36374 1859 36430
rect 1927 36374 1983 36430
rect 2051 36374 2107 36430
rect 315 36250 371 36306
rect 439 36250 495 36306
rect 563 36250 619 36306
rect 687 36250 743 36306
rect 811 36250 867 36306
rect 935 36250 991 36306
rect 1059 36250 1115 36306
rect 1183 36250 1239 36306
rect 1307 36250 1363 36306
rect 1431 36250 1487 36306
rect 1555 36250 1611 36306
rect 1679 36250 1735 36306
rect 1803 36250 1859 36306
rect 1927 36250 1983 36306
rect 2051 36250 2107 36306
rect 315 36126 371 36182
rect 439 36126 495 36182
rect 563 36126 619 36182
rect 687 36126 743 36182
rect 811 36126 867 36182
rect 935 36126 991 36182
rect 1059 36126 1115 36182
rect 1183 36126 1239 36182
rect 1307 36126 1363 36182
rect 1431 36126 1487 36182
rect 1555 36126 1611 36182
rect 1679 36126 1735 36182
rect 1803 36126 1859 36182
rect 1927 36126 1983 36182
rect 2051 36126 2107 36182
rect 315 36002 371 36058
rect 439 36002 495 36058
rect 563 36002 619 36058
rect 687 36002 743 36058
rect 811 36002 867 36058
rect 935 36002 991 36058
rect 1059 36002 1115 36058
rect 1183 36002 1239 36058
rect 1307 36002 1363 36058
rect 1431 36002 1487 36058
rect 1555 36002 1611 36058
rect 1679 36002 1735 36058
rect 1803 36002 1859 36058
rect 1927 36002 1983 36058
rect 2051 36002 2107 36058
rect 315 35878 371 35934
rect 439 35878 495 35934
rect 563 35878 619 35934
rect 687 35878 743 35934
rect 811 35878 867 35934
rect 935 35878 991 35934
rect 1059 35878 1115 35934
rect 1183 35878 1239 35934
rect 1307 35878 1363 35934
rect 1431 35878 1487 35934
rect 1555 35878 1611 35934
rect 1679 35878 1735 35934
rect 1803 35878 1859 35934
rect 1927 35878 1983 35934
rect 2051 35878 2107 35934
rect 315 35754 371 35810
rect 439 35754 495 35810
rect 563 35754 619 35810
rect 687 35754 743 35810
rect 811 35754 867 35810
rect 935 35754 991 35810
rect 1059 35754 1115 35810
rect 1183 35754 1239 35810
rect 1307 35754 1363 35810
rect 1431 35754 1487 35810
rect 1555 35754 1611 35810
rect 1679 35754 1735 35810
rect 1803 35754 1859 35810
rect 1927 35754 1983 35810
rect 2051 35754 2107 35810
rect 315 35630 371 35686
rect 439 35630 495 35686
rect 563 35630 619 35686
rect 687 35630 743 35686
rect 811 35630 867 35686
rect 935 35630 991 35686
rect 1059 35630 1115 35686
rect 1183 35630 1239 35686
rect 1307 35630 1363 35686
rect 1431 35630 1487 35686
rect 1555 35630 1611 35686
rect 1679 35630 1735 35686
rect 1803 35630 1859 35686
rect 1927 35630 1983 35686
rect 2051 35630 2107 35686
rect 315 35506 371 35562
rect 439 35506 495 35562
rect 563 35506 619 35562
rect 687 35506 743 35562
rect 811 35506 867 35562
rect 935 35506 991 35562
rect 1059 35506 1115 35562
rect 1183 35506 1239 35562
rect 1307 35506 1363 35562
rect 1431 35506 1487 35562
rect 1555 35506 1611 35562
rect 1679 35506 1735 35562
rect 1803 35506 1859 35562
rect 1927 35506 1983 35562
rect 2051 35506 2107 35562
rect 315 35382 371 35438
rect 439 35382 495 35438
rect 563 35382 619 35438
rect 687 35382 743 35438
rect 811 35382 867 35438
rect 935 35382 991 35438
rect 1059 35382 1115 35438
rect 1183 35382 1239 35438
rect 1307 35382 1363 35438
rect 1431 35382 1487 35438
rect 1555 35382 1611 35438
rect 1679 35382 1735 35438
rect 1803 35382 1859 35438
rect 1927 35382 1983 35438
rect 2051 35382 2107 35438
rect 315 35258 371 35314
rect 439 35258 495 35314
rect 563 35258 619 35314
rect 687 35258 743 35314
rect 811 35258 867 35314
rect 935 35258 991 35314
rect 1059 35258 1115 35314
rect 1183 35258 1239 35314
rect 1307 35258 1363 35314
rect 1431 35258 1487 35314
rect 1555 35258 1611 35314
rect 1679 35258 1735 35314
rect 1803 35258 1859 35314
rect 1927 35258 1983 35314
rect 2051 35258 2107 35314
rect 315 35134 371 35190
rect 439 35134 495 35190
rect 563 35134 619 35190
rect 687 35134 743 35190
rect 811 35134 867 35190
rect 935 35134 991 35190
rect 1059 35134 1115 35190
rect 1183 35134 1239 35190
rect 1307 35134 1363 35190
rect 1431 35134 1487 35190
rect 1555 35134 1611 35190
rect 1679 35134 1735 35190
rect 1803 35134 1859 35190
rect 1927 35134 1983 35190
rect 2051 35134 2107 35190
rect 315 35010 371 35066
rect 439 35010 495 35066
rect 563 35010 619 35066
rect 687 35010 743 35066
rect 811 35010 867 35066
rect 935 35010 991 35066
rect 1059 35010 1115 35066
rect 1183 35010 1239 35066
rect 1307 35010 1363 35066
rect 1431 35010 1487 35066
rect 1555 35010 1611 35066
rect 1679 35010 1735 35066
rect 1803 35010 1859 35066
rect 1927 35010 1983 35066
rect 2051 35010 2107 35066
rect 315 34886 371 34942
rect 439 34886 495 34942
rect 563 34886 619 34942
rect 687 34886 743 34942
rect 811 34886 867 34942
rect 935 34886 991 34942
rect 1059 34886 1115 34942
rect 1183 34886 1239 34942
rect 1307 34886 1363 34942
rect 1431 34886 1487 34942
rect 1555 34886 1611 34942
rect 1679 34886 1735 34942
rect 1803 34886 1859 34942
rect 1927 34886 1983 34942
rect 2051 34886 2107 34942
rect 315 34762 371 34818
rect 439 34762 495 34818
rect 563 34762 619 34818
rect 687 34762 743 34818
rect 811 34762 867 34818
rect 935 34762 991 34818
rect 1059 34762 1115 34818
rect 1183 34762 1239 34818
rect 1307 34762 1363 34818
rect 1431 34762 1487 34818
rect 1555 34762 1611 34818
rect 1679 34762 1735 34818
rect 1803 34762 1859 34818
rect 1927 34762 1983 34818
rect 2051 34762 2107 34818
rect 315 34638 371 34694
rect 439 34638 495 34694
rect 563 34638 619 34694
rect 687 34638 743 34694
rect 811 34638 867 34694
rect 935 34638 991 34694
rect 1059 34638 1115 34694
rect 1183 34638 1239 34694
rect 1307 34638 1363 34694
rect 1431 34638 1487 34694
rect 1555 34638 1611 34694
rect 1679 34638 1735 34694
rect 1803 34638 1859 34694
rect 1927 34638 1983 34694
rect 2051 34638 2107 34694
rect 315 34514 371 34570
rect 439 34514 495 34570
rect 563 34514 619 34570
rect 687 34514 743 34570
rect 811 34514 867 34570
rect 935 34514 991 34570
rect 1059 34514 1115 34570
rect 1183 34514 1239 34570
rect 1307 34514 1363 34570
rect 1431 34514 1487 34570
rect 1555 34514 1611 34570
rect 1679 34514 1735 34570
rect 1803 34514 1859 34570
rect 1927 34514 1983 34570
rect 2051 34514 2107 34570
rect 315 34390 371 34446
rect 439 34390 495 34446
rect 563 34390 619 34446
rect 687 34390 743 34446
rect 811 34390 867 34446
rect 935 34390 991 34446
rect 1059 34390 1115 34446
rect 1183 34390 1239 34446
rect 1307 34390 1363 34446
rect 1431 34390 1487 34446
rect 1555 34390 1611 34446
rect 1679 34390 1735 34446
rect 1803 34390 1859 34446
rect 1927 34390 1983 34446
rect 2051 34390 2107 34446
rect 315 34266 371 34322
rect 439 34266 495 34322
rect 563 34266 619 34322
rect 687 34266 743 34322
rect 811 34266 867 34322
rect 935 34266 991 34322
rect 1059 34266 1115 34322
rect 1183 34266 1239 34322
rect 1307 34266 1363 34322
rect 1431 34266 1487 34322
rect 1555 34266 1611 34322
rect 1679 34266 1735 34322
rect 1803 34266 1859 34322
rect 1927 34266 1983 34322
rect 2051 34266 2107 34322
rect 315 34142 371 34198
rect 439 34142 495 34198
rect 563 34142 619 34198
rect 687 34142 743 34198
rect 811 34142 867 34198
rect 935 34142 991 34198
rect 1059 34142 1115 34198
rect 1183 34142 1239 34198
rect 1307 34142 1363 34198
rect 1431 34142 1487 34198
rect 1555 34142 1611 34198
rect 1679 34142 1735 34198
rect 1803 34142 1859 34198
rect 1927 34142 1983 34198
rect 2051 34142 2107 34198
rect 315 34018 371 34074
rect 439 34018 495 34074
rect 563 34018 619 34074
rect 687 34018 743 34074
rect 811 34018 867 34074
rect 935 34018 991 34074
rect 1059 34018 1115 34074
rect 1183 34018 1239 34074
rect 1307 34018 1363 34074
rect 1431 34018 1487 34074
rect 1555 34018 1611 34074
rect 1679 34018 1735 34074
rect 1803 34018 1859 34074
rect 1927 34018 1983 34074
rect 2051 34018 2107 34074
rect 315 33894 371 33950
rect 439 33894 495 33950
rect 563 33894 619 33950
rect 687 33894 743 33950
rect 811 33894 867 33950
rect 935 33894 991 33950
rect 1059 33894 1115 33950
rect 1183 33894 1239 33950
rect 1307 33894 1363 33950
rect 1431 33894 1487 33950
rect 1555 33894 1611 33950
rect 1679 33894 1735 33950
rect 1803 33894 1859 33950
rect 1927 33894 1983 33950
rect 2051 33894 2107 33950
rect 315 33770 371 33826
rect 439 33770 495 33826
rect 563 33770 619 33826
rect 687 33770 743 33826
rect 811 33770 867 33826
rect 935 33770 991 33826
rect 1059 33770 1115 33826
rect 1183 33770 1239 33826
rect 1307 33770 1363 33826
rect 1431 33770 1487 33826
rect 1555 33770 1611 33826
rect 1679 33770 1735 33826
rect 1803 33770 1859 33826
rect 1927 33770 1983 33826
rect 2051 33770 2107 33826
rect 315 33646 371 33702
rect 439 33646 495 33702
rect 563 33646 619 33702
rect 687 33646 743 33702
rect 811 33646 867 33702
rect 935 33646 991 33702
rect 1059 33646 1115 33702
rect 1183 33646 1239 33702
rect 1307 33646 1363 33702
rect 1431 33646 1487 33702
rect 1555 33646 1611 33702
rect 1679 33646 1735 33702
rect 1803 33646 1859 33702
rect 1927 33646 1983 33702
rect 2051 33646 2107 33702
rect 2808 36498 2864 36554
rect 2932 36498 2988 36554
rect 3056 36498 3112 36554
rect 3180 36498 3236 36554
rect 3304 36498 3360 36554
rect 3428 36498 3484 36554
rect 3552 36498 3608 36554
rect 3676 36498 3732 36554
rect 3800 36498 3856 36554
rect 3924 36498 3980 36554
rect 4048 36498 4104 36554
rect 4172 36498 4228 36554
rect 4296 36498 4352 36554
rect 4420 36498 4476 36554
rect 4544 36498 4600 36554
rect 4668 36498 4724 36554
rect 2808 36374 2864 36430
rect 2932 36374 2988 36430
rect 3056 36374 3112 36430
rect 3180 36374 3236 36430
rect 3304 36374 3360 36430
rect 3428 36374 3484 36430
rect 3552 36374 3608 36430
rect 3676 36374 3732 36430
rect 3800 36374 3856 36430
rect 3924 36374 3980 36430
rect 4048 36374 4104 36430
rect 4172 36374 4228 36430
rect 4296 36374 4352 36430
rect 4420 36374 4476 36430
rect 4544 36374 4600 36430
rect 4668 36374 4724 36430
rect 2808 36250 2864 36306
rect 2932 36250 2988 36306
rect 3056 36250 3112 36306
rect 3180 36250 3236 36306
rect 3304 36250 3360 36306
rect 3428 36250 3484 36306
rect 3552 36250 3608 36306
rect 3676 36250 3732 36306
rect 3800 36250 3856 36306
rect 3924 36250 3980 36306
rect 4048 36250 4104 36306
rect 4172 36250 4228 36306
rect 4296 36250 4352 36306
rect 4420 36250 4476 36306
rect 4544 36250 4600 36306
rect 4668 36250 4724 36306
rect 2808 36126 2864 36182
rect 2932 36126 2988 36182
rect 3056 36126 3112 36182
rect 3180 36126 3236 36182
rect 3304 36126 3360 36182
rect 3428 36126 3484 36182
rect 3552 36126 3608 36182
rect 3676 36126 3732 36182
rect 3800 36126 3856 36182
rect 3924 36126 3980 36182
rect 4048 36126 4104 36182
rect 4172 36126 4228 36182
rect 4296 36126 4352 36182
rect 4420 36126 4476 36182
rect 4544 36126 4600 36182
rect 4668 36126 4724 36182
rect 2808 36002 2864 36058
rect 2932 36002 2988 36058
rect 3056 36002 3112 36058
rect 3180 36002 3236 36058
rect 3304 36002 3360 36058
rect 3428 36002 3484 36058
rect 3552 36002 3608 36058
rect 3676 36002 3732 36058
rect 3800 36002 3856 36058
rect 3924 36002 3980 36058
rect 4048 36002 4104 36058
rect 4172 36002 4228 36058
rect 4296 36002 4352 36058
rect 4420 36002 4476 36058
rect 4544 36002 4600 36058
rect 4668 36002 4724 36058
rect 2808 35878 2864 35934
rect 2932 35878 2988 35934
rect 3056 35878 3112 35934
rect 3180 35878 3236 35934
rect 3304 35878 3360 35934
rect 3428 35878 3484 35934
rect 3552 35878 3608 35934
rect 3676 35878 3732 35934
rect 3800 35878 3856 35934
rect 3924 35878 3980 35934
rect 4048 35878 4104 35934
rect 4172 35878 4228 35934
rect 4296 35878 4352 35934
rect 4420 35878 4476 35934
rect 4544 35878 4600 35934
rect 4668 35878 4724 35934
rect 2808 35754 2864 35810
rect 2932 35754 2988 35810
rect 3056 35754 3112 35810
rect 3180 35754 3236 35810
rect 3304 35754 3360 35810
rect 3428 35754 3484 35810
rect 3552 35754 3608 35810
rect 3676 35754 3732 35810
rect 3800 35754 3856 35810
rect 3924 35754 3980 35810
rect 4048 35754 4104 35810
rect 4172 35754 4228 35810
rect 4296 35754 4352 35810
rect 4420 35754 4476 35810
rect 4544 35754 4600 35810
rect 4668 35754 4724 35810
rect 2808 35630 2864 35686
rect 2932 35630 2988 35686
rect 3056 35630 3112 35686
rect 3180 35630 3236 35686
rect 3304 35630 3360 35686
rect 3428 35630 3484 35686
rect 3552 35630 3608 35686
rect 3676 35630 3732 35686
rect 3800 35630 3856 35686
rect 3924 35630 3980 35686
rect 4048 35630 4104 35686
rect 4172 35630 4228 35686
rect 4296 35630 4352 35686
rect 4420 35630 4476 35686
rect 4544 35630 4600 35686
rect 4668 35630 4724 35686
rect 2808 35506 2864 35562
rect 2932 35506 2988 35562
rect 3056 35506 3112 35562
rect 3180 35506 3236 35562
rect 3304 35506 3360 35562
rect 3428 35506 3484 35562
rect 3552 35506 3608 35562
rect 3676 35506 3732 35562
rect 3800 35506 3856 35562
rect 3924 35506 3980 35562
rect 4048 35506 4104 35562
rect 4172 35506 4228 35562
rect 4296 35506 4352 35562
rect 4420 35506 4476 35562
rect 4544 35506 4600 35562
rect 4668 35506 4724 35562
rect 2808 35382 2864 35438
rect 2932 35382 2988 35438
rect 3056 35382 3112 35438
rect 3180 35382 3236 35438
rect 3304 35382 3360 35438
rect 3428 35382 3484 35438
rect 3552 35382 3608 35438
rect 3676 35382 3732 35438
rect 3800 35382 3856 35438
rect 3924 35382 3980 35438
rect 4048 35382 4104 35438
rect 4172 35382 4228 35438
rect 4296 35382 4352 35438
rect 4420 35382 4476 35438
rect 4544 35382 4600 35438
rect 4668 35382 4724 35438
rect 2808 35258 2864 35314
rect 2932 35258 2988 35314
rect 3056 35258 3112 35314
rect 3180 35258 3236 35314
rect 3304 35258 3360 35314
rect 3428 35258 3484 35314
rect 3552 35258 3608 35314
rect 3676 35258 3732 35314
rect 3800 35258 3856 35314
rect 3924 35258 3980 35314
rect 4048 35258 4104 35314
rect 4172 35258 4228 35314
rect 4296 35258 4352 35314
rect 4420 35258 4476 35314
rect 4544 35258 4600 35314
rect 4668 35258 4724 35314
rect 2808 35134 2864 35190
rect 2932 35134 2988 35190
rect 3056 35134 3112 35190
rect 3180 35134 3236 35190
rect 3304 35134 3360 35190
rect 3428 35134 3484 35190
rect 3552 35134 3608 35190
rect 3676 35134 3732 35190
rect 3800 35134 3856 35190
rect 3924 35134 3980 35190
rect 4048 35134 4104 35190
rect 4172 35134 4228 35190
rect 4296 35134 4352 35190
rect 4420 35134 4476 35190
rect 4544 35134 4600 35190
rect 4668 35134 4724 35190
rect 2808 35010 2864 35066
rect 2932 35010 2988 35066
rect 3056 35010 3112 35066
rect 3180 35010 3236 35066
rect 3304 35010 3360 35066
rect 3428 35010 3484 35066
rect 3552 35010 3608 35066
rect 3676 35010 3732 35066
rect 3800 35010 3856 35066
rect 3924 35010 3980 35066
rect 4048 35010 4104 35066
rect 4172 35010 4228 35066
rect 4296 35010 4352 35066
rect 4420 35010 4476 35066
rect 4544 35010 4600 35066
rect 4668 35010 4724 35066
rect 2808 34886 2864 34942
rect 2932 34886 2988 34942
rect 3056 34886 3112 34942
rect 3180 34886 3236 34942
rect 3304 34886 3360 34942
rect 3428 34886 3484 34942
rect 3552 34886 3608 34942
rect 3676 34886 3732 34942
rect 3800 34886 3856 34942
rect 3924 34886 3980 34942
rect 4048 34886 4104 34942
rect 4172 34886 4228 34942
rect 4296 34886 4352 34942
rect 4420 34886 4476 34942
rect 4544 34886 4600 34942
rect 4668 34886 4724 34942
rect 2808 34762 2864 34818
rect 2932 34762 2988 34818
rect 3056 34762 3112 34818
rect 3180 34762 3236 34818
rect 3304 34762 3360 34818
rect 3428 34762 3484 34818
rect 3552 34762 3608 34818
rect 3676 34762 3732 34818
rect 3800 34762 3856 34818
rect 3924 34762 3980 34818
rect 4048 34762 4104 34818
rect 4172 34762 4228 34818
rect 4296 34762 4352 34818
rect 4420 34762 4476 34818
rect 4544 34762 4600 34818
rect 4668 34762 4724 34818
rect 2808 34638 2864 34694
rect 2932 34638 2988 34694
rect 3056 34638 3112 34694
rect 3180 34638 3236 34694
rect 3304 34638 3360 34694
rect 3428 34638 3484 34694
rect 3552 34638 3608 34694
rect 3676 34638 3732 34694
rect 3800 34638 3856 34694
rect 3924 34638 3980 34694
rect 4048 34638 4104 34694
rect 4172 34638 4228 34694
rect 4296 34638 4352 34694
rect 4420 34638 4476 34694
rect 4544 34638 4600 34694
rect 4668 34638 4724 34694
rect 2808 34514 2864 34570
rect 2932 34514 2988 34570
rect 3056 34514 3112 34570
rect 3180 34514 3236 34570
rect 3304 34514 3360 34570
rect 3428 34514 3484 34570
rect 3552 34514 3608 34570
rect 3676 34514 3732 34570
rect 3800 34514 3856 34570
rect 3924 34514 3980 34570
rect 4048 34514 4104 34570
rect 4172 34514 4228 34570
rect 4296 34514 4352 34570
rect 4420 34514 4476 34570
rect 4544 34514 4600 34570
rect 4668 34514 4724 34570
rect 2808 34390 2864 34446
rect 2932 34390 2988 34446
rect 3056 34390 3112 34446
rect 3180 34390 3236 34446
rect 3304 34390 3360 34446
rect 3428 34390 3484 34446
rect 3552 34390 3608 34446
rect 3676 34390 3732 34446
rect 3800 34390 3856 34446
rect 3924 34390 3980 34446
rect 4048 34390 4104 34446
rect 4172 34390 4228 34446
rect 4296 34390 4352 34446
rect 4420 34390 4476 34446
rect 4544 34390 4600 34446
rect 4668 34390 4724 34446
rect 2808 34266 2864 34322
rect 2932 34266 2988 34322
rect 3056 34266 3112 34322
rect 3180 34266 3236 34322
rect 3304 34266 3360 34322
rect 3428 34266 3484 34322
rect 3552 34266 3608 34322
rect 3676 34266 3732 34322
rect 3800 34266 3856 34322
rect 3924 34266 3980 34322
rect 4048 34266 4104 34322
rect 4172 34266 4228 34322
rect 4296 34266 4352 34322
rect 4420 34266 4476 34322
rect 4544 34266 4600 34322
rect 4668 34266 4724 34322
rect 2808 34142 2864 34198
rect 2932 34142 2988 34198
rect 3056 34142 3112 34198
rect 3180 34142 3236 34198
rect 3304 34142 3360 34198
rect 3428 34142 3484 34198
rect 3552 34142 3608 34198
rect 3676 34142 3732 34198
rect 3800 34142 3856 34198
rect 3924 34142 3980 34198
rect 4048 34142 4104 34198
rect 4172 34142 4228 34198
rect 4296 34142 4352 34198
rect 4420 34142 4476 34198
rect 4544 34142 4600 34198
rect 4668 34142 4724 34198
rect 2808 34018 2864 34074
rect 2932 34018 2988 34074
rect 3056 34018 3112 34074
rect 3180 34018 3236 34074
rect 3304 34018 3360 34074
rect 3428 34018 3484 34074
rect 3552 34018 3608 34074
rect 3676 34018 3732 34074
rect 3800 34018 3856 34074
rect 3924 34018 3980 34074
rect 4048 34018 4104 34074
rect 4172 34018 4228 34074
rect 4296 34018 4352 34074
rect 4420 34018 4476 34074
rect 4544 34018 4600 34074
rect 4668 34018 4724 34074
rect 2808 33894 2864 33950
rect 2932 33894 2988 33950
rect 3056 33894 3112 33950
rect 3180 33894 3236 33950
rect 3304 33894 3360 33950
rect 3428 33894 3484 33950
rect 3552 33894 3608 33950
rect 3676 33894 3732 33950
rect 3800 33894 3856 33950
rect 3924 33894 3980 33950
rect 4048 33894 4104 33950
rect 4172 33894 4228 33950
rect 4296 33894 4352 33950
rect 4420 33894 4476 33950
rect 4544 33894 4600 33950
rect 4668 33894 4724 33950
rect 2808 33770 2864 33826
rect 2932 33770 2988 33826
rect 3056 33770 3112 33826
rect 3180 33770 3236 33826
rect 3304 33770 3360 33826
rect 3428 33770 3484 33826
rect 3552 33770 3608 33826
rect 3676 33770 3732 33826
rect 3800 33770 3856 33826
rect 3924 33770 3980 33826
rect 4048 33770 4104 33826
rect 4172 33770 4228 33826
rect 4296 33770 4352 33826
rect 4420 33770 4476 33826
rect 4544 33770 4600 33826
rect 4668 33770 4724 33826
rect 2808 33646 2864 33702
rect 2932 33646 2988 33702
rect 3056 33646 3112 33702
rect 3180 33646 3236 33702
rect 3304 33646 3360 33702
rect 3428 33646 3484 33702
rect 3552 33646 3608 33702
rect 3676 33646 3732 33702
rect 3800 33646 3856 33702
rect 3924 33646 3980 33702
rect 4048 33646 4104 33702
rect 4172 33646 4228 33702
rect 4296 33646 4352 33702
rect 4420 33646 4476 33702
rect 4544 33646 4600 33702
rect 4668 33646 4724 33702
rect 5178 36498 5234 36554
rect 5302 36498 5358 36554
rect 5426 36498 5482 36554
rect 5550 36498 5606 36554
rect 5674 36498 5730 36554
rect 5798 36498 5854 36554
rect 5922 36498 5978 36554
rect 6046 36498 6102 36554
rect 6170 36498 6226 36554
rect 6294 36498 6350 36554
rect 6418 36498 6474 36554
rect 6542 36498 6598 36554
rect 6666 36498 6722 36554
rect 6790 36498 6846 36554
rect 6914 36498 6970 36554
rect 7038 36498 7094 36554
rect 5178 36374 5234 36430
rect 5302 36374 5358 36430
rect 5426 36374 5482 36430
rect 5550 36374 5606 36430
rect 5674 36374 5730 36430
rect 5798 36374 5854 36430
rect 5922 36374 5978 36430
rect 6046 36374 6102 36430
rect 6170 36374 6226 36430
rect 6294 36374 6350 36430
rect 6418 36374 6474 36430
rect 6542 36374 6598 36430
rect 6666 36374 6722 36430
rect 6790 36374 6846 36430
rect 6914 36374 6970 36430
rect 7038 36374 7094 36430
rect 5178 36250 5234 36306
rect 5302 36250 5358 36306
rect 5426 36250 5482 36306
rect 5550 36250 5606 36306
rect 5674 36250 5730 36306
rect 5798 36250 5854 36306
rect 5922 36250 5978 36306
rect 6046 36250 6102 36306
rect 6170 36250 6226 36306
rect 6294 36250 6350 36306
rect 6418 36250 6474 36306
rect 6542 36250 6598 36306
rect 6666 36250 6722 36306
rect 6790 36250 6846 36306
rect 6914 36250 6970 36306
rect 7038 36250 7094 36306
rect 5178 36126 5234 36182
rect 5302 36126 5358 36182
rect 5426 36126 5482 36182
rect 5550 36126 5606 36182
rect 5674 36126 5730 36182
rect 5798 36126 5854 36182
rect 5922 36126 5978 36182
rect 6046 36126 6102 36182
rect 6170 36126 6226 36182
rect 6294 36126 6350 36182
rect 6418 36126 6474 36182
rect 6542 36126 6598 36182
rect 6666 36126 6722 36182
rect 6790 36126 6846 36182
rect 6914 36126 6970 36182
rect 7038 36126 7094 36182
rect 5178 36002 5234 36058
rect 5302 36002 5358 36058
rect 5426 36002 5482 36058
rect 5550 36002 5606 36058
rect 5674 36002 5730 36058
rect 5798 36002 5854 36058
rect 5922 36002 5978 36058
rect 6046 36002 6102 36058
rect 6170 36002 6226 36058
rect 6294 36002 6350 36058
rect 6418 36002 6474 36058
rect 6542 36002 6598 36058
rect 6666 36002 6722 36058
rect 6790 36002 6846 36058
rect 6914 36002 6970 36058
rect 7038 36002 7094 36058
rect 5178 35878 5234 35934
rect 5302 35878 5358 35934
rect 5426 35878 5482 35934
rect 5550 35878 5606 35934
rect 5674 35878 5730 35934
rect 5798 35878 5854 35934
rect 5922 35878 5978 35934
rect 6046 35878 6102 35934
rect 6170 35878 6226 35934
rect 6294 35878 6350 35934
rect 6418 35878 6474 35934
rect 6542 35878 6598 35934
rect 6666 35878 6722 35934
rect 6790 35878 6846 35934
rect 6914 35878 6970 35934
rect 7038 35878 7094 35934
rect 5178 35754 5234 35810
rect 5302 35754 5358 35810
rect 5426 35754 5482 35810
rect 5550 35754 5606 35810
rect 5674 35754 5730 35810
rect 5798 35754 5854 35810
rect 5922 35754 5978 35810
rect 6046 35754 6102 35810
rect 6170 35754 6226 35810
rect 6294 35754 6350 35810
rect 6418 35754 6474 35810
rect 6542 35754 6598 35810
rect 6666 35754 6722 35810
rect 6790 35754 6846 35810
rect 6914 35754 6970 35810
rect 7038 35754 7094 35810
rect 5178 35630 5234 35686
rect 5302 35630 5358 35686
rect 5426 35630 5482 35686
rect 5550 35630 5606 35686
rect 5674 35630 5730 35686
rect 5798 35630 5854 35686
rect 5922 35630 5978 35686
rect 6046 35630 6102 35686
rect 6170 35630 6226 35686
rect 6294 35630 6350 35686
rect 6418 35630 6474 35686
rect 6542 35630 6598 35686
rect 6666 35630 6722 35686
rect 6790 35630 6846 35686
rect 6914 35630 6970 35686
rect 7038 35630 7094 35686
rect 5178 35506 5234 35562
rect 5302 35506 5358 35562
rect 5426 35506 5482 35562
rect 5550 35506 5606 35562
rect 5674 35506 5730 35562
rect 5798 35506 5854 35562
rect 5922 35506 5978 35562
rect 6046 35506 6102 35562
rect 6170 35506 6226 35562
rect 6294 35506 6350 35562
rect 6418 35506 6474 35562
rect 6542 35506 6598 35562
rect 6666 35506 6722 35562
rect 6790 35506 6846 35562
rect 6914 35506 6970 35562
rect 7038 35506 7094 35562
rect 5178 35382 5234 35438
rect 5302 35382 5358 35438
rect 5426 35382 5482 35438
rect 5550 35382 5606 35438
rect 5674 35382 5730 35438
rect 5798 35382 5854 35438
rect 5922 35382 5978 35438
rect 6046 35382 6102 35438
rect 6170 35382 6226 35438
rect 6294 35382 6350 35438
rect 6418 35382 6474 35438
rect 6542 35382 6598 35438
rect 6666 35382 6722 35438
rect 6790 35382 6846 35438
rect 6914 35382 6970 35438
rect 7038 35382 7094 35438
rect 5178 35258 5234 35314
rect 5302 35258 5358 35314
rect 5426 35258 5482 35314
rect 5550 35258 5606 35314
rect 5674 35258 5730 35314
rect 5798 35258 5854 35314
rect 5922 35258 5978 35314
rect 6046 35258 6102 35314
rect 6170 35258 6226 35314
rect 6294 35258 6350 35314
rect 6418 35258 6474 35314
rect 6542 35258 6598 35314
rect 6666 35258 6722 35314
rect 6790 35258 6846 35314
rect 6914 35258 6970 35314
rect 7038 35258 7094 35314
rect 5178 35134 5234 35190
rect 5302 35134 5358 35190
rect 5426 35134 5482 35190
rect 5550 35134 5606 35190
rect 5674 35134 5730 35190
rect 5798 35134 5854 35190
rect 5922 35134 5978 35190
rect 6046 35134 6102 35190
rect 6170 35134 6226 35190
rect 6294 35134 6350 35190
rect 6418 35134 6474 35190
rect 6542 35134 6598 35190
rect 6666 35134 6722 35190
rect 6790 35134 6846 35190
rect 6914 35134 6970 35190
rect 7038 35134 7094 35190
rect 5178 35010 5234 35066
rect 5302 35010 5358 35066
rect 5426 35010 5482 35066
rect 5550 35010 5606 35066
rect 5674 35010 5730 35066
rect 5798 35010 5854 35066
rect 5922 35010 5978 35066
rect 6046 35010 6102 35066
rect 6170 35010 6226 35066
rect 6294 35010 6350 35066
rect 6418 35010 6474 35066
rect 6542 35010 6598 35066
rect 6666 35010 6722 35066
rect 6790 35010 6846 35066
rect 6914 35010 6970 35066
rect 7038 35010 7094 35066
rect 5178 34886 5234 34942
rect 5302 34886 5358 34942
rect 5426 34886 5482 34942
rect 5550 34886 5606 34942
rect 5674 34886 5730 34942
rect 5798 34886 5854 34942
rect 5922 34886 5978 34942
rect 6046 34886 6102 34942
rect 6170 34886 6226 34942
rect 6294 34886 6350 34942
rect 6418 34886 6474 34942
rect 6542 34886 6598 34942
rect 6666 34886 6722 34942
rect 6790 34886 6846 34942
rect 6914 34886 6970 34942
rect 7038 34886 7094 34942
rect 5178 34762 5234 34818
rect 5302 34762 5358 34818
rect 5426 34762 5482 34818
rect 5550 34762 5606 34818
rect 5674 34762 5730 34818
rect 5798 34762 5854 34818
rect 5922 34762 5978 34818
rect 6046 34762 6102 34818
rect 6170 34762 6226 34818
rect 6294 34762 6350 34818
rect 6418 34762 6474 34818
rect 6542 34762 6598 34818
rect 6666 34762 6722 34818
rect 6790 34762 6846 34818
rect 6914 34762 6970 34818
rect 7038 34762 7094 34818
rect 5178 34638 5234 34694
rect 5302 34638 5358 34694
rect 5426 34638 5482 34694
rect 5550 34638 5606 34694
rect 5674 34638 5730 34694
rect 5798 34638 5854 34694
rect 5922 34638 5978 34694
rect 6046 34638 6102 34694
rect 6170 34638 6226 34694
rect 6294 34638 6350 34694
rect 6418 34638 6474 34694
rect 6542 34638 6598 34694
rect 6666 34638 6722 34694
rect 6790 34638 6846 34694
rect 6914 34638 6970 34694
rect 7038 34638 7094 34694
rect 5178 34514 5234 34570
rect 5302 34514 5358 34570
rect 5426 34514 5482 34570
rect 5550 34514 5606 34570
rect 5674 34514 5730 34570
rect 5798 34514 5854 34570
rect 5922 34514 5978 34570
rect 6046 34514 6102 34570
rect 6170 34514 6226 34570
rect 6294 34514 6350 34570
rect 6418 34514 6474 34570
rect 6542 34514 6598 34570
rect 6666 34514 6722 34570
rect 6790 34514 6846 34570
rect 6914 34514 6970 34570
rect 7038 34514 7094 34570
rect 5178 34390 5234 34446
rect 5302 34390 5358 34446
rect 5426 34390 5482 34446
rect 5550 34390 5606 34446
rect 5674 34390 5730 34446
rect 5798 34390 5854 34446
rect 5922 34390 5978 34446
rect 6046 34390 6102 34446
rect 6170 34390 6226 34446
rect 6294 34390 6350 34446
rect 6418 34390 6474 34446
rect 6542 34390 6598 34446
rect 6666 34390 6722 34446
rect 6790 34390 6846 34446
rect 6914 34390 6970 34446
rect 7038 34390 7094 34446
rect 5178 34266 5234 34322
rect 5302 34266 5358 34322
rect 5426 34266 5482 34322
rect 5550 34266 5606 34322
rect 5674 34266 5730 34322
rect 5798 34266 5854 34322
rect 5922 34266 5978 34322
rect 6046 34266 6102 34322
rect 6170 34266 6226 34322
rect 6294 34266 6350 34322
rect 6418 34266 6474 34322
rect 6542 34266 6598 34322
rect 6666 34266 6722 34322
rect 6790 34266 6846 34322
rect 6914 34266 6970 34322
rect 7038 34266 7094 34322
rect 5178 34142 5234 34198
rect 5302 34142 5358 34198
rect 5426 34142 5482 34198
rect 5550 34142 5606 34198
rect 5674 34142 5730 34198
rect 5798 34142 5854 34198
rect 5922 34142 5978 34198
rect 6046 34142 6102 34198
rect 6170 34142 6226 34198
rect 6294 34142 6350 34198
rect 6418 34142 6474 34198
rect 6542 34142 6598 34198
rect 6666 34142 6722 34198
rect 6790 34142 6846 34198
rect 6914 34142 6970 34198
rect 7038 34142 7094 34198
rect 5178 34018 5234 34074
rect 5302 34018 5358 34074
rect 5426 34018 5482 34074
rect 5550 34018 5606 34074
rect 5674 34018 5730 34074
rect 5798 34018 5854 34074
rect 5922 34018 5978 34074
rect 6046 34018 6102 34074
rect 6170 34018 6226 34074
rect 6294 34018 6350 34074
rect 6418 34018 6474 34074
rect 6542 34018 6598 34074
rect 6666 34018 6722 34074
rect 6790 34018 6846 34074
rect 6914 34018 6970 34074
rect 7038 34018 7094 34074
rect 5178 33894 5234 33950
rect 5302 33894 5358 33950
rect 5426 33894 5482 33950
rect 5550 33894 5606 33950
rect 5674 33894 5730 33950
rect 5798 33894 5854 33950
rect 5922 33894 5978 33950
rect 6046 33894 6102 33950
rect 6170 33894 6226 33950
rect 6294 33894 6350 33950
rect 6418 33894 6474 33950
rect 6542 33894 6598 33950
rect 6666 33894 6722 33950
rect 6790 33894 6846 33950
rect 6914 33894 6970 33950
rect 7038 33894 7094 33950
rect 5178 33770 5234 33826
rect 5302 33770 5358 33826
rect 5426 33770 5482 33826
rect 5550 33770 5606 33826
rect 5674 33770 5730 33826
rect 5798 33770 5854 33826
rect 5922 33770 5978 33826
rect 6046 33770 6102 33826
rect 6170 33770 6226 33826
rect 6294 33770 6350 33826
rect 6418 33770 6474 33826
rect 6542 33770 6598 33826
rect 6666 33770 6722 33826
rect 6790 33770 6846 33826
rect 6914 33770 6970 33826
rect 7038 33770 7094 33826
rect 5178 33646 5234 33702
rect 5302 33646 5358 33702
rect 5426 33646 5482 33702
rect 5550 33646 5606 33702
rect 5674 33646 5730 33702
rect 5798 33646 5854 33702
rect 5922 33646 5978 33702
rect 6046 33646 6102 33702
rect 6170 33646 6226 33702
rect 6294 33646 6350 33702
rect 6418 33646 6474 33702
rect 6542 33646 6598 33702
rect 6666 33646 6722 33702
rect 6790 33646 6846 33702
rect 6914 33646 6970 33702
rect 7038 33646 7094 33702
rect 7884 36498 7940 36554
rect 8008 36498 8064 36554
rect 8132 36498 8188 36554
rect 8256 36498 8312 36554
rect 8380 36498 8436 36554
rect 8504 36498 8560 36554
rect 8628 36498 8684 36554
rect 8752 36498 8808 36554
rect 8876 36498 8932 36554
rect 9000 36498 9056 36554
rect 9124 36498 9180 36554
rect 9248 36498 9304 36554
rect 9372 36498 9428 36554
rect 9496 36498 9552 36554
rect 9620 36498 9676 36554
rect 9744 36498 9800 36554
rect 7884 36374 7940 36430
rect 8008 36374 8064 36430
rect 8132 36374 8188 36430
rect 8256 36374 8312 36430
rect 8380 36374 8436 36430
rect 8504 36374 8560 36430
rect 8628 36374 8684 36430
rect 8752 36374 8808 36430
rect 8876 36374 8932 36430
rect 9000 36374 9056 36430
rect 9124 36374 9180 36430
rect 9248 36374 9304 36430
rect 9372 36374 9428 36430
rect 9496 36374 9552 36430
rect 9620 36374 9676 36430
rect 9744 36374 9800 36430
rect 7884 36250 7940 36306
rect 8008 36250 8064 36306
rect 8132 36250 8188 36306
rect 8256 36250 8312 36306
rect 8380 36250 8436 36306
rect 8504 36250 8560 36306
rect 8628 36250 8684 36306
rect 8752 36250 8808 36306
rect 8876 36250 8932 36306
rect 9000 36250 9056 36306
rect 9124 36250 9180 36306
rect 9248 36250 9304 36306
rect 9372 36250 9428 36306
rect 9496 36250 9552 36306
rect 9620 36250 9676 36306
rect 9744 36250 9800 36306
rect 7884 36126 7940 36182
rect 8008 36126 8064 36182
rect 8132 36126 8188 36182
rect 8256 36126 8312 36182
rect 8380 36126 8436 36182
rect 8504 36126 8560 36182
rect 8628 36126 8684 36182
rect 8752 36126 8808 36182
rect 8876 36126 8932 36182
rect 9000 36126 9056 36182
rect 9124 36126 9180 36182
rect 9248 36126 9304 36182
rect 9372 36126 9428 36182
rect 9496 36126 9552 36182
rect 9620 36126 9676 36182
rect 9744 36126 9800 36182
rect 7884 36002 7940 36058
rect 8008 36002 8064 36058
rect 8132 36002 8188 36058
rect 8256 36002 8312 36058
rect 8380 36002 8436 36058
rect 8504 36002 8560 36058
rect 8628 36002 8684 36058
rect 8752 36002 8808 36058
rect 8876 36002 8932 36058
rect 9000 36002 9056 36058
rect 9124 36002 9180 36058
rect 9248 36002 9304 36058
rect 9372 36002 9428 36058
rect 9496 36002 9552 36058
rect 9620 36002 9676 36058
rect 9744 36002 9800 36058
rect 7884 35878 7940 35934
rect 8008 35878 8064 35934
rect 8132 35878 8188 35934
rect 8256 35878 8312 35934
rect 8380 35878 8436 35934
rect 8504 35878 8560 35934
rect 8628 35878 8684 35934
rect 8752 35878 8808 35934
rect 8876 35878 8932 35934
rect 9000 35878 9056 35934
rect 9124 35878 9180 35934
rect 9248 35878 9304 35934
rect 9372 35878 9428 35934
rect 9496 35878 9552 35934
rect 9620 35878 9676 35934
rect 9744 35878 9800 35934
rect 7884 35754 7940 35810
rect 8008 35754 8064 35810
rect 8132 35754 8188 35810
rect 8256 35754 8312 35810
rect 8380 35754 8436 35810
rect 8504 35754 8560 35810
rect 8628 35754 8684 35810
rect 8752 35754 8808 35810
rect 8876 35754 8932 35810
rect 9000 35754 9056 35810
rect 9124 35754 9180 35810
rect 9248 35754 9304 35810
rect 9372 35754 9428 35810
rect 9496 35754 9552 35810
rect 9620 35754 9676 35810
rect 9744 35754 9800 35810
rect 7884 35630 7940 35686
rect 8008 35630 8064 35686
rect 8132 35630 8188 35686
rect 8256 35630 8312 35686
rect 8380 35630 8436 35686
rect 8504 35630 8560 35686
rect 8628 35630 8684 35686
rect 8752 35630 8808 35686
rect 8876 35630 8932 35686
rect 9000 35630 9056 35686
rect 9124 35630 9180 35686
rect 9248 35630 9304 35686
rect 9372 35630 9428 35686
rect 9496 35630 9552 35686
rect 9620 35630 9676 35686
rect 9744 35630 9800 35686
rect 7884 35506 7940 35562
rect 8008 35506 8064 35562
rect 8132 35506 8188 35562
rect 8256 35506 8312 35562
rect 8380 35506 8436 35562
rect 8504 35506 8560 35562
rect 8628 35506 8684 35562
rect 8752 35506 8808 35562
rect 8876 35506 8932 35562
rect 9000 35506 9056 35562
rect 9124 35506 9180 35562
rect 9248 35506 9304 35562
rect 9372 35506 9428 35562
rect 9496 35506 9552 35562
rect 9620 35506 9676 35562
rect 9744 35506 9800 35562
rect 7884 35382 7940 35438
rect 8008 35382 8064 35438
rect 8132 35382 8188 35438
rect 8256 35382 8312 35438
rect 8380 35382 8436 35438
rect 8504 35382 8560 35438
rect 8628 35382 8684 35438
rect 8752 35382 8808 35438
rect 8876 35382 8932 35438
rect 9000 35382 9056 35438
rect 9124 35382 9180 35438
rect 9248 35382 9304 35438
rect 9372 35382 9428 35438
rect 9496 35382 9552 35438
rect 9620 35382 9676 35438
rect 9744 35382 9800 35438
rect 7884 35258 7940 35314
rect 8008 35258 8064 35314
rect 8132 35258 8188 35314
rect 8256 35258 8312 35314
rect 8380 35258 8436 35314
rect 8504 35258 8560 35314
rect 8628 35258 8684 35314
rect 8752 35258 8808 35314
rect 8876 35258 8932 35314
rect 9000 35258 9056 35314
rect 9124 35258 9180 35314
rect 9248 35258 9304 35314
rect 9372 35258 9428 35314
rect 9496 35258 9552 35314
rect 9620 35258 9676 35314
rect 9744 35258 9800 35314
rect 7884 35134 7940 35190
rect 8008 35134 8064 35190
rect 8132 35134 8188 35190
rect 8256 35134 8312 35190
rect 8380 35134 8436 35190
rect 8504 35134 8560 35190
rect 8628 35134 8684 35190
rect 8752 35134 8808 35190
rect 8876 35134 8932 35190
rect 9000 35134 9056 35190
rect 9124 35134 9180 35190
rect 9248 35134 9304 35190
rect 9372 35134 9428 35190
rect 9496 35134 9552 35190
rect 9620 35134 9676 35190
rect 9744 35134 9800 35190
rect 7884 35010 7940 35066
rect 8008 35010 8064 35066
rect 8132 35010 8188 35066
rect 8256 35010 8312 35066
rect 8380 35010 8436 35066
rect 8504 35010 8560 35066
rect 8628 35010 8684 35066
rect 8752 35010 8808 35066
rect 8876 35010 8932 35066
rect 9000 35010 9056 35066
rect 9124 35010 9180 35066
rect 9248 35010 9304 35066
rect 9372 35010 9428 35066
rect 9496 35010 9552 35066
rect 9620 35010 9676 35066
rect 9744 35010 9800 35066
rect 7884 34886 7940 34942
rect 8008 34886 8064 34942
rect 8132 34886 8188 34942
rect 8256 34886 8312 34942
rect 8380 34886 8436 34942
rect 8504 34886 8560 34942
rect 8628 34886 8684 34942
rect 8752 34886 8808 34942
rect 8876 34886 8932 34942
rect 9000 34886 9056 34942
rect 9124 34886 9180 34942
rect 9248 34886 9304 34942
rect 9372 34886 9428 34942
rect 9496 34886 9552 34942
rect 9620 34886 9676 34942
rect 9744 34886 9800 34942
rect 7884 34762 7940 34818
rect 8008 34762 8064 34818
rect 8132 34762 8188 34818
rect 8256 34762 8312 34818
rect 8380 34762 8436 34818
rect 8504 34762 8560 34818
rect 8628 34762 8684 34818
rect 8752 34762 8808 34818
rect 8876 34762 8932 34818
rect 9000 34762 9056 34818
rect 9124 34762 9180 34818
rect 9248 34762 9304 34818
rect 9372 34762 9428 34818
rect 9496 34762 9552 34818
rect 9620 34762 9676 34818
rect 9744 34762 9800 34818
rect 7884 34638 7940 34694
rect 8008 34638 8064 34694
rect 8132 34638 8188 34694
rect 8256 34638 8312 34694
rect 8380 34638 8436 34694
rect 8504 34638 8560 34694
rect 8628 34638 8684 34694
rect 8752 34638 8808 34694
rect 8876 34638 8932 34694
rect 9000 34638 9056 34694
rect 9124 34638 9180 34694
rect 9248 34638 9304 34694
rect 9372 34638 9428 34694
rect 9496 34638 9552 34694
rect 9620 34638 9676 34694
rect 9744 34638 9800 34694
rect 7884 34514 7940 34570
rect 8008 34514 8064 34570
rect 8132 34514 8188 34570
rect 8256 34514 8312 34570
rect 8380 34514 8436 34570
rect 8504 34514 8560 34570
rect 8628 34514 8684 34570
rect 8752 34514 8808 34570
rect 8876 34514 8932 34570
rect 9000 34514 9056 34570
rect 9124 34514 9180 34570
rect 9248 34514 9304 34570
rect 9372 34514 9428 34570
rect 9496 34514 9552 34570
rect 9620 34514 9676 34570
rect 9744 34514 9800 34570
rect 7884 34390 7940 34446
rect 8008 34390 8064 34446
rect 8132 34390 8188 34446
rect 8256 34390 8312 34446
rect 8380 34390 8436 34446
rect 8504 34390 8560 34446
rect 8628 34390 8684 34446
rect 8752 34390 8808 34446
rect 8876 34390 8932 34446
rect 9000 34390 9056 34446
rect 9124 34390 9180 34446
rect 9248 34390 9304 34446
rect 9372 34390 9428 34446
rect 9496 34390 9552 34446
rect 9620 34390 9676 34446
rect 9744 34390 9800 34446
rect 7884 34266 7940 34322
rect 8008 34266 8064 34322
rect 8132 34266 8188 34322
rect 8256 34266 8312 34322
rect 8380 34266 8436 34322
rect 8504 34266 8560 34322
rect 8628 34266 8684 34322
rect 8752 34266 8808 34322
rect 8876 34266 8932 34322
rect 9000 34266 9056 34322
rect 9124 34266 9180 34322
rect 9248 34266 9304 34322
rect 9372 34266 9428 34322
rect 9496 34266 9552 34322
rect 9620 34266 9676 34322
rect 9744 34266 9800 34322
rect 7884 34142 7940 34198
rect 8008 34142 8064 34198
rect 8132 34142 8188 34198
rect 8256 34142 8312 34198
rect 8380 34142 8436 34198
rect 8504 34142 8560 34198
rect 8628 34142 8684 34198
rect 8752 34142 8808 34198
rect 8876 34142 8932 34198
rect 9000 34142 9056 34198
rect 9124 34142 9180 34198
rect 9248 34142 9304 34198
rect 9372 34142 9428 34198
rect 9496 34142 9552 34198
rect 9620 34142 9676 34198
rect 9744 34142 9800 34198
rect 7884 34018 7940 34074
rect 8008 34018 8064 34074
rect 8132 34018 8188 34074
rect 8256 34018 8312 34074
rect 8380 34018 8436 34074
rect 8504 34018 8560 34074
rect 8628 34018 8684 34074
rect 8752 34018 8808 34074
rect 8876 34018 8932 34074
rect 9000 34018 9056 34074
rect 9124 34018 9180 34074
rect 9248 34018 9304 34074
rect 9372 34018 9428 34074
rect 9496 34018 9552 34074
rect 9620 34018 9676 34074
rect 9744 34018 9800 34074
rect 7884 33894 7940 33950
rect 8008 33894 8064 33950
rect 8132 33894 8188 33950
rect 8256 33894 8312 33950
rect 8380 33894 8436 33950
rect 8504 33894 8560 33950
rect 8628 33894 8684 33950
rect 8752 33894 8808 33950
rect 8876 33894 8932 33950
rect 9000 33894 9056 33950
rect 9124 33894 9180 33950
rect 9248 33894 9304 33950
rect 9372 33894 9428 33950
rect 9496 33894 9552 33950
rect 9620 33894 9676 33950
rect 9744 33894 9800 33950
rect 7884 33770 7940 33826
rect 8008 33770 8064 33826
rect 8132 33770 8188 33826
rect 8256 33770 8312 33826
rect 8380 33770 8436 33826
rect 8504 33770 8560 33826
rect 8628 33770 8684 33826
rect 8752 33770 8808 33826
rect 8876 33770 8932 33826
rect 9000 33770 9056 33826
rect 9124 33770 9180 33826
rect 9248 33770 9304 33826
rect 9372 33770 9428 33826
rect 9496 33770 9552 33826
rect 9620 33770 9676 33826
rect 9744 33770 9800 33826
rect 7884 33646 7940 33702
rect 8008 33646 8064 33702
rect 8132 33646 8188 33702
rect 8256 33646 8312 33702
rect 8380 33646 8436 33702
rect 8504 33646 8560 33702
rect 8628 33646 8684 33702
rect 8752 33646 8808 33702
rect 8876 33646 8932 33702
rect 9000 33646 9056 33702
rect 9124 33646 9180 33702
rect 9248 33646 9304 33702
rect 9372 33646 9428 33702
rect 9496 33646 9552 33702
rect 9620 33646 9676 33702
rect 9744 33646 9800 33702
rect 10254 36498 10310 36554
rect 10378 36498 10434 36554
rect 10502 36498 10558 36554
rect 10626 36498 10682 36554
rect 10750 36498 10806 36554
rect 10874 36498 10930 36554
rect 10998 36498 11054 36554
rect 11122 36498 11178 36554
rect 11246 36498 11302 36554
rect 11370 36498 11426 36554
rect 11494 36498 11550 36554
rect 11618 36498 11674 36554
rect 11742 36498 11798 36554
rect 11866 36498 11922 36554
rect 11990 36498 12046 36554
rect 12114 36498 12170 36554
rect 10254 36374 10310 36430
rect 10378 36374 10434 36430
rect 10502 36374 10558 36430
rect 10626 36374 10682 36430
rect 10750 36374 10806 36430
rect 10874 36374 10930 36430
rect 10998 36374 11054 36430
rect 11122 36374 11178 36430
rect 11246 36374 11302 36430
rect 11370 36374 11426 36430
rect 11494 36374 11550 36430
rect 11618 36374 11674 36430
rect 11742 36374 11798 36430
rect 11866 36374 11922 36430
rect 11990 36374 12046 36430
rect 12114 36374 12170 36430
rect 10254 36250 10310 36306
rect 10378 36250 10434 36306
rect 10502 36250 10558 36306
rect 10626 36250 10682 36306
rect 10750 36250 10806 36306
rect 10874 36250 10930 36306
rect 10998 36250 11054 36306
rect 11122 36250 11178 36306
rect 11246 36250 11302 36306
rect 11370 36250 11426 36306
rect 11494 36250 11550 36306
rect 11618 36250 11674 36306
rect 11742 36250 11798 36306
rect 11866 36250 11922 36306
rect 11990 36250 12046 36306
rect 12114 36250 12170 36306
rect 10254 36126 10310 36182
rect 10378 36126 10434 36182
rect 10502 36126 10558 36182
rect 10626 36126 10682 36182
rect 10750 36126 10806 36182
rect 10874 36126 10930 36182
rect 10998 36126 11054 36182
rect 11122 36126 11178 36182
rect 11246 36126 11302 36182
rect 11370 36126 11426 36182
rect 11494 36126 11550 36182
rect 11618 36126 11674 36182
rect 11742 36126 11798 36182
rect 11866 36126 11922 36182
rect 11990 36126 12046 36182
rect 12114 36126 12170 36182
rect 10254 36002 10310 36058
rect 10378 36002 10434 36058
rect 10502 36002 10558 36058
rect 10626 36002 10682 36058
rect 10750 36002 10806 36058
rect 10874 36002 10930 36058
rect 10998 36002 11054 36058
rect 11122 36002 11178 36058
rect 11246 36002 11302 36058
rect 11370 36002 11426 36058
rect 11494 36002 11550 36058
rect 11618 36002 11674 36058
rect 11742 36002 11798 36058
rect 11866 36002 11922 36058
rect 11990 36002 12046 36058
rect 12114 36002 12170 36058
rect 10254 35878 10310 35934
rect 10378 35878 10434 35934
rect 10502 35878 10558 35934
rect 10626 35878 10682 35934
rect 10750 35878 10806 35934
rect 10874 35878 10930 35934
rect 10998 35878 11054 35934
rect 11122 35878 11178 35934
rect 11246 35878 11302 35934
rect 11370 35878 11426 35934
rect 11494 35878 11550 35934
rect 11618 35878 11674 35934
rect 11742 35878 11798 35934
rect 11866 35878 11922 35934
rect 11990 35878 12046 35934
rect 12114 35878 12170 35934
rect 10254 35754 10310 35810
rect 10378 35754 10434 35810
rect 10502 35754 10558 35810
rect 10626 35754 10682 35810
rect 10750 35754 10806 35810
rect 10874 35754 10930 35810
rect 10998 35754 11054 35810
rect 11122 35754 11178 35810
rect 11246 35754 11302 35810
rect 11370 35754 11426 35810
rect 11494 35754 11550 35810
rect 11618 35754 11674 35810
rect 11742 35754 11798 35810
rect 11866 35754 11922 35810
rect 11990 35754 12046 35810
rect 12114 35754 12170 35810
rect 10254 35630 10310 35686
rect 10378 35630 10434 35686
rect 10502 35630 10558 35686
rect 10626 35630 10682 35686
rect 10750 35630 10806 35686
rect 10874 35630 10930 35686
rect 10998 35630 11054 35686
rect 11122 35630 11178 35686
rect 11246 35630 11302 35686
rect 11370 35630 11426 35686
rect 11494 35630 11550 35686
rect 11618 35630 11674 35686
rect 11742 35630 11798 35686
rect 11866 35630 11922 35686
rect 11990 35630 12046 35686
rect 12114 35630 12170 35686
rect 10254 35506 10310 35562
rect 10378 35506 10434 35562
rect 10502 35506 10558 35562
rect 10626 35506 10682 35562
rect 10750 35506 10806 35562
rect 10874 35506 10930 35562
rect 10998 35506 11054 35562
rect 11122 35506 11178 35562
rect 11246 35506 11302 35562
rect 11370 35506 11426 35562
rect 11494 35506 11550 35562
rect 11618 35506 11674 35562
rect 11742 35506 11798 35562
rect 11866 35506 11922 35562
rect 11990 35506 12046 35562
rect 12114 35506 12170 35562
rect 10254 35382 10310 35438
rect 10378 35382 10434 35438
rect 10502 35382 10558 35438
rect 10626 35382 10682 35438
rect 10750 35382 10806 35438
rect 10874 35382 10930 35438
rect 10998 35382 11054 35438
rect 11122 35382 11178 35438
rect 11246 35382 11302 35438
rect 11370 35382 11426 35438
rect 11494 35382 11550 35438
rect 11618 35382 11674 35438
rect 11742 35382 11798 35438
rect 11866 35382 11922 35438
rect 11990 35382 12046 35438
rect 12114 35382 12170 35438
rect 10254 35258 10310 35314
rect 10378 35258 10434 35314
rect 10502 35258 10558 35314
rect 10626 35258 10682 35314
rect 10750 35258 10806 35314
rect 10874 35258 10930 35314
rect 10998 35258 11054 35314
rect 11122 35258 11178 35314
rect 11246 35258 11302 35314
rect 11370 35258 11426 35314
rect 11494 35258 11550 35314
rect 11618 35258 11674 35314
rect 11742 35258 11798 35314
rect 11866 35258 11922 35314
rect 11990 35258 12046 35314
rect 12114 35258 12170 35314
rect 10254 35134 10310 35190
rect 10378 35134 10434 35190
rect 10502 35134 10558 35190
rect 10626 35134 10682 35190
rect 10750 35134 10806 35190
rect 10874 35134 10930 35190
rect 10998 35134 11054 35190
rect 11122 35134 11178 35190
rect 11246 35134 11302 35190
rect 11370 35134 11426 35190
rect 11494 35134 11550 35190
rect 11618 35134 11674 35190
rect 11742 35134 11798 35190
rect 11866 35134 11922 35190
rect 11990 35134 12046 35190
rect 12114 35134 12170 35190
rect 10254 35010 10310 35066
rect 10378 35010 10434 35066
rect 10502 35010 10558 35066
rect 10626 35010 10682 35066
rect 10750 35010 10806 35066
rect 10874 35010 10930 35066
rect 10998 35010 11054 35066
rect 11122 35010 11178 35066
rect 11246 35010 11302 35066
rect 11370 35010 11426 35066
rect 11494 35010 11550 35066
rect 11618 35010 11674 35066
rect 11742 35010 11798 35066
rect 11866 35010 11922 35066
rect 11990 35010 12046 35066
rect 12114 35010 12170 35066
rect 10254 34886 10310 34942
rect 10378 34886 10434 34942
rect 10502 34886 10558 34942
rect 10626 34886 10682 34942
rect 10750 34886 10806 34942
rect 10874 34886 10930 34942
rect 10998 34886 11054 34942
rect 11122 34886 11178 34942
rect 11246 34886 11302 34942
rect 11370 34886 11426 34942
rect 11494 34886 11550 34942
rect 11618 34886 11674 34942
rect 11742 34886 11798 34942
rect 11866 34886 11922 34942
rect 11990 34886 12046 34942
rect 12114 34886 12170 34942
rect 10254 34762 10310 34818
rect 10378 34762 10434 34818
rect 10502 34762 10558 34818
rect 10626 34762 10682 34818
rect 10750 34762 10806 34818
rect 10874 34762 10930 34818
rect 10998 34762 11054 34818
rect 11122 34762 11178 34818
rect 11246 34762 11302 34818
rect 11370 34762 11426 34818
rect 11494 34762 11550 34818
rect 11618 34762 11674 34818
rect 11742 34762 11798 34818
rect 11866 34762 11922 34818
rect 11990 34762 12046 34818
rect 12114 34762 12170 34818
rect 10254 34638 10310 34694
rect 10378 34638 10434 34694
rect 10502 34638 10558 34694
rect 10626 34638 10682 34694
rect 10750 34638 10806 34694
rect 10874 34638 10930 34694
rect 10998 34638 11054 34694
rect 11122 34638 11178 34694
rect 11246 34638 11302 34694
rect 11370 34638 11426 34694
rect 11494 34638 11550 34694
rect 11618 34638 11674 34694
rect 11742 34638 11798 34694
rect 11866 34638 11922 34694
rect 11990 34638 12046 34694
rect 12114 34638 12170 34694
rect 10254 34514 10310 34570
rect 10378 34514 10434 34570
rect 10502 34514 10558 34570
rect 10626 34514 10682 34570
rect 10750 34514 10806 34570
rect 10874 34514 10930 34570
rect 10998 34514 11054 34570
rect 11122 34514 11178 34570
rect 11246 34514 11302 34570
rect 11370 34514 11426 34570
rect 11494 34514 11550 34570
rect 11618 34514 11674 34570
rect 11742 34514 11798 34570
rect 11866 34514 11922 34570
rect 11990 34514 12046 34570
rect 12114 34514 12170 34570
rect 10254 34390 10310 34446
rect 10378 34390 10434 34446
rect 10502 34390 10558 34446
rect 10626 34390 10682 34446
rect 10750 34390 10806 34446
rect 10874 34390 10930 34446
rect 10998 34390 11054 34446
rect 11122 34390 11178 34446
rect 11246 34390 11302 34446
rect 11370 34390 11426 34446
rect 11494 34390 11550 34446
rect 11618 34390 11674 34446
rect 11742 34390 11798 34446
rect 11866 34390 11922 34446
rect 11990 34390 12046 34446
rect 12114 34390 12170 34446
rect 10254 34266 10310 34322
rect 10378 34266 10434 34322
rect 10502 34266 10558 34322
rect 10626 34266 10682 34322
rect 10750 34266 10806 34322
rect 10874 34266 10930 34322
rect 10998 34266 11054 34322
rect 11122 34266 11178 34322
rect 11246 34266 11302 34322
rect 11370 34266 11426 34322
rect 11494 34266 11550 34322
rect 11618 34266 11674 34322
rect 11742 34266 11798 34322
rect 11866 34266 11922 34322
rect 11990 34266 12046 34322
rect 12114 34266 12170 34322
rect 10254 34142 10310 34198
rect 10378 34142 10434 34198
rect 10502 34142 10558 34198
rect 10626 34142 10682 34198
rect 10750 34142 10806 34198
rect 10874 34142 10930 34198
rect 10998 34142 11054 34198
rect 11122 34142 11178 34198
rect 11246 34142 11302 34198
rect 11370 34142 11426 34198
rect 11494 34142 11550 34198
rect 11618 34142 11674 34198
rect 11742 34142 11798 34198
rect 11866 34142 11922 34198
rect 11990 34142 12046 34198
rect 12114 34142 12170 34198
rect 10254 34018 10310 34074
rect 10378 34018 10434 34074
rect 10502 34018 10558 34074
rect 10626 34018 10682 34074
rect 10750 34018 10806 34074
rect 10874 34018 10930 34074
rect 10998 34018 11054 34074
rect 11122 34018 11178 34074
rect 11246 34018 11302 34074
rect 11370 34018 11426 34074
rect 11494 34018 11550 34074
rect 11618 34018 11674 34074
rect 11742 34018 11798 34074
rect 11866 34018 11922 34074
rect 11990 34018 12046 34074
rect 12114 34018 12170 34074
rect 10254 33894 10310 33950
rect 10378 33894 10434 33950
rect 10502 33894 10558 33950
rect 10626 33894 10682 33950
rect 10750 33894 10806 33950
rect 10874 33894 10930 33950
rect 10998 33894 11054 33950
rect 11122 33894 11178 33950
rect 11246 33894 11302 33950
rect 11370 33894 11426 33950
rect 11494 33894 11550 33950
rect 11618 33894 11674 33950
rect 11742 33894 11798 33950
rect 11866 33894 11922 33950
rect 11990 33894 12046 33950
rect 12114 33894 12170 33950
rect 10254 33770 10310 33826
rect 10378 33770 10434 33826
rect 10502 33770 10558 33826
rect 10626 33770 10682 33826
rect 10750 33770 10806 33826
rect 10874 33770 10930 33826
rect 10998 33770 11054 33826
rect 11122 33770 11178 33826
rect 11246 33770 11302 33826
rect 11370 33770 11426 33826
rect 11494 33770 11550 33826
rect 11618 33770 11674 33826
rect 11742 33770 11798 33826
rect 11866 33770 11922 33826
rect 11990 33770 12046 33826
rect 12114 33770 12170 33826
rect 10254 33646 10310 33702
rect 10378 33646 10434 33702
rect 10502 33646 10558 33702
rect 10626 33646 10682 33702
rect 10750 33646 10806 33702
rect 10874 33646 10930 33702
rect 10998 33646 11054 33702
rect 11122 33646 11178 33702
rect 11246 33646 11302 33702
rect 11370 33646 11426 33702
rect 11494 33646 11550 33702
rect 11618 33646 11674 33702
rect 11742 33646 11798 33702
rect 11866 33646 11922 33702
rect 11990 33646 12046 33702
rect 12114 33646 12170 33702
rect 12871 36498 12927 36554
rect 12995 36498 13051 36554
rect 13119 36498 13175 36554
rect 13243 36498 13299 36554
rect 13367 36498 13423 36554
rect 13491 36498 13547 36554
rect 13615 36498 13671 36554
rect 13739 36498 13795 36554
rect 13863 36498 13919 36554
rect 13987 36498 14043 36554
rect 14111 36498 14167 36554
rect 14235 36498 14291 36554
rect 14359 36498 14415 36554
rect 14483 36498 14539 36554
rect 14607 36498 14663 36554
rect 12871 36374 12927 36430
rect 12995 36374 13051 36430
rect 13119 36374 13175 36430
rect 13243 36374 13299 36430
rect 13367 36374 13423 36430
rect 13491 36374 13547 36430
rect 13615 36374 13671 36430
rect 13739 36374 13795 36430
rect 13863 36374 13919 36430
rect 13987 36374 14043 36430
rect 14111 36374 14167 36430
rect 14235 36374 14291 36430
rect 14359 36374 14415 36430
rect 14483 36374 14539 36430
rect 14607 36374 14663 36430
rect 12871 36250 12927 36306
rect 12995 36250 13051 36306
rect 13119 36250 13175 36306
rect 13243 36250 13299 36306
rect 13367 36250 13423 36306
rect 13491 36250 13547 36306
rect 13615 36250 13671 36306
rect 13739 36250 13795 36306
rect 13863 36250 13919 36306
rect 13987 36250 14043 36306
rect 14111 36250 14167 36306
rect 14235 36250 14291 36306
rect 14359 36250 14415 36306
rect 14483 36250 14539 36306
rect 14607 36250 14663 36306
rect 12871 36126 12927 36182
rect 12995 36126 13051 36182
rect 13119 36126 13175 36182
rect 13243 36126 13299 36182
rect 13367 36126 13423 36182
rect 13491 36126 13547 36182
rect 13615 36126 13671 36182
rect 13739 36126 13795 36182
rect 13863 36126 13919 36182
rect 13987 36126 14043 36182
rect 14111 36126 14167 36182
rect 14235 36126 14291 36182
rect 14359 36126 14415 36182
rect 14483 36126 14539 36182
rect 14607 36126 14663 36182
rect 12871 36002 12927 36058
rect 12995 36002 13051 36058
rect 13119 36002 13175 36058
rect 13243 36002 13299 36058
rect 13367 36002 13423 36058
rect 13491 36002 13547 36058
rect 13615 36002 13671 36058
rect 13739 36002 13795 36058
rect 13863 36002 13919 36058
rect 13987 36002 14043 36058
rect 14111 36002 14167 36058
rect 14235 36002 14291 36058
rect 14359 36002 14415 36058
rect 14483 36002 14539 36058
rect 14607 36002 14663 36058
rect 12871 35878 12927 35934
rect 12995 35878 13051 35934
rect 13119 35878 13175 35934
rect 13243 35878 13299 35934
rect 13367 35878 13423 35934
rect 13491 35878 13547 35934
rect 13615 35878 13671 35934
rect 13739 35878 13795 35934
rect 13863 35878 13919 35934
rect 13987 35878 14043 35934
rect 14111 35878 14167 35934
rect 14235 35878 14291 35934
rect 14359 35878 14415 35934
rect 14483 35878 14539 35934
rect 14607 35878 14663 35934
rect 12871 35754 12927 35810
rect 12995 35754 13051 35810
rect 13119 35754 13175 35810
rect 13243 35754 13299 35810
rect 13367 35754 13423 35810
rect 13491 35754 13547 35810
rect 13615 35754 13671 35810
rect 13739 35754 13795 35810
rect 13863 35754 13919 35810
rect 13987 35754 14043 35810
rect 14111 35754 14167 35810
rect 14235 35754 14291 35810
rect 14359 35754 14415 35810
rect 14483 35754 14539 35810
rect 14607 35754 14663 35810
rect 12871 35630 12927 35686
rect 12995 35630 13051 35686
rect 13119 35630 13175 35686
rect 13243 35630 13299 35686
rect 13367 35630 13423 35686
rect 13491 35630 13547 35686
rect 13615 35630 13671 35686
rect 13739 35630 13795 35686
rect 13863 35630 13919 35686
rect 13987 35630 14043 35686
rect 14111 35630 14167 35686
rect 14235 35630 14291 35686
rect 14359 35630 14415 35686
rect 14483 35630 14539 35686
rect 14607 35630 14663 35686
rect 12871 35506 12927 35562
rect 12995 35506 13051 35562
rect 13119 35506 13175 35562
rect 13243 35506 13299 35562
rect 13367 35506 13423 35562
rect 13491 35506 13547 35562
rect 13615 35506 13671 35562
rect 13739 35506 13795 35562
rect 13863 35506 13919 35562
rect 13987 35506 14043 35562
rect 14111 35506 14167 35562
rect 14235 35506 14291 35562
rect 14359 35506 14415 35562
rect 14483 35506 14539 35562
rect 14607 35506 14663 35562
rect 12871 35382 12927 35438
rect 12995 35382 13051 35438
rect 13119 35382 13175 35438
rect 13243 35382 13299 35438
rect 13367 35382 13423 35438
rect 13491 35382 13547 35438
rect 13615 35382 13671 35438
rect 13739 35382 13795 35438
rect 13863 35382 13919 35438
rect 13987 35382 14043 35438
rect 14111 35382 14167 35438
rect 14235 35382 14291 35438
rect 14359 35382 14415 35438
rect 14483 35382 14539 35438
rect 14607 35382 14663 35438
rect 12871 35258 12927 35314
rect 12995 35258 13051 35314
rect 13119 35258 13175 35314
rect 13243 35258 13299 35314
rect 13367 35258 13423 35314
rect 13491 35258 13547 35314
rect 13615 35258 13671 35314
rect 13739 35258 13795 35314
rect 13863 35258 13919 35314
rect 13987 35258 14043 35314
rect 14111 35258 14167 35314
rect 14235 35258 14291 35314
rect 14359 35258 14415 35314
rect 14483 35258 14539 35314
rect 14607 35258 14663 35314
rect 12871 35134 12927 35190
rect 12995 35134 13051 35190
rect 13119 35134 13175 35190
rect 13243 35134 13299 35190
rect 13367 35134 13423 35190
rect 13491 35134 13547 35190
rect 13615 35134 13671 35190
rect 13739 35134 13795 35190
rect 13863 35134 13919 35190
rect 13987 35134 14043 35190
rect 14111 35134 14167 35190
rect 14235 35134 14291 35190
rect 14359 35134 14415 35190
rect 14483 35134 14539 35190
rect 14607 35134 14663 35190
rect 12871 35010 12927 35066
rect 12995 35010 13051 35066
rect 13119 35010 13175 35066
rect 13243 35010 13299 35066
rect 13367 35010 13423 35066
rect 13491 35010 13547 35066
rect 13615 35010 13671 35066
rect 13739 35010 13795 35066
rect 13863 35010 13919 35066
rect 13987 35010 14043 35066
rect 14111 35010 14167 35066
rect 14235 35010 14291 35066
rect 14359 35010 14415 35066
rect 14483 35010 14539 35066
rect 14607 35010 14663 35066
rect 12871 34886 12927 34942
rect 12995 34886 13051 34942
rect 13119 34886 13175 34942
rect 13243 34886 13299 34942
rect 13367 34886 13423 34942
rect 13491 34886 13547 34942
rect 13615 34886 13671 34942
rect 13739 34886 13795 34942
rect 13863 34886 13919 34942
rect 13987 34886 14043 34942
rect 14111 34886 14167 34942
rect 14235 34886 14291 34942
rect 14359 34886 14415 34942
rect 14483 34886 14539 34942
rect 14607 34886 14663 34942
rect 12871 34762 12927 34818
rect 12995 34762 13051 34818
rect 13119 34762 13175 34818
rect 13243 34762 13299 34818
rect 13367 34762 13423 34818
rect 13491 34762 13547 34818
rect 13615 34762 13671 34818
rect 13739 34762 13795 34818
rect 13863 34762 13919 34818
rect 13987 34762 14043 34818
rect 14111 34762 14167 34818
rect 14235 34762 14291 34818
rect 14359 34762 14415 34818
rect 14483 34762 14539 34818
rect 14607 34762 14663 34818
rect 12871 34638 12927 34694
rect 12995 34638 13051 34694
rect 13119 34638 13175 34694
rect 13243 34638 13299 34694
rect 13367 34638 13423 34694
rect 13491 34638 13547 34694
rect 13615 34638 13671 34694
rect 13739 34638 13795 34694
rect 13863 34638 13919 34694
rect 13987 34638 14043 34694
rect 14111 34638 14167 34694
rect 14235 34638 14291 34694
rect 14359 34638 14415 34694
rect 14483 34638 14539 34694
rect 14607 34638 14663 34694
rect 12871 34514 12927 34570
rect 12995 34514 13051 34570
rect 13119 34514 13175 34570
rect 13243 34514 13299 34570
rect 13367 34514 13423 34570
rect 13491 34514 13547 34570
rect 13615 34514 13671 34570
rect 13739 34514 13795 34570
rect 13863 34514 13919 34570
rect 13987 34514 14043 34570
rect 14111 34514 14167 34570
rect 14235 34514 14291 34570
rect 14359 34514 14415 34570
rect 14483 34514 14539 34570
rect 14607 34514 14663 34570
rect 12871 34390 12927 34446
rect 12995 34390 13051 34446
rect 13119 34390 13175 34446
rect 13243 34390 13299 34446
rect 13367 34390 13423 34446
rect 13491 34390 13547 34446
rect 13615 34390 13671 34446
rect 13739 34390 13795 34446
rect 13863 34390 13919 34446
rect 13987 34390 14043 34446
rect 14111 34390 14167 34446
rect 14235 34390 14291 34446
rect 14359 34390 14415 34446
rect 14483 34390 14539 34446
rect 14607 34390 14663 34446
rect 12871 34266 12927 34322
rect 12995 34266 13051 34322
rect 13119 34266 13175 34322
rect 13243 34266 13299 34322
rect 13367 34266 13423 34322
rect 13491 34266 13547 34322
rect 13615 34266 13671 34322
rect 13739 34266 13795 34322
rect 13863 34266 13919 34322
rect 13987 34266 14043 34322
rect 14111 34266 14167 34322
rect 14235 34266 14291 34322
rect 14359 34266 14415 34322
rect 14483 34266 14539 34322
rect 14607 34266 14663 34322
rect 12871 34142 12927 34198
rect 12995 34142 13051 34198
rect 13119 34142 13175 34198
rect 13243 34142 13299 34198
rect 13367 34142 13423 34198
rect 13491 34142 13547 34198
rect 13615 34142 13671 34198
rect 13739 34142 13795 34198
rect 13863 34142 13919 34198
rect 13987 34142 14043 34198
rect 14111 34142 14167 34198
rect 14235 34142 14291 34198
rect 14359 34142 14415 34198
rect 14483 34142 14539 34198
rect 14607 34142 14663 34198
rect 12871 34018 12927 34074
rect 12995 34018 13051 34074
rect 13119 34018 13175 34074
rect 13243 34018 13299 34074
rect 13367 34018 13423 34074
rect 13491 34018 13547 34074
rect 13615 34018 13671 34074
rect 13739 34018 13795 34074
rect 13863 34018 13919 34074
rect 13987 34018 14043 34074
rect 14111 34018 14167 34074
rect 14235 34018 14291 34074
rect 14359 34018 14415 34074
rect 14483 34018 14539 34074
rect 14607 34018 14663 34074
rect 12871 33894 12927 33950
rect 12995 33894 13051 33950
rect 13119 33894 13175 33950
rect 13243 33894 13299 33950
rect 13367 33894 13423 33950
rect 13491 33894 13547 33950
rect 13615 33894 13671 33950
rect 13739 33894 13795 33950
rect 13863 33894 13919 33950
rect 13987 33894 14043 33950
rect 14111 33894 14167 33950
rect 14235 33894 14291 33950
rect 14359 33894 14415 33950
rect 14483 33894 14539 33950
rect 14607 33894 14663 33950
rect 12871 33770 12927 33826
rect 12995 33770 13051 33826
rect 13119 33770 13175 33826
rect 13243 33770 13299 33826
rect 13367 33770 13423 33826
rect 13491 33770 13547 33826
rect 13615 33770 13671 33826
rect 13739 33770 13795 33826
rect 13863 33770 13919 33826
rect 13987 33770 14043 33826
rect 14111 33770 14167 33826
rect 14235 33770 14291 33826
rect 14359 33770 14415 33826
rect 14483 33770 14539 33826
rect 14607 33770 14663 33826
rect 12871 33646 12927 33702
rect 12995 33646 13051 33702
rect 13119 33646 13175 33702
rect 13243 33646 13299 33702
rect 13367 33646 13423 33702
rect 13491 33646 13547 33702
rect 13615 33646 13671 33702
rect 13739 33646 13795 33702
rect 13863 33646 13919 33702
rect 13987 33646 14043 33702
rect 14111 33646 14167 33702
rect 14235 33646 14291 33702
rect 14359 33646 14415 33702
rect 14483 33646 14539 33702
rect 14607 33646 14663 33702
rect 14902 36584 14958 36586
rect 14902 36532 14904 36584
rect 14904 36532 14956 36584
rect 14956 36532 14958 36584
rect 14902 36476 14958 36532
rect 14902 36424 14904 36476
rect 14904 36424 14956 36476
rect 14956 36424 14958 36476
rect 14902 36368 14958 36424
rect 14902 36316 14904 36368
rect 14904 36316 14956 36368
rect 14956 36316 14958 36368
rect 14902 36260 14958 36316
rect 14902 36208 14904 36260
rect 14904 36208 14956 36260
rect 14956 36208 14958 36260
rect 14902 36152 14958 36208
rect 14902 36100 14904 36152
rect 14904 36100 14956 36152
rect 14956 36100 14958 36152
rect 14902 36044 14958 36100
rect 14902 35992 14904 36044
rect 14904 35992 14956 36044
rect 14956 35992 14958 36044
rect 14902 35936 14958 35992
rect 14902 35884 14904 35936
rect 14904 35884 14956 35936
rect 14956 35884 14958 35936
rect 14902 35828 14958 35884
rect 14902 35776 14904 35828
rect 14904 35776 14956 35828
rect 14956 35776 14958 35828
rect 14902 35720 14958 35776
rect 14902 35668 14904 35720
rect 14904 35668 14956 35720
rect 14956 35668 14958 35720
rect 14902 35612 14958 35668
rect 14902 35560 14904 35612
rect 14904 35560 14956 35612
rect 14956 35560 14958 35612
rect 14902 35504 14958 35560
rect 14902 35452 14904 35504
rect 14904 35452 14956 35504
rect 14956 35452 14958 35504
rect 14902 35396 14958 35452
rect 14902 35344 14904 35396
rect 14904 35344 14956 35396
rect 14956 35344 14958 35396
rect 14902 35288 14958 35344
rect 14902 35236 14904 35288
rect 14904 35236 14956 35288
rect 14956 35236 14958 35288
rect 14902 35180 14958 35236
rect 14902 35128 14904 35180
rect 14904 35128 14956 35180
rect 14956 35128 14958 35180
rect 14902 35072 14958 35128
rect 14902 35020 14904 35072
rect 14904 35020 14956 35072
rect 14956 35020 14958 35072
rect 14902 34964 14958 35020
rect 14902 34912 14904 34964
rect 14904 34912 14956 34964
rect 14956 34912 14958 34964
rect 14902 34856 14958 34912
rect 14902 34804 14904 34856
rect 14904 34804 14956 34856
rect 14956 34804 14958 34856
rect 14902 34748 14958 34804
rect 14902 34696 14904 34748
rect 14904 34696 14956 34748
rect 14956 34696 14958 34748
rect 14902 34640 14958 34696
rect 14902 34588 14904 34640
rect 14904 34588 14956 34640
rect 14956 34588 14958 34640
rect 14902 34532 14958 34588
rect 14902 34480 14904 34532
rect 14904 34480 14956 34532
rect 14956 34480 14958 34532
rect 14902 34424 14958 34480
rect 14902 34372 14904 34424
rect 14904 34372 14956 34424
rect 14956 34372 14958 34424
rect 14902 34316 14958 34372
rect 14902 34264 14904 34316
rect 14904 34264 14956 34316
rect 14956 34264 14958 34316
rect 14902 34208 14958 34264
rect 14902 34156 14904 34208
rect 14904 34156 14956 34208
rect 14956 34156 14958 34208
rect 14902 34100 14958 34156
rect 14902 34048 14904 34100
rect 14904 34048 14956 34100
rect 14956 34048 14958 34100
rect 14902 33992 14958 34048
rect 14902 33940 14904 33992
rect 14904 33940 14956 33992
rect 14956 33940 14958 33992
rect 14902 33884 14958 33940
rect 14902 33832 14904 33884
rect 14904 33832 14956 33884
rect 14956 33832 14958 33884
rect 14902 33776 14958 33832
rect 14902 33724 14904 33776
rect 14904 33724 14956 33776
rect 14956 33724 14958 33776
rect 14902 33668 14958 33724
rect 14902 33616 14904 33668
rect 14904 33616 14956 33668
rect 14956 33616 14958 33668
rect 14902 33614 14958 33616
rect 2491 33298 2547 33354
rect 2615 33298 2671 33354
rect 2491 33174 2547 33230
rect 2615 33174 2671 33230
rect 2491 33050 2547 33106
rect 2615 33050 2671 33106
rect 2491 32926 2547 32982
rect 2615 32926 2671 32982
rect 2491 32802 2547 32858
rect 2615 32802 2671 32858
rect 2491 32678 2547 32734
rect 2615 32678 2671 32734
rect 2491 32554 2547 32610
rect 2615 32554 2671 32610
rect 2491 32430 2547 32486
rect 2615 32430 2671 32486
rect 2491 32306 2547 32362
rect 2615 32306 2671 32362
rect 2491 32182 2547 32238
rect 2615 32182 2671 32238
rect 2491 32058 2547 32114
rect 2615 32058 2671 32114
rect 2491 31934 2547 31990
rect 2615 31934 2671 31990
rect 2491 31810 2547 31866
rect 2615 31810 2671 31866
rect 2491 31686 2547 31742
rect 2615 31686 2671 31742
rect 2491 31562 2547 31618
rect 2615 31562 2671 31618
rect 2491 31438 2547 31494
rect 2615 31438 2671 31494
rect 2491 31314 2547 31370
rect 2615 31314 2671 31370
rect 2491 31190 2547 31246
rect 2615 31190 2671 31246
rect 2491 31066 2547 31122
rect 2615 31066 2671 31122
rect 2491 30942 2547 30998
rect 2615 30942 2671 30998
rect 2491 30818 2547 30874
rect 2615 30818 2671 30874
rect 2491 30694 2547 30750
rect 2615 30694 2671 30750
rect 2491 30570 2547 30626
rect 2615 30570 2671 30626
rect 2491 30446 2547 30502
rect 2615 30446 2671 30502
rect 4861 33298 4917 33354
rect 4985 33298 5041 33354
rect 4861 33174 4917 33230
rect 4985 33174 5041 33230
rect 4861 33050 4917 33106
rect 4985 33050 5041 33106
rect 4861 32926 4917 32982
rect 4985 32926 5041 32982
rect 4861 32802 4917 32858
rect 4985 32802 5041 32858
rect 4861 32678 4917 32734
rect 4985 32678 5041 32734
rect 4861 32554 4917 32610
rect 4985 32554 5041 32610
rect 4861 32430 4917 32486
rect 4985 32430 5041 32486
rect 4861 32306 4917 32362
rect 4985 32306 5041 32362
rect 4861 32182 4917 32238
rect 4985 32182 5041 32238
rect 4861 32058 4917 32114
rect 4985 32058 5041 32114
rect 4861 31934 4917 31990
rect 4985 31934 5041 31990
rect 4861 31810 4917 31866
rect 4985 31810 5041 31866
rect 4861 31686 4917 31742
rect 4985 31686 5041 31742
rect 4861 31562 4917 31618
rect 4985 31562 5041 31618
rect 4861 31438 4917 31494
rect 4985 31438 5041 31494
rect 4861 31314 4917 31370
rect 4985 31314 5041 31370
rect 4861 31190 4917 31246
rect 4985 31190 5041 31246
rect 4861 31066 4917 31122
rect 4985 31066 5041 31122
rect 4861 30942 4917 30998
rect 4985 30942 5041 30998
rect 4861 30818 4917 30874
rect 4985 30818 5041 30874
rect 4861 30694 4917 30750
rect 4985 30694 5041 30750
rect 4861 30570 4917 30626
rect 4985 30570 5041 30626
rect 4861 30446 4917 30502
rect 4985 30446 5041 30502
rect 7275 33298 7331 33354
rect 7399 33298 7455 33354
rect 7523 33298 7579 33354
rect 7647 33298 7703 33354
rect 7275 33174 7331 33230
rect 7399 33174 7455 33230
rect 7523 33174 7579 33230
rect 7647 33174 7703 33230
rect 7275 33050 7331 33106
rect 7399 33050 7455 33106
rect 7523 33050 7579 33106
rect 7647 33050 7703 33106
rect 7275 32926 7331 32982
rect 7399 32926 7455 32982
rect 7523 32926 7579 32982
rect 7647 32926 7703 32982
rect 7275 32802 7331 32858
rect 7399 32802 7455 32858
rect 7523 32802 7579 32858
rect 7647 32802 7703 32858
rect 7275 32678 7331 32734
rect 7399 32678 7455 32734
rect 7523 32678 7579 32734
rect 7647 32678 7703 32734
rect 7275 32554 7331 32610
rect 7399 32554 7455 32610
rect 7523 32554 7579 32610
rect 7647 32554 7703 32610
rect 7275 32430 7331 32486
rect 7399 32430 7455 32486
rect 7523 32430 7579 32486
rect 7647 32430 7703 32486
rect 7275 32306 7331 32362
rect 7399 32306 7455 32362
rect 7523 32306 7579 32362
rect 7647 32306 7703 32362
rect 7275 32182 7331 32238
rect 7399 32182 7455 32238
rect 7523 32182 7579 32238
rect 7647 32182 7703 32238
rect 7275 32058 7331 32114
rect 7399 32058 7455 32114
rect 7523 32058 7579 32114
rect 7647 32058 7703 32114
rect 7275 31934 7331 31990
rect 7399 31934 7455 31990
rect 7523 31934 7579 31990
rect 7647 31934 7703 31990
rect 7275 31810 7331 31866
rect 7399 31810 7455 31866
rect 7523 31810 7579 31866
rect 7647 31810 7703 31866
rect 7275 31686 7331 31742
rect 7399 31686 7455 31742
rect 7523 31686 7579 31742
rect 7647 31686 7703 31742
rect 7275 31562 7331 31618
rect 7399 31562 7455 31618
rect 7523 31562 7579 31618
rect 7647 31562 7703 31618
rect 7275 31438 7331 31494
rect 7399 31438 7455 31494
rect 7523 31438 7579 31494
rect 7647 31438 7703 31494
rect 7275 31314 7331 31370
rect 7399 31314 7455 31370
rect 7523 31314 7579 31370
rect 7647 31314 7703 31370
rect 7275 31190 7331 31246
rect 7399 31190 7455 31246
rect 7523 31190 7579 31246
rect 7647 31190 7703 31246
rect 7275 31066 7331 31122
rect 7399 31066 7455 31122
rect 7523 31066 7579 31122
rect 7647 31066 7703 31122
rect 7275 30942 7331 30998
rect 7399 30942 7455 30998
rect 7523 30942 7579 30998
rect 7647 30942 7703 30998
rect 7275 30818 7331 30874
rect 7399 30818 7455 30874
rect 7523 30818 7579 30874
rect 7647 30818 7703 30874
rect 7275 30694 7331 30750
rect 7399 30694 7455 30750
rect 7523 30694 7579 30750
rect 7647 30694 7703 30750
rect 7275 30570 7331 30626
rect 7399 30570 7455 30626
rect 7523 30570 7579 30626
rect 7647 30570 7703 30626
rect 7275 30446 7331 30502
rect 7399 30446 7455 30502
rect 7523 30446 7579 30502
rect 7647 30446 7703 30502
rect 9937 33298 9993 33354
rect 10061 33298 10117 33354
rect 9937 33174 9993 33230
rect 10061 33174 10117 33230
rect 9937 33050 9993 33106
rect 10061 33050 10117 33106
rect 9937 32926 9993 32982
rect 10061 32926 10117 32982
rect 9937 32802 9993 32858
rect 10061 32802 10117 32858
rect 9937 32678 9993 32734
rect 10061 32678 10117 32734
rect 9937 32554 9993 32610
rect 10061 32554 10117 32610
rect 9937 32430 9993 32486
rect 10061 32430 10117 32486
rect 9937 32306 9993 32362
rect 10061 32306 10117 32362
rect 9937 32182 9993 32238
rect 10061 32182 10117 32238
rect 9937 32058 9993 32114
rect 10061 32058 10117 32114
rect 9937 31934 9993 31990
rect 10061 31934 10117 31990
rect 9937 31810 9993 31866
rect 10061 31810 10117 31866
rect 9937 31686 9993 31742
rect 10061 31686 10117 31742
rect 9937 31562 9993 31618
rect 10061 31562 10117 31618
rect 9937 31438 9993 31494
rect 10061 31438 10117 31494
rect 9937 31314 9993 31370
rect 10061 31314 10117 31370
rect 9937 31190 9993 31246
rect 10061 31190 10117 31246
rect 9937 31066 9993 31122
rect 10061 31066 10117 31122
rect 9937 30942 9993 30998
rect 10061 30942 10117 30998
rect 9937 30818 9993 30874
rect 10061 30818 10117 30874
rect 9937 30694 9993 30750
rect 10061 30694 10117 30750
rect 9937 30570 9993 30626
rect 10061 30570 10117 30626
rect 9937 30446 9993 30502
rect 10061 30446 10117 30502
rect 12307 33298 12363 33354
rect 12431 33298 12487 33354
rect 12307 33174 12363 33230
rect 12431 33174 12487 33230
rect 12307 33050 12363 33106
rect 12431 33050 12487 33106
rect 12307 32926 12363 32982
rect 12431 32926 12487 32982
rect 12307 32802 12363 32858
rect 12431 32802 12487 32858
rect 12307 32678 12363 32734
rect 12431 32678 12487 32734
rect 12307 32554 12363 32610
rect 12431 32554 12487 32610
rect 12307 32430 12363 32486
rect 12431 32430 12487 32486
rect 12307 32306 12363 32362
rect 12431 32306 12487 32362
rect 12307 32182 12363 32238
rect 12431 32182 12487 32238
rect 12307 32058 12363 32114
rect 12431 32058 12487 32114
rect 12307 31934 12363 31990
rect 12431 31934 12487 31990
rect 12307 31810 12363 31866
rect 12431 31810 12487 31866
rect 12307 31686 12363 31742
rect 12431 31686 12487 31742
rect 12307 31562 12363 31618
rect 12431 31562 12487 31618
rect 12307 31438 12363 31494
rect 12431 31438 12487 31494
rect 12307 31314 12363 31370
rect 12431 31314 12487 31370
rect 12307 31190 12363 31246
rect 12431 31190 12487 31246
rect 12307 31066 12363 31122
rect 12431 31066 12487 31122
rect 12307 30942 12363 30998
rect 12431 30942 12487 30998
rect 12307 30818 12363 30874
rect 12431 30818 12487 30874
rect 12307 30694 12363 30750
rect 12431 30694 12487 30750
rect 12307 30570 12363 30626
rect 12431 30570 12487 30626
rect 12307 30446 12363 30502
rect 12431 30446 12487 30502
rect 2491 30092 2547 30148
rect 2615 30092 2671 30148
rect 2491 29968 2547 30024
rect 2615 29968 2671 30024
rect 2491 29844 2547 29900
rect 2615 29844 2671 29900
rect 2491 29720 2547 29776
rect 2615 29720 2671 29776
rect 2491 29596 2547 29652
rect 2615 29596 2671 29652
rect 2491 29472 2547 29528
rect 2615 29472 2671 29528
rect 2491 29348 2547 29404
rect 2615 29348 2671 29404
rect 2491 29224 2547 29280
rect 2615 29224 2671 29280
rect 2491 29100 2547 29156
rect 2615 29100 2671 29156
rect 2491 28976 2547 29032
rect 2615 28976 2671 29032
rect 2491 28852 2547 28908
rect 2615 28852 2671 28908
rect 4861 30092 4917 30148
rect 4985 30092 5041 30148
rect 4861 29968 4917 30024
rect 4985 29968 5041 30024
rect 4861 29844 4917 29900
rect 4985 29844 5041 29900
rect 4861 29720 4917 29776
rect 4985 29720 5041 29776
rect 4861 29596 4917 29652
rect 4985 29596 5041 29652
rect 4861 29472 4917 29528
rect 4985 29472 5041 29528
rect 4861 29348 4917 29404
rect 4985 29348 5041 29404
rect 4861 29224 4917 29280
rect 4985 29224 5041 29280
rect 4861 29100 4917 29156
rect 4985 29100 5041 29156
rect 4861 28976 4917 29032
rect 4985 28976 5041 29032
rect 4861 28852 4917 28908
rect 4985 28852 5041 28908
rect 7275 30092 7331 30148
rect 7399 30092 7455 30148
rect 7523 30092 7579 30148
rect 7647 30092 7703 30148
rect 7275 29968 7331 30024
rect 7399 29968 7455 30024
rect 7523 29968 7579 30024
rect 7647 29968 7703 30024
rect 7275 29844 7331 29900
rect 7399 29844 7455 29900
rect 7523 29844 7579 29900
rect 7647 29844 7703 29900
rect 7275 29720 7331 29776
rect 7399 29720 7455 29776
rect 7523 29720 7579 29776
rect 7647 29720 7703 29776
rect 7275 29596 7331 29652
rect 7399 29596 7455 29652
rect 7523 29596 7579 29652
rect 7647 29596 7703 29652
rect 7275 29472 7331 29528
rect 7399 29472 7455 29528
rect 7523 29472 7579 29528
rect 7647 29472 7703 29528
rect 7275 29348 7331 29404
rect 7399 29348 7455 29404
rect 7523 29348 7579 29404
rect 7647 29348 7703 29404
rect 7275 29224 7331 29280
rect 7399 29224 7455 29280
rect 7523 29224 7579 29280
rect 7647 29224 7703 29280
rect 7275 29100 7331 29156
rect 7399 29100 7455 29156
rect 7523 29100 7579 29156
rect 7647 29100 7703 29156
rect 7275 28976 7331 29032
rect 7399 28976 7455 29032
rect 7523 28976 7579 29032
rect 7647 28976 7703 29032
rect 7275 28852 7331 28908
rect 7399 28852 7455 28908
rect 7523 28852 7579 28908
rect 7647 28852 7703 28908
rect 9937 30092 9993 30148
rect 10061 30092 10117 30148
rect 9937 29968 9993 30024
rect 10061 29968 10117 30024
rect 9937 29844 9993 29900
rect 10061 29844 10117 29900
rect 9937 29720 9993 29776
rect 10061 29720 10117 29776
rect 9937 29596 9993 29652
rect 10061 29596 10117 29652
rect 9937 29472 9993 29528
rect 10061 29472 10117 29528
rect 9937 29348 9993 29404
rect 10061 29348 10117 29404
rect 9937 29224 9993 29280
rect 10061 29224 10117 29280
rect 9937 29100 9993 29156
rect 10061 29100 10117 29156
rect 9937 28976 9993 29032
rect 10061 28976 10117 29032
rect 9937 28852 9993 28908
rect 10061 28852 10117 28908
rect 12307 30092 12363 30148
rect 12431 30092 12487 30148
rect 12307 29968 12363 30024
rect 12431 29968 12487 30024
rect 12307 29844 12363 29900
rect 12431 29844 12487 29900
rect 12307 29720 12363 29776
rect 12431 29720 12487 29776
rect 12307 29596 12363 29652
rect 12431 29596 12487 29652
rect 12307 29472 12363 29528
rect 12431 29472 12487 29528
rect 12307 29348 12363 29404
rect 12431 29348 12487 29404
rect 12307 29224 12363 29280
rect 12431 29224 12487 29280
rect 12307 29100 12363 29156
rect 12431 29100 12487 29156
rect 12307 28976 12363 29032
rect 12431 28976 12487 29032
rect 12307 28852 12363 28908
rect 12431 28852 12487 28908
rect 20 28574 76 28576
rect 20 28522 22 28574
rect 22 28522 74 28574
rect 74 28522 76 28574
rect 20 28466 76 28522
rect 20 28414 22 28466
rect 22 28414 74 28466
rect 74 28414 76 28466
rect 20 28358 76 28414
rect 20 28306 22 28358
rect 22 28306 74 28358
rect 74 28306 76 28358
rect 20 28250 76 28306
rect 20 28198 22 28250
rect 22 28198 74 28250
rect 74 28198 76 28250
rect 20 28142 76 28198
rect 20 28090 22 28142
rect 22 28090 74 28142
rect 74 28090 76 28142
rect 20 28034 76 28090
rect 20 27982 22 28034
rect 22 27982 74 28034
rect 74 27982 76 28034
rect 20 27926 76 27982
rect 20 27874 22 27926
rect 22 27874 74 27926
rect 74 27874 76 27926
rect 20 27818 76 27874
rect 20 27766 22 27818
rect 22 27766 74 27818
rect 74 27766 76 27818
rect 20 27710 76 27766
rect 20 27658 22 27710
rect 22 27658 74 27710
rect 74 27658 76 27710
rect 20 27602 76 27658
rect 20 27550 22 27602
rect 22 27550 74 27602
rect 74 27550 76 27602
rect 20 27494 76 27550
rect 20 27442 22 27494
rect 22 27442 74 27494
rect 74 27442 76 27494
rect 20 27386 76 27442
rect 20 27334 22 27386
rect 22 27334 74 27386
rect 74 27334 76 27386
rect 20 27278 76 27334
rect 20 27226 22 27278
rect 22 27226 74 27278
rect 74 27226 76 27278
rect 20 27224 76 27226
rect 315 28492 371 28548
rect 439 28492 495 28548
rect 563 28492 619 28548
rect 687 28492 743 28548
rect 811 28492 867 28548
rect 935 28492 991 28548
rect 1059 28492 1115 28548
rect 1183 28492 1239 28548
rect 1307 28492 1363 28548
rect 1431 28492 1487 28548
rect 1555 28492 1611 28548
rect 1679 28492 1735 28548
rect 1803 28492 1859 28548
rect 1927 28492 1983 28548
rect 2051 28492 2107 28548
rect 315 28368 371 28424
rect 439 28368 495 28424
rect 563 28368 619 28424
rect 687 28368 743 28424
rect 811 28368 867 28424
rect 935 28368 991 28424
rect 1059 28368 1115 28424
rect 1183 28368 1239 28424
rect 1307 28368 1363 28424
rect 1431 28368 1487 28424
rect 1555 28368 1611 28424
rect 1679 28368 1735 28424
rect 1803 28368 1859 28424
rect 1927 28368 1983 28424
rect 2051 28368 2107 28424
rect 315 28244 371 28300
rect 439 28244 495 28300
rect 563 28244 619 28300
rect 687 28244 743 28300
rect 811 28244 867 28300
rect 935 28244 991 28300
rect 1059 28244 1115 28300
rect 1183 28244 1239 28300
rect 1307 28244 1363 28300
rect 1431 28244 1487 28300
rect 1555 28244 1611 28300
rect 1679 28244 1735 28300
rect 1803 28244 1859 28300
rect 1927 28244 1983 28300
rect 2051 28244 2107 28300
rect 315 28120 371 28176
rect 439 28120 495 28176
rect 563 28120 619 28176
rect 687 28120 743 28176
rect 811 28120 867 28176
rect 935 28120 991 28176
rect 1059 28120 1115 28176
rect 1183 28120 1239 28176
rect 1307 28120 1363 28176
rect 1431 28120 1487 28176
rect 1555 28120 1611 28176
rect 1679 28120 1735 28176
rect 1803 28120 1859 28176
rect 1927 28120 1983 28176
rect 2051 28120 2107 28176
rect 315 27996 371 28052
rect 439 27996 495 28052
rect 563 27996 619 28052
rect 687 27996 743 28052
rect 811 27996 867 28052
rect 935 27996 991 28052
rect 1059 27996 1115 28052
rect 1183 27996 1239 28052
rect 1307 27996 1363 28052
rect 1431 27996 1487 28052
rect 1555 27996 1611 28052
rect 1679 27996 1735 28052
rect 1803 27996 1859 28052
rect 1927 27996 1983 28052
rect 2051 27996 2107 28052
rect 315 27872 371 27928
rect 439 27872 495 27928
rect 563 27872 619 27928
rect 687 27872 743 27928
rect 811 27872 867 27928
rect 935 27872 991 27928
rect 1059 27872 1115 27928
rect 1183 27872 1239 27928
rect 1307 27872 1363 27928
rect 1431 27872 1487 27928
rect 1555 27872 1611 27928
rect 1679 27872 1735 27928
rect 1803 27872 1859 27928
rect 1927 27872 1983 27928
rect 2051 27872 2107 27928
rect 315 27748 371 27804
rect 439 27748 495 27804
rect 563 27748 619 27804
rect 687 27748 743 27804
rect 811 27748 867 27804
rect 935 27748 991 27804
rect 1059 27748 1115 27804
rect 1183 27748 1239 27804
rect 1307 27748 1363 27804
rect 1431 27748 1487 27804
rect 1555 27748 1611 27804
rect 1679 27748 1735 27804
rect 1803 27748 1859 27804
rect 1927 27748 1983 27804
rect 2051 27748 2107 27804
rect 315 27624 371 27680
rect 439 27624 495 27680
rect 563 27624 619 27680
rect 687 27624 743 27680
rect 811 27624 867 27680
rect 935 27624 991 27680
rect 1059 27624 1115 27680
rect 1183 27624 1239 27680
rect 1307 27624 1363 27680
rect 1431 27624 1487 27680
rect 1555 27624 1611 27680
rect 1679 27624 1735 27680
rect 1803 27624 1859 27680
rect 1927 27624 1983 27680
rect 2051 27624 2107 27680
rect 315 27500 371 27556
rect 439 27500 495 27556
rect 563 27500 619 27556
rect 687 27500 743 27556
rect 811 27500 867 27556
rect 935 27500 991 27556
rect 1059 27500 1115 27556
rect 1183 27500 1239 27556
rect 1307 27500 1363 27556
rect 1431 27500 1487 27556
rect 1555 27500 1611 27556
rect 1679 27500 1735 27556
rect 1803 27500 1859 27556
rect 1927 27500 1983 27556
rect 2051 27500 2107 27556
rect 315 27376 371 27432
rect 439 27376 495 27432
rect 563 27376 619 27432
rect 687 27376 743 27432
rect 811 27376 867 27432
rect 935 27376 991 27432
rect 1059 27376 1115 27432
rect 1183 27376 1239 27432
rect 1307 27376 1363 27432
rect 1431 27376 1487 27432
rect 1555 27376 1611 27432
rect 1679 27376 1735 27432
rect 1803 27376 1859 27432
rect 1927 27376 1983 27432
rect 2051 27376 2107 27432
rect 315 27252 371 27308
rect 439 27252 495 27308
rect 563 27252 619 27308
rect 687 27252 743 27308
rect 811 27252 867 27308
rect 935 27252 991 27308
rect 1059 27252 1115 27308
rect 1183 27252 1239 27308
rect 1307 27252 1363 27308
rect 1431 27252 1487 27308
rect 1555 27252 1611 27308
rect 1679 27252 1735 27308
rect 1803 27252 1859 27308
rect 1927 27252 1983 27308
rect 2051 27252 2107 27308
rect 2808 28492 2864 28548
rect 2932 28492 2988 28548
rect 3056 28492 3112 28548
rect 3180 28492 3236 28548
rect 3304 28492 3360 28548
rect 3428 28492 3484 28548
rect 3552 28492 3608 28548
rect 3676 28492 3732 28548
rect 3800 28492 3856 28548
rect 3924 28492 3980 28548
rect 4048 28492 4104 28548
rect 4172 28492 4228 28548
rect 4296 28492 4352 28548
rect 4420 28492 4476 28548
rect 4544 28492 4600 28548
rect 4668 28492 4724 28548
rect 2808 28368 2864 28424
rect 2932 28368 2988 28424
rect 3056 28368 3112 28424
rect 3180 28368 3236 28424
rect 3304 28368 3360 28424
rect 3428 28368 3484 28424
rect 3552 28368 3608 28424
rect 3676 28368 3732 28424
rect 3800 28368 3856 28424
rect 3924 28368 3980 28424
rect 4048 28368 4104 28424
rect 4172 28368 4228 28424
rect 4296 28368 4352 28424
rect 4420 28368 4476 28424
rect 4544 28368 4600 28424
rect 4668 28368 4724 28424
rect 2808 28244 2864 28300
rect 2932 28244 2988 28300
rect 3056 28244 3112 28300
rect 3180 28244 3236 28300
rect 3304 28244 3360 28300
rect 3428 28244 3484 28300
rect 3552 28244 3608 28300
rect 3676 28244 3732 28300
rect 3800 28244 3856 28300
rect 3924 28244 3980 28300
rect 4048 28244 4104 28300
rect 4172 28244 4228 28300
rect 4296 28244 4352 28300
rect 4420 28244 4476 28300
rect 4544 28244 4600 28300
rect 4668 28244 4724 28300
rect 2808 28120 2864 28176
rect 2932 28120 2988 28176
rect 3056 28120 3112 28176
rect 3180 28120 3236 28176
rect 3304 28120 3360 28176
rect 3428 28120 3484 28176
rect 3552 28120 3608 28176
rect 3676 28120 3732 28176
rect 3800 28120 3856 28176
rect 3924 28120 3980 28176
rect 4048 28120 4104 28176
rect 4172 28120 4228 28176
rect 4296 28120 4352 28176
rect 4420 28120 4476 28176
rect 4544 28120 4600 28176
rect 4668 28120 4724 28176
rect 2808 27996 2864 28052
rect 2932 27996 2988 28052
rect 3056 27996 3112 28052
rect 3180 27996 3236 28052
rect 3304 27996 3360 28052
rect 3428 27996 3484 28052
rect 3552 27996 3608 28052
rect 3676 27996 3732 28052
rect 3800 27996 3856 28052
rect 3924 27996 3980 28052
rect 4048 27996 4104 28052
rect 4172 27996 4228 28052
rect 4296 27996 4352 28052
rect 4420 27996 4476 28052
rect 4544 27996 4600 28052
rect 4668 27996 4724 28052
rect 2808 27872 2864 27928
rect 2932 27872 2988 27928
rect 3056 27872 3112 27928
rect 3180 27872 3236 27928
rect 3304 27872 3360 27928
rect 3428 27872 3484 27928
rect 3552 27872 3608 27928
rect 3676 27872 3732 27928
rect 3800 27872 3856 27928
rect 3924 27872 3980 27928
rect 4048 27872 4104 27928
rect 4172 27872 4228 27928
rect 4296 27872 4352 27928
rect 4420 27872 4476 27928
rect 4544 27872 4600 27928
rect 4668 27872 4724 27928
rect 2808 27748 2864 27804
rect 2932 27748 2988 27804
rect 3056 27748 3112 27804
rect 3180 27748 3236 27804
rect 3304 27748 3360 27804
rect 3428 27748 3484 27804
rect 3552 27748 3608 27804
rect 3676 27748 3732 27804
rect 3800 27748 3856 27804
rect 3924 27748 3980 27804
rect 4048 27748 4104 27804
rect 4172 27748 4228 27804
rect 4296 27748 4352 27804
rect 4420 27748 4476 27804
rect 4544 27748 4600 27804
rect 4668 27748 4724 27804
rect 2808 27624 2864 27680
rect 2932 27624 2988 27680
rect 3056 27624 3112 27680
rect 3180 27624 3236 27680
rect 3304 27624 3360 27680
rect 3428 27624 3484 27680
rect 3552 27624 3608 27680
rect 3676 27624 3732 27680
rect 3800 27624 3856 27680
rect 3924 27624 3980 27680
rect 4048 27624 4104 27680
rect 4172 27624 4228 27680
rect 4296 27624 4352 27680
rect 4420 27624 4476 27680
rect 4544 27624 4600 27680
rect 4668 27624 4724 27680
rect 2808 27500 2864 27556
rect 2932 27500 2988 27556
rect 3056 27500 3112 27556
rect 3180 27500 3236 27556
rect 3304 27500 3360 27556
rect 3428 27500 3484 27556
rect 3552 27500 3608 27556
rect 3676 27500 3732 27556
rect 3800 27500 3856 27556
rect 3924 27500 3980 27556
rect 4048 27500 4104 27556
rect 4172 27500 4228 27556
rect 4296 27500 4352 27556
rect 4420 27500 4476 27556
rect 4544 27500 4600 27556
rect 4668 27500 4724 27556
rect 2808 27376 2864 27432
rect 2932 27376 2988 27432
rect 3056 27376 3112 27432
rect 3180 27376 3236 27432
rect 3304 27376 3360 27432
rect 3428 27376 3484 27432
rect 3552 27376 3608 27432
rect 3676 27376 3732 27432
rect 3800 27376 3856 27432
rect 3924 27376 3980 27432
rect 4048 27376 4104 27432
rect 4172 27376 4228 27432
rect 4296 27376 4352 27432
rect 4420 27376 4476 27432
rect 4544 27376 4600 27432
rect 4668 27376 4724 27432
rect 2808 27252 2864 27308
rect 2932 27252 2988 27308
rect 3056 27252 3112 27308
rect 3180 27252 3236 27308
rect 3304 27252 3360 27308
rect 3428 27252 3484 27308
rect 3552 27252 3608 27308
rect 3676 27252 3732 27308
rect 3800 27252 3856 27308
rect 3924 27252 3980 27308
rect 4048 27252 4104 27308
rect 4172 27252 4228 27308
rect 4296 27252 4352 27308
rect 4420 27252 4476 27308
rect 4544 27252 4600 27308
rect 4668 27252 4724 27308
rect 5178 28492 5234 28548
rect 5302 28492 5358 28548
rect 5426 28492 5482 28548
rect 5550 28492 5606 28548
rect 5674 28492 5730 28548
rect 5798 28492 5854 28548
rect 5922 28492 5978 28548
rect 6046 28492 6102 28548
rect 6170 28492 6226 28548
rect 6294 28492 6350 28548
rect 6418 28492 6474 28548
rect 6542 28492 6598 28548
rect 6666 28492 6722 28548
rect 6790 28492 6846 28548
rect 6914 28492 6970 28548
rect 7038 28492 7094 28548
rect 5178 28368 5234 28424
rect 5302 28368 5358 28424
rect 5426 28368 5482 28424
rect 5550 28368 5606 28424
rect 5674 28368 5730 28424
rect 5798 28368 5854 28424
rect 5922 28368 5978 28424
rect 6046 28368 6102 28424
rect 6170 28368 6226 28424
rect 6294 28368 6350 28424
rect 6418 28368 6474 28424
rect 6542 28368 6598 28424
rect 6666 28368 6722 28424
rect 6790 28368 6846 28424
rect 6914 28368 6970 28424
rect 7038 28368 7094 28424
rect 5178 28244 5234 28300
rect 5302 28244 5358 28300
rect 5426 28244 5482 28300
rect 5550 28244 5606 28300
rect 5674 28244 5730 28300
rect 5798 28244 5854 28300
rect 5922 28244 5978 28300
rect 6046 28244 6102 28300
rect 6170 28244 6226 28300
rect 6294 28244 6350 28300
rect 6418 28244 6474 28300
rect 6542 28244 6598 28300
rect 6666 28244 6722 28300
rect 6790 28244 6846 28300
rect 6914 28244 6970 28300
rect 7038 28244 7094 28300
rect 5178 28120 5234 28176
rect 5302 28120 5358 28176
rect 5426 28120 5482 28176
rect 5550 28120 5606 28176
rect 5674 28120 5730 28176
rect 5798 28120 5854 28176
rect 5922 28120 5978 28176
rect 6046 28120 6102 28176
rect 6170 28120 6226 28176
rect 6294 28120 6350 28176
rect 6418 28120 6474 28176
rect 6542 28120 6598 28176
rect 6666 28120 6722 28176
rect 6790 28120 6846 28176
rect 6914 28120 6970 28176
rect 7038 28120 7094 28176
rect 5178 27996 5234 28052
rect 5302 27996 5358 28052
rect 5426 27996 5482 28052
rect 5550 27996 5606 28052
rect 5674 27996 5730 28052
rect 5798 27996 5854 28052
rect 5922 27996 5978 28052
rect 6046 27996 6102 28052
rect 6170 27996 6226 28052
rect 6294 27996 6350 28052
rect 6418 27996 6474 28052
rect 6542 27996 6598 28052
rect 6666 27996 6722 28052
rect 6790 27996 6846 28052
rect 6914 27996 6970 28052
rect 7038 27996 7094 28052
rect 5178 27872 5234 27928
rect 5302 27872 5358 27928
rect 5426 27872 5482 27928
rect 5550 27872 5606 27928
rect 5674 27872 5730 27928
rect 5798 27872 5854 27928
rect 5922 27872 5978 27928
rect 6046 27872 6102 27928
rect 6170 27872 6226 27928
rect 6294 27872 6350 27928
rect 6418 27872 6474 27928
rect 6542 27872 6598 27928
rect 6666 27872 6722 27928
rect 6790 27872 6846 27928
rect 6914 27872 6970 27928
rect 7038 27872 7094 27928
rect 5178 27748 5234 27804
rect 5302 27748 5358 27804
rect 5426 27748 5482 27804
rect 5550 27748 5606 27804
rect 5674 27748 5730 27804
rect 5798 27748 5854 27804
rect 5922 27748 5978 27804
rect 6046 27748 6102 27804
rect 6170 27748 6226 27804
rect 6294 27748 6350 27804
rect 6418 27748 6474 27804
rect 6542 27748 6598 27804
rect 6666 27748 6722 27804
rect 6790 27748 6846 27804
rect 6914 27748 6970 27804
rect 7038 27748 7094 27804
rect 5178 27624 5234 27680
rect 5302 27624 5358 27680
rect 5426 27624 5482 27680
rect 5550 27624 5606 27680
rect 5674 27624 5730 27680
rect 5798 27624 5854 27680
rect 5922 27624 5978 27680
rect 6046 27624 6102 27680
rect 6170 27624 6226 27680
rect 6294 27624 6350 27680
rect 6418 27624 6474 27680
rect 6542 27624 6598 27680
rect 6666 27624 6722 27680
rect 6790 27624 6846 27680
rect 6914 27624 6970 27680
rect 7038 27624 7094 27680
rect 5178 27500 5234 27556
rect 5302 27500 5358 27556
rect 5426 27500 5482 27556
rect 5550 27500 5606 27556
rect 5674 27500 5730 27556
rect 5798 27500 5854 27556
rect 5922 27500 5978 27556
rect 6046 27500 6102 27556
rect 6170 27500 6226 27556
rect 6294 27500 6350 27556
rect 6418 27500 6474 27556
rect 6542 27500 6598 27556
rect 6666 27500 6722 27556
rect 6790 27500 6846 27556
rect 6914 27500 6970 27556
rect 7038 27500 7094 27556
rect 5178 27376 5234 27432
rect 5302 27376 5358 27432
rect 5426 27376 5482 27432
rect 5550 27376 5606 27432
rect 5674 27376 5730 27432
rect 5798 27376 5854 27432
rect 5922 27376 5978 27432
rect 6046 27376 6102 27432
rect 6170 27376 6226 27432
rect 6294 27376 6350 27432
rect 6418 27376 6474 27432
rect 6542 27376 6598 27432
rect 6666 27376 6722 27432
rect 6790 27376 6846 27432
rect 6914 27376 6970 27432
rect 7038 27376 7094 27432
rect 5178 27252 5234 27308
rect 5302 27252 5358 27308
rect 5426 27252 5482 27308
rect 5550 27252 5606 27308
rect 5674 27252 5730 27308
rect 5798 27252 5854 27308
rect 5922 27252 5978 27308
rect 6046 27252 6102 27308
rect 6170 27252 6226 27308
rect 6294 27252 6350 27308
rect 6418 27252 6474 27308
rect 6542 27252 6598 27308
rect 6666 27252 6722 27308
rect 6790 27252 6846 27308
rect 6914 27252 6970 27308
rect 7038 27252 7094 27308
rect 7884 28492 7940 28548
rect 8008 28492 8064 28548
rect 8132 28492 8188 28548
rect 8256 28492 8312 28548
rect 8380 28492 8436 28548
rect 8504 28492 8560 28548
rect 8628 28492 8684 28548
rect 8752 28492 8808 28548
rect 8876 28492 8932 28548
rect 9000 28492 9056 28548
rect 9124 28492 9180 28548
rect 9248 28492 9304 28548
rect 9372 28492 9428 28548
rect 9496 28492 9552 28548
rect 9620 28492 9676 28548
rect 9744 28492 9800 28548
rect 7884 28368 7940 28424
rect 8008 28368 8064 28424
rect 8132 28368 8188 28424
rect 8256 28368 8312 28424
rect 8380 28368 8436 28424
rect 8504 28368 8560 28424
rect 8628 28368 8684 28424
rect 8752 28368 8808 28424
rect 8876 28368 8932 28424
rect 9000 28368 9056 28424
rect 9124 28368 9180 28424
rect 9248 28368 9304 28424
rect 9372 28368 9428 28424
rect 9496 28368 9552 28424
rect 9620 28368 9676 28424
rect 9744 28368 9800 28424
rect 7884 28244 7940 28300
rect 8008 28244 8064 28300
rect 8132 28244 8188 28300
rect 8256 28244 8312 28300
rect 8380 28244 8436 28300
rect 8504 28244 8560 28300
rect 8628 28244 8684 28300
rect 8752 28244 8808 28300
rect 8876 28244 8932 28300
rect 9000 28244 9056 28300
rect 9124 28244 9180 28300
rect 9248 28244 9304 28300
rect 9372 28244 9428 28300
rect 9496 28244 9552 28300
rect 9620 28244 9676 28300
rect 9744 28244 9800 28300
rect 7884 28120 7940 28176
rect 8008 28120 8064 28176
rect 8132 28120 8188 28176
rect 8256 28120 8312 28176
rect 8380 28120 8436 28176
rect 8504 28120 8560 28176
rect 8628 28120 8684 28176
rect 8752 28120 8808 28176
rect 8876 28120 8932 28176
rect 9000 28120 9056 28176
rect 9124 28120 9180 28176
rect 9248 28120 9304 28176
rect 9372 28120 9428 28176
rect 9496 28120 9552 28176
rect 9620 28120 9676 28176
rect 9744 28120 9800 28176
rect 7884 27996 7940 28052
rect 8008 27996 8064 28052
rect 8132 27996 8188 28052
rect 8256 27996 8312 28052
rect 8380 27996 8436 28052
rect 8504 27996 8560 28052
rect 8628 27996 8684 28052
rect 8752 27996 8808 28052
rect 8876 27996 8932 28052
rect 9000 27996 9056 28052
rect 9124 27996 9180 28052
rect 9248 27996 9304 28052
rect 9372 27996 9428 28052
rect 9496 27996 9552 28052
rect 9620 27996 9676 28052
rect 9744 27996 9800 28052
rect 7884 27872 7940 27928
rect 8008 27872 8064 27928
rect 8132 27872 8188 27928
rect 8256 27872 8312 27928
rect 8380 27872 8436 27928
rect 8504 27872 8560 27928
rect 8628 27872 8684 27928
rect 8752 27872 8808 27928
rect 8876 27872 8932 27928
rect 9000 27872 9056 27928
rect 9124 27872 9180 27928
rect 9248 27872 9304 27928
rect 9372 27872 9428 27928
rect 9496 27872 9552 27928
rect 9620 27872 9676 27928
rect 9744 27872 9800 27928
rect 7884 27748 7940 27804
rect 8008 27748 8064 27804
rect 8132 27748 8188 27804
rect 8256 27748 8312 27804
rect 8380 27748 8436 27804
rect 8504 27748 8560 27804
rect 8628 27748 8684 27804
rect 8752 27748 8808 27804
rect 8876 27748 8932 27804
rect 9000 27748 9056 27804
rect 9124 27748 9180 27804
rect 9248 27748 9304 27804
rect 9372 27748 9428 27804
rect 9496 27748 9552 27804
rect 9620 27748 9676 27804
rect 9744 27748 9800 27804
rect 7884 27624 7940 27680
rect 8008 27624 8064 27680
rect 8132 27624 8188 27680
rect 8256 27624 8312 27680
rect 8380 27624 8436 27680
rect 8504 27624 8560 27680
rect 8628 27624 8684 27680
rect 8752 27624 8808 27680
rect 8876 27624 8932 27680
rect 9000 27624 9056 27680
rect 9124 27624 9180 27680
rect 9248 27624 9304 27680
rect 9372 27624 9428 27680
rect 9496 27624 9552 27680
rect 9620 27624 9676 27680
rect 9744 27624 9800 27680
rect 7884 27500 7940 27556
rect 8008 27500 8064 27556
rect 8132 27500 8188 27556
rect 8256 27500 8312 27556
rect 8380 27500 8436 27556
rect 8504 27500 8560 27556
rect 8628 27500 8684 27556
rect 8752 27500 8808 27556
rect 8876 27500 8932 27556
rect 9000 27500 9056 27556
rect 9124 27500 9180 27556
rect 9248 27500 9304 27556
rect 9372 27500 9428 27556
rect 9496 27500 9552 27556
rect 9620 27500 9676 27556
rect 9744 27500 9800 27556
rect 7884 27376 7940 27432
rect 8008 27376 8064 27432
rect 8132 27376 8188 27432
rect 8256 27376 8312 27432
rect 8380 27376 8436 27432
rect 8504 27376 8560 27432
rect 8628 27376 8684 27432
rect 8752 27376 8808 27432
rect 8876 27376 8932 27432
rect 9000 27376 9056 27432
rect 9124 27376 9180 27432
rect 9248 27376 9304 27432
rect 9372 27376 9428 27432
rect 9496 27376 9552 27432
rect 9620 27376 9676 27432
rect 9744 27376 9800 27432
rect 7884 27252 7940 27308
rect 8008 27252 8064 27308
rect 8132 27252 8188 27308
rect 8256 27252 8312 27308
rect 8380 27252 8436 27308
rect 8504 27252 8560 27308
rect 8628 27252 8684 27308
rect 8752 27252 8808 27308
rect 8876 27252 8932 27308
rect 9000 27252 9056 27308
rect 9124 27252 9180 27308
rect 9248 27252 9304 27308
rect 9372 27252 9428 27308
rect 9496 27252 9552 27308
rect 9620 27252 9676 27308
rect 9744 27252 9800 27308
rect 10254 28492 10310 28548
rect 10378 28492 10434 28548
rect 10502 28492 10558 28548
rect 10626 28492 10682 28548
rect 10750 28492 10806 28548
rect 10874 28492 10930 28548
rect 10998 28492 11054 28548
rect 11122 28492 11178 28548
rect 11246 28492 11302 28548
rect 11370 28492 11426 28548
rect 11494 28492 11550 28548
rect 11618 28492 11674 28548
rect 11742 28492 11798 28548
rect 11866 28492 11922 28548
rect 11990 28492 12046 28548
rect 12114 28492 12170 28548
rect 10254 28368 10310 28424
rect 10378 28368 10434 28424
rect 10502 28368 10558 28424
rect 10626 28368 10682 28424
rect 10750 28368 10806 28424
rect 10874 28368 10930 28424
rect 10998 28368 11054 28424
rect 11122 28368 11178 28424
rect 11246 28368 11302 28424
rect 11370 28368 11426 28424
rect 11494 28368 11550 28424
rect 11618 28368 11674 28424
rect 11742 28368 11798 28424
rect 11866 28368 11922 28424
rect 11990 28368 12046 28424
rect 12114 28368 12170 28424
rect 10254 28244 10310 28300
rect 10378 28244 10434 28300
rect 10502 28244 10558 28300
rect 10626 28244 10682 28300
rect 10750 28244 10806 28300
rect 10874 28244 10930 28300
rect 10998 28244 11054 28300
rect 11122 28244 11178 28300
rect 11246 28244 11302 28300
rect 11370 28244 11426 28300
rect 11494 28244 11550 28300
rect 11618 28244 11674 28300
rect 11742 28244 11798 28300
rect 11866 28244 11922 28300
rect 11990 28244 12046 28300
rect 12114 28244 12170 28300
rect 10254 28120 10310 28176
rect 10378 28120 10434 28176
rect 10502 28120 10558 28176
rect 10626 28120 10682 28176
rect 10750 28120 10806 28176
rect 10874 28120 10930 28176
rect 10998 28120 11054 28176
rect 11122 28120 11178 28176
rect 11246 28120 11302 28176
rect 11370 28120 11426 28176
rect 11494 28120 11550 28176
rect 11618 28120 11674 28176
rect 11742 28120 11798 28176
rect 11866 28120 11922 28176
rect 11990 28120 12046 28176
rect 12114 28120 12170 28176
rect 10254 27996 10310 28052
rect 10378 27996 10434 28052
rect 10502 27996 10558 28052
rect 10626 27996 10682 28052
rect 10750 27996 10806 28052
rect 10874 27996 10930 28052
rect 10998 27996 11054 28052
rect 11122 27996 11178 28052
rect 11246 27996 11302 28052
rect 11370 27996 11426 28052
rect 11494 27996 11550 28052
rect 11618 27996 11674 28052
rect 11742 27996 11798 28052
rect 11866 27996 11922 28052
rect 11990 27996 12046 28052
rect 12114 27996 12170 28052
rect 10254 27872 10310 27928
rect 10378 27872 10434 27928
rect 10502 27872 10558 27928
rect 10626 27872 10682 27928
rect 10750 27872 10806 27928
rect 10874 27872 10930 27928
rect 10998 27872 11054 27928
rect 11122 27872 11178 27928
rect 11246 27872 11302 27928
rect 11370 27872 11426 27928
rect 11494 27872 11550 27928
rect 11618 27872 11674 27928
rect 11742 27872 11798 27928
rect 11866 27872 11922 27928
rect 11990 27872 12046 27928
rect 12114 27872 12170 27928
rect 10254 27748 10310 27804
rect 10378 27748 10434 27804
rect 10502 27748 10558 27804
rect 10626 27748 10682 27804
rect 10750 27748 10806 27804
rect 10874 27748 10930 27804
rect 10998 27748 11054 27804
rect 11122 27748 11178 27804
rect 11246 27748 11302 27804
rect 11370 27748 11426 27804
rect 11494 27748 11550 27804
rect 11618 27748 11674 27804
rect 11742 27748 11798 27804
rect 11866 27748 11922 27804
rect 11990 27748 12046 27804
rect 12114 27748 12170 27804
rect 10254 27624 10310 27680
rect 10378 27624 10434 27680
rect 10502 27624 10558 27680
rect 10626 27624 10682 27680
rect 10750 27624 10806 27680
rect 10874 27624 10930 27680
rect 10998 27624 11054 27680
rect 11122 27624 11178 27680
rect 11246 27624 11302 27680
rect 11370 27624 11426 27680
rect 11494 27624 11550 27680
rect 11618 27624 11674 27680
rect 11742 27624 11798 27680
rect 11866 27624 11922 27680
rect 11990 27624 12046 27680
rect 12114 27624 12170 27680
rect 10254 27500 10310 27556
rect 10378 27500 10434 27556
rect 10502 27500 10558 27556
rect 10626 27500 10682 27556
rect 10750 27500 10806 27556
rect 10874 27500 10930 27556
rect 10998 27500 11054 27556
rect 11122 27500 11178 27556
rect 11246 27500 11302 27556
rect 11370 27500 11426 27556
rect 11494 27500 11550 27556
rect 11618 27500 11674 27556
rect 11742 27500 11798 27556
rect 11866 27500 11922 27556
rect 11990 27500 12046 27556
rect 12114 27500 12170 27556
rect 10254 27376 10310 27432
rect 10378 27376 10434 27432
rect 10502 27376 10558 27432
rect 10626 27376 10682 27432
rect 10750 27376 10806 27432
rect 10874 27376 10930 27432
rect 10998 27376 11054 27432
rect 11122 27376 11178 27432
rect 11246 27376 11302 27432
rect 11370 27376 11426 27432
rect 11494 27376 11550 27432
rect 11618 27376 11674 27432
rect 11742 27376 11798 27432
rect 11866 27376 11922 27432
rect 11990 27376 12046 27432
rect 12114 27376 12170 27432
rect 10254 27252 10310 27308
rect 10378 27252 10434 27308
rect 10502 27252 10558 27308
rect 10626 27252 10682 27308
rect 10750 27252 10806 27308
rect 10874 27252 10930 27308
rect 10998 27252 11054 27308
rect 11122 27252 11178 27308
rect 11246 27252 11302 27308
rect 11370 27252 11426 27308
rect 11494 27252 11550 27308
rect 11618 27252 11674 27308
rect 11742 27252 11798 27308
rect 11866 27252 11922 27308
rect 11990 27252 12046 27308
rect 12114 27252 12170 27308
rect 12871 28492 12927 28548
rect 12995 28492 13051 28548
rect 13119 28492 13175 28548
rect 13243 28492 13299 28548
rect 13367 28492 13423 28548
rect 13491 28492 13547 28548
rect 13615 28492 13671 28548
rect 13739 28492 13795 28548
rect 13863 28492 13919 28548
rect 13987 28492 14043 28548
rect 14111 28492 14167 28548
rect 14235 28492 14291 28548
rect 14359 28492 14415 28548
rect 14483 28492 14539 28548
rect 14607 28492 14663 28548
rect 12871 28368 12927 28424
rect 12995 28368 13051 28424
rect 13119 28368 13175 28424
rect 13243 28368 13299 28424
rect 13367 28368 13423 28424
rect 13491 28368 13547 28424
rect 13615 28368 13671 28424
rect 13739 28368 13795 28424
rect 13863 28368 13919 28424
rect 13987 28368 14043 28424
rect 14111 28368 14167 28424
rect 14235 28368 14291 28424
rect 14359 28368 14415 28424
rect 14483 28368 14539 28424
rect 14607 28368 14663 28424
rect 12871 28244 12927 28300
rect 12995 28244 13051 28300
rect 13119 28244 13175 28300
rect 13243 28244 13299 28300
rect 13367 28244 13423 28300
rect 13491 28244 13547 28300
rect 13615 28244 13671 28300
rect 13739 28244 13795 28300
rect 13863 28244 13919 28300
rect 13987 28244 14043 28300
rect 14111 28244 14167 28300
rect 14235 28244 14291 28300
rect 14359 28244 14415 28300
rect 14483 28244 14539 28300
rect 14607 28244 14663 28300
rect 12871 28120 12927 28176
rect 12995 28120 13051 28176
rect 13119 28120 13175 28176
rect 13243 28120 13299 28176
rect 13367 28120 13423 28176
rect 13491 28120 13547 28176
rect 13615 28120 13671 28176
rect 13739 28120 13795 28176
rect 13863 28120 13919 28176
rect 13987 28120 14043 28176
rect 14111 28120 14167 28176
rect 14235 28120 14291 28176
rect 14359 28120 14415 28176
rect 14483 28120 14539 28176
rect 14607 28120 14663 28176
rect 12871 27996 12927 28052
rect 12995 27996 13051 28052
rect 13119 27996 13175 28052
rect 13243 27996 13299 28052
rect 13367 27996 13423 28052
rect 13491 27996 13547 28052
rect 13615 27996 13671 28052
rect 13739 27996 13795 28052
rect 13863 27996 13919 28052
rect 13987 27996 14043 28052
rect 14111 27996 14167 28052
rect 14235 27996 14291 28052
rect 14359 27996 14415 28052
rect 14483 27996 14539 28052
rect 14607 27996 14663 28052
rect 12871 27872 12927 27928
rect 12995 27872 13051 27928
rect 13119 27872 13175 27928
rect 13243 27872 13299 27928
rect 13367 27872 13423 27928
rect 13491 27872 13547 27928
rect 13615 27872 13671 27928
rect 13739 27872 13795 27928
rect 13863 27872 13919 27928
rect 13987 27872 14043 27928
rect 14111 27872 14167 27928
rect 14235 27872 14291 27928
rect 14359 27872 14415 27928
rect 14483 27872 14539 27928
rect 14607 27872 14663 27928
rect 12871 27748 12927 27804
rect 12995 27748 13051 27804
rect 13119 27748 13175 27804
rect 13243 27748 13299 27804
rect 13367 27748 13423 27804
rect 13491 27748 13547 27804
rect 13615 27748 13671 27804
rect 13739 27748 13795 27804
rect 13863 27748 13919 27804
rect 13987 27748 14043 27804
rect 14111 27748 14167 27804
rect 14235 27748 14291 27804
rect 14359 27748 14415 27804
rect 14483 27748 14539 27804
rect 14607 27748 14663 27804
rect 12871 27624 12927 27680
rect 12995 27624 13051 27680
rect 13119 27624 13175 27680
rect 13243 27624 13299 27680
rect 13367 27624 13423 27680
rect 13491 27624 13547 27680
rect 13615 27624 13671 27680
rect 13739 27624 13795 27680
rect 13863 27624 13919 27680
rect 13987 27624 14043 27680
rect 14111 27624 14167 27680
rect 14235 27624 14291 27680
rect 14359 27624 14415 27680
rect 14483 27624 14539 27680
rect 14607 27624 14663 27680
rect 12871 27500 12927 27556
rect 12995 27500 13051 27556
rect 13119 27500 13175 27556
rect 13243 27500 13299 27556
rect 13367 27500 13423 27556
rect 13491 27500 13547 27556
rect 13615 27500 13671 27556
rect 13739 27500 13795 27556
rect 13863 27500 13919 27556
rect 13987 27500 14043 27556
rect 14111 27500 14167 27556
rect 14235 27500 14291 27556
rect 14359 27500 14415 27556
rect 14483 27500 14539 27556
rect 14607 27500 14663 27556
rect 12871 27376 12927 27432
rect 12995 27376 13051 27432
rect 13119 27376 13175 27432
rect 13243 27376 13299 27432
rect 13367 27376 13423 27432
rect 13491 27376 13547 27432
rect 13615 27376 13671 27432
rect 13739 27376 13795 27432
rect 13863 27376 13919 27432
rect 13987 27376 14043 27432
rect 14111 27376 14167 27432
rect 14235 27376 14291 27432
rect 14359 27376 14415 27432
rect 14483 27376 14539 27432
rect 14607 27376 14663 27432
rect 12871 27252 12927 27308
rect 12995 27252 13051 27308
rect 13119 27252 13175 27308
rect 13243 27252 13299 27308
rect 13367 27252 13423 27308
rect 13491 27252 13547 27308
rect 13615 27252 13671 27308
rect 13739 27252 13795 27308
rect 13863 27252 13919 27308
rect 13987 27252 14043 27308
rect 14111 27252 14167 27308
rect 14235 27252 14291 27308
rect 14359 27252 14415 27308
rect 14483 27252 14539 27308
rect 14607 27252 14663 27308
rect 14902 28574 14958 28576
rect 14902 28522 14904 28574
rect 14904 28522 14956 28574
rect 14956 28522 14958 28574
rect 14902 28466 14958 28522
rect 14902 28414 14904 28466
rect 14904 28414 14956 28466
rect 14956 28414 14958 28466
rect 14902 28358 14958 28414
rect 14902 28306 14904 28358
rect 14904 28306 14956 28358
rect 14956 28306 14958 28358
rect 14902 28250 14958 28306
rect 14902 28198 14904 28250
rect 14904 28198 14956 28250
rect 14956 28198 14958 28250
rect 14902 28142 14958 28198
rect 14902 28090 14904 28142
rect 14904 28090 14956 28142
rect 14956 28090 14958 28142
rect 14902 28034 14958 28090
rect 14902 27982 14904 28034
rect 14904 27982 14956 28034
rect 14956 27982 14958 28034
rect 14902 27926 14958 27982
rect 14902 27874 14904 27926
rect 14904 27874 14956 27926
rect 14956 27874 14958 27926
rect 14902 27818 14958 27874
rect 14902 27766 14904 27818
rect 14904 27766 14956 27818
rect 14956 27766 14958 27818
rect 14902 27710 14958 27766
rect 14902 27658 14904 27710
rect 14904 27658 14956 27710
rect 14956 27658 14958 27710
rect 14902 27602 14958 27658
rect 14902 27550 14904 27602
rect 14904 27550 14956 27602
rect 14956 27550 14958 27602
rect 14902 27494 14958 27550
rect 14902 27442 14904 27494
rect 14904 27442 14956 27494
rect 14956 27442 14958 27494
rect 14902 27386 14958 27442
rect 14902 27334 14904 27386
rect 14904 27334 14956 27386
rect 14956 27334 14958 27386
rect 14902 27278 14958 27334
rect 14902 27226 14904 27278
rect 14904 27226 14956 27278
rect 14956 27226 14958 27278
rect 14902 27224 14958 27226
rect 2491 26898 2547 26954
rect 2615 26898 2671 26954
rect 2491 26774 2547 26830
rect 2615 26774 2671 26830
rect 2491 26650 2547 26706
rect 2615 26650 2671 26706
rect 2491 26526 2547 26582
rect 2615 26526 2671 26582
rect 2491 26402 2547 26458
rect 2615 26402 2671 26458
rect 2491 26278 2547 26334
rect 2615 26278 2671 26334
rect 2491 26154 2547 26210
rect 2615 26154 2671 26210
rect 2491 26030 2547 26086
rect 2615 26030 2671 26086
rect 2491 25906 2547 25962
rect 2615 25906 2671 25962
rect 2491 25782 2547 25838
rect 2615 25782 2671 25838
rect 2491 25658 2547 25714
rect 2615 25658 2671 25714
rect 2491 25534 2547 25590
rect 2615 25534 2671 25590
rect 2491 25410 2547 25466
rect 2615 25410 2671 25466
rect 2491 25286 2547 25342
rect 2615 25286 2671 25342
rect 2491 25162 2547 25218
rect 2615 25162 2671 25218
rect 2491 25038 2547 25094
rect 2615 25038 2671 25094
rect 2491 24914 2547 24970
rect 2615 24914 2671 24970
rect 2491 24790 2547 24846
rect 2615 24790 2671 24846
rect 2491 24666 2547 24722
rect 2615 24666 2671 24722
rect 2491 24542 2547 24598
rect 2615 24542 2671 24598
rect 2491 24418 2547 24474
rect 2615 24418 2671 24474
rect 2491 24294 2547 24350
rect 2615 24294 2671 24350
rect 2491 24170 2547 24226
rect 2615 24170 2671 24226
rect 2491 24046 2547 24102
rect 2615 24046 2671 24102
rect 4861 26898 4917 26954
rect 4985 26898 5041 26954
rect 4861 26774 4917 26830
rect 4985 26774 5041 26830
rect 4861 26650 4917 26706
rect 4985 26650 5041 26706
rect 4861 26526 4917 26582
rect 4985 26526 5041 26582
rect 4861 26402 4917 26458
rect 4985 26402 5041 26458
rect 4861 26278 4917 26334
rect 4985 26278 5041 26334
rect 4861 26154 4917 26210
rect 4985 26154 5041 26210
rect 4861 26030 4917 26086
rect 4985 26030 5041 26086
rect 4861 25906 4917 25962
rect 4985 25906 5041 25962
rect 4861 25782 4917 25838
rect 4985 25782 5041 25838
rect 4861 25658 4917 25714
rect 4985 25658 5041 25714
rect 4861 25534 4917 25590
rect 4985 25534 5041 25590
rect 4861 25410 4917 25466
rect 4985 25410 5041 25466
rect 4861 25286 4917 25342
rect 4985 25286 5041 25342
rect 4861 25162 4917 25218
rect 4985 25162 5041 25218
rect 4861 25038 4917 25094
rect 4985 25038 5041 25094
rect 4861 24914 4917 24970
rect 4985 24914 5041 24970
rect 4861 24790 4917 24846
rect 4985 24790 5041 24846
rect 4861 24666 4917 24722
rect 4985 24666 5041 24722
rect 4861 24542 4917 24598
rect 4985 24542 5041 24598
rect 4861 24418 4917 24474
rect 4985 24418 5041 24474
rect 4861 24294 4917 24350
rect 4985 24294 5041 24350
rect 4861 24170 4917 24226
rect 4985 24170 5041 24226
rect 4861 24046 4917 24102
rect 4985 24046 5041 24102
rect 7275 26898 7331 26954
rect 7399 26898 7455 26954
rect 7523 26898 7579 26954
rect 7647 26898 7703 26954
rect 7275 26774 7331 26830
rect 7399 26774 7455 26830
rect 7523 26774 7579 26830
rect 7647 26774 7703 26830
rect 7275 26650 7331 26706
rect 7399 26650 7455 26706
rect 7523 26650 7579 26706
rect 7647 26650 7703 26706
rect 7275 26526 7331 26582
rect 7399 26526 7455 26582
rect 7523 26526 7579 26582
rect 7647 26526 7703 26582
rect 7275 26402 7331 26458
rect 7399 26402 7455 26458
rect 7523 26402 7579 26458
rect 7647 26402 7703 26458
rect 7275 26278 7331 26334
rect 7399 26278 7455 26334
rect 7523 26278 7579 26334
rect 7647 26278 7703 26334
rect 7275 26154 7331 26210
rect 7399 26154 7455 26210
rect 7523 26154 7579 26210
rect 7647 26154 7703 26210
rect 7275 26030 7331 26086
rect 7399 26030 7455 26086
rect 7523 26030 7579 26086
rect 7647 26030 7703 26086
rect 7275 25906 7331 25962
rect 7399 25906 7455 25962
rect 7523 25906 7579 25962
rect 7647 25906 7703 25962
rect 7275 25782 7331 25838
rect 7399 25782 7455 25838
rect 7523 25782 7579 25838
rect 7647 25782 7703 25838
rect 7275 25658 7331 25714
rect 7399 25658 7455 25714
rect 7523 25658 7579 25714
rect 7647 25658 7703 25714
rect 7275 25534 7331 25590
rect 7399 25534 7455 25590
rect 7523 25534 7579 25590
rect 7647 25534 7703 25590
rect 7275 25410 7331 25466
rect 7399 25410 7455 25466
rect 7523 25410 7579 25466
rect 7647 25410 7703 25466
rect 7275 25286 7331 25342
rect 7399 25286 7455 25342
rect 7523 25286 7579 25342
rect 7647 25286 7703 25342
rect 7275 25162 7331 25218
rect 7399 25162 7455 25218
rect 7523 25162 7579 25218
rect 7647 25162 7703 25218
rect 7275 25038 7331 25094
rect 7399 25038 7455 25094
rect 7523 25038 7579 25094
rect 7647 25038 7703 25094
rect 7275 24914 7331 24970
rect 7399 24914 7455 24970
rect 7523 24914 7579 24970
rect 7647 24914 7703 24970
rect 7275 24790 7331 24846
rect 7399 24790 7455 24846
rect 7523 24790 7579 24846
rect 7647 24790 7703 24846
rect 7275 24666 7331 24722
rect 7399 24666 7455 24722
rect 7523 24666 7579 24722
rect 7647 24666 7703 24722
rect 7275 24542 7331 24598
rect 7399 24542 7455 24598
rect 7523 24542 7579 24598
rect 7647 24542 7703 24598
rect 7275 24418 7331 24474
rect 7399 24418 7455 24474
rect 7523 24418 7579 24474
rect 7647 24418 7703 24474
rect 7275 24294 7331 24350
rect 7399 24294 7455 24350
rect 7523 24294 7579 24350
rect 7647 24294 7703 24350
rect 7275 24170 7331 24226
rect 7399 24170 7455 24226
rect 7523 24170 7579 24226
rect 7647 24170 7703 24226
rect 7275 24046 7331 24102
rect 7399 24046 7455 24102
rect 7523 24046 7579 24102
rect 7647 24046 7703 24102
rect 9937 26898 9993 26954
rect 10061 26898 10117 26954
rect 9937 26774 9993 26830
rect 10061 26774 10117 26830
rect 9937 26650 9993 26706
rect 10061 26650 10117 26706
rect 9937 26526 9993 26582
rect 10061 26526 10117 26582
rect 9937 26402 9993 26458
rect 10061 26402 10117 26458
rect 9937 26278 9993 26334
rect 10061 26278 10117 26334
rect 9937 26154 9993 26210
rect 10061 26154 10117 26210
rect 9937 26030 9993 26086
rect 10061 26030 10117 26086
rect 9937 25906 9993 25962
rect 10061 25906 10117 25962
rect 9937 25782 9993 25838
rect 10061 25782 10117 25838
rect 9937 25658 9993 25714
rect 10061 25658 10117 25714
rect 9937 25534 9993 25590
rect 10061 25534 10117 25590
rect 9937 25410 9993 25466
rect 10061 25410 10117 25466
rect 9937 25286 9993 25342
rect 10061 25286 10117 25342
rect 9937 25162 9993 25218
rect 10061 25162 10117 25218
rect 9937 25038 9993 25094
rect 10061 25038 10117 25094
rect 9937 24914 9993 24970
rect 10061 24914 10117 24970
rect 9937 24790 9993 24846
rect 10061 24790 10117 24846
rect 9937 24666 9993 24722
rect 10061 24666 10117 24722
rect 9937 24542 9993 24598
rect 10061 24542 10117 24598
rect 9937 24418 9993 24474
rect 10061 24418 10117 24474
rect 9937 24294 9993 24350
rect 10061 24294 10117 24350
rect 9937 24170 9993 24226
rect 10061 24170 10117 24226
rect 9937 24046 9993 24102
rect 10061 24046 10117 24102
rect 12307 26898 12363 26954
rect 12431 26898 12487 26954
rect 12307 26774 12363 26830
rect 12431 26774 12487 26830
rect 12307 26650 12363 26706
rect 12431 26650 12487 26706
rect 12307 26526 12363 26582
rect 12431 26526 12487 26582
rect 12307 26402 12363 26458
rect 12431 26402 12487 26458
rect 12307 26278 12363 26334
rect 12431 26278 12487 26334
rect 12307 26154 12363 26210
rect 12431 26154 12487 26210
rect 12307 26030 12363 26086
rect 12431 26030 12487 26086
rect 12307 25906 12363 25962
rect 12431 25906 12487 25962
rect 12307 25782 12363 25838
rect 12431 25782 12487 25838
rect 12307 25658 12363 25714
rect 12431 25658 12487 25714
rect 12307 25534 12363 25590
rect 12431 25534 12487 25590
rect 12307 25410 12363 25466
rect 12431 25410 12487 25466
rect 12307 25286 12363 25342
rect 12431 25286 12487 25342
rect 12307 25162 12363 25218
rect 12431 25162 12487 25218
rect 12307 25038 12363 25094
rect 12431 25038 12487 25094
rect 12307 24914 12363 24970
rect 12431 24914 12487 24970
rect 12307 24790 12363 24846
rect 12431 24790 12487 24846
rect 12307 24666 12363 24722
rect 12431 24666 12487 24722
rect 12307 24542 12363 24598
rect 12431 24542 12487 24598
rect 12307 24418 12363 24474
rect 12431 24418 12487 24474
rect 12307 24294 12363 24350
rect 12431 24294 12487 24350
rect 12307 24170 12363 24226
rect 12431 24170 12487 24226
rect 12307 24046 12363 24102
rect 12431 24046 12487 24102
rect 2491 23698 2547 23754
rect 2615 23698 2671 23754
rect 2491 23574 2547 23630
rect 2615 23574 2671 23630
rect 2491 23450 2547 23506
rect 2615 23450 2671 23506
rect 2491 23326 2547 23382
rect 2615 23326 2671 23382
rect 2491 23202 2547 23258
rect 2615 23202 2671 23258
rect 2491 23078 2547 23134
rect 2615 23078 2671 23134
rect 2491 22954 2547 23010
rect 2615 22954 2671 23010
rect 2491 22830 2547 22886
rect 2615 22830 2671 22886
rect 2491 22706 2547 22762
rect 2615 22706 2671 22762
rect 2491 22582 2547 22638
rect 2615 22582 2671 22638
rect 2491 22458 2547 22514
rect 2615 22458 2671 22514
rect 2491 22334 2547 22390
rect 2615 22334 2671 22390
rect 2491 22210 2547 22266
rect 2615 22210 2671 22266
rect 2491 22086 2547 22142
rect 2615 22086 2671 22142
rect 2491 21962 2547 22018
rect 2615 21962 2671 22018
rect 2491 21838 2547 21894
rect 2615 21838 2671 21894
rect 2491 21714 2547 21770
rect 2615 21714 2671 21770
rect 2491 21590 2547 21646
rect 2615 21590 2671 21646
rect 2491 21466 2547 21522
rect 2615 21466 2671 21522
rect 2491 21342 2547 21398
rect 2615 21342 2671 21398
rect 2491 21218 2547 21274
rect 2615 21218 2671 21274
rect 2491 21094 2547 21150
rect 2615 21094 2671 21150
rect 2491 20970 2547 21026
rect 2615 20970 2671 21026
rect 2491 20846 2547 20902
rect 2615 20846 2671 20902
rect 4861 23698 4917 23754
rect 4985 23698 5041 23754
rect 4861 23574 4917 23630
rect 4985 23574 5041 23630
rect 4861 23450 4917 23506
rect 4985 23450 5041 23506
rect 4861 23326 4917 23382
rect 4985 23326 5041 23382
rect 4861 23202 4917 23258
rect 4985 23202 5041 23258
rect 4861 23078 4917 23134
rect 4985 23078 5041 23134
rect 4861 22954 4917 23010
rect 4985 22954 5041 23010
rect 4861 22830 4917 22886
rect 4985 22830 5041 22886
rect 4861 22706 4917 22762
rect 4985 22706 5041 22762
rect 4861 22582 4917 22638
rect 4985 22582 5041 22638
rect 4861 22458 4917 22514
rect 4985 22458 5041 22514
rect 4861 22334 4917 22390
rect 4985 22334 5041 22390
rect 4861 22210 4917 22266
rect 4985 22210 5041 22266
rect 4861 22086 4917 22142
rect 4985 22086 5041 22142
rect 4861 21962 4917 22018
rect 4985 21962 5041 22018
rect 4861 21838 4917 21894
rect 4985 21838 5041 21894
rect 4861 21714 4917 21770
rect 4985 21714 5041 21770
rect 4861 21590 4917 21646
rect 4985 21590 5041 21646
rect 4861 21466 4917 21522
rect 4985 21466 5041 21522
rect 4861 21342 4917 21398
rect 4985 21342 5041 21398
rect 4861 21218 4917 21274
rect 4985 21218 5041 21274
rect 4861 21094 4917 21150
rect 4985 21094 5041 21150
rect 4861 20970 4917 21026
rect 4985 20970 5041 21026
rect 4861 20846 4917 20902
rect 4985 20846 5041 20902
rect 7275 23698 7331 23754
rect 7399 23698 7455 23754
rect 7523 23698 7579 23754
rect 7647 23698 7703 23754
rect 7275 23574 7331 23630
rect 7399 23574 7455 23630
rect 7523 23574 7579 23630
rect 7647 23574 7703 23630
rect 7275 23450 7331 23506
rect 7399 23450 7455 23506
rect 7523 23450 7579 23506
rect 7647 23450 7703 23506
rect 7275 23326 7331 23382
rect 7399 23326 7455 23382
rect 7523 23326 7579 23382
rect 7647 23326 7703 23382
rect 7275 23202 7331 23258
rect 7399 23202 7455 23258
rect 7523 23202 7579 23258
rect 7647 23202 7703 23258
rect 7275 23078 7331 23134
rect 7399 23078 7455 23134
rect 7523 23078 7579 23134
rect 7647 23078 7703 23134
rect 7275 22954 7331 23010
rect 7399 22954 7455 23010
rect 7523 22954 7579 23010
rect 7647 22954 7703 23010
rect 7275 22830 7331 22886
rect 7399 22830 7455 22886
rect 7523 22830 7579 22886
rect 7647 22830 7703 22886
rect 7275 22706 7331 22762
rect 7399 22706 7455 22762
rect 7523 22706 7579 22762
rect 7647 22706 7703 22762
rect 7275 22582 7331 22638
rect 7399 22582 7455 22638
rect 7523 22582 7579 22638
rect 7647 22582 7703 22638
rect 7275 22458 7331 22514
rect 7399 22458 7455 22514
rect 7523 22458 7579 22514
rect 7647 22458 7703 22514
rect 7275 22334 7331 22390
rect 7399 22334 7455 22390
rect 7523 22334 7579 22390
rect 7647 22334 7703 22390
rect 7275 22210 7331 22266
rect 7399 22210 7455 22266
rect 7523 22210 7579 22266
rect 7647 22210 7703 22266
rect 7275 22086 7331 22142
rect 7399 22086 7455 22142
rect 7523 22086 7579 22142
rect 7647 22086 7703 22142
rect 7275 21962 7331 22018
rect 7399 21962 7455 22018
rect 7523 21962 7579 22018
rect 7647 21962 7703 22018
rect 7275 21838 7331 21894
rect 7399 21838 7455 21894
rect 7523 21838 7579 21894
rect 7647 21838 7703 21894
rect 7275 21714 7331 21770
rect 7399 21714 7455 21770
rect 7523 21714 7579 21770
rect 7647 21714 7703 21770
rect 7275 21590 7331 21646
rect 7399 21590 7455 21646
rect 7523 21590 7579 21646
rect 7647 21590 7703 21646
rect 7275 21466 7331 21522
rect 7399 21466 7455 21522
rect 7523 21466 7579 21522
rect 7647 21466 7703 21522
rect 7275 21342 7331 21398
rect 7399 21342 7455 21398
rect 7523 21342 7579 21398
rect 7647 21342 7703 21398
rect 7275 21218 7331 21274
rect 7399 21218 7455 21274
rect 7523 21218 7579 21274
rect 7647 21218 7703 21274
rect 7275 21094 7331 21150
rect 7399 21094 7455 21150
rect 7523 21094 7579 21150
rect 7647 21094 7703 21150
rect 7275 20970 7331 21026
rect 7399 20970 7455 21026
rect 7523 20970 7579 21026
rect 7647 20970 7703 21026
rect 7275 20846 7331 20902
rect 7399 20846 7455 20902
rect 7523 20846 7579 20902
rect 7647 20846 7703 20902
rect 9937 23698 9993 23754
rect 10061 23698 10117 23754
rect 9937 23574 9993 23630
rect 10061 23574 10117 23630
rect 9937 23450 9993 23506
rect 10061 23450 10117 23506
rect 9937 23326 9993 23382
rect 10061 23326 10117 23382
rect 9937 23202 9993 23258
rect 10061 23202 10117 23258
rect 9937 23078 9993 23134
rect 10061 23078 10117 23134
rect 9937 22954 9993 23010
rect 10061 22954 10117 23010
rect 9937 22830 9993 22886
rect 10061 22830 10117 22886
rect 9937 22706 9993 22762
rect 10061 22706 10117 22762
rect 9937 22582 9993 22638
rect 10061 22582 10117 22638
rect 9937 22458 9993 22514
rect 10061 22458 10117 22514
rect 9937 22334 9993 22390
rect 10061 22334 10117 22390
rect 9937 22210 9993 22266
rect 10061 22210 10117 22266
rect 9937 22086 9993 22142
rect 10061 22086 10117 22142
rect 9937 21962 9993 22018
rect 10061 21962 10117 22018
rect 9937 21838 9993 21894
rect 10061 21838 10117 21894
rect 9937 21714 9993 21770
rect 10061 21714 10117 21770
rect 9937 21590 9993 21646
rect 10061 21590 10117 21646
rect 9937 21466 9993 21522
rect 10061 21466 10117 21522
rect 9937 21342 9993 21398
rect 10061 21342 10117 21398
rect 9937 21218 9993 21274
rect 10061 21218 10117 21274
rect 9937 21094 9993 21150
rect 10061 21094 10117 21150
rect 9937 20970 9993 21026
rect 10061 20970 10117 21026
rect 9937 20846 9993 20902
rect 10061 20846 10117 20902
rect 12307 23698 12363 23754
rect 12431 23698 12487 23754
rect 12307 23574 12363 23630
rect 12431 23574 12487 23630
rect 12307 23450 12363 23506
rect 12431 23450 12487 23506
rect 12307 23326 12363 23382
rect 12431 23326 12487 23382
rect 12307 23202 12363 23258
rect 12431 23202 12487 23258
rect 12307 23078 12363 23134
rect 12431 23078 12487 23134
rect 12307 22954 12363 23010
rect 12431 22954 12487 23010
rect 12307 22830 12363 22886
rect 12431 22830 12487 22886
rect 12307 22706 12363 22762
rect 12431 22706 12487 22762
rect 12307 22582 12363 22638
rect 12431 22582 12487 22638
rect 12307 22458 12363 22514
rect 12431 22458 12487 22514
rect 12307 22334 12363 22390
rect 12431 22334 12487 22390
rect 12307 22210 12363 22266
rect 12431 22210 12487 22266
rect 12307 22086 12363 22142
rect 12431 22086 12487 22142
rect 12307 21962 12363 22018
rect 12431 21962 12487 22018
rect 12307 21838 12363 21894
rect 12431 21838 12487 21894
rect 12307 21714 12363 21770
rect 12431 21714 12487 21770
rect 12307 21590 12363 21646
rect 12431 21590 12487 21646
rect 12307 21466 12363 21522
rect 12431 21466 12487 21522
rect 12307 21342 12363 21398
rect 12431 21342 12487 21398
rect 12307 21218 12363 21274
rect 12431 21218 12487 21274
rect 12307 21094 12363 21150
rect 12431 21094 12487 21150
rect 12307 20970 12363 21026
rect 12431 20970 12487 21026
rect 12307 20846 12363 20902
rect 12431 20846 12487 20902
rect 2491 20498 2547 20554
rect 2615 20498 2671 20554
rect 2491 20374 2547 20430
rect 2615 20374 2671 20430
rect 2491 20250 2547 20306
rect 2615 20250 2671 20306
rect 2491 20126 2547 20182
rect 2615 20126 2671 20182
rect 2491 20002 2547 20058
rect 2615 20002 2671 20058
rect 2491 19878 2547 19934
rect 2615 19878 2671 19934
rect 2491 19754 2547 19810
rect 2615 19754 2671 19810
rect 2491 19630 2547 19686
rect 2615 19630 2671 19686
rect 2491 19506 2547 19562
rect 2615 19506 2671 19562
rect 2491 19382 2547 19438
rect 2615 19382 2671 19438
rect 2491 19258 2547 19314
rect 2615 19258 2671 19314
rect 2491 19134 2547 19190
rect 2615 19134 2671 19190
rect 2491 19010 2547 19066
rect 2615 19010 2671 19066
rect 2491 18886 2547 18942
rect 2615 18886 2671 18942
rect 2491 18762 2547 18818
rect 2615 18762 2671 18818
rect 2491 18638 2547 18694
rect 2615 18638 2671 18694
rect 2491 18514 2547 18570
rect 2615 18514 2671 18570
rect 2491 18390 2547 18446
rect 2615 18390 2671 18446
rect 2491 18266 2547 18322
rect 2615 18266 2671 18322
rect 2491 18142 2547 18198
rect 2615 18142 2671 18198
rect 2491 18018 2547 18074
rect 2615 18018 2671 18074
rect 2491 17894 2547 17950
rect 2615 17894 2671 17950
rect 2491 17770 2547 17826
rect 2615 17770 2671 17826
rect 2491 17646 2547 17702
rect 2615 17646 2671 17702
rect 4861 20498 4917 20554
rect 4985 20498 5041 20554
rect 4861 20374 4917 20430
rect 4985 20374 5041 20430
rect 4861 20250 4917 20306
rect 4985 20250 5041 20306
rect 4861 20126 4917 20182
rect 4985 20126 5041 20182
rect 4861 20002 4917 20058
rect 4985 20002 5041 20058
rect 4861 19878 4917 19934
rect 4985 19878 5041 19934
rect 4861 19754 4917 19810
rect 4985 19754 5041 19810
rect 4861 19630 4917 19686
rect 4985 19630 5041 19686
rect 4861 19506 4917 19562
rect 4985 19506 5041 19562
rect 4861 19382 4917 19438
rect 4985 19382 5041 19438
rect 4861 19258 4917 19314
rect 4985 19258 5041 19314
rect 4861 19134 4917 19190
rect 4985 19134 5041 19190
rect 4861 19010 4917 19066
rect 4985 19010 5041 19066
rect 4861 18886 4917 18942
rect 4985 18886 5041 18942
rect 4861 18762 4917 18818
rect 4985 18762 5041 18818
rect 4861 18638 4917 18694
rect 4985 18638 5041 18694
rect 4861 18514 4917 18570
rect 4985 18514 5041 18570
rect 4861 18390 4917 18446
rect 4985 18390 5041 18446
rect 4861 18266 4917 18322
rect 4985 18266 5041 18322
rect 4861 18142 4917 18198
rect 4985 18142 5041 18198
rect 4861 18018 4917 18074
rect 4985 18018 5041 18074
rect 4861 17894 4917 17950
rect 4985 17894 5041 17950
rect 4861 17770 4917 17826
rect 4985 17770 5041 17826
rect 4861 17646 4917 17702
rect 4985 17646 5041 17702
rect 7275 20498 7331 20554
rect 7399 20498 7455 20554
rect 7523 20498 7579 20554
rect 7647 20498 7703 20554
rect 7275 20374 7331 20430
rect 7399 20374 7455 20430
rect 7523 20374 7579 20430
rect 7647 20374 7703 20430
rect 7275 20250 7331 20306
rect 7399 20250 7455 20306
rect 7523 20250 7579 20306
rect 7647 20250 7703 20306
rect 7275 20126 7331 20182
rect 7399 20126 7455 20182
rect 7523 20126 7579 20182
rect 7647 20126 7703 20182
rect 7275 20002 7331 20058
rect 7399 20002 7455 20058
rect 7523 20002 7579 20058
rect 7647 20002 7703 20058
rect 7275 19878 7331 19934
rect 7399 19878 7455 19934
rect 7523 19878 7579 19934
rect 7647 19878 7703 19934
rect 7275 19754 7331 19810
rect 7399 19754 7455 19810
rect 7523 19754 7579 19810
rect 7647 19754 7703 19810
rect 7275 19630 7331 19686
rect 7399 19630 7455 19686
rect 7523 19630 7579 19686
rect 7647 19630 7703 19686
rect 7275 19506 7331 19562
rect 7399 19506 7455 19562
rect 7523 19506 7579 19562
rect 7647 19506 7703 19562
rect 7275 19382 7331 19438
rect 7399 19382 7455 19438
rect 7523 19382 7579 19438
rect 7647 19382 7703 19438
rect 7275 19258 7331 19314
rect 7399 19258 7455 19314
rect 7523 19258 7579 19314
rect 7647 19258 7703 19314
rect 7275 19134 7331 19190
rect 7399 19134 7455 19190
rect 7523 19134 7579 19190
rect 7647 19134 7703 19190
rect 7275 19010 7331 19066
rect 7399 19010 7455 19066
rect 7523 19010 7579 19066
rect 7647 19010 7703 19066
rect 7275 18886 7331 18942
rect 7399 18886 7455 18942
rect 7523 18886 7579 18942
rect 7647 18886 7703 18942
rect 7275 18762 7331 18818
rect 7399 18762 7455 18818
rect 7523 18762 7579 18818
rect 7647 18762 7703 18818
rect 7275 18638 7331 18694
rect 7399 18638 7455 18694
rect 7523 18638 7579 18694
rect 7647 18638 7703 18694
rect 7275 18514 7331 18570
rect 7399 18514 7455 18570
rect 7523 18514 7579 18570
rect 7647 18514 7703 18570
rect 7275 18390 7331 18446
rect 7399 18390 7455 18446
rect 7523 18390 7579 18446
rect 7647 18390 7703 18446
rect 7275 18266 7331 18322
rect 7399 18266 7455 18322
rect 7523 18266 7579 18322
rect 7647 18266 7703 18322
rect 7275 18142 7331 18198
rect 7399 18142 7455 18198
rect 7523 18142 7579 18198
rect 7647 18142 7703 18198
rect 7275 18018 7331 18074
rect 7399 18018 7455 18074
rect 7523 18018 7579 18074
rect 7647 18018 7703 18074
rect 7275 17894 7331 17950
rect 7399 17894 7455 17950
rect 7523 17894 7579 17950
rect 7647 17894 7703 17950
rect 7275 17770 7331 17826
rect 7399 17770 7455 17826
rect 7523 17770 7579 17826
rect 7647 17770 7703 17826
rect 7275 17646 7331 17702
rect 7399 17646 7455 17702
rect 7523 17646 7579 17702
rect 7647 17646 7703 17702
rect 9937 20498 9993 20554
rect 10061 20498 10117 20554
rect 9937 20374 9993 20430
rect 10061 20374 10117 20430
rect 9937 20250 9993 20306
rect 10061 20250 10117 20306
rect 9937 20126 9993 20182
rect 10061 20126 10117 20182
rect 9937 20002 9993 20058
rect 10061 20002 10117 20058
rect 9937 19878 9993 19934
rect 10061 19878 10117 19934
rect 9937 19754 9993 19810
rect 10061 19754 10117 19810
rect 9937 19630 9993 19686
rect 10061 19630 10117 19686
rect 9937 19506 9993 19562
rect 10061 19506 10117 19562
rect 9937 19382 9993 19438
rect 10061 19382 10117 19438
rect 9937 19258 9993 19314
rect 10061 19258 10117 19314
rect 9937 19134 9993 19190
rect 10061 19134 10117 19190
rect 9937 19010 9993 19066
rect 10061 19010 10117 19066
rect 9937 18886 9993 18942
rect 10061 18886 10117 18942
rect 9937 18762 9993 18818
rect 10061 18762 10117 18818
rect 9937 18638 9993 18694
rect 10061 18638 10117 18694
rect 9937 18514 9993 18570
rect 10061 18514 10117 18570
rect 9937 18390 9993 18446
rect 10061 18390 10117 18446
rect 9937 18266 9993 18322
rect 10061 18266 10117 18322
rect 9937 18142 9993 18198
rect 10061 18142 10117 18198
rect 9937 18018 9993 18074
rect 10061 18018 10117 18074
rect 9937 17894 9993 17950
rect 10061 17894 10117 17950
rect 9937 17770 9993 17826
rect 10061 17770 10117 17826
rect 9937 17646 9993 17702
rect 10061 17646 10117 17702
rect 12307 20498 12363 20554
rect 12431 20498 12487 20554
rect 12307 20374 12363 20430
rect 12431 20374 12487 20430
rect 12307 20250 12363 20306
rect 12431 20250 12487 20306
rect 12307 20126 12363 20182
rect 12431 20126 12487 20182
rect 12307 20002 12363 20058
rect 12431 20002 12487 20058
rect 12307 19878 12363 19934
rect 12431 19878 12487 19934
rect 12307 19754 12363 19810
rect 12431 19754 12487 19810
rect 12307 19630 12363 19686
rect 12431 19630 12487 19686
rect 12307 19506 12363 19562
rect 12431 19506 12487 19562
rect 12307 19382 12363 19438
rect 12431 19382 12487 19438
rect 12307 19258 12363 19314
rect 12431 19258 12487 19314
rect 12307 19134 12363 19190
rect 12431 19134 12487 19190
rect 12307 19010 12363 19066
rect 12431 19010 12487 19066
rect 12307 18886 12363 18942
rect 12431 18886 12487 18942
rect 12307 18762 12363 18818
rect 12431 18762 12487 18818
rect 12307 18638 12363 18694
rect 12431 18638 12487 18694
rect 12307 18514 12363 18570
rect 12431 18514 12487 18570
rect 12307 18390 12363 18446
rect 12431 18390 12487 18446
rect 12307 18266 12363 18322
rect 12431 18266 12487 18322
rect 12307 18142 12363 18198
rect 12431 18142 12487 18198
rect 12307 18018 12363 18074
rect 12431 18018 12487 18074
rect 12307 17894 12363 17950
rect 12431 17894 12487 17950
rect 12307 17770 12363 17826
rect 12431 17770 12487 17826
rect 12307 17646 12363 17702
rect 12431 17646 12487 17702
rect 2491 17298 2547 17354
rect 2615 17298 2671 17354
rect 2491 17174 2547 17230
rect 2615 17174 2671 17230
rect 2491 17050 2547 17106
rect 2615 17050 2671 17106
rect 2491 16926 2547 16982
rect 2615 16926 2671 16982
rect 2491 16802 2547 16858
rect 2615 16802 2671 16858
rect 2491 16678 2547 16734
rect 2615 16678 2671 16734
rect 2491 16554 2547 16610
rect 2615 16554 2671 16610
rect 2491 16430 2547 16486
rect 2615 16430 2671 16486
rect 2491 16306 2547 16362
rect 2615 16306 2671 16362
rect 2491 16182 2547 16238
rect 2615 16182 2671 16238
rect 2491 16058 2547 16114
rect 2615 16058 2671 16114
rect 2491 15934 2547 15990
rect 2615 15934 2671 15990
rect 2491 15810 2547 15866
rect 2615 15810 2671 15866
rect 2491 15686 2547 15742
rect 2615 15686 2671 15742
rect 2491 15562 2547 15618
rect 2615 15562 2671 15618
rect 2491 15438 2547 15494
rect 2615 15438 2671 15494
rect 2491 15314 2547 15370
rect 2615 15314 2671 15370
rect 2491 15190 2547 15246
rect 2615 15190 2671 15246
rect 2491 15066 2547 15122
rect 2615 15066 2671 15122
rect 2491 14942 2547 14998
rect 2615 14942 2671 14998
rect 2491 14818 2547 14874
rect 2615 14818 2671 14874
rect 2491 14694 2547 14750
rect 2615 14694 2671 14750
rect 2491 14570 2547 14626
rect 2615 14570 2671 14626
rect 2491 14446 2547 14502
rect 2615 14446 2671 14502
rect 4861 17298 4917 17354
rect 4985 17298 5041 17354
rect 4861 17174 4917 17230
rect 4985 17174 5041 17230
rect 4861 17050 4917 17106
rect 4985 17050 5041 17106
rect 4861 16926 4917 16982
rect 4985 16926 5041 16982
rect 4861 16802 4917 16858
rect 4985 16802 5041 16858
rect 4861 16678 4917 16734
rect 4985 16678 5041 16734
rect 4861 16554 4917 16610
rect 4985 16554 5041 16610
rect 4861 16430 4917 16486
rect 4985 16430 5041 16486
rect 4861 16306 4917 16362
rect 4985 16306 5041 16362
rect 4861 16182 4917 16238
rect 4985 16182 5041 16238
rect 4861 16058 4917 16114
rect 4985 16058 5041 16114
rect 4861 15934 4917 15990
rect 4985 15934 5041 15990
rect 4861 15810 4917 15866
rect 4985 15810 5041 15866
rect 4861 15686 4917 15742
rect 4985 15686 5041 15742
rect 4861 15562 4917 15618
rect 4985 15562 5041 15618
rect 4861 15438 4917 15494
rect 4985 15438 5041 15494
rect 4861 15314 4917 15370
rect 4985 15314 5041 15370
rect 4861 15190 4917 15246
rect 4985 15190 5041 15246
rect 4861 15066 4917 15122
rect 4985 15066 5041 15122
rect 4861 14942 4917 14998
rect 4985 14942 5041 14998
rect 4861 14818 4917 14874
rect 4985 14818 5041 14874
rect 4861 14694 4917 14750
rect 4985 14694 5041 14750
rect 4861 14570 4917 14626
rect 4985 14570 5041 14626
rect 4861 14446 4917 14502
rect 4985 14446 5041 14502
rect 7275 17298 7331 17354
rect 7399 17298 7455 17354
rect 7523 17298 7579 17354
rect 7647 17298 7703 17354
rect 7275 17174 7331 17230
rect 7399 17174 7455 17230
rect 7523 17174 7579 17230
rect 7647 17174 7703 17230
rect 7275 17050 7331 17106
rect 7399 17050 7455 17106
rect 7523 17050 7579 17106
rect 7647 17050 7703 17106
rect 7275 16926 7331 16982
rect 7399 16926 7455 16982
rect 7523 16926 7579 16982
rect 7647 16926 7703 16982
rect 7275 16802 7331 16858
rect 7399 16802 7455 16858
rect 7523 16802 7579 16858
rect 7647 16802 7703 16858
rect 7275 16678 7331 16734
rect 7399 16678 7455 16734
rect 7523 16678 7579 16734
rect 7647 16678 7703 16734
rect 7275 16554 7331 16610
rect 7399 16554 7455 16610
rect 7523 16554 7579 16610
rect 7647 16554 7703 16610
rect 7275 16430 7331 16486
rect 7399 16430 7455 16486
rect 7523 16430 7579 16486
rect 7647 16430 7703 16486
rect 7275 16306 7331 16362
rect 7399 16306 7455 16362
rect 7523 16306 7579 16362
rect 7647 16306 7703 16362
rect 7275 16182 7331 16238
rect 7399 16182 7455 16238
rect 7523 16182 7579 16238
rect 7647 16182 7703 16238
rect 7275 16058 7331 16114
rect 7399 16058 7455 16114
rect 7523 16058 7579 16114
rect 7647 16058 7703 16114
rect 7275 15934 7331 15990
rect 7399 15934 7455 15990
rect 7523 15934 7579 15990
rect 7647 15934 7703 15990
rect 7275 15810 7331 15866
rect 7399 15810 7455 15866
rect 7523 15810 7579 15866
rect 7647 15810 7703 15866
rect 7275 15686 7331 15742
rect 7399 15686 7455 15742
rect 7523 15686 7579 15742
rect 7647 15686 7703 15742
rect 7275 15562 7331 15618
rect 7399 15562 7455 15618
rect 7523 15562 7579 15618
rect 7647 15562 7703 15618
rect 7275 15438 7331 15494
rect 7399 15438 7455 15494
rect 7523 15438 7579 15494
rect 7647 15438 7703 15494
rect 7275 15314 7331 15370
rect 7399 15314 7455 15370
rect 7523 15314 7579 15370
rect 7647 15314 7703 15370
rect 7275 15190 7331 15246
rect 7399 15190 7455 15246
rect 7523 15190 7579 15246
rect 7647 15190 7703 15246
rect 7275 15066 7331 15122
rect 7399 15066 7455 15122
rect 7523 15066 7579 15122
rect 7647 15066 7703 15122
rect 7275 14942 7331 14998
rect 7399 14942 7455 14998
rect 7523 14942 7579 14998
rect 7647 14942 7703 14998
rect 7275 14818 7331 14874
rect 7399 14818 7455 14874
rect 7523 14818 7579 14874
rect 7647 14818 7703 14874
rect 7275 14694 7331 14750
rect 7399 14694 7455 14750
rect 7523 14694 7579 14750
rect 7647 14694 7703 14750
rect 7275 14570 7331 14626
rect 7399 14570 7455 14626
rect 7523 14570 7579 14626
rect 7647 14570 7703 14626
rect 7275 14446 7331 14502
rect 7399 14446 7455 14502
rect 7523 14446 7579 14502
rect 7647 14446 7703 14502
rect 9937 17298 9993 17354
rect 10061 17298 10117 17354
rect 9937 17174 9993 17230
rect 10061 17174 10117 17230
rect 9937 17050 9993 17106
rect 10061 17050 10117 17106
rect 9937 16926 9993 16982
rect 10061 16926 10117 16982
rect 9937 16802 9993 16858
rect 10061 16802 10117 16858
rect 9937 16678 9993 16734
rect 10061 16678 10117 16734
rect 9937 16554 9993 16610
rect 10061 16554 10117 16610
rect 9937 16430 9993 16486
rect 10061 16430 10117 16486
rect 9937 16306 9993 16362
rect 10061 16306 10117 16362
rect 9937 16182 9993 16238
rect 10061 16182 10117 16238
rect 9937 16058 9993 16114
rect 10061 16058 10117 16114
rect 9937 15934 9993 15990
rect 10061 15934 10117 15990
rect 9937 15810 9993 15866
rect 10061 15810 10117 15866
rect 9937 15686 9993 15742
rect 10061 15686 10117 15742
rect 9937 15562 9993 15618
rect 10061 15562 10117 15618
rect 9937 15438 9993 15494
rect 10061 15438 10117 15494
rect 9937 15314 9993 15370
rect 10061 15314 10117 15370
rect 9937 15190 9993 15246
rect 10061 15190 10117 15246
rect 9937 15066 9993 15122
rect 10061 15066 10117 15122
rect 9937 14942 9993 14998
rect 10061 14942 10117 14998
rect 9937 14818 9993 14874
rect 10061 14818 10117 14874
rect 9937 14694 9993 14750
rect 10061 14694 10117 14750
rect 9937 14570 9993 14626
rect 10061 14570 10117 14626
rect 9937 14446 9993 14502
rect 10061 14446 10117 14502
rect 12307 17298 12363 17354
rect 12431 17298 12487 17354
rect 12307 17174 12363 17230
rect 12431 17174 12487 17230
rect 12307 17050 12363 17106
rect 12431 17050 12487 17106
rect 12307 16926 12363 16982
rect 12431 16926 12487 16982
rect 12307 16802 12363 16858
rect 12431 16802 12487 16858
rect 12307 16678 12363 16734
rect 12431 16678 12487 16734
rect 12307 16554 12363 16610
rect 12431 16554 12487 16610
rect 12307 16430 12363 16486
rect 12431 16430 12487 16486
rect 12307 16306 12363 16362
rect 12431 16306 12487 16362
rect 12307 16182 12363 16238
rect 12431 16182 12487 16238
rect 12307 16058 12363 16114
rect 12431 16058 12487 16114
rect 12307 15934 12363 15990
rect 12431 15934 12487 15990
rect 12307 15810 12363 15866
rect 12431 15810 12487 15866
rect 12307 15686 12363 15742
rect 12431 15686 12487 15742
rect 12307 15562 12363 15618
rect 12431 15562 12487 15618
rect 12307 15438 12363 15494
rect 12431 15438 12487 15494
rect 12307 15314 12363 15370
rect 12431 15314 12487 15370
rect 12307 15190 12363 15246
rect 12431 15190 12487 15246
rect 12307 15066 12363 15122
rect 12431 15066 12487 15122
rect 12307 14942 12363 14998
rect 12431 14942 12487 14998
rect 12307 14818 12363 14874
rect 12431 14818 12487 14874
rect 12307 14694 12363 14750
rect 12431 14694 12487 14750
rect 12307 14570 12363 14626
rect 12431 14570 12487 14626
rect 12307 14446 12363 14502
rect 12431 14446 12487 14502
rect 20 14174 76 14176
rect 20 14122 22 14174
rect 22 14122 74 14174
rect 74 14122 76 14174
rect 20 14066 76 14122
rect 20 14014 22 14066
rect 22 14014 74 14066
rect 74 14014 76 14066
rect 20 13958 76 14014
rect 20 13906 22 13958
rect 22 13906 74 13958
rect 74 13906 76 13958
rect 20 13850 76 13906
rect 20 13798 22 13850
rect 22 13798 74 13850
rect 74 13798 76 13850
rect 20 13742 76 13798
rect 20 13690 22 13742
rect 22 13690 74 13742
rect 74 13690 76 13742
rect 20 13634 76 13690
rect 20 13582 22 13634
rect 22 13582 74 13634
rect 74 13582 76 13634
rect 20 13526 76 13582
rect 20 13474 22 13526
rect 22 13474 74 13526
rect 74 13474 76 13526
rect 20 13418 76 13474
rect 20 13366 22 13418
rect 22 13366 74 13418
rect 74 13366 76 13418
rect 20 13310 76 13366
rect 20 13258 22 13310
rect 22 13258 74 13310
rect 74 13258 76 13310
rect 20 13202 76 13258
rect 20 13150 22 13202
rect 22 13150 74 13202
rect 74 13150 76 13202
rect 20 13094 76 13150
rect 20 13042 22 13094
rect 22 13042 74 13094
rect 74 13042 76 13094
rect 20 12986 76 13042
rect 20 12934 22 12986
rect 22 12934 74 12986
rect 74 12934 76 12986
rect 20 12878 76 12934
rect 20 12826 22 12878
rect 22 12826 74 12878
rect 74 12826 76 12878
rect 20 12824 76 12826
rect 315 14092 371 14148
rect 439 14092 495 14148
rect 563 14092 619 14148
rect 687 14092 743 14148
rect 811 14092 867 14148
rect 935 14092 991 14148
rect 1059 14092 1115 14148
rect 1183 14092 1239 14148
rect 1307 14092 1363 14148
rect 1431 14092 1487 14148
rect 1555 14092 1611 14148
rect 1679 14092 1735 14148
rect 1803 14092 1859 14148
rect 1927 14092 1983 14148
rect 2051 14092 2107 14148
rect 315 13968 371 14024
rect 439 13968 495 14024
rect 563 13968 619 14024
rect 687 13968 743 14024
rect 811 13968 867 14024
rect 935 13968 991 14024
rect 1059 13968 1115 14024
rect 1183 13968 1239 14024
rect 1307 13968 1363 14024
rect 1431 13968 1487 14024
rect 1555 13968 1611 14024
rect 1679 13968 1735 14024
rect 1803 13968 1859 14024
rect 1927 13968 1983 14024
rect 2051 13968 2107 14024
rect 315 13844 371 13900
rect 439 13844 495 13900
rect 563 13844 619 13900
rect 687 13844 743 13900
rect 811 13844 867 13900
rect 935 13844 991 13900
rect 1059 13844 1115 13900
rect 1183 13844 1239 13900
rect 1307 13844 1363 13900
rect 1431 13844 1487 13900
rect 1555 13844 1611 13900
rect 1679 13844 1735 13900
rect 1803 13844 1859 13900
rect 1927 13844 1983 13900
rect 2051 13844 2107 13900
rect 315 13720 371 13776
rect 439 13720 495 13776
rect 563 13720 619 13776
rect 687 13720 743 13776
rect 811 13720 867 13776
rect 935 13720 991 13776
rect 1059 13720 1115 13776
rect 1183 13720 1239 13776
rect 1307 13720 1363 13776
rect 1431 13720 1487 13776
rect 1555 13720 1611 13776
rect 1679 13720 1735 13776
rect 1803 13720 1859 13776
rect 1927 13720 1983 13776
rect 2051 13720 2107 13776
rect 315 13596 371 13652
rect 439 13596 495 13652
rect 563 13596 619 13652
rect 687 13596 743 13652
rect 811 13596 867 13652
rect 935 13596 991 13652
rect 1059 13596 1115 13652
rect 1183 13596 1239 13652
rect 1307 13596 1363 13652
rect 1431 13596 1487 13652
rect 1555 13596 1611 13652
rect 1679 13596 1735 13652
rect 1803 13596 1859 13652
rect 1927 13596 1983 13652
rect 2051 13596 2107 13652
rect 315 13472 371 13528
rect 439 13472 495 13528
rect 563 13472 619 13528
rect 687 13472 743 13528
rect 811 13472 867 13528
rect 935 13472 991 13528
rect 1059 13472 1115 13528
rect 1183 13472 1239 13528
rect 1307 13472 1363 13528
rect 1431 13472 1487 13528
rect 1555 13472 1611 13528
rect 1679 13472 1735 13528
rect 1803 13472 1859 13528
rect 1927 13472 1983 13528
rect 2051 13472 2107 13528
rect 315 13348 371 13404
rect 439 13348 495 13404
rect 563 13348 619 13404
rect 687 13348 743 13404
rect 811 13348 867 13404
rect 935 13348 991 13404
rect 1059 13348 1115 13404
rect 1183 13348 1239 13404
rect 1307 13348 1363 13404
rect 1431 13348 1487 13404
rect 1555 13348 1611 13404
rect 1679 13348 1735 13404
rect 1803 13348 1859 13404
rect 1927 13348 1983 13404
rect 2051 13348 2107 13404
rect 315 13224 371 13280
rect 439 13224 495 13280
rect 563 13224 619 13280
rect 687 13224 743 13280
rect 811 13224 867 13280
rect 935 13224 991 13280
rect 1059 13224 1115 13280
rect 1183 13224 1239 13280
rect 1307 13224 1363 13280
rect 1431 13224 1487 13280
rect 1555 13224 1611 13280
rect 1679 13224 1735 13280
rect 1803 13224 1859 13280
rect 1927 13224 1983 13280
rect 2051 13224 2107 13280
rect 315 13100 371 13156
rect 439 13100 495 13156
rect 563 13100 619 13156
rect 687 13100 743 13156
rect 811 13100 867 13156
rect 935 13100 991 13156
rect 1059 13100 1115 13156
rect 1183 13100 1239 13156
rect 1307 13100 1363 13156
rect 1431 13100 1487 13156
rect 1555 13100 1611 13156
rect 1679 13100 1735 13156
rect 1803 13100 1859 13156
rect 1927 13100 1983 13156
rect 2051 13100 2107 13156
rect 315 12976 371 13032
rect 439 12976 495 13032
rect 563 12976 619 13032
rect 687 12976 743 13032
rect 811 12976 867 13032
rect 935 12976 991 13032
rect 1059 12976 1115 13032
rect 1183 12976 1239 13032
rect 1307 12976 1363 13032
rect 1431 12976 1487 13032
rect 1555 12976 1611 13032
rect 1679 12976 1735 13032
rect 1803 12976 1859 13032
rect 1927 12976 1983 13032
rect 2051 12976 2107 13032
rect 315 12852 371 12908
rect 439 12852 495 12908
rect 563 12852 619 12908
rect 687 12852 743 12908
rect 811 12852 867 12908
rect 935 12852 991 12908
rect 1059 12852 1115 12908
rect 1183 12852 1239 12908
rect 1307 12852 1363 12908
rect 1431 12852 1487 12908
rect 1555 12852 1611 12908
rect 1679 12852 1735 12908
rect 1803 12852 1859 12908
rect 1927 12852 1983 12908
rect 2051 12852 2107 12908
rect 2808 14092 2864 14148
rect 2932 14092 2988 14148
rect 3056 14092 3112 14148
rect 3180 14092 3236 14148
rect 3304 14092 3360 14148
rect 3428 14092 3484 14148
rect 3552 14092 3608 14148
rect 3676 14092 3732 14148
rect 3800 14092 3856 14148
rect 3924 14092 3980 14148
rect 4048 14092 4104 14148
rect 4172 14092 4228 14148
rect 4296 14092 4352 14148
rect 4420 14092 4476 14148
rect 4544 14092 4600 14148
rect 4668 14092 4724 14148
rect 2808 13968 2864 14024
rect 2932 13968 2988 14024
rect 3056 13968 3112 14024
rect 3180 13968 3236 14024
rect 3304 13968 3360 14024
rect 3428 13968 3484 14024
rect 3552 13968 3608 14024
rect 3676 13968 3732 14024
rect 3800 13968 3856 14024
rect 3924 13968 3980 14024
rect 4048 13968 4104 14024
rect 4172 13968 4228 14024
rect 4296 13968 4352 14024
rect 4420 13968 4476 14024
rect 4544 13968 4600 14024
rect 4668 13968 4724 14024
rect 2808 13844 2864 13900
rect 2932 13844 2988 13900
rect 3056 13844 3112 13900
rect 3180 13844 3236 13900
rect 3304 13844 3360 13900
rect 3428 13844 3484 13900
rect 3552 13844 3608 13900
rect 3676 13844 3732 13900
rect 3800 13844 3856 13900
rect 3924 13844 3980 13900
rect 4048 13844 4104 13900
rect 4172 13844 4228 13900
rect 4296 13844 4352 13900
rect 4420 13844 4476 13900
rect 4544 13844 4600 13900
rect 4668 13844 4724 13900
rect 2808 13720 2864 13776
rect 2932 13720 2988 13776
rect 3056 13720 3112 13776
rect 3180 13720 3236 13776
rect 3304 13720 3360 13776
rect 3428 13720 3484 13776
rect 3552 13720 3608 13776
rect 3676 13720 3732 13776
rect 3800 13720 3856 13776
rect 3924 13720 3980 13776
rect 4048 13720 4104 13776
rect 4172 13720 4228 13776
rect 4296 13720 4352 13776
rect 4420 13720 4476 13776
rect 4544 13720 4600 13776
rect 4668 13720 4724 13776
rect 2808 13596 2864 13652
rect 2932 13596 2988 13652
rect 3056 13596 3112 13652
rect 3180 13596 3236 13652
rect 3304 13596 3360 13652
rect 3428 13596 3484 13652
rect 3552 13596 3608 13652
rect 3676 13596 3732 13652
rect 3800 13596 3856 13652
rect 3924 13596 3980 13652
rect 4048 13596 4104 13652
rect 4172 13596 4228 13652
rect 4296 13596 4352 13652
rect 4420 13596 4476 13652
rect 4544 13596 4600 13652
rect 4668 13596 4724 13652
rect 2808 13472 2864 13528
rect 2932 13472 2988 13528
rect 3056 13472 3112 13528
rect 3180 13472 3236 13528
rect 3304 13472 3360 13528
rect 3428 13472 3484 13528
rect 3552 13472 3608 13528
rect 3676 13472 3732 13528
rect 3800 13472 3856 13528
rect 3924 13472 3980 13528
rect 4048 13472 4104 13528
rect 4172 13472 4228 13528
rect 4296 13472 4352 13528
rect 4420 13472 4476 13528
rect 4544 13472 4600 13528
rect 4668 13472 4724 13528
rect 2808 13348 2864 13404
rect 2932 13348 2988 13404
rect 3056 13348 3112 13404
rect 3180 13348 3236 13404
rect 3304 13348 3360 13404
rect 3428 13348 3484 13404
rect 3552 13348 3608 13404
rect 3676 13348 3732 13404
rect 3800 13348 3856 13404
rect 3924 13348 3980 13404
rect 4048 13348 4104 13404
rect 4172 13348 4228 13404
rect 4296 13348 4352 13404
rect 4420 13348 4476 13404
rect 4544 13348 4600 13404
rect 4668 13348 4724 13404
rect 2808 13224 2864 13280
rect 2932 13224 2988 13280
rect 3056 13224 3112 13280
rect 3180 13224 3236 13280
rect 3304 13224 3360 13280
rect 3428 13224 3484 13280
rect 3552 13224 3608 13280
rect 3676 13224 3732 13280
rect 3800 13224 3856 13280
rect 3924 13224 3980 13280
rect 4048 13224 4104 13280
rect 4172 13224 4228 13280
rect 4296 13224 4352 13280
rect 4420 13224 4476 13280
rect 4544 13224 4600 13280
rect 4668 13224 4724 13280
rect 2808 13100 2864 13156
rect 2932 13100 2988 13156
rect 3056 13100 3112 13156
rect 3180 13100 3236 13156
rect 3304 13100 3360 13156
rect 3428 13100 3484 13156
rect 3552 13100 3608 13156
rect 3676 13100 3732 13156
rect 3800 13100 3856 13156
rect 3924 13100 3980 13156
rect 4048 13100 4104 13156
rect 4172 13100 4228 13156
rect 4296 13100 4352 13156
rect 4420 13100 4476 13156
rect 4544 13100 4600 13156
rect 4668 13100 4724 13156
rect 2808 12976 2864 13032
rect 2932 12976 2988 13032
rect 3056 12976 3112 13032
rect 3180 12976 3236 13032
rect 3304 12976 3360 13032
rect 3428 12976 3484 13032
rect 3552 12976 3608 13032
rect 3676 12976 3732 13032
rect 3800 12976 3856 13032
rect 3924 12976 3980 13032
rect 4048 12976 4104 13032
rect 4172 12976 4228 13032
rect 4296 12976 4352 13032
rect 4420 12976 4476 13032
rect 4544 12976 4600 13032
rect 4668 12976 4724 13032
rect 2808 12852 2864 12908
rect 2932 12852 2988 12908
rect 3056 12852 3112 12908
rect 3180 12852 3236 12908
rect 3304 12852 3360 12908
rect 3428 12852 3484 12908
rect 3552 12852 3608 12908
rect 3676 12852 3732 12908
rect 3800 12852 3856 12908
rect 3924 12852 3980 12908
rect 4048 12852 4104 12908
rect 4172 12852 4228 12908
rect 4296 12852 4352 12908
rect 4420 12852 4476 12908
rect 4544 12852 4600 12908
rect 4668 12852 4724 12908
rect 5178 14092 5234 14148
rect 5302 14092 5358 14148
rect 5426 14092 5482 14148
rect 5550 14092 5606 14148
rect 5674 14092 5730 14148
rect 5798 14092 5854 14148
rect 5922 14092 5978 14148
rect 6046 14092 6102 14148
rect 6170 14092 6226 14148
rect 6294 14092 6350 14148
rect 6418 14092 6474 14148
rect 6542 14092 6598 14148
rect 6666 14092 6722 14148
rect 6790 14092 6846 14148
rect 6914 14092 6970 14148
rect 7038 14092 7094 14148
rect 5178 13968 5234 14024
rect 5302 13968 5358 14024
rect 5426 13968 5482 14024
rect 5550 13968 5606 14024
rect 5674 13968 5730 14024
rect 5798 13968 5854 14024
rect 5922 13968 5978 14024
rect 6046 13968 6102 14024
rect 6170 13968 6226 14024
rect 6294 13968 6350 14024
rect 6418 13968 6474 14024
rect 6542 13968 6598 14024
rect 6666 13968 6722 14024
rect 6790 13968 6846 14024
rect 6914 13968 6970 14024
rect 7038 13968 7094 14024
rect 5178 13844 5234 13900
rect 5302 13844 5358 13900
rect 5426 13844 5482 13900
rect 5550 13844 5606 13900
rect 5674 13844 5730 13900
rect 5798 13844 5854 13900
rect 5922 13844 5978 13900
rect 6046 13844 6102 13900
rect 6170 13844 6226 13900
rect 6294 13844 6350 13900
rect 6418 13844 6474 13900
rect 6542 13844 6598 13900
rect 6666 13844 6722 13900
rect 6790 13844 6846 13900
rect 6914 13844 6970 13900
rect 7038 13844 7094 13900
rect 5178 13720 5234 13776
rect 5302 13720 5358 13776
rect 5426 13720 5482 13776
rect 5550 13720 5606 13776
rect 5674 13720 5730 13776
rect 5798 13720 5854 13776
rect 5922 13720 5978 13776
rect 6046 13720 6102 13776
rect 6170 13720 6226 13776
rect 6294 13720 6350 13776
rect 6418 13720 6474 13776
rect 6542 13720 6598 13776
rect 6666 13720 6722 13776
rect 6790 13720 6846 13776
rect 6914 13720 6970 13776
rect 7038 13720 7094 13776
rect 5178 13596 5234 13652
rect 5302 13596 5358 13652
rect 5426 13596 5482 13652
rect 5550 13596 5606 13652
rect 5674 13596 5730 13652
rect 5798 13596 5854 13652
rect 5922 13596 5978 13652
rect 6046 13596 6102 13652
rect 6170 13596 6226 13652
rect 6294 13596 6350 13652
rect 6418 13596 6474 13652
rect 6542 13596 6598 13652
rect 6666 13596 6722 13652
rect 6790 13596 6846 13652
rect 6914 13596 6970 13652
rect 7038 13596 7094 13652
rect 5178 13472 5234 13528
rect 5302 13472 5358 13528
rect 5426 13472 5482 13528
rect 5550 13472 5606 13528
rect 5674 13472 5730 13528
rect 5798 13472 5854 13528
rect 5922 13472 5978 13528
rect 6046 13472 6102 13528
rect 6170 13472 6226 13528
rect 6294 13472 6350 13528
rect 6418 13472 6474 13528
rect 6542 13472 6598 13528
rect 6666 13472 6722 13528
rect 6790 13472 6846 13528
rect 6914 13472 6970 13528
rect 7038 13472 7094 13528
rect 5178 13348 5234 13404
rect 5302 13348 5358 13404
rect 5426 13348 5482 13404
rect 5550 13348 5606 13404
rect 5674 13348 5730 13404
rect 5798 13348 5854 13404
rect 5922 13348 5978 13404
rect 6046 13348 6102 13404
rect 6170 13348 6226 13404
rect 6294 13348 6350 13404
rect 6418 13348 6474 13404
rect 6542 13348 6598 13404
rect 6666 13348 6722 13404
rect 6790 13348 6846 13404
rect 6914 13348 6970 13404
rect 7038 13348 7094 13404
rect 5178 13224 5234 13280
rect 5302 13224 5358 13280
rect 5426 13224 5482 13280
rect 5550 13224 5606 13280
rect 5674 13224 5730 13280
rect 5798 13224 5854 13280
rect 5922 13224 5978 13280
rect 6046 13224 6102 13280
rect 6170 13224 6226 13280
rect 6294 13224 6350 13280
rect 6418 13224 6474 13280
rect 6542 13224 6598 13280
rect 6666 13224 6722 13280
rect 6790 13224 6846 13280
rect 6914 13224 6970 13280
rect 7038 13224 7094 13280
rect 5178 13100 5234 13156
rect 5302 13100 5358 13156
rect 5426 13100 5482 13156
rect 5550 13100 5606 13156
rect 5674 13100 5730 13156
rect 5798 13100 5854 13156
rect 5922 13100 5978 13156
rect 6046 13100 6102 13156
rect 6170 13100 6226 13156
rect 6294 13100 6350 13156
rect 6418 13100 6474 13156
rect 6542 13100 6598 13156
rect 6666 13100 6722 13156
rect 6790 13100 6846 13156
rect 6914 13100 6970 13156
rect 7038 13100 7094 13156
rect 5178 12976 5234 13032
rect 5302 12976 5358 13032
rect 5426 12976 5482 13032
rect 5550 12976 5606 13032
rect 5674 12976 5730 13032
rect 5798 12976 5854 13032
rect 5922 12976 5978 13032
rect 6046 12976 6102 13032
rect 6170 12976 6226 13032
rect 6294 12976 6350 13032
rect 6418 12976 6474 13032
rect 6542 12976 6598 13032
rect 6666 12976 6722 13032
rect 6790 12976 6846 13032
rect 6914 12976 6970 13032
rect 7038 12976 7094 13032
rect 5178 12852 5234 12908
rect 5302 12852 5358 12908
rect 5426 12852 5482 12908
rect 5550 12852 5606 12908
rect 5674 12852 5730 12908
rect 5798 12852 5854 12908
rect 5922 12852 5978 12908
rect 6046 12852 6102 12908
rect 6170 12852 6226 12908
rect 6294 12852 6350 12908
rect 6418 12852 6474 12908
rect 6542 12852 6598 12908
rect 6666 12852 6722 12908
rect 6790 12852 6846 12908
rect 6914 12852 6970 12908
rect 7038 12852 7094 12908
rect 7884 14092 7940 14148
rect 8008 14092 8064 14148
rect 8132 14092 8188 14148
rect 8256 14092 8312 14148
rect 8380 14092 8436 14148
rect 8504 14092 8560 14148
rect 8628 14092 8684 14148
rect 8752 14092 8808 14148
rect 8876 14092 8932 14148
rect 9000 14092 9056 14148
rect 9124 14092 9180 14148
rect 9248 14092 9304 14148
rect 9372 14092 9428 14148
rect 9496 14092 9552 14148
rect 9620 14092 9676 14148
rect 9744 14092 9800 14148
rect 7884 13968 7940 14024
rect 8008 13968 8064 14024
rect 8132 13968 8188 14024
rect 8256 13968 8312 14024
rect 8380 13968 8436 14024
rect 8504 13968 8560 14024
rect 8628 13968 8684 14024
rect 8752 13968 8808 14024
rect 8876 13968 8932 14024
rect 9000 13968 9056 14024
rect 9124 13968 9180 14024
rect 9248 13968 9304 14024
rect 9372 13968 9428 14024
rect 9496 13968 9552 14024
rect 9620 13968 9676 14024
rect 9744 13968 9800 14024
rect 7884 13844 7940 13900
rect 8008 13844 8064 13900
rect 8132 13844 8188 13900
rect 8256 13844 8312 13900
rect 8380 13844 8436 13900
rect 8504 13844 8560 13900
rect 8628 13844 8684 13900
rect 8752 13844 8808 13900
rect 8876 13844 8932 13900
rect 9000 13844 9056 13900
rect 9124 13844 9180 13900
rect 9248 13844 9304 13900
rect 9372 13844 9428 13900
rect 9496 13844 9552 13900
rect 9620 13844 9676 13900
rect 9744 13844 9800 13900
rect 7884 13720 7940 13776
rect 8008 13720 8064 13776
rect 8132 13720 8188 13776
rect 8256 13720 8312 13776
rect 8380 13720 8436 13776
rect 8504 13720 8560 13776
rect 8628 13720 8684 13776
rect 8752 13720 8808 13776
rect 8876 13720 8932 13776
rect 9000 13720 9056 13776
rect 9124 13720 9180 13776
rect 9248 13720 9304 13776
rect 9372 13720 9428 13776
rect 9496 13720 9552 13776
rect 9620 13720 9676 13776
rect 9744 13720 9800 13776
rect 7884 13596 7940 13652
rect 8008 13596 8064 13652
rect 8132 13596 8188 13652
rect 8256 13596 8312 13652
rect 8380 13596 8436 13652
rect 8504 13596 8560 13652
rect 8628 13596 8684 13652
rect 8752 13596 8808 13652
rect 8876 13596 8932 13652
rect 9000 13596 9056 13652
rect 9124 13596 9180 13652
rect 9248 13596 9304 13652
rect 9372 13596 9428 13652
rect 9496 13596 9552 13652
rect 9620 13596 9676 13652
rect 9744 13596 9800 13652
rect 7884 13472 7940 13528
rect 8008 13472 8064 13528
rect 8132 13472 8188 13528
rect 8256 13472 8312 13528
rect 8380 13472 8436 13528
rect 8504 13472 8560 13528
rect 8628 13472 8684 13528
rect 8752 13472 8808 13528
rect 8876 13472 8932 13528
rect 9000 13472 9056 13528
rect 9124 13472 9180 13528
rect 9248 13472 9304 13528
rect 9372 13472 9428 13528
rect 9496 13472 9552 13528
rect 9620 13472 9676 13528
rect 9744 13472 9800 13528
rect 7884 13348 7940 13404
rect 8008 13348 8064 13404
rect 8132 13348 8188 13404
rect 8256 13348 8312 13404
rect 8380 13348 8436 13404
rect 8504 13348 8560 13404
rect 8628 13348 8684 13404
rect 8752 13348 8808 13404
rect 8876 13348 8932 13404
rect 9000 13348 9056 13404
rect 9124 13348 9180 13404
rect 9248 13348 9304 13404
rect 9372 13348 9428 13404
rect 9496 13348 9552 13404
rect 9620 13348 9676 13404
rect 9744 13348 9800 13404
rect 7884 13224 7940 13280
rect 8008 13224 8064 13280
rect 8132 13224 8188 13280
rect 8256 13224 8312 13280
rect 8380 13224 8436 13280
rect 8504 13224 8560 13280
rect 8628 13224 8684 13280
rect 8752 13224 8808 13280
rect 8876 13224 8932 13280
rect 9000 13224 9056 13280
rect 9124 13224 9180 13280
rect 9248 13224 9304 13280
rect 9372 13224 9428 13280
rect 9496 13224 9552 13280
rect 9620 13224 9676 13280
rect 9744 13224 9800 13280
rect 7884 13100 7940 13156
rect 8008 13100 8064 13156
rect 8132 13100 8188 13156
rect 8256 13100 8312 13156
rect 8380 13100 8436 13156
rect 8504 13100 8560 13156
rect 8628 13100 8684 13156
rect 8752 13100 8808 13156
rect 8876 13100 8932 13156
rect 9000 13100 9056 13156
rect 9124 13100 9180 13156
rect 9248 13100 9304 13156
rect 9372 13100 9428 13156
rect 9496 13100 9552 13156
rect 9620 13100 9676 13156
rect 9744 13100 9800 13156
rect 7884 12976 7940 13032
rect 8008 12976 8064 13032
rect 8132 12976 8188 13032
rect 8256 12976 8312 13032
rect 8380 12976 8436 13032
rect 8504 12976 8560 13032
rect 8628 12976 8684 13032
rect 8752 12976 8808 13032
rect 8876 12976 8932 13032
rect 9000 12976 9056 13032
rect 9124 12976 9180 13032
rect 9248 12976 9304 13032
rect 9372 12976 9428 13032
rect 9496 12976 9552 13032
rect 9620 12976 9676 13032
rect 9744 12976 9800 13032
rect 7884 12852 7940 12908
rect 8008 12852 8064 12908
rect 8132 12852 8188 12908
rect 8256 12852 8312 12908
rect 8380 12852 8436 12908
rect 8504 12852 8560 12908
rect 8628 12852 8684 12908
rect 8752 12852 8808 12908
rect 8876 12852 8932 12908
rect 9000 12852 9056 12908
rect 9124 12852 9180 12908
rect 9248 12852 9304 12908
rect 9372 12852 9428 12908
rect 9496 12852 9552 12908
rect 9620 12852 9676 12908
rect 9744 12852 9800 12908
rect 10254 14092 10310 14148
rect 10378 14092 10434 14148
rect 10502 14092 10558 14148
rect 10626 14092 10682 14148
rect 10750 14092 10806 14148
rect 10874 14092 10930 14148
rect 10998 14092 11054 14148
rect 11122 14092 11178 14148
rect 11246 14092 11302 14148
rect 11370 14092 11426 14148
rect 11494 14092 11550 14148
rect 11618 14092 11674 14148
rect 11742 14092 11798 14148
rect 11866 14092 11922 14148
rect 11990 14092 12046 14148
rect 12114 14092 12170 14148
rect 10254 13968 10310 14024
rect 10378 13968 10434 14024
rect 10502 13968 10558 14024
rect 10626 13968 10682 14024
rect 10750 13968 10806 14024
rect 10874 13968 10930 14024
rect 10998 13968 11054 14024
rect 11122 13968 11178 14024
rect 11246 13968 11302 14024
rect 11370 13968 11426 14024
rect 11494 13968 11550 14024
rect 11618 13968 11674 14024
rect 11742 13968 11798 14024
rect 11866 13968 11922 14024
rect 11990 13968 12046 14024
rect 12114 13968 12170 14024
rect 10254 13844 10310 13900
rect 10378 13844 10434 13900
rect 10502 13844 10558 13900
rect 10626 13844 10682 13900
rect 10750 13844 10806 13900
rect 10874 13844 10930 13900
rect 10998 13844 11054 13900
rect 11122 13844 11178 13900
rect 11246 13844 11302 13900
rect 11370 13844 11426 13900
rect 11494 13844 11550 13900
rect 11618 13844 11674 13900
rect 11742 13844 11798 13900
rect 11866 13844 11922 13900
rect 11990 13844 12046 13900
rect 12114 13844 12170 13900
rect 10254 13720 10310 13776
rect 10378 13720 10434 13776
rect 10502 13720 10558 13776
rect 10626 13720 10682 13776
rect 10750 13720 10806 13776
rect 10874 13720 10930 13776
rect 10998 13720 11054 13776
rect 11122 13720 11178 13776
rect 11246 13720 11302 13776
rect 11370 13720 11426 13776
rect 11494 13720 11550 13776
rect 11618 13720 11674 13776
rect 11742 13720 11798 13776
rect 11866 13720 11922 13776
rect 11990 13720 12046 13776
rect 12114 13720 12170 13776
rect 10254 13596 10310 13652
rect 10378 13596 10434 13652
rect 10502 13596 10558 13652
rect 10626 13596 10682 13652
rect 10750 13596 10806 13652
rect 10874 13596 10930 13652
rect 10998 13596 11054 13652
rect 11122 13596 11178 13652
rect 11246 13596 11302 13652
rect 11370 13596 11426 13652
rect 11494 13596 11550 13652
rect 11618 13596 11674 13652
rect 11742 13596 11798 13652
rect 11866 13596 11922 13652
rect 11990 13596 12046 13652
rect 12114 13596 12170 13652
rect 10254 13472 10310 13528
rect 10378 13472 10434 13528
rect 10502 13472 10558 13528
rect 10626 13472 10682 13528
rect 10750 13472 10806 13528
rect 10874 13472 10930 13528
rect 10998 13472 11054 13528
rect 11122 13472 11178 13528
rect 11246 13472 11302 13528
rect 11370 13472 11426 13528
rect 11494 13472 11550 13528
rect 11618 13472 11674 13528
rect 11742 13472 11798 13528
rect 11866 13472 11922 13528
rect 11990 13472 12046 13528
rect 12114 13472 12170 13528
rect 10254 13348 10310 13404
rect 10378 13348 10434 13404
rect 10502 13348 10558 13404
rect 10626 13348 10682 13404
rect 10750 13348 10806 13404
rect 10874 13348 10930 13404
rect 10998 13348 11054 13404
rect 11122 13348 11178 13404
rect 11246 13348 11302 13404
rect 11370 13348 11426 13404
rect 11494 13348 11550 13404
rect 11618 13348 11674 13404
rect 11742 13348 11798 13404
rect 11866 13348 11922 13404
rect 11990 13348 12046 13404
rect 12114 13348 12170 13404
rect 10254 13224 10310 13280
rect 10378 13224 10434 13280
rect 10502 13224 10558 13280
rect 10626 13224 10682 13280
rect 10750 13224 10806 13280
rect 10874 13224 10930 13280
rect 10998 13224 11054 13280
rect 11122 13224 11178 13280
rect 11246 13224 11302 13280
rect 11370 13224 11426 13280
rect 11494 13224 11550 13280
rect 11618 13224 11674 13280
rect 11742 13224 11798 13280
rect 11866 13224 11922 13280
rect 11990 13224 12046 13280
rect 12114 13224 12170 13280
rect 10254 13100 10310 13156
rect 10378 13100 10434 13156
rect 10502 13100 10558 13156
rect 10626 13100 10682 13156
rect 10750 13100 10806 13156
rect 10874 13100 10930 13156
rect 10998 13100 11054 13156
rect 11122 13100 11178 13156
rect 11246 13100 11302 13156
rect 11370 13100 11426 13156
rect 11494 13100 11550 13156
rect 11618 13100 11674 13156
rect 11742 13100 11798 13156
rect 11866 13100 11922 13156
rect 11990 13100 12046 13156
rect 12114 13100 12170 13156
rect 10254 12976 10310 13032
rect 10378 12976 10434 13032
rect 10502 12976 10558 13032
rect 10626 12976 10682 13032
rect 10750 12976 10806 13032
rect 10874 12976 10930 13032
rect 10998 12976 11054 13032
rect 11122 12976 11178 13032
rect 11246 12976 11302 13032
rect 11370 12976 11426 13032
rect 11494 12976 11550 13032
rect 11618 12976 11674 13032
rect 11742 12976 11798 13032
rect 11866 12976 11922 13032
rect 11990 12976 12046 13032
rect 12114 12976 12170 13032
rect 10254 12852 10310 12908
rect 10378 12852 10434 12908
rect 10502 12852 10558 12908
rect 10626 12852 10682 12908
rect 10750 12852 10806 12908
rect 10874 12852 10930 12908
rect 10998 12852 11054 12908
rect 11122 12852 11178 12908
rect 11246 12852 11302 12908
rect 11370 12852 11426 12908
rect 11494 12852 11550 12908
rect 11618 12852 11674 12908
rect 11742 12852 11798 12908
rect 11866 12852 11922 12908
rect 11990 12852 12046 12908
rect 12114 12852 12170 12908
rect 12871 14092 12927 14148
rect 12995 14092 13051 14148
rect 13119 14092 13175 14148
rect 13243 14092 13299 14148
rect 13367 14092 13423 14148
rect 13491 14092 13547 14148
rect 13615 14092 13671 14148
rect 13739 14092 13795 14148
rect 13863 14092 13919 14148
rect 13987 14092 14043 14148
rect 14111 14092 14167 14148
rect 14235 14092 14291 14148
rect 14359 14092 14415 14148
rect 14483 14092 14539 14148
rect 14607 14092 14663 14148
rect 12871 13968 12927 14024
rect 12995 13968 13051 14024
rect 13119 13968 13175 14024
rect 13243 13968 13299 14024
rect 13367 13968 13423 14024
rect 13491 13968 13547 14024
rect 13615 13968 13671 14024
rect 13739 13968 13795 14024
rect 13863 13968 13919 14024
rect 13987 13968 14043 14024
rect 14111 13968 14167 14024
rect 14235 13968 14291 14024
rect 14359 13968 14415 14024
rect 14483 13968 14539 14024
rect 14607 13968 14663 14024
rect 12871 13844 12927 13900
rect 12995 13844 13051 13900
rect 13119 13844 13175 13900
rect 13243 13844 13299 13900
rect 13367 13844 13423 13900
rect 13491 13844 13547 13900
rect 13615 13844 13671 13900
rect 13739 13844 13795 13900
rect 13863 13844 13919 13900
rect 13987 13844 14043 13900
rect 14111 13844 14167 13900
rect 14235 13844 14291 13900
rect 14359 13844 14415 13900
rect 14483 13844 14539 13900
rect 14607 13844 14663 13900
rect 12871 13720 12927 13776
rect 12995 13720 13051 13776
rect 13119 13720 13175 13776
rect 13243 13720 13299 13776
rect 13367 13720 13423 13776
rect 13491 13720 13547 13776
rect 13615 13720 13671 13776
rect 13739 13720 13795 13776
rect 13863 13720 13919 13776
rect 13987 13720 14043 13776
rect 14111 13720 14167 13776
rect 14235 13720 14291 13776
rect 14359 13720 14415 13776
rect 14483 13720 14539 13776
rect 14607 13720 14663 13776
rect 12871 13596 12927 13652
rect 12995 13596 13051 13652
rect 13119 13596 13175 13652
rect 13243 13596 13299 13652
rect 13367 13596 13423 13652
rect 13491 13596 13547 13652
rect 13615 13596 13671 13652
rect 13739 13596 13795 13652
rect 13863 13596 13919 13652
rect 13987 13596 14043 13652
rect 14111 13596 14167 13652
rect 14235 13596 14291 13652
rect 14359 13596 14415 13652
rect 14483 13596 14539 13652
rect 14607 13596 14663 13652
rect 12871 13472 12927 13528
rect 12995 13472 13051 13528
rect 13119 13472 13175 13528
rect 13243 13472 13299 13528
rect 13367 13472 13423 13528
rect 13491 13472 13547 13528
rect 13615 13472 13671 13528
rect 13739 13472 13795 13528
rect 13863 13472 13919 13528
rect 13987 13472 14043 13528
rect 14111 13472 14167 13528
rect 14235 13472 14291 13528
rect 14359 13472 14415 13528
rect 14483 13472 14539 13528
rect 14607 13472 14663 13528
rect 12871 13348 12927 13404
rect 12995 13348 13051 13404
rect 13119 13348 13175 13404
rect 13243 13348 13299 13404
rect 13367 13348 13423 13404
rect 13491 13348 13547 13404
rect 13615 13348 13671 13404
rect 13739 13348 13795 13404
rect 13863 13348 13919 13404
rect 13987 13348 14043 13404
rect 14111 13348 14167 13404
rect 14235 13348 14291 13404
rect 14359 13348 14415 13404
rect 14483 13348 14539 13404
rect 14607 13348 14663 13404
rect 12871 13224 12927 13280
rect 12995 13224 13051 13280
rect 13119 13224 13175 13280
rect 13243 13224 13299 13280
rect 13367 13224 13423 13280
rect 13491 13224 13547 13280
rect 13615 13224 13671 13280
rect 13739 13224 13795 13280
rect 13863 13224 13919 13280
rect 13987 13224 14043 13280
rect 14111 13224 14167 13280
rect 14235 13224 14291 13280
rect 14359 13224 14415 13280
rect 14483 13224 14539 13280
rect 14607 13224 14663 13280
rect 12871 13100 12927 13156
rect 12995 13100 13051 13156
rect 13119 13100 13175 13156
rect 13243 13100 13299 13156
rect 13367 13100 13423 13156
rect 13491 13100 13547 13156
rect 13615 13100 13671 13156
rect 13739 13100 13795 13156
rect 13863 13100 13919 13156
rect 13987 13100 14043 13156
rect 14111 13100 14167 13156
rect 14235 13100 14291 13156
rect 14359 13100 14415 13156
rect 14483 13100 14539 13156
rect 14607 13100 14663 13156
rect 12871 12976 12927 13032
rect 12995 12976 13051 13032
rect 13119 12976 13175 13032
rect 13243 12976 13299 13032
rect 13367 12976 13423 13032
rect 13491 12976 13547 13032
rect 13615 12976 13671 13032
rect 13739 12976 13795 13032
rect 13863 12976 13919 13032
rect 13987 12976 14043 13032
rect 14111 12976 14167 13032
rect 14235 12976 14291 13032
rect 14359 12976 14415 13032
rect 14483 12976 14539 13032
rect 14607 12976 14663 13032
rect 12871 12852 12927 12908
rect 12995 12852 13051 12908
rect 13119 12852 13175 12908
rect 13243 12852 13299 12908
rect 13367 12852 13423 12908
rect 13491 12852 13547 12908
rect 13615 12852 13671 12908
rect 13739 12852 13795 12908
rect 13863 12852 13919 12908
rect 13987 12852 14043 12908
rect 14111 12852 14167 12908
rect 14235 12852 14291 12908
rect 14359 12852 14415 12908
rect 14483 12852 14539 12908
rect 14607 12852 14663 12908
rect 14902 14174 14958 14176
rect 14902 14122 14904 14174
rect 14904 14122 14956 14174
rect 14956 14122 14958 14174
rect 14902 14066 14958 14122
rect 14902 14014 14904 14066
rect 14904 14014 14956 14066
rect 14956 14014 14958 14066
rect 14902 13958 14958 14014
rect 14902 13906 14904 13958
rect 14904 13906 14956 13958
rect 14956 13906 14958 13958
rect 14902 13850 14958 13906
rect 14902 13798 14904 13850
rect 14904 13798 14956 13850
rect 14956 13798 14958 13850
rect 14902 13742 14958 13798
rect 14902 13690 14904 13742
rect 14904 13690 14956 13742
rect 14956 13690 14958 13742
rect 14902 13634 14958 13690
rect 14902 13582 14904 13634
rect 14904 13582 14956 13634
rect 14956 13582 14958 13634
rect 14902 13526 14958 13582
rect 14902 13474 14904 13526
rect 14904 13474 14956 13526
rect 14956 13474 14958 13526
rect 14902 13418 14958 13474
rect 14902 13366 14904 13418
rect 14904 13366 14956 13418
rect 14956 13366 14958 13418
rect 14902 13310 14958 13366
rect 14902 13258 14904 13310
rect 14904 13258 14956 13310
rect 14956 13258 14958 13310
rect 14902 13202 14958 13258
rect 14902 13150 14904 13202
rect 14904 13150 14956 13202
rect 14956 13150 14958 13202
rect 14902 13094 14958 13150
rect 14902 13042 14904 13094
rect 14904 13042 14956 13094
rect 14956 13042 14958 13094
rect 14902 12986 14958 13042
rect 14902 12934 14904 12986
rect 14904 12934 14956 12986
rect 14956 12934 14958 12986
rect 14902 12878 14958 12934
rect 14902 12826 14904 12878
rect 14904 12826 14956 12878
rect 14956 12826 14958 12878
rect 14902 12824 14958 12826
rect 2491 12492 2547 12548
rect 2615 12492 2671 12548
rect 2491 12368 2547 12424
rect 2615 12368 2671 12424
rect 2491 12244 2547 12300
rect 2615 12244 2671 12300
rect 2491 12120 2547 12176
rect 2615 12120 2671 12176
rect 2491 11996 2547 12052
rect 2615 11996 2671 12052
rect 2491 11872 2547 11928
rect 2615 11872 2671 11928
rect 2491 11748 2547 11804
rect 2615 11748 2671 11804
rect 2491 11624 2547 11680
rect 2615 11624 2671 11680
rect 2491 11500 2547 11556
rect 2615 11500 2671 11556
rect 2491 11376 2547 11432
rect 2615 11376 2671 11432
rect 2491 11252 2547 11308
rect 2615 11252 2671 11308
rect 4861 12492 4917 12548
rect 4985 12492 5041 12548
rect 4861 12368 4917 12424
rect 4985 12368 5041 12424
rect 4861 12244 4917 12300
rect 4985 12244 5041 12300
rect 4861 12120 4917 12176
rect 4985 12120 5041 12176
rect 4861 11996 4917 12052
rect 4985 11996 5041 12052
rect 4861 11872 4917 11928
rect 4985 11872 5041 11928
rect 4861 11748 4917 11804
rect 4985 11748 5041 11804
rect 4861 11624 4917 11680
rect 4985 11624 5041 11680
rect 4861 11500 4917 11556
rect 4985 11500 5041 11556
rect 4861 11376 4917 11432
rect 4985 11376 5041 11432
rect 4861 11252 4917 11308
rect 4985 11252 5041 11308
rect 7275 12492 7331 12548
rect 7399 12492 7455 12548
rect 7523 12492 7579 12548
rect 7647 12492 7703 12548
rect 7275 12368 7331 12424
rect 7399 12368 7455 12424
rect 7523 12368 7579 12424
rect 7647 12368 7703 12424
rect 7275 12244 7331 12300
rect 7399 12244 7455 12300
rect 7523 12244 7579 12300
rect 7647 12244 7703 12300
rect 7275 12120 7331 12176
rect 7399 12120 7455 12176
rect 7523 12120 7579 12176
rect 7647 12120 7703 12176
rect 7275 11996 7331 12052
rect 7399 11996 7455 12052
rect 7523 11996 7579 12052
rect 7647 11996 7703 12052
rect 7275 11872 7331 11928
rect 7399 11872 7455 11928
rect 7523 11872 7579 11928
rect 7647 11872 7703 11928
rect 7275 11748 7331 11804
rect 7399 11748 7455 11804
rect 7523 11748 7579 11804
rect 7647 11748 7703 11804
rect 7275 11624 7331 11680
rect 7399 11624 7455 11680
rect 7523 11624 7579 11680
rect 7647 11624 7703 11680
rect 7275 11500 7331 11556
rect 7399 11500 7455 11556
rect 7523 11500 7579 11556
rect 7647 11500 7703 11556
rect 7275 11376 7331 11432
rect 7399 11376 7455 11432
rect 7523 11376 7579 11432
rect 7647 11376 7703 11432
rect 7275 11252 7331 11308
rect 7399 11252 7455 11308
rect 7523 11252 7579 11308
rect 7647 11252 7703 11308
rect 9937 12492 9993 12548
rect 10061 12492 10117 12548
rect 9937 12368 9993 12424
rect 10061 12368 10117 12424
rect 9937 12244 9993 12300
rect 10061 12244 10117 12300
rect 9937 12120 9993 12176
rect 10061 12120 10117 12176
rect 9937 11996 9993 12052
rect 10061 11996 10117 12052
rect 9937 11872 9993 11928
rect 10061 11872 10117 11928
rect 9937 11748 9993 11804
rect 10061 11748 10117 11804
rect 9937 11624 9993 11680
rect 10061 11624 10117 11680
rect 9937 11500 9993 11556
rect 10061 11500 10117 11556
rect 9937 11376 9993 11432
rect 10061 11376 10117 11432
rect 9937 11252 9993 11308
rect 10061 11252 10117 11308
rect 12307 12492 12363 12548
rect 12431 12492 12487 12548
rect 12307 12368 12363 12424
rect 12431 12368 12487 12424
rect 12307 12244 12363 12300
rect 12431 12244 12487 12300
rect 12307 12120 12363 12176
rect 12431 12120 12487 12176
rect 12307 11996 12363 12052
rect 12431 11996 12487 12052
rect 12307 11872 12363 11928
rect 12431 11872 12487 11928
rect 12307 11748 12363 11804
rect 12431 11748 12487 11804
rect 12307 11624 12363 11680
rect 12431 11624 12487 11680
rect 12307 11500 12363 11556
rect 12431 11500 12487 11556
rect 12307 11376 12363 11432
rect 12431 11376 12487 11432
rect 12307 11252 12363 11308
rect 12431 11252 12487 11308
rect 20 10984 76 10986
rect 20 10932 22 10984
rect 22 10932 74 10984
rect 74 10932 76 10984
rect 20 10876 76 10932
rect 20 10824 22 10876
rect 22 10824 74 10876
rect 74 10824 76 10876
rect 20 10768 76 10824
rect 20 10716 22 10768
rect 22 10716 74 10768
rect 74 10716 76 10768
rect 20 10660 76 10716
rect 20 10608 22 10660
rect 22 10608 74 10660
rect 74 10608 76 10660
rect 20 10552 76 10608
rect 20 10500 22 10552
rect 22 10500 74 10552
rect 74 10500 76 10552
rect 20 10444 76 10500
rect 20 10392 22 10444
rect 22 10392 74 10444
rect 74 10392 76 10444
rect 20 10336 76 10392
rect 20 10284 22 10336
rect 22 10284 74 10336
rect 74 10284 76 10336
rect 20 10228 76 10284
rect 20 10176 22 10228
rect 22 10176 74 10228
rect 74 10176 76 10228
rect 20 10120 76 10176
rect 20 10068 22 10120
rect 22 10068 74 10120
rect 74 10068 76 10120
rect 20 10012 76 10068
rect 20 9960 22 10012
rect 22 9960 74 10012
rect 74 9960 76 10012
rect 20 9904 76 9960
rect 20 9852 22 9904
rect 22 9852 74 9904
rect 74 9852 76 9904
rect 20 9796 76 9852
rect 20 9744 22 9796
rect 22 9744 74 9796
rect 74 9744 76 9796
rect 20 9688 76 9744
rect 20 9636 22 9688
rect 22 9636 74 9688
rect 74 9636 76 9688
rect 20 9580 76 9636
rect 20 9528 22 9580
rect 22 9528 74 9580
rect 74 9528 76 9580
rect 20 9472 76 9528
rect 20 9420 22 9472
rect 22 9420 74 9472
rect 74 9420 76 9472
rect 20 9364 76 9420
rect 20 9312 22 9364
rect 22 9312 74 9364
rect 74 9312 76 9364
rect 20 9256 76 9312
rect 20 9204 22 9256
rect 22 9204 74 9256
rect 74 9204 76 9256
rect 20 9148 76 9204
rect 20 9096 22 9148
rect 22 9096 74 9148
rect 74 9096 76 9148
rect 20 9040 76 9096
rect 20 8988 22 9040
rect 22 8988 74 9040
rect 74 8988 76 9040
rect 20 8932 76 8988
rect 20 8880 22 8932
rect 22 8880 74 8932
rect 74 8880 76 8932
rect 20 8824 76 8880
rect 20 8772 22 8824
rect 22 8772 74 8824
rect 74 8772 76 8824
rect 20 8716 76 8772
rect 20 8664 22 8716
rect 22 8664 74 8716
rect 74 8664 76 8716
rect 20 8608 76 8664
rect 20 8556 22 8608
rect 22 8556 74 8608
rect 74 8556 76 8608
rect 20 8500 76 8556
rect 20 8448 22 8500
rect 22 8448 74 8500
rect 74 8448 76 8500
rect 20 8392 76 8448
rect 20 8340 22 8392
rect 22 8340 74 8392
rect 74 8340 76 8392
rect 20 8284 76 8340
rect 20 8232 22 8284
rect 22 8232 74 8284
rect 74 8232 76 8284
rect 20 8176 76 8232
rect 20 8124 22 8176
rect 22 8124 74 8176
rect 74 8124 76 8176
rect 20 8068 76 8124
rect 20 8016 22 8068
rect 22 8016 74 8068
rect 74 8016 76 8068
rect 20 8014 76 8016
rect 315 10898 371 10954
rect 439 10898 495 10954
rect 563 10898 619 10954
rect 687 10898 743 10954
rect 811 10898 867 10954
rect 935 10898 991 10954
rect 1059 10898 1115 10954
rect 1183 10898 1239 10954
rect 1307 10898 1363 10954
rect 1431 10898 1487 10954
rect 1555 10898 1611 10954
rect 1679 10898 1735 10954
rect 1803 10898 1859 10954
rect 1927 10898 1983 10954
rect 2051 10898 2107 10954
rect 315 10774 371 10830
rect 439 10774 495 10830
rect 563 10774 619 10830
rect 687 10774 743 10830
rect 811 10774 867 10830
rect 935 10774 991 10830
rect 1059 10774 1115 10830
rect 1183 10774 1239 10830
rect 1307 10774 1363 10830
rect 1431 10774 1487 10830
rect 1555 10774 1611 10830
rect 1679 10774 1735 10830
rect 1803 10774 1859 10830
rect 1927 10774 1983 10830
rect 2051 10774 2107 10830
rect 315 10650 371 10706
rect 439 10650 495 10706
rect 563 10650 619 10706
rect 687 10650 743 10706
rect 811 10650 867 10706
rect 935 10650 991 10706
rect 1059 10650 1115 10706
rect 1183 10650 1239 10706
rect 1307 10650 1363 10706
rect 1431 10650 1487 10706
rect 1555 10650 1611 10706
rect 1679 10650 1735 10706
rect 1803 10650 1859 10706
rect 1927 10650 1983 10706
rect 2051 10650 2107 10706
rect 315 10526 371 10582
rect 439 10526 495 10582
rect 563 10526 619 10582
rect 687 10526 743 10582
rect 811 10526 867 10582
rect 935 10526 991 10582
rect 1059 10526 1115 10582
rect 1183 10526 1239 10582
rect 1307 10526 1363 10582
rect 1431 10526 1487 10582
rect 1555 10526 1611 10582
rect 1679 10526 1735 10582
rect 1803 10526 1859 10582
rect 1927 10526 1983 10582
rect 2051 10526 2107 10582
rect 315 10402 371 10458
rect 439 10402 495 10458
rect 563 10402 619 10458
rect 687 10402 743 10458
rect 811 10402 867 10458
rect 935 10402 991 10458
rect 1059 10402 1115 10458
rect 1183 10402 1239 10458
rect 1307 10402 1363 10458
rect 1431 10402 1487 10458
rect 1555 10402 1611 10458
rect 1679 10402 1735 10458
rect 1803 10402 1859 10458
rect 1927 10402 1983 10458
rect 2051 10402 2107 10458
rect 315 10278 371 10334
rect 439 10278 495 10334
rect 563 10278 619 10334
rect 687 10278 743 10334
rect 811 10278 867 10334
rect 935 10278 991 10334
rect 1059 10278 1115 10334
rect 1183 10278 1239 10334
rect 1307 10278 1363 10334
rect 1431 10278 1487 10334
rect 1555 10278 1611 10334
rect 1679 10278 1735 10334
rect 1803 10278 1859 10334
rect 1927 10278 1983 10334
rect 2051 10278 2107 10334
rect 315 10154 371 10210
rect 439 10154 495 10210
rect 563 10154 619 10210
rect 687 10154 743 10210
rect 811 10154 867 10210
rect 935 10154 991 10210
rect 1059 10154 1115 10210
rect 1183 10154 1239 10210
rect 1307 10154 1363 10210
rect 1431 10154 1487 10210
rect 1555 10154 1611 10210
rect 1679 10154 1735 10210
rect 1803 10154 1859 10210
rect 1927 10154 1983 10210
rect 2051 10154 2107 10210
rect 315 10030 371 10086
rect 439 10030 495 10086
rect 563 10030 619 10086
rect 687 10030 743 10086
rect 811 10030 867 10086
rect 935 10030 991 10086
rect 1059 10030 1115 10086
rect 1183 10030 1239 10086
rect 1307 10030 1363 10086
rect 1431 10030 1487 10086
rect 1555 10030 1611 10086
rect 1679 10030 1735 10086
rect 1803 10030 1859 10086
rect 1927 10030 1983 10086
rect 2051 10030 2107 10086
rect 315 9906 371 9962
rect 439 9906 495 9962
rect 563 9906 619 9962
rect 687 9906 743 9962
rect 811 9906 867 9962
rect 935 9906 991 9962
rect 1059 9906 1115 9962
rect 1183 9906 1239 9962
rect 1307 9906 1363 9962
rect 1431 9906 1487 9962
rect 1555 9906 1611 9962
rect 1679 9906 1735 9962
rect 1803 9906 1859 9962
rect 1927 9906 1983 9962
rect 2051 9906 2107 9962
rect 315 9782 371 9838
rect 439 9782 495 9838
rect 563 9782 619 9838
rect 687 9782 743 9838
rect 811 9782 867 9838
rect 935 9782 991 9838
rect 1059 9782 1115 9838
rect 1183 9782 1239 9838
rect 1307 9782 1363 9838
rect 1431 9782 1487 9838
rect 1555 9782 1611 9838
rect 1679 9782 1735 9838
rect 1803 9782 1859 9838
rect 1927 9782 1983 9838
rect 2051 9782 2107 9838
rect 315 9658 371 9714
rect 439 9658 495 9714
rect 563 9658 619 9714
rect 687 9658 743 9714
rect 811 9658 867 9714
rect 935 9658 991 9714
rect 1059 9658 1115 9714
rect 1183 9658 1239 9714
rect 1307 9658 1363 9714
rect 1431 9658 1487 9714
rect 1555 9658 1611 9714
rect 1679 9658 1735 9714
rect 1803 9658 1859 9714
rect 1927 9658 1983 9714
rect 2051 9658 2107 9714
rect 315 9534 371 9590
rect 439 9534 495 9590
rect 563 9534 619 9590
rect 687 9534 743 9590
rect 811 9534 867 9590
rect 935 9534 991 9590
rect 1059 9534 1115 9590
rect 1183 9534 1239 9590
rect 1307 9534 1363 9590
rect 1431 9534 1487 9590
rect 1555 9534 1611 9590
rect 1679 9534 1735 9590
rect 1803 9534 1859 9590
rect 1927 9534 1983 9590
rect 2051 9534 2107 9590
rect 315 9410 371 9466
rect 439 9410 495 9466
rect 563 9410 619 9466
rect 687 9410 743 9466
rect 811 9410 867 9466
rect 935 9410 991 9466
rect 1059 9410 1115 9466
rect 1183 9410 1239 9466
rect 1307 9410 1363 9466
rect 1431 9410 1487 9466
rect 1555 9410 1611 9466
rect 1679 9410 1735 9466
rect 1803 9410 1859 9466
rect 1927 9410 1983 9466
rect 2051 9410 2107 9466
rect 315 9286 371 9342
rect 439 9286 495 9342
rect 563 9286 619 9342
rect 687 9286 743 9342
rect 811 9286 867 9342
rect 935 9286 991 9342
rect 1059 9286 1115 9342
rect 1183 9286 1239 9342
rect 1307 9286 1363 9342
rect 1431 9286 1487 9342
rect 1555 9286 1611 9342
rect 1679 9286 1735 9342
rect 1803 9286 1859 9342
rect 1927 9286 1983 9342
rect 2051 9286 2107 9342
rect 315 9162 371 9218
rect 439 9162 495 9218
rect 563 9162 619 9218
rect 687 9162 743 9218
rect 811 9162 867 9218
rect 935 9162 991 9218
rect 1059 9162 1115 9218
rect 1183 9162 1239 9218
rect 1307 9162 1363 9218
rect 1431 9162 1487 9218
rect 1555 9162 1611 9218
rect 1679 9162 1735 9218
rect 1803 9162 1859 9218
rect 1927 9162 1983 9218
rect 2051 9162 2107 9218
rect 315 9038 371 9094
rect 439 9038 495 9094
rect 563 9038 619 9094
rect 687 9038 743 9094
rect 811 9038 867 9094
rect 935 9038 991 9094
rect 1059 9038 1115 9094
rect 1183 9038 1239 9094
rect 1307 9038 1363 9094
rect 1431 9038 1487 9094
rect 1555 9038 1611 9094
rect 1679 9038 1735 9094
rect 1803 9038 1859 9094
rect 1927 9038 1983 9094
rect 2051 9038 2107 9094
rect 315 8914 371 8970
rect 439 8914 495 8970
rect 563 8914 619 8970
rect 687 8914 743 8970
rect 811 8914 867 8970
rect 935 8914 991 8970
rect 1059 8914 1115 8970
rect 1183 8914 1239 8970
rect 1307 8914 1363 8970
rect 1431 8914 1487 8970
rect 1555 8914 1611 8970
rect 1679 8914 1735 8970
rect 1803 8914 1859 8970
rect 1927 8914 1983 8970
rect 2051 8914 2107 8970
rect 315 8790 371 8846
rect 439 8790 495 8846
rect 563 8790 619 8846
rect 687 8790 743 8846
rect 811 8790 867 8846
rect 935 8790 991 8846
rect 1059 8790 1115 8846
rect 1183 8790 1239 8846
rect 1307 8790 1363 8846
rect 1431 8790 1487 8846
rect 1555 8790 1611 8846
rect 1679 8790 1735 8846
rect 1803 8790 1859 8846
rect 1927 8790 1983 8846
rect 2051 8790 2107 8846
rect 315 8666 371 8722
rect 439 8666 495 8722
rect 563 8666 619 8722
rect 687 8666 743 8722
rect 811 8666 867 8722
rect 935 8666 991 8722
rect 1059 8666 1115 8722
rect 1183 8666 1239 8722
rect 1307 8666 1363 8722
rect 1431 8666 1487 8722
rect 1555 8666 1611 8722
rect 1679 8666 1735 8722
rect 1803 8666 1859 8722
rect 1927 8666 1983 8722
rect 2051 8666 2107 8722
rect 315 8542 371 8598
rect 439 8542 495 8598
rect 563 8542 619 8598
rect 687 8542 743 8598
rect 811 8542 867 8598
rect 935 8542 991 8598
rect 1059 8542 1115 8598
rect 1183 8542 1239 8598
rect 1307 8542 1363 8598
rect 1431 8542 1487 8598
rect 1555 8542 1611 8598
rect 1679 8542 1735 8598
rect 1803 8542 1859 8598
rect 1927 8542 1983 8598
rect 2051 8542 2107 8598
rect 315 8418 371 8474
rect 439 8418 495 8474
rect 563 8418 619 8474
rect 687 8418 743 8474
rect 811 8418 867 8474
rect 935 8418 991 8474
rect 1059 8418 1115 8474
rect 1183 8418 1239 8474
rect 1307 8418 1363 8474
rect 1431 8418 1487 8474
rect 1555 8418 1611 8474
rect 1679 8418 1735 8474
rect 1803 8418 1859 8474
rect 1927 8418 1983 8474
rect 2051 8418 2107 8474
rect 315 8294 371 8350
rect 439 8294 495 8350
rect 563 8294 619 8350
rect 687 8294 743 8350
rect 811 8294 867 8350
rect 935 8294 991 8350
rect 1059 8294 1115 8350
rect 1183 8294 1239 8350
rect 1307 8294 1363 8350
rect 1431 8294 1487 8350
rect 1555 8294 1611 8350
rect 1679 8294 1735 8350
rect 1803 8294 1859 8350
rect 1927 8294 1983 8350
rect 2051 8294 2107 8350
rect 315 8170 371 8226
rect 439 8170 495 8226
rect 563 8170 619 8226
rect 687 8170 743 8226
rect 811 8170 867 8226
rect 935 8170 991 8226
rect 1059 8170 1115 8226
rect 1183 8170 1239 8226
rect 1307 8170 1363 8226
rect 1431 8170 1487 8226
rect 1555 8170 1611 8226
rect 1679 8170 1735 8226
rect 1803 8170 1859 8226
rect 1927 8170 1983 8226
rect 2051 8170 2107 8226
rect 315 8046 371 8102
rect 439 8046 495 8102
rect 563 8046 619 8102
rect 687 8046 743 8102
rect 811 8046 867 8102
rect 935 8046 991 8102
rect 1059 8046 1115 8102
rect 1183 8046 1239 8102
rect 1307 8046 1363 8102
rect 1431 8046 1487 8102
rect 1555 8046 1611 8102
rect 1679 8046 1735 8102
rect 1803 8046 1859 8102
rect 1927 8046 1983 8102
rect 2051 8046 2107 8102
rect 2808 10898 2864 10954
rect 2932 10898 2988 10954
rect 3056 10898 3112 10954
rect 3180 10898 3236 10954
rect 3304 10898 3360 10954
rect 3428 10898 3484 10954
rect 3552 10898 3608 10954
rect 3676 10898 3732 10954
rect 3800 10898 3856 10954
rect 3924 10898 3980 10954
rect 4048 10898 4104 10954
rect 4172 10898 4228 10954
rect 4296 10898 4352 10954
rect 4420 10898 4476 10954
rect 4544 10898 4600 10954
rect 4668 10898 4724 10954
rect 2808 10774 2864 10830
rect 2932 10774 2988 10830
rect 3056 10774 3112 10830
rect 3180 10774 3236 10830
rect 3304 10774 3360 10830
rect 3428 10774 3484 10830
rect 3552 10774 3608 10830
rect 3676 10774 3732 10830
rect 3800 10774 3856 10830
rect 3924 10774 3980 10830
rect 4048 10774 4104 10830
rect 4172 10774 4228 10830
rect 4296 10774 4352 10830
rect 4420 10774 4476 10830
rect 4544 10774 4600 10830
rect 4668 10774 4724 10830
rect 2808 10650 2864 10706
rect 2932 10650 2988 10706
rect 3056 10650 3112 10706
rect 3180 10650 3236 10706
rect 3304 10650 3360 10706
rect 3428 10650 3484 10706
rect 3552 10650 3608 10706
rect 3676 10650 3732 10706
rect 3800 10650 3856 10706
rect 3924 10650 3980 10706
rect 4048 10650 4104 10706
rect 4172 10650 4228 10706
rect 4296 10650 4352 10706
rect 4420 10650 4476 10706
rect 4544 10650 4600 10706
rect 4668 10650 4724 10706
rect 2808 10526 2864 10582
rect 2932 10526 2988 10582
rect 3056 10526 3112 10582
rect 3180 10526 3236 10582
rect 3304 10526 3360 10582
rect 3428 10526 3484 10582
rect 3552 10526 3608 10582
rect 3676 10526 3732 10582
rect 3800 10526 3856 10582
rect 3924 10526 3980 10582
rect 4048 10526 4104 10582
rect 4172 10526 4228 10582
rect 4296 10526 4352 10582
rect 4420 10526 4476 10582
rect 4544 10526 4600 10582
rect 4668 10526 4724 10582
rect 2808 10402 2864 10458
rect 2932 10402 2988 10458
rect 3056 10402 3112 10458
rect 3180 10402 3236 10458
rect 3304 10402 3360 10458
rect 3428 10402 3484 10458
rect 3552 10402 3608 10458
rect 3676 10402 3732 10458
rect 3800 10402 3856 10458
rect 3924 10402 3980 10458
rect 4048 10402 4104 10458
rect 4172 10402 4228 10458
rect 4296 10402 4352 10458
rect 4420 10402 4476 10458
rect 4544 10402 4600 10458
rect 4668 10402 4724 10458
rect 2808 10278 2864 10334
rect 2932 10278 2988 10334
rect 3056 10278 3112 10334
rect 3180 10278 3236 10334
rect 3304 10278 3360 10334
rect 3428 10278 3484 10334
rect 3552 10278 3608 10334
rect 3676 10278 3732 10334
rect 3800 10278 3856 10334
rect 3924 10278 3980 10334
rect 4048 10278 4104 10334
rect 4172 10278 4228 10334
rect 4296 10278 4352 10334
rect 4420 10278 4476 10334
rect 4544 10278 4600 10334
rect 4668 10278 4724 10334
rect 2808 10154 2864 10210
rect 2932 10154 2988 10210
rect 3056 10154 3112 10210
rect 3180 10154 3236 10210
rect 3304 10154 3360 10210
rect 3428 10154 3484 10210
rect 3552 10154 3608 10210
rect 3676 10154 3732 10210
rect 3800 10154 3856 10210
rect 3924 10154 3980 10210
rect 4048 10154 4104 10210
rect 4172 10154 4228 10210
rect 4296 10154 4352 10210
rect 4420 10154 4476 10210
rect 4544 10154 4600 10210
rect 4668 10154 4724 10210
rect 2808 10030 2864 10086
rect 2932 10030 2988 10086
rect 3056 10030 3112 10086
rect 3180 10030 3236 10086
rect 3304 10030 3360 10086
rect 3428 10030 3484 10086
rect 3552 10030 3608 10086
rect 3676 10030 3732 10086
rect 3800 10030 3856 10086
rect 3924 10030 3980 10086
rect 4048 10030 4104 10086
rect 4172 10030 4228 10086
rect 4296 10030 4352 10086
rect 4420 10030 4476 10086
rect 4544 10030 4600 10086
rect 4668 10030 4724 10086
rect 2808 9906 2864 9962
rect 2932 9906 2988 9962
rect 3056 9906 3112 9962
rect 3180 9906 3236 9962
rect 3304 9906 3360 9962
rect 3428 9906 3484 9962
rect 3552 9906 3608 9962
rect 3676 9906 3732 9962
rect 3800 9906 3856 9962
rect 3924 9906 3980 9962
rect 4048 9906 4104 9962
rect 4172 9906 4228 9962
rect 4296 9906 4352 9962
rect 4420 9906 4476 9962
rect 4544 9906 4600 9962
rect 4668 9906 4724 9962
rect 2808 9782 2864 9838
rect 2932 9782 2988 9838
rect 3056 9782 3112 9838
rect 3180 9782 3236 9838
rect 3304 9782 3360 9838
rect 3428 9782 3484 9838
rect 3552 9782 3608 9838
rect 3676 9782 3732 9838
rect 3800 9782 3856 9838
rect 3924 9782 3980 9838
rect 4048 9782 4104 9838
rect 4172 9782 4228 9838
rect 4296 9782 4352 9838
rect 4420 9782 4476 9838
rect 4544 9782 4600 9838
rect 4668 9782 4724 9838
rect 2808 9658 2864 9714
rect 2932 9658 2988 9714
rect 3056 9658 3112 9714
rect 3180 9658 3236 9714
rect 3304 9658 3360 9714
rect 3428 9658 3484 9714
rect 3552 9658 3608 9714
rect 3676 9658 3732 9714
rect 3800 9658 3856 9714
rect 3924 9658 3980 9714
rect 4048 9658 4104 9714
rect 4172 9658 4228 9714
rect 4296 9658 4352 9714
rect 4420 9658 4476 9714
rect 4544 9658 4600 9714
rect 4668 9658 4724 9714
rect 2808 9534 2864 9590
rect 2932 9534 2988 9590
rect 3056 9534 3112 9590
rect 3180 9534 3236 9590
rect 3304 9534 3360 9590
rect 3428 9534 3484 9590
rect 3552 9534 3608 9590
rect 3676 9534 3732 9590
rect 3800 9534 3856 9590
rect 3924 9534 3980 9590
rect 4048 9534 4104 9590
rect 4172 9534 4228 9590
rect 4296 9534 4352 9590
rect 4420 9534 4476 9590
rect 4544 9534 4600 9590
rect 4668 9534 4724 9590
rect 2808 9410 2864 9466
rect 2932 9410 2988 9466
rect 3056 9410 3112 9466
rect 3180 9410 3236 9466
rect 3304 9410 3360 9466
rect 3428 9410 3484 9466
rect 3552 9410 3608 9466
rect 3676 9410 3732 9466
rect 3800 9410 3856 9466
rect 3924 9410 3980 9466
rect 4048 9410 4104 9466
rect 4172 9410 4228 9466
rect 4296 9410 4352 9466
rect 4420 9410 4476 9466
rect 4544 9410 4600 9466
rect 4668 9410 4724 9466
rect 2808 9286 2864 9342
rect 2932 9286 2988 9342
rect 3056 9286 3112 9342
rect 3180 9286 3236 9342
rect 3304 9286 3360 9342
rect 3428 9286 3484 9342
rect 3552 9286 3608 9342
rect 3676 9286 3732 9342
rect 3800 9286 3856 9342
rect 3924 9286 3980 9342
rect 4048 9286 4104 9342
rect 4172 9286 4228 9342
rect 4296 9286 4352 9342
rect 4420 9286 4476 9342
rect 4544 9286 4600 9342
rect 4668 9286 4724 9342
rect 2808 9162 2864 9218
rect 2932 9162 2988 9218
rect 3056 9162 3112 9218
rect 3180 9162 3236 9218
rect 3304 9162 3360 9218
rect 3428 9162 3484 9218
rect 3552 9162 3608 9218
rect 3676 9162 3732 9218
rect 3800 9162 3856 9218
rect 3924 9162 3980 9218
rect 4048 9162 4104 9218
rect 4172 9162 4228 9218
rect 4296 9162 4352 9218
rect 4420 9162 4476 9218
rect 4544 9162 4600 9218
rect 4668 9162 4724 9218
rect 2808 9038 2864 9094
rect 2932 9038 2988 9094
rect 3056 9038 3112 9094
rect 3180 9038 3236 9094
rect 3304 9038 3360 9094
rect 3428 9038 3484 9094
rect 3552 9038 3608 9094
rect 3676 9038 3732 9094
rect 3800 9038 3856 9094
rect 3924 9038 3980 9094
rect 4048 9038 4104 9094
rect 4172 9038 4228 9094
rect 4296 9038 4352 9094
rect 4420 9038 4476 9094
rect 4544 9038 4600 9094
rect 4668 9038 4724 9094
rect 2808 8914 2864 8970
rect 2932 8914 2988 8970
rect 3056 8914 3112 8970
rect 3180 8914 3236 8970
rect 3304 8914 3360 8970
rect 3428 8914 3484 8970
rect 3552 8914 3608 8970
rect 3676 8914 3732 8970
rect 3800 8914 3856 8970
rect 3924 8914 3980 8970
rect 4048 8914 4104 8970
rect 4172 8914 4228 8970
rect 4296 8914 4352 8970
rect 4420 8914 4476 8970
rect 4544 8914 4600 8970
rect 4668 8914 4724 8970
rect 2808 8790 2864 8846
rect 2932 8790 2988 8846
rect 3056 8790 3112 8846
rect 3180 8790 3236 8846
rect 3304 8790 3360 8846
rect 3428 8790 3484 8846
rect 3552 8790 3608 8846
rect 3676 8790 3732 8846
rect 3800 8790 3856 8846
rect 3924 8790 3980 8846
rect 4048 8790 4104 8846
rect 4172 8790 4228 8846
rect 4296 8790 4352 8846
rect 4420 8790 4476 8846
rect 4544 8790 4600 8846
rect 4668 8790 4724 8846
rect 2808 8666 2864 8722
rect 2932 8666 2988 8722
rect 3056 8666 3112 8722
rect 3180 8666 3236 8722
rect 3304 8666 3360 8722
rect 3428 8666 3484 8722
rect 3552 8666 3608 8722
rect 3676 8666 3732 8722
rect 3800 8666 3856 8722
rect 3924 8666 3980 8722
rect 4048 8666 4104 8722
rect 4172 8666 4228 8722
rect 4296 8666 4352 8722
rect 4420 8666 4476 8722
rect 4544 8666 4600 8722
rect 4668 8666 4724 8722
rect 2808 8542 2864 8598
rect 2932 8542 2988 8598
rect 3056 8542 3112 8598
rect 3180 8542 3236 8598
rect 3304 8542 3360 8598
rect 3428 8542 3484 8598
rect 3552 8542 3608 8598
rect 3676 8542 3732 8598
rect 3800 8542 3856 8598
rect 3924 8542 3980 8598
rect 4048 8542 4104 8598
rect 4172 8542 4228 8598
rect 4296 8542 4352 8598
rect 4420 8542 4476 8598
rect 4544 8542 4600 8598
rect 4668 8542 4724 8598
rect 2808 8418 2864 8474
rect 2932 8418 2988 8474
rect 3056 8418 3112 8474
rect 3180 8418 3236 8474
rect 3304 8418 3360 8474
rect 3428 8418 3484 8474
rect 3552 8418 3608 8474
rect 3676 8418 3732 8474
rect 3800 8418 3856 8474
rect 3924 8418 3980 8474
rect 4048 8418 4104 8474
rect 4172 8418 4228 8474
rect 4296 8418 4352 8474
rect 4420 8418 4476 8474
rect 4544 8418 4600 8474
rect 4668 8418 4724 8474
rect 2808 8294 2864 8350
rect 2932 8294 2988 8350
rect 3056 8294 3112 8350
rect 3180 8294 3236 8350
rect 3304 8294 3360 8350
rect 3428 8294 3484 8350
rect 3552 8294 3608 8350
rect 3676 8294 3732 8350
rect 3800 8294 3856 8350
rect 3924 8294 3980 8350
rect 4048 8294 4104 8350
rect 4172 8294 4228 8350
rect 4296 8294 4352 8350
rect 4420 8294 4476 8350
rect 4544 8294 4600 8350
rect 4668 8294 4724 8350
rect 2808 8170 2864 8226
rect 2932 8170 2988 8226
rect 3056 8170 3112 8226
rect 3180 8170 3236 8226
rect 3304 8170 3360 8226
rect 3428 8170 3484 8226
rect 3552 8170 3608 8226
rect 3676 8170 3732 8226
rect 3800 8170 3856 8226
rect 3924 8170 3980 8226
rect 4048 8170 4104 8226
rect 4172 8170 4228 8226
rect 4296 8170 4352 8226
rect 4420 8170 4476 8226
rect 4544 8170 4600 8226
rect 4668 8170 4724 8226
rect 2808 8046 2864 8102
rect 2932 8046 2988 8102
rect 3056 8046 3112 8102
rect 3180 8046 3236 8102
rect 3304 8046 3360 8102
rect 3428 8046 3484 8102
rect 3552 8046 3608 8102
rect 3676 8046 3732 8102
rect 3800 8046 3856 8102
rect 3924 8046 3980 8102
rect 4048 8046 4104 8102
rect 4172 8046 4228 8102
rect 4296 8046 4352 8102
rect 4420 8046 4476 8102
rect 4544 8046 4600 8102
rect 4668 8046 4724 8102
rect 5178 10898 5234 10954
rect 5302 10898 5358 10954
rect 5426 10898 5482 10954
rect 5550 10898 5606 10954
rect 5674 10898 5730 10954
rect 5798 10898 5854 10954
rect 5922 10898 5978 10954
rect 6046 10898 6102 10954
rect 6170 10898 6226 10954
rect 6294 10898 6350 10954
rect 6418 10898 6474 10954
rect 6542 10898 6598 10954
rect 6666 10898 6722 10954
rect 6790 10898 6846 10954
rect 6914 10898 6970 10954
rect 7038 10898 7094 10954
rect 5178 10774 5234 10830
rect 5302 10774 5358 10830
rect 5426 10774 5482 10830
rect 5550 10774 5606 10830
rect 5674 10774 5730 10830
rect 5798 10774 5854 10830
rect 5922 10774 5978 10830
rect 6046 10774 6102 10830
rect 6170 10774 6226 10830
rect 6294 10774 6350 10830
rect 6418 10774 6474 10830
rect 6542 10774 6598 10830
rect 6666 10774 6722 10830
rect 6790 10774 6846 10830
rect 6914 10774 6970 10830
rect 7038 10774 7094 10830
rect 5178 10650 5234 10706
rect 5302 10650 5358 10706
rect 5426 10650 5482 10706
rect 5550 10650 5606 10706
rect 5674 10650 5730 10706
rect 5798 10650 5854 10706
rect 5922 10650 5978 10706
rect 6046 10650 6102 10706
rect 6170 10650 6226 10706
rect 6294 10650 6350 10706
rect 6418 10650 6474 10706
rect 6542 10650 6598 10706
rect 6666 10650 6722 10706
rect 6790 10650 6846 10706
rect 6914 10650 6970 10706
rect 7038 10650 7094 10706
rect 5178 10526 5234 10582
rect 5302 10526 5358 10582
rect 5426 10526 5482 10582
rect 5550 10526 5606 10582
rect 5674 10526 5730 10582
rect 5798 10526 5854 10582
rect 5922 10526 5978 10582
rect 6046 10526 6102 10582
rect 6170 10526 6226 10582
rect 6294 10526 6350 10582
rect 6418 10526 6474 10582
rect 6542 10526 6598 10582
rect 6666 10526 6722 10582
rect 6790 10526 6846 10582
rect 6914 10526 6970 10582
rect 7038 10526 7094 10582
rect 5178 10402 5234 10458
rect 5302 10402 5358 10458
rect 5426 10402 5482 10458
rect 5550 10402 5606 10458
rect 5674 10402 5730 10458
rect 5798 10402 5854 10458
rect 5922 10402 5978 10458
rect 6046 10402 6102 10458
rect 6170 10402 6226 10458
rect 6294 10402 6350 10458
rect 6418 10402 6474 10458
rect 6542 10402 6598 10458
rect 6666 10402 6722 10458
rect 6790 10402 6846 10458
rect 6914 10402 6970 10458
rect 7038 10402 7094 10458
rect 5178 10278 5234 10334
rect 5302 10278 5358 10334
rect 5426 10278 5482 10334
rect 5550 10278 5606 10334
rect 5674 10278 5730 10334
rect 5798 10278 5854 10334
rect 5922 10278 5978 10334
rect 6046 10278 6102 10334
rect 6170 10278 6226 10334
rect 6294 10278 6350 10334
rect 6418 10278 6474 10334
rect 6542 10278 6598 10334
rect 6666 10278 6722 10334
rect 6790 10278 6846 10334
rect 6914 10278 6970 10334
rect 7038 10278 7094 10334
rect 5178 10154 5234 10210
rect 5302 10154 5358 10210
rect 5426 10154 5482 10210
rect 5550 10154 5606 10210
rect 5674 10154 5730 10210
rect 5798 10154 5854 10210
rect 5922 10154 5978 10210
rect 6046 10154 6102 10210
rect 6170 10154 6226 10210
rect 6294 10154 6350 10210
rect 6418 10154 6474 10210
rect 6542 10154 6598 10210
rect 6666 10154 6722 10210
rect 6790 10154 6846 10210
rect 6914 10154 6970 10210
rect 7038 10154 7094 10210
rect 5178 10030 5234 10086
rect 5302 10030 5358 10086
rect 5426 10030 5482 10086
rect 5550 10030 5606 10086
rect 5674 10030 5730 10086
rect 5798 10030 5854 10086
rect 5922 10030 5978 10086
rect 6046 10030 6102 10086
rect 6170 10030 6226 10086
rect 6294 10030 6350 10086
rect 6418 10030 6474 10086
rect 6542 10030 6598 10086
rect 6666 10030 6722 10086
rect 6790 10030 6846 10086
rect 6914 10030 6970 10086
rect 7038 10030 7094 10086
rect 5178 9906 5234 9962
rect 5302 9906 5358 9962
rect 5426 9906 5482 9962
rect 5550 9906 5606 9962
rect 5674 9906 5730 9962
rect 5798 9906 5854 9962
rect 5922 9906 5978 9962
rect 6046 9906 6102 9962
rect 6170 9906 6226 9962
rect 6294 9906 6350 9962
rect 6418 9906 6474 9962
rect 6542 9906 6598 9962
rect 6666 9906 6722 9962
rect 6790 9906 6846 9962
rect 6914 9906 6970 9962
rect 7038 9906 7094 9962
rect 5178 9782 5234 9838
rect 5302 9782 5358 9838
rect 5426 9782 5482 9838
rect 5550 9782 5606 9838
rect 5674 9782 5730 9838
rect 5798 9782 5854 9838
rect 5922 9782 5978 9838
rect 6046 9782 6102 9838
rect 6170 9782 6226 9838
rect 6294 9782 6350 9838
rect 6418 9782 6474 9838
rect 6542 9782 6598 9838
rect 6666 9782 6722 9838
rect 6790 9782 6846 9838
rect 6914 9782 6970 9838
rect 7038 9782 7094 9838
rect 5178 9658 5234 9714
rect 5302 9658 5358 9714
rect 5426 9658 5482 9714
rect 5550 9658 5606 9714
rect 5674 9658 5730 9714
rect 5798 9658 5854 9714
rect 5922 9658 5978 9714
rect 6046 9658 6102 9714
rect 6170 9658 6226 9714
rect 6294 9658 6350 9714
rect 6418 9658 6474 9714
rect 6542 9658 6598 9714
rect 6666 9658 6722 9714
rect 6790 9658 6846 9714
rect 6914 9658 6970 9714
rect 7038 9658 7094 9714
rect 5178 9534 5234 9590
rect 5302 9534 5358 9590
rect 5426 9534 5482 9590
rect 5550 9534 5606 9590
rect 5674 9534 5730 9590
rect 5798 9534 5854 9590
rect 5922 9534 5978 9590
rect 6046 9534 6102 9590
rect 6170 9534 6226 9590
rect 6294 9534 6350 9590
rect 6418 9534 6474 9590
rect 6542 9534 6598 9590
rect 6666 9534 6722 9590
rect 6790 9534 6846 9590
rect 6914 9534 6970 9590
rect 7038 9534 7094 9590
rect 5178 9410 5234 9466
rect 5302 9410 5358 9466
rect 5426 9410 5482 9466
rect 5550 9410 5606 9466
rect 5674 9410 5730 9466
rect 5798 9410 5854 9466
rect 5922 9410 5978 9466
rect 6046 9410 6102 9466
rect 6170 9410 6226 9466
rect 6294 9410 6350 9466
rect 6418 9410 6474 9466
rect 6542 9410 6598 9466
rect 6666 9410 6722 9466
rect 6790 9410 6846 9466
rect 6914 9410 6970 9466
rect 7038 9410 7094 9466
rect 5178 9286 5234 9342
rect 5302 9286 5358 9342
rect 5426 9286 5482 9342
rect 5550 9286 5606 9342
rect 5674 9286 5730 9342
rect 5798 9286 5854 9342
rect 5922 9286 5978 9342
rect 6046 9286 6102 9342
rect 6170 9286 6226 9342
rect 6294 9286 6350 9342
rect 6418 9286 6474 9342
rect 6542 9286 6598 9342
rect 6666 9286 6722 9342
rect 6790 9286 6846 9342
rect 6914 9286 6970 9342
rect 7038 9286 7094 9342
rect 5178 9162 5234 9218
rect 5302 9162 5358 9218
rect 5426 9162 5482 9218
rect 5550 9162 5606 9218
rect 5674 9162 5730 9218
rect 5798 9162 5854 9218
rect 5922 9162 5978 9218
rect 6046 9162 6102 9218
rect 6170 9162 6226 9218
rect 6294 9162 6350 9218
rect 6418 9162 6474 9218
rect 6542 9162 6598 9218
rect 6666 9162 6722 9218
rect 6790 9162 6846 9218
rect 6914 9162 6970 9218
rect 7038 9162 7094 9218
rect 5178 9038 5234 9094
rect 5302 9038 5358 9094
rect 5426 9038 5482 9094
rect 5550 9038 5606 9094
rect 5674 9038 5730 9094
rect 5798 9038 5854 9094
rect 5922 9038 5978 9094
rect 6046 9038 6102 9094
rect 6170 9038 6226 9094
rect 6294 9038 6350 9094
rect 6418 9038 6474 9094
rect 6542 9038 6598 9094
rect 6666 9038 6722 9094
rect 6790 9038 6846 9094
rect 6914 9038 6970 9094
rect 7038 9038 7094 9094
rect 5178 8914 5234 8970
rect 5302 8914 5358 8970
rect 5426 8914 5482 8970
rect 5550 8914 5606 8970
rect 5674 8914 5730 8970
rect 5798 8914 5854 8970
rect 5922 8914 5978 8970
rect 6046 8914 6102 8970
rect 6170 8914 6226 8970
rect 6294 8914 6350 8970
rect 6418 8914 6474 8970
rect 6542 8914 6598 8970
rect 6666 8914 6722 8970
rect 6790 8914 6846 8970
rect 6914 8914 6970 8970
rect 7038 8914 7094 8970
rect 5178 8790 5234 8846
rect 5302 8790 5358 8846
rect 5426 8790 5482 8846
rect 5550 8790 5606 8846
rect 5674 8790 5730 8846
rect 5798 8790 5854 8846
rect 5922 8790 5978 8846
rect 6046 8790 6102 8846
rect 6170 8790 6226 8846
rect 6294 8790 6350 8846
rect 6418 8790 6474 8846
rect 6542 8790 6598 8846
rect 6666 8790 6722 8846
rect 6790 8790 6846 8846
rect 6914 8790 6970 8846
rect 7038 8790 7094 8846
rect 5178 8666 5234 8722
rect 5302 8666 5358 8722
rect 5426 8666 5482 8722
rect 5550 8666 5606 8722
rect 5674 8666 5730 8722
rect 5798 8666 5854 8722
rect 5922 8666 5978 8722
rect 6046 8666 6102 8722
rect 6170 8666 6226 8722
rect 6294 8666 6350 8722
rect 6418 8666 6474 8722
rect 6542 8666 6598 8722
rect 6666 8666 6722 8722
rect 6790 8666 6846 8722
rect 6914 8666 6970 8722
rect 7038 8666 7094 8722
rect 5178 8542 5234 8598
rect 5302 8542 5358 8598
rect 5426 8542 5482 8598
rect 5550 8542 5606 8598
rect 5674 8542 5730 8598
rect 5798 8542 5854 8598
rect 5922 8542 5978 8598
rect 6046 8542 6102 8598
rect 6170 8542 6226 8598
rect 6294 8542 6350 8598
rect 6418 8542 6474 8598
rect 6542 8542 6598 8598
rect 6666 8542 6722 8598
rect 6790 8542 6846 8598
rect 6914 8542 6970 8598
rect 7038 8542 7094 8598
rect 5178 8418 5234 8474
rect 5302 8418 5358 8474
rect 5426 8418 5482 8474
rect 5550 8418 5606 8474
rect 5674 8418 5730 8474
rect 5798 8418 5854 8474
rect 5922 8418 5978 8474
rect 6046 8418 6102 8474
rect 6170 8418 6226 8474
rect 6294 8418 6350 8474
rect 6418 8418 6474 8474
rect 6542 8418 6598 8474
rect 6666 8418 6722 8474
rect 6790 8418 6846 8474
rect 6914 8418 6970 8474
rect 7038 8418 7094 8474
rect 5178 8294 5234 8350
rect 5302 8294 5358 8350
rect 5426 8294 5482 8350
rect 5550 8294 5606 8350
rect 5674 8294 5730 8350
rect 5798 8294 5854 8350
rect 5922 8294 5978 8350
rect 6046 8294 6102 8350
rect 6170 8294 6226 8350
rect 6294 8294 6350 8350
rect 6418 8294 6474 8350
rect 6542 8294 6598 8350
rect 6666 8294 6722 8350
rect 6790 8294 6846 8350
rect 6914 8294 6970 8350
rect 7038 8294 7094 8350
rect 5178 8170 5234 8226
rect 5302 8170 5358 8226
rect 5426 8170 5482 8226
rect 5550 8170 5606 8226
rect 5674 8170 5730 8226
rect 5798 8170 5854 8226
rect 5922 8170 5978 8226
rect 6046 8170 6102 8226
rect 6170 8170 6226 8226
rect 6294 8170 6350 8226
rect 6418 8170 6474 8226
rect 6542 8170 6598 8226
rect 6666 8170 6722 8226
rect 6790 8170 6846 8226
rect 6914 8170 6970 8226
rect 7038 8170 7094 8226
rect 5178 8046 5234 8102
rect 5302 8046 5358 8102
rect 5426 8046 5482 8102
rect 5550 8046 5606 8102
rect 5674 8046 5730 8102
rect 5798 8046 5854 8102
rect 5922 8046 5978 8102
rect 6046 8046 6102 8102
rect 6170 8046 6226 8102
rect 6294 8046 6350 8102
rect 6418 8046 6474 8102
rect 6542 8046 6598 8102
rect 6666 8046 6722 8102
rect 6790 8046 6846 8102
rect 6914 8046 6970 8102
rect 7038 8046 7094 8102
rect 7884 10898 7940 10954
rect 8008 10898 8064 10954
rect 8132 10898 8188 10954
rect 8256 10898 8312 10954
rect 8380 10898 8436 10954
rect 8504 10898 8560 10954
rect 8628 10898 8684 10954
rect 8752 10898 8808 10954
rect 8876 10898 8932 10954
rect 9000 10898 9056 10954
rect 9124 10898 9180 10954
rect 9248 10898 9304 10954
rect 9372 10898 9428 10954
rect 9496 10898 9552 10954
rect 9620 10898 9676 10954
rect 9744 10898 9800 10954
rect 7884 10774 7940 10830
rect 8008 10774 8064 10830
rect 8132 10774 8188 10830
rect 8256 10774 8312 10830
rect 8380 10774 8436 10830
rect 8504 10774 8560 10830
rect 8628 10774 8684 10830
rect 8752 10774 8808 10830
rect 8876 10774 8932 10830
rect 9000 10774 9056 10830
rect 9124 10774 9180 10830
rect 9248 10774 9304 10830
rect 9372 10774 9428 10830
rect 9496 10774 9552 10830
rect 9620 10774 9676 10830
rect 9744 10774 9800 10830
rect 7884 10650 7940 10706
rect 8008 10650 8064 10706
rect 8132 10650 8188 10706
rect 8256 10650 8312 10706
rect 8380 10650 8436 10706
rect 8504 10650 8560 10706
rect 8628 10650 8684 10706
rect 8752 10650 8808 10706
rect 8876 10650 8932 10706
rect 9000 10650 9056 10706
rect 9124 10650 9180 10706
rect 9248 10650 9304 10706
rect 9372 10650 9428 10706
rect 9496 10650 9552 10706
rect 9620 10650 9676 10706
rect 9744 10650 9800 10706
rect 7884 10526 7940 10582
rect 8008 10526 8064 10582
rect 8132 10526 8188 10582
rect 8256 10526 8312 10582
rect 8380 10526 8436 10582
rect 8504 10526 8560 10582
rect 8628 10526 8684 10582
rect 8752 10526 8808 10582
rect 8876 10526 8932 10582
rect 9000 10526 9056 10582
rect 9124 10526 9180 10582
rect 9248 10526 9304 10582
rect 9372 10526 9428 10582
rect 9496 10526 9552 10582
rect 9620 10526 9676 10582
rect 9744 10526 9800 10582
rect 7884 10402 7940 10458
rect 8008 10402 8064 10458
rect 8132 10402 8188 10458
rect 8256 10402 8312 10458
rect 8380 10402 8436 10458
rect 8504 10402 8560 10458
rect 8628 10402 8684 10458
rect 8752 10402 8808 10458
rect 8876 10402 8932 10458
rect 9000 10402 9056 10458
rect 9124 10402 9180 10458
rect 9248 10402 9304 10458
rect 9372 10402 9428 10458
rect 9496 10402 9552 10458
rect 9620 10402 9676 10458
rect 9744 10402 9800 10458
rect 7884 10278 7940 10334
rect 8008 10278 8064 10334
rect 8132 10278 8188 10334
rect 8256 10278 8312 10334
rect 8380 10278 8436 10334
rect 8504 10278 8560 10334
rect 8628 10278 8684 10334
rect 8752 10278 8808 10334
rect 8876 10278 8932 10334
rect 9000 10278 9056 10334
rect 9124 10278 9180 10334
rect 9248 10278 9304 10334
rect 9372 10278 9428 10334
rect 9496 10278 9552 10334
rect 9620 10278 9676 10334
rect 9744 10278 9800 10334
rect 7884 10154 7940 10210
rect 8008 10154 8064 10210
rect 8132 10154 8188 10210
rect 8256 10154 8312 10210
rect 8380 10154 8436 10210
rect 8504 10154 8560 10210
rect 8628 10154 8684 10210
rect 8752 10154 8808 10210
rect 8876 10154 8932 10210
rect 9000 10154 9056 10210
rect 9124 10154 9180 10210
rect 9248 10154 9304 10210
rect 9372 10154 9428 10210
rect 9496 10154 9552 10210
rect 9620 10154 9676 10210
rect 9744 10154 9800 10210
rect 7884 10030 7940 10086
rect 8008 10030 8064 10086
rect 8132 10030 8188 10086
rect 8256 10030 8312 10086
rect 8380 10030 8436 10086
rect 8504 10030 8560 10086
rect 8628 10030 8684 10086
rect 8752 10030 8808 10086
rect 8876 10030 8932 10086
rect 9000 10030 9056 10086
rect 9124 10030 9180 10086
rect 9248 10030 9304 10086
rect 9372 10030 9428 10086
rect 9496 10030 9552 10086
rect 9620 10030 9676 10086
rect 9744 10030 9800 10086
rect 7884 9906 7940 9962
rect 8008 9906 8064 9962
rect 8132 9906 8188 9962
rect 8256 9906 8312 9962
rect 8380 9906 8436 9962
rect 8504 9906 8560 9962
rect 8628 9906 8684 9962
rect 8752 9906 8808 9962
rect 8876 9906 8932 9962
rect 9000 9906 9056 9962
rect 9124 9906 9180 9962
rect 9248 9906 9304 9962
rect 9372 9906 9428 9962
rect 9496 9906 9552 9962
rect 9620 9906 9676 9962
rect 9744 9906 9800 9962
rect 7884 9782 7940 9838
rect 8008 9782 8064 9838
rect 8132 9782 8188 9838
rect 8256 9782 8312 9838
rect 8380 9782 8436 9838
rect 8504 9782 8560 9838
rect 8628 9782 8684 9838
rect 8752 9782 8808 9838
rect 8876 9782 8932 9838
rect 9000 9782 9056 9838
rect 9124 9782 9180 9838
rect 9248 9782 9304 9838
rect 9372 9782 9428 9838
rect 9496 9782 9552 9838
rect 9620 9782 9676 9838
rect 9744 9782 9800 9838
rect 7884 9658 7940 9714
rect 8008 9658 8064 9714
rect 8132 9658 8188 9714
rect 8256 9658 8312 9714
rect 8380 9658 8436 9714
rect 8504 9658 8560 9714
rect 8628 9658 8684 9714
rect 8752 9658 8808 9714
rect 8876 9658 8932 9714
rect 9000 9658 9056 9714
rect 9124 9658 9180 9714
rect 9248 9658 9304 9714
rect 9372 9658 9428 9714
rect 9496 9658 9552 9714
rect 9620 9658 9676 9714
rect 9744 9658 9800 9714
rect 7884 9534 7940 9590
rect 8008 9534 8064 9590
rect 8132 9534 8188 9590
rect 8256 9534 8312 9590
rect 8380 9534 8436 9590
rect 8504 9534 8560 9590
rect 8628 9534 8684 9590
rect 8752 9534 8808 9590
rect 8876 9534 8932 9590
rect 9000 9534 9056 9590
rect 9124 9534 9180 9590
rect 9248 9534 9304 9590
rect 9372 9534 9428 9590
rect 9496 9534 9552 9590
rect 9620 9534 9676 9590
rect 9744 9534 9800 9590
rect 7884 9410 7940 9466
rect 8008 9410 8064 9466
rect 8132 9410 8188 9466
rect 8256 9410 8312 9466
rect 8380 9410 8436 9466
rect 8504 9410 8560 9466
rect 8628 9410 8684 9466
rect 8752 9410 8808 9466
rect 8876 9410 8932 9466
rect 9000 9410 9056 9466
rect 9124 9410 9180 9466
rect 9248 9410 9304 9466
rect 9372 9410 9428 9466
rect 9496 9410 9552 9466
rect 9620 9410 9676 9466
rect 9744 9410 9800 9466
rect 7884 9286 7940 9342
rect 8008 9286 8064 9342
rect 8132 9286 8188 9342
rect 8256 9286 8312 9342
rect 8380 9286 8436 9342
rect 8504 9286 8560 9342
rect 8628 9286 8684 9342
rect 8752 9286 8808 9342
rect 8876 9286 8932 9342
rect 9000 9286 9056 9342
rect 9124 9286 9180 9342
rect 9248 9286 9304 9342
rect 9372 9286 9428 9342
rect 9496 9286 9552 9342
rect 9620 9286 9676 9342
rect 9744 9286 9800 9342
rect 7884 9162 7940 9218
rect 8008 9162 8064 9218
rect 8132 9162 8188 9218
rect 8256 9162 8312 9218
rect 8380 9162 8436 9218
rect 8504 9162 8560 9218
rect 8628 9162 8684 9218
rect 8752 9162 8808 9218
rect 8876 9162 8932 9218
rect 9000 9162 9056 9218
rect 9124 9162 9180 9218
rect 9248 9162 9304 9218
rect 9372 9162 9428 9218
rect 9496 9162 9552 9218
rect 9620 9162 9676 9218
rect 9744 9162 9800 9218
rect 7884 9038 7940 9094
rect 8008 9038 8064 9094
rect 8132 9038 8188 9094
rect 8256 9038 8312 9094
rect 8380 9038 8436 9094
rect 8504 9038 8560 9094
rect 8628 9038 8684 9094
rect 8752 9038 8808 9094
rect 8876 9038 8932 9094
rect 9000 9038 9056 9094
rect 9124 9038 9180 9094
rect 9248 9038 9304 9094
rect 9372 9038 9428 9094
rect 9496 9038 9552 9094
rect 9620 9038 9676 9094
rect 9744 9038 9800 9094
rect 7884 8914 7940 8970
rect 8008 8914 8064 8970
rect 8132 8914 8188 8970
rect 8256 8914 8312 8970
rect 8380 8914 8436 8970
rect 8504 8914 8560 8970
rect 8628 8914 8684 8970
rect 8752 8914 8808 8970
rect 8876 8914 8932 8970
rect 9000 8914 9056 8970
rect 9124 8914 9180 8970
rect 9248 8914 9304 8970
rect 9372 8914 9428 8970
rect 9496 8914 9552 8970
rect 9620 8914 9676 8970
rect 9744 8914 9800 8970
rect 7884 8790 7940 8846
rect 8008 8790 8064 8846
rect 8132 8790 8188 8846
rect 8256 8790 8312 8846
rect 8380 8790 8436 8846
rect 8504 8790 8560 8846
rect 8628 8790 8684 8846
rect 8752 8790 8808 8846
rect 8876 8790 8932 8846
rect 9000 8790 9056 8846
rect 9124 8790 9180 8846
rect 9248 8790 9304 8846
rect 9372 8790 9428 8846
rect 9496 8790 9552 8846
rect 9620 8790 9676 8846
rect 9744 8790 9800 8846
rect 7884 8666 7940 8722
rect 8008 8666 8064 8722
rect 8132 8666 8188 8722
rect 8256 8666 8312 8722
rect 8380 8666 8436 8722
rect 8504 8666 8560 8722
rect 8628 8666 8684 8722
rect 8752 8666 8808 8722
rect 8876 8666 8932 8722
rect 9000 8666 9056 8722
rect 9124 8666 9180 8722
rect 9248 8666 9304 8722
rect 9372 8666 9428 8722
rect 9496 8666 9552 8722
rect 9620 8666 9676 8722
rect 9744 8666 9800 8722
rect 7884 8542 7940 8598
rect 8008 8542 8064 8598
rect 8132 8542 8188 8598
rect 8256 8542 8312 8598
rect 8380 8542 8436 8598
rect 8504 8542 8560 8598
rect 8628 8542 8684 8598
rect 8752 8542 8808 8598
rect 8876 8542 8932 8598
rect 9000 8542 9056 8598
rect 9124 8542 9180 8598
rect 9248 8542 9304 8598
rect 9372 8542 9428 8598
rect 9496 8542 9552 8598
rect 9620 8542 9676 8598
rect 9744 8542 9800 8598
rect 7884 8418 7940 8474
rect 8008 8418 8064 8474
rect 8132 8418 8188 8474
rect 8256 8418 8312 8474
rect 8380 8418 8436 8474
rect 8504 8418 8560 8474
rect 8628 8418 8684 8474
rect 8752 8418 8808 8474
rect 8876 8418 8932 8474
rect 9000 8418 9056 8474
rect 9124 8418 9180 8474
rect 9248 8418 9304 8474
rect 9372 8418 9428 8474
rect 9496 8418 9552 8474
rect 9620 8418 9676 8474
rect 9744 8418 9800 8474
rect 7884 8294 7940 8350
rect 8008 8294 8064 8350
rect 8132 8294 8188 8350
rect 8256 8294 8312 8350
rect 8380 8294 8436 8350
rect 8504 8294 8560 8350
rect 8628 8294 8684 8350
rect 8752 8294 8808 8350
rect 8876 8294 8932 8350
rect 9000 8294 9056 8350
rect 9124 8294 9180 8350
rect 9248 8294 9304 8350
rect 9372 8294 9428 8350
rect 9496 8294 9552 8350
rect 9620 8294 9676 8350
rect 9744 8294 9800 8350
rect 7884 8170 7940 8226
rect 8008 8170 8064 8226
rect 8132 8170 8188 8226
rect 8256 8170 8312 8226
rect 8380 8170 8436 8226
rect 8504 8170 8560 8226
rect 8628 8170 8684 8226
rect 8752 8170 8808 8226
rect 8876 8170 8932 8226
rect 9000 8170 9056 8226
rect 9124 8170 9180 8226
rect 9248 8170 9304 8226
rect 9372 8170 9428 8226
rect 9496 8170 9552 8226
rect 9620 8170 9676 8226
rect 9744 8170 9800 8226
rect 7884 8046 7940 8102
rect 8008 8046 8064 8102
rect 8132 8046 8188 8102
rect 8256 8046 8312 8102
rect 8380 8046 8436 8102
rect 8504 8046 8560 8102
rect 8628 8046 8684 8102
rect 8752 8046 8808 8102
rect 8876 8046 8932 8102
rect 9000 8046 9056 8102
rect 9124 8046 9180 8102
rect 9248 8046 9304 8102
rect 9372 8046 9428 8102
rect 9496 8046 9552 8102
rect 9620 8046 9676 8102
rect 9744 8046 9800 8102
rect 10254 10898 10310 10954
rect 10378 10898 10434 10954
rect 10502 10898 10558 10954
rect 10626 10898 10682 10954
rect 10750 10898 10806 10954
rect 10874 10898 10930 10954
rect 10998 10898 11054 10954
rect 11122 10898 11178 10954
rect 11246 10898 11302 10954
rect 11370 10898 11426 10954
rect 11494 10898 11550 10954
rect 11618 10898 11674 10954
rect 11742 10898 11798 10954
rect 11866 10898 11922 10954
rect 11990 10898 12046 10954
rect 12114 10898 12170 10954
rect 10254 10774 10310 10830
rect 10378 10774 10434 10830
rect 10502 10774 10558 10830
rect 10626 10774 10682 10830
rect 10750 10774 10806 10830
rect 10874 10774 10930 10830
rect 10998 10774 11054 10830
rect 11122 10774 11178 10830
rect 11246 10774 11302 10830
rect 11370 10774 11426 10830
rect 11494 10774 11550 10830
rect 11618 10774 11674 10830
rect 11742 10774 11798 10830
rect 11866 10774 11922 10830
rect 11990 10774 12046 10830
rect 12114 10774 12170 10830
rect 10254 10650 10310 10706
rect 10378 10650 10434 10706
rect 10502 10650 10558 10706
rect 10626 10650 10682 10706
rect 10750 10650 10806 10706
rect 10874 10650 10930 10706
rect 10998 10650 11054 10706
rect 11122 10650 11178 10706
rect 11246 10650 11302 10706
rect 11370 10650 11426 10706
rect 11494 10650 11550 10706
rect 11618 10650 11674 10706
rect 11742 10650 11798 10706
rect 11866 10650 11922 10706
rect 11990 10650 12046 10706
rect 12114 10650 12170 10706
rect 10254 10526 10310 10582
rect 10378 10526 10434 10582
rect 10502 10526 10558 10582
rect 10626 10526 10682 10582
rect 10750 10526 10806 10582
rect 10874 10526 10930 10582
rect 10998 10526 11054 10582
rect 11122 10526 11178 10582
rect 11246 10526 11302 10582
rect 11370 10526 11426 10582
rect 11494 10526 11550 10582
rect 11618 10526 11674 10582
rect 11742 10526 11798 10582
rect 11866 10526 11922 10582
rect 11990 10526 12046 10582
rect 12114 10526 12170 10582
rect 10254 10402 10310 10458
rect 10378 10402 10434 10458
rect 10502 10402 10558 10458
rect 10626 10402 10682 10458
rect 10750 10402 10806 10458
rect 10874 10402 10930 10458
rect 10998 10402 11054 10458
rect 11122 10402 11178 10458
rect 11246 10402 11302 10458
rect 11370 10402 11426 10458
rect 11494 10402 11550 10458
rect 11618 10402 11674 10458
rect 11742 10402 11798 10458
rect 11866 10402 11922 10458
rect 11990 10402 12046 10458
rect 12114 10402 12170 10458
rect 10254 10278 10310 10334
rect 10378 10278 10434 10334
rect 10502 10278 10558 10334
rect 10626 10278 10682 10334
rect 10750 10278 10806 10334
rect 10874 10278 10930 10334
rect 10998 10278 11054 10334
rect 11122 10278 11178 10334
rect 11246 10278 11302 10334
rect 11370 10278 11426 10334
rect 11494 10278 11550 10334
rect 11618 10278 11674 10334
rect 11742 10278 11798 10334
rect 11866 10278 11922 10334
rect 11990 10278 12046 10334
rect 12114 10278 12170 10334
rect 10254 10154 10310 10210
rect 10378 10154 10434 10210
rect 10502 10154 10558 10210
rect 10626 10154 10682 10210
rect 10750 10154 10806 10210
rect 10874 10154 10930 10210
rect 10998 10154 11054 10210
rect 11122 10154 11178 10210
rect 11246 10154 11302 10210
rect 11370 10154 11426 10210
rect 11494 10154 11550 10210
rect 11618 10154 11674 10210
rect 11742 10154 11798 10210
rect 11866 10154 11922 10210
rect 11990 10154 12046 10210
rect 12114 10154 12170 10210
rect 10254 10030 10310 10086
rect 10378 10030 10434 10086
rect 10502 10030 10558 10086
rect 10626 10030 10682 10086
rect 10750 10030 10806 10086
rect 10874 10030 10930 10086
rect 10998 10030 11054 10086
rect 11122 10030 11178 10086
rect 11246 10030 11302 10086
rect 11370 10030 11426 10086
rect 11494 10030 11550 10086
rect 11618 10030 11674 10086
rect 11742 10030 11798 10086
rect 11866 10030 11922 10086
rect 11990 10030 12046 10086
rect 12114 10030 12170 10086
rect 10254 9906 10310 9962
rect 10378 9906 10434 9962
rect 10502 9906 10558 9962
rect 10626 9906 10682 9962
rect 10750 9906 10806 9962
rect 10874 9906 10930 9962
rect 10998 9906 11054 9962
rect 11122 9906 11178 9962
rect 11246 9906 11302 9962
rect 11370 9906 11426 9962
rect 11494 9906 11550 9962
rect 11618 9906 11674 9962
rect 11742 9906 11798 9962
rect 11866 9906 11922 9962
rect 11990 9906 12046 9962
rect 12114 9906 12170 9962
rect 10254 9782 10310 9838
rect 10378 9782 10434 9838
rect 10502 9782 10558 9838
rect 10626 9782 10682 9838
rect 10750 9782 10806 9838
rect 10874 9782 10930 9838
rect 10998 9782 11054 9838
rect 11122 9782 11178 9838
rect 11246 9782 11302 9838
rect 11370 9782 11426 9838
rect 11494 9782 11550 9838
rect 11618 9782 11674 9838
rect 11742 9782 11798 9838
rect 11866 9782 11922 9838
rect 11990 9782 12046 9838
rect 12114 9782 12170 9838
rect 10254 9658 10310 9714
rect 10378 9658 10434 9714
rect 10502 9658 10558 9714
rect 10626 9658 10682 9714
rect 10750 9658 10806 9714
rect 10874 9658 10930 9714
rect 10998 9658 11054 9714
rect 11122 9658 11178 9714
rect 11246 9658 11302 9714
rect 11370 9658 11426 9714
rect 11494 9658 11550 9714
rect 11618 9658 11674 9714
rect 11742 9658 11798 9714
rect 11866 9658 11922 9714
rect 11990 9658 12046 9714
rect 12114 9658 12170 9714
rect 10254 9534 10310 9590
rect 10378 9534 10434 9590
rect 10502 9534 10558 9590
rect 10626 9534 10682 9590
rect 10750 9534 10806 9590
rect 10874 9534 10930 9590
rect 10998 9534 11054 9590
rect 11122 9534 11178 9590
rect 11246 9534 11302 9590
rect 11370 9534 11426 9590
rect 11494 9534 11550 9590
rect 11618 9534 11674 9590
rect 11742 9534 11798 9590
rect 11866 9534 11922 9590
rect 11990 9534 12046 9590
rect 12114 9534 12170 9590
rect 10254 9410 10310 9466
rect 10378 9410 10434 9466
rect 10502 9410 10558 9466
rect 10626 9410 10682 9466
rect 10750 9410 10806 9466
rect 10874 9410 10930 9466
rect 10998 9410 11054 9466
rect 11122 9410 11178 9466
rect 11246 9410 11302 9466
rect 11370 9410 11426 9466
rect 11494 9410 11550 9466
rect 11618 9410 11674 9466
rect 11742 9410 11798 9466
rect 11866 9410 11922 9466
rect 11990 9410 12046 9466
rect 12114 9410 12170 9466
rect 10254 9286 10310 9342
rect 10378 9286 10434 9342
rect 10502 9286 10558 9342
rect 10626 9286 10682 9342
rect 10750 9286 10806 9342
rect 10874 9286 10930 9342
rect 10998 9286 11054 9342
rect 11122 9286 11178 9342
rect 11246 9286 11302 9342
rect 11370 9286 11426 9342
rect 11494 9286 11550 9342
rect 11618 9286 11674 9342
rect 11742 9286 11798 9342
rect 11866 9286 11922 9342
rect 11990 9286 12046 9342
rect 12114 9286 12170 9342
rect 10254 9162 10310 9218
rect 10378 9162 10434 9218
rect 10502 9162 10558 9218
rect 10626 9162 10682 9218
rect 10750 9162 10806 9218
rect 10874 9162 10930 9218
rect 10998 9162 11054 9218
rect 11122 9162 11178 9218
rect 11246 9162 11302 9218
rect 11370 9162 11426 9218
rect 11494 9162 11550 9218
rect 11618 9162 11674 9218
rect 11742 9162 11798 9218
rect 11866 9162 11922 9218
rect 11990 9162 12046 9218
rect 12114 9162 12170 9218
rect 10254 9038 10310 9094
rect 10378 9038 10434 9094
rect 10502 9038 10558 9094
rect 10626 9038 10682 9094
rect 10750 9038 10806 9094
rect 10874 9038 10930 9094
rect 10998 9038 11054 9094
rect 11122 9038 11178 9094
rect 11246 9038 11302 9094
rect 11370 9038 11426 9094
rect 11494 9038 11550 9094
rect 11618 9038 11674 9094
rect 11742 9038 11798 9094
rect 11866 9038 11922 9094
rect 11990 9038 12046 9094
rect 12114 9038 12170 9094
rect 10254 8914 10310 8970
rect 10378 8914 10434 8970
rect 10502 8914 10558 8970
rect 10626 8914 10682 8970
rect 10750 8914 10806 8970
rect 10874 8914 10930 8970
rect 10998 8914 11054 8970
rect 11122 8914 11178 8970
rect 11246 8914 11302 8970
rect 11370 8914 11426 8970
rect 11494 8914 11550 8970
rect 11618 8914 11674 8970
rect 11742 8914 11798 8970
rect 11866 8914 11922 8970
rect 11990 8914 12046 8970
rect 12114 8914 12170 8970
rect 10254 8790 10310 8846
rect 10378 8790 10434 8846
rect 10502 8790 10558 8846
rect 10626 8790 10682 8846
rect 10750 8790 10806 8846
rect 10874 8790 10930 8846
rect 10998 8790 11054 8846
rect 11122 8790 11178 8846
rect 11246 8790 11302 8846
rect 11370 8790 11426 8846
rect 11494 8790 11550 8846
rect 11618 8790 11674 8846
rect 11742 8790 11798 8846
rect 11866 8790 11922 8846
rect 11990 8790 12046 8846
rect 12114 8790 12170 8846
rect 10254 8666 10310 8722
rect 10378 8666 10434 8722
rect 10502 8666 10558 8722
rect 10626 8666 10682 8722
rect 10750 8666 10806 8722
rect 10874 8666 10930 8722
rect 10998 8666 11054 8722
rect 11122 8666 11178 8722
rect 11246 8666 11302 8722
rect 11370 8666 11426 8722
rect 11494 8666 11550 8722
rect 11618 8666 11674 8722
rect 11742 8666 11798 8722
rect 11866 8666 11922 8722
rect 11990 8666 12046 8722
rect 12114 8666 12170 8722
rect 10254 8542 10310 8598
rect 10378 8542 10434 8598
rect 10502 8542 10558 8598
rect 10626 8542 10682 8598
rect 10750 8542 10806 8598
rect 10874 8542 10930 8598
rect 10998 8542 11054 8598
rect 11122 8542 11178 8598
rect 11246 8542 11302 8598
rect 11370 8542 11426 8598
rect 11494 8542 11550 8598
rect 11618 8542 11674 8598
rect 11742 8542 11798 8598
rect 11866 8542 11922 8598
rect 11990 8542 12046 8598
rect 12114 8542 12170 8598
rect 10254 8418 10310 8474
rect 10378 8418 10434 8474
rect 10502 8418 10558 8474
rect 10626 8418 10682 8474
rect 10750 8418 10806 8474
rect 10874 8418 10930 8474
rect 10998 8418 11054 8474
rect 11122 8418 11178 8474
rect 11246 8418 11302 8474
rect 11370 8418 11426 8474
rect 11494 8418 11550 8474
rect 11618 8418 11674 8474
rect 11742 8418 11798 8474
rect 11866 8418 11922 8474
rect 11990 8418 12046 8474
rect 12114 8418 12170 8474
rect 10254 8294 10310 8350
rect 10378 8294 10434 8350
rect 10502 8294 10558 8350
rect 10626 8294 10682 8350
rect 10750 8294 10806 8350
rect 10874 8294 10930 8350
rect 10998 8294 11054 8350
rect 11122 8294 11178 8350
rect 11246 8294 11302 8350
rect 11370 8294 11426 8350
rect 11494 8294 11550 8350
rect 11618 8294 11674 8350
rect 11742 8294 11798 8350
rect 11866 8294 11922 8350
rect 11990 8294 12046 8350
rect 12114 8294 12170 8350
rect 10254 8170 10310 8226
rect 10378 8170 10434 8226
rect 10502 8170 10558 8226
rect 10626 8170 10682 8226
rect 10750 8170 10806 8226
rect 10874 8170 10930 8226
rect 10998 8170 11054 8226
rect 11122 8170 11178 8226
rect 11246 8170 11302 8226
rect 11370 8170 11426 8226
rect 11494 8170 11550 8226
rect 11618 8170 11674 8226
rect 11742 8170 11798 8226
rect 11866 8170 11922 8226
rect 11990 8170 12046 8226
rect 12114 8170 12170 8226
rect 10254 8046 10310 8102
rect 10378 8046 10434 8102
rect 10502 8046 10558 8102
rect 10626 8046 10682 8102
rect 10750 8046 10806 8102
rect 10874 8046 10930 8102
rect 10998 8046 11054 8102
rect 11122 8046 11178 8102
rect 11246 8046 11302 8102
rect 11370 8046 11426 8102
rect 11494 8046 11550 8102
rect 11618 8046 11674 8102
rect 11742 8046 11798 8102
rect 11866 8046 11922 8102
rect 11990 8046 12046 8102
rect 12114 8046 12170 8102
rect 12871 10898 12927 10954
rect 12995 10898 13051 10954
rect 13119 10898 13175 10954
rect 13243 10898 13299 10954
rect 13367 10898 13423 10954
rect 13491 10898 13547 10954
rect 13615 10898 13671 10954
rect 13739 10898 13795 10954
rect 13863 10898 13919 10954
rect 13987 10898 14043 10954
rect 14111 10898 14167 10954
rect 14235 10898 14291 10954
rect 14359 10898 14415 10954
rect 14483 10898 14539 10954
rect 14607 10898 14663 10954
rect 12871 10774 12927 10830
rect 12995 10774 13051 10830
rect 13119 10774 13175 10830
rect 13243 10774 13299 10830
rect 13367 10774 13423 10830
rect 13491 10774 13547 10830
rect 13615 10774 13671 10830
rect 13739 10774 13795 10830
rect 13863 10774 13919 10830
rect 13987 10774 14043 10830
rect 14111 10774 14167 10830
rect 14235 10774 14291 10830
rect 14359 10774 14415 10830
rect 14483 10774 14539 10830
rect 14607 10774 14663 10830
rect 12871 10650 12927 10706
rect 12995 10650 13051 10706
rect 13119 10650 13175 10706
rect 13243 10650 13299 10706
rect 13367 10650 13423 10706
rect 13491 10650 13547 10706
rect 13615 10650 13671 10706
rect 13739 10650 13795 10706
rect 13863 10650 13919 10706
rect 13987 10650 14043 10706
rect 14111 10650 14167 10706
rect 14235 10650 14291 10706
rect 14359 10650 14415 10706
rect 14483 10650 14539 10706
rect 14607 10650 14663 10706
rect 12871 10526 12927 10582
rect 12995 10526 13051 10582
rect 13119 10526 13175 10582
rect 13243 10526 13299 10582
rect 13367 10526 13423 10582
rect 13491 10526 13547 10582
rect 13615 10526 13671 10582
rect 13739 10526 13795 10582
rect 13863 10526 13919 10582
rect 13987 10526 14043 10582
rect 14111 10526 14167 10582
rect 14235 10526 14291 10582
rect 14359 10526 14415 10582
rect 14483 10526 14539 10582
rect 14607 10526 14663 10582
rect 12871 10402 12927 10458
rect 12995 10402 13051 10458
rect 13119 10402 13175 10458
rect 13243 10402 13299 10458
rect 13367 10402 13423 10458
rect 13491 10402 13547 10458
rect 13615 10402 13671 10458
rect 13739 10402 13795 10458
rect 13863 10402 13919 10458
rect 13987 10402 14043 10458
rect 14111 10402 14167 10458
rect 14235 10402 14291 10458
rect 14359 10402 14415 10458
rect 14483 10402 14539 10458
rect 14607 10402 14663 10458
rect 12871 10278 12927 10334
rect 12995 10278 13051 10334
rect 13119 10278 13175 10334
rect 13243 10278 13299 10334
rect 13367 10278 13423 10334
rect 13491 10278 13547 10334
rect 13615 10278 13671 10334
rect 13739 10278 13795 10334
rect 13863 10278 13919 10334
rect 13987 10278 14043 10334
rect 14111 10278 14167 10334
rect 14235 10278 14291 10334
rect 14359 10278 14415 10334
rect 14483 10278 14539 10334
rect 14607 10278 14663 10334
rect 12871 10154 12927 10210
rect 12995 10154 13051 10210
rect 13119 10154 13175 10210
rect 13243 10154 13299 10210
rect 13367 10154 13423 10210
rect 13491 10154 13547 10210
rect 13615 10154 13671 10210
rect 13739 10154 13795 10210
rect 13863 10154 13919 10210
rect 13987 10154 14043 10210
rect 14111 10154 14167 10210
rect 14235 10154 14291 10210
rect 14359 10154 14415 10210
rect 14483 10154 14539 10210
rect 14607 10154 14663 10210
rect 12871 10030 12927 10086
rect 12995 10030 13051 10086
rect 13119 10030 13175 10086
rect 13243 10030 13299 10086
rect 13367 10030 13423 10086
rect 13491 10030 13547 10086
rect 13615 10030 13671 10086
rect 13739 10030 13795 10086
rect 13863 10030 13919 10086
rect 13987 10030 14043 10086
rect 14111 10030 14167 10086
rect 14235 10030 14291 10086
rect 14359 10030 14415 10086
rect 14483 10030 14539 10086
rect 14607 10030 14663 10086
rect 12871 9906 12927 9962
rect 12995 9906 13051 9962
rect 13119 9906 13175 9962
rect 13243 9906 13299 9962
rect 13367 9906 13423 9962
rect 13491 9906 13547 9962
rect 13615 9906 13671 9962
rect 13739 9906 13795 9962
rect 13863 9906 13919 9962
rect 13987 9906 14043 9962
rect 14111 9906 14167 9962
rect 14235 9906 14291 9962
rect 14359 9906 14415 9962
rect 14483 9906 14539 9962
rect 14607 9906 14663 9962
rect 12871 9782 12927 9838
rect 12995 9782 13051 9838
rect 13119 9782 13175 9838
rect 13243 9782 13299 9838
rect 13367 9782 13423 9838
rect 13491 9782 13547 9838
rect 13615 9782 13671 9838
rect 13739 9782 13795 9838
rect 13863 9782 13919 9838
rect 13987 9782 14043 9838
rect 14111 9782 14167 9838
rect 14235 9782 14291 9838
rect 14359 9782 14415 9838
rect 14483 9782 14539 9838
rect 14607 9782 14663 9838
rect 12871 9658 12927 9714
rect 12995 9658 13051 9714
rect 13119 9658 13175 9714
rect 13243 9658 13299 9714
rect 13367 9658 13423 9714
rect 13491 9658 13547 9714
rect 13615 9658 13671 9714
rect 13739 9658 13795 9714
rect 13863 9658 13919 9714
rect 13987 9658 14043 9714
rect 14111 9658 14167 9714
rect 14235 9658 14291 9714
rect 14359 9658 14415 9714
rect 14483 9658 14539 9714
rect 14607 9658 14663 9714
rect 12871 9534 12927 9590
rect 12995 9534 13051 9590
rect 13119 9534 13175 9590
rect 13243 9534 13299 9590
rect 13367 9534 13423 9590
rect 13491 9534 13547 9590
rect 13615 9534 13671 9590
rect 13739 9534 13795 9590
rect 13863 9534 13919 9590
rect 13987 9534 14043 9590
rect 14111 9534 14167 9590
rect 14235 9534 14291 9590
rect 14359 9534 14415 9590
rect 14483 9534 14539 9590
rect 14607 9534 14663 9590
rect 12871 9410 12927 9466
rect 12995 9410 13051 9466
rect 13119 9410 13175 9466
rect 13243 9410 13299 9466
rect 13367 9410 13423 9466
rect 13491 9410 13547 9466
rect 13615 9410 13671 9466
rect 13739 9410 13795 9466
rect 13863 9410 13919 9466
rect 13987 9410 14043 9466
rect 14111 9410 14167 9466
rect 14235 9410 14291 9466
rect 14359 9410 14415 9466
rect 14483 9410 14539 9466
rect 14607 9410 14663 9466
rect 12871 9286 12927 9342
rect 12995 9286 13051 9342
rect 13119 9286 13175 9342
rect 13243 9286 13299 9342
rect 13367 9286 13423 9342
rect 13491 9286 13547 9342
rect 13615 9286 13671 9342
rect 13739 9286 13795 9342
rect 13863 9286 13919 9342
rect 13987 9286 14043 9342
rect 14111 9286 14167 9342
rect 14235 9286 14291 9342
rect 14359 9286 14415 9342
rect 14483 9286 14539 9342
rect 14607 9286 14663 9342
rect 12871 9162 12927 9218
rect 12995 9162 13051 9218
rect 13119 9162 13175 9218
rect 13243 9162 13299 9218
rect 13367 9162 13423 9218
rect 13491 9162 13547 9218
rect 13615 9162 13671 9218
rect 13739 9162 13795 9218
rect 13863 9162 13919 9218
rect 13987 9162 14043 9218
rect 14111 9162 14167 9218
rect 14235 9162 14291 9218
rect 14359 9162 14415 9218
rect 14483 9162 14539 9218
rect 14607 9162 14663 9218
rect 12871 9038 12927 9094
rect 12995 9038 13051 9094
rect 13119 9038 13175 9094
rect 13243 9038 13299 9094
rect 13367 9038 13423 9094
rect 13491 9038 13547 9094
rect 13615 9038 13671 9094
rect 13739 9038 13795 9094
rect 13863 9038 13919 9094
rect 13987 9038 14043 9094
rect 14111 9038 14167 9094
rect 14235 9038 14291 9094
rect 14359 9038 14415 9094
rect 14483 9038 14539 9094
rect 14607 9038 14663 9094
rect 12871 8914 12927 8970
rect 12995 8914 13051 8970
rect 13119 8914 13175 8970
rect 13243 8914 13299 8970
rect 13367 8914 13423 8970
rect 13491 8914 13547 8970
rect 13615 8914 13671 8970
rect 13739 8914 13795 8970
rect 13863 8914 13919 8970
rect 13987 8914 14043 8970
rect 14111 8914 14167 8970
rect 14235 8914 14291 8970
rect 14359 8914 14415 8970
rect 14483 8914 14539 8970
rect 14607 8914 14663 8970
rect 12871 8790 12927 8846
rect 12995 8790 13051 8846
rect 13119 8790 13175 8846
rect 13243 8790 13299 8846
rect 13367 8790 13423 8846
rect 13491 8790 13547 8846
rect 13615 8790 13671 8846
rect 13739 8790 13795 8846
rect 13863 8790 13919 8846
rect 13987 8790 14043 8846
rect 14111 8790 14167 8846
rect 14235 8790 14291 8846
rect 14359 8790 14415 8846
rect 14483 8790 14539 8846
rect 14607 8790 14663 8846
rect 12871 8666 12927 8722
rect 12995 8666 13051 8722
rect 13119 8666 13175 8722
rect 13243 8666 13299 8722
rect 13367 8666 13423 8722
rect 13491 8666 13547 8722
rect 13615 8666 13671 8722
rect 13739 8666 13795 8722
rect 13863 8666 13919 8722
rect 13987 8666 14043 8722
rect 14111 8666 14167 8722
rect 14235 8666 14291 8722
rect 14359 8666 14415 8722
rect 14483 8666 14539 8722
rect 14607 8666 14663 8722
rect 12871 8542 12927 8598
rect 12995 8542 13051 8598
rect 13119 8542 13175 8598
rect 13243 8542 13299 8598
rect 13367 8542 13423 8598
rect 13491 8542 13547 8598
rect 13615 8542 13671 8598
rect 13739 8542 13795 8598
rect 13863 8542 13919 8598
rect 13987 8542 14043 8598
rect 14111 8542 14167 8598
rect 14235 8542 14291 8598
rect 14359 8542 14415 8598
rect 14483 8542 14539 8598
rect 14607 8542 14663 8598
rect 12871 8418 12927 8474
rect 12995 8418 13051 8474
rect 13119 8418 13175 8474
rect 13243 8418 13299 8474
rect 13367 8418 13423 8474
rect 13491 8418 13547 8474
rect 13615 8418 13671 8474
rect 13739 8418 13795 8474
rect 13863 8418 13919 8474
rect 13987 8418 14043 8474
rect 14111 8418 14167 8474
rect 14235 8418 14291 8474
rect 14359 8418 14415 8474
rect 14483 8418 14539 8474
rect 14607 8418 14663 8474
rect 12871 8294 12927 8350
rect 12995 8294 13051 8350
rect 13119 8294 13175 8350
rect 13243 8294 13299 8350
rect 13367 8294 13423 8350
rect 13491 8294 13547 8350
rect 13615 8294 13671 8350
rect 13739 8294 13795 8350
rect 13863 8294 13919 8350
rect 13987 8294 14043 8350
rect 14111 8294 14167 8350
rect 14235 8294 14291 8350
rect 14359 8294 14415 8350
rect 14483 8294 14539 8350
rect 14607 8294 14663 8350
rect 12871 8170 12927 8226
rect 12995 8170 13051 8226
rect 13119 8170 13175 8226
rect 13243 8170 13299 8226
rect 13367 8170 13423 8226
rect 13491 8170 13547 8226
rect 13615 8170 13671 8226
rect 13739 8170 13795 8226
rect 13863 8170 13919 8226
rect 13987 8170 14043 8226
rect 14111 8170 14167 8226
rect 14235 8170 14291 8226
rect 14359 8170 14415 8226
rect 14483 8170 14539 8226
rect 14607 8170 14663 8226
rect 12871 8046 12927 8102
rect 12995 8046 13051 8102
rect 13119 8046 13175 8102
rect 13243 8046 13299 8102
rect 13367 8046 13423 8102
rect 13491 8046 13547 8102
rect 13615 8046 13671 8102
rect 13739 8046 13795 8102
rect 13863 8046 13919 8102
rect 13987 8046 14043 8102
rect 14111 8046 14167 8102
rect 14235 8046 14291 8102
rect 14359 8046 14415 8102
rect 14483 8046 14539 8102
rect 14607 8046 14663 8102
rect 14902 10984 14958 10986
rect 14902 10932 14904 10984
rect 14904 10932 14956 10984
rect 14956 10932 14958 10984
rect 14902 10876 14958 10932
rect 14902 10824 14904 10876
rect 14904 10824 14956 10876
rect 14956 10824 14958 10876
rect 14902 10768 14958 10824
rect 14902 10716 14904 10768
rect 14904 10716 14956 10768
rect 14956 10716 14958 10768
rect 14902 10660 14958 10716
rect 14902 10608 14904 10660
rect 14904 10608 14956 10660
rect 14956 10608 14958 10660
rect 14902 10552 14958 10608
rect 14902 10500 14904 10552
rect 14904 10500 14956 10552
rect 14956 10500 14958 10552
rect 14902 10444 14958 10500
rect 14902 10392 14904 10444
rect 14904 10392 14956 10444
rect 14956 10392 14958 10444
rect 14902 10336 14958 10392
rect 14902 10284 14904 10336
rect 14904 10284 14956 10336
rect 14956 10284 14958 10336
rect 14902 10228 14958 10284
rect 14902 10176 14904 10228
rect 14904 10176 14956 10228
rect 14956 10176 14958 10228
rect 14902 10120 14958 10176
rect 14902 10068 14904 10120
rect 14904 10068 14956 10120
rect 14956 10068 14958 10120
rect 14902 10012 14958 10068
rect 14902 9960 14904 10012
rect 14904 9960 14956 10012
rect 14956 9960 14958 10012
rect 14902 9904 14958 9960
rect 14902 9852 14904 9904
rect 14904 9852 14956 9904
rect 14956 9852 14958 9904
rect 14902 9796 14958 9852
rect 14902 9744 14904 9796
rect 14904 9744 14956 9796
rect 14956 9744 14958 9796
rect 14902 9688 14958 9744
rect 14902 9636 14904 9688
rect 14904 9636 14956 9688
rect 14956 9636 14958 9688
rect 14902 9580 14958 9636
rect 14902 9528 14904 9580
rect 14904 9528 14956 9580
rect 14956 9528 14958 9580
rect 14902 9472 14958 9528
rect 14902 9420 14904 9472
rect 14904 9420 14956 9472
rect 14956 9420 14958 9472
rect 14902 9364 14958 9420
rect 14902 9312 14904 9364
rect 14904 9312 14956 9364
rect 14956 9312 14958 9364
rect 14902 9256 14958 9312
rect 14902 9204 14904 9256
rect 14904 9204 14956 9256
rect 14956 9204 14958 9256
rect 14902 9148 14958 9204
rect 14902 9096 14904 9148
rect 14904 9096 14956 9148
rect 14956 9096 14958 9148
rect 14902 9040 14958 9096
rect 14902 8988 14904 9040
rect 14904 8988 14956 9040
rect 14956 8988 14958 9040
rect 14902 8932 14958 8988
rect 14902 8880 14904 8932
rect 14904 8880 14956 8932
rect 14956 8880 14958 8932
rect 14902 8824 14958 8880
rect 14902 8772 14904 8824
rect 14904 8772 14956 8824
rect 14956 8772 14958 8824
rect 14902 8716 14958 8772
rect 14902 8664 14904 8716
rect 14904 8664 14956 8716
rect 14956 8664 14958 8716
rect 14902 8608 14958 8664
rect 14902 8556 14904 8608
rect 14904 8556 14956 8608
rect 14956 8556 14958 8608
rect 14902 8500 14958 8556
rect 14902 8448 14904 8500
rect 14904 8448 14956 8500
rect 14956 8448 14958 8500
rect 14902 8392 14958 8448
rect 14902 8340 14904 8392
rect 14904 8340 14956 8392
rect 14956 8340 14958 8392
rect 14902 8284 14958 8340
rect 14902 8232 14904 8284
rect 14904 8232 14956 8284
rect 14956 8232 14958 8284
rect 14902 8176 14958 8232
rect 14902 8124 14904 8176
rect 14904 8124 14956 8176
rect 14956 8124 14958 8176
rect 14902 8068 14958 8124
rect 14902 8016 14904 8068
rect 14904 8016 14956 8068
rect 14956 8016 14958 8068
rect 14902 8014 14958 8016
rect 20 7784 76 7786
rect 20 7732 22 7784
rect 22 7732 74 7784
rect 74 7732 76 7784
rect 20 7676 76 7732
rect 20 7624 22 7676
rect 22 7624 74 7676
rect 74 7624 76 7676
rect 20 7568 76 7624
rect 20 7516 22 7568
rect 22 7516 74 7568
rect 74 7516 76 7568
rect 20 7460 76 7516
rect 20 7408 22 7460
rect 22 7408 74 7460
rect 74 7408 76 7460
rect 20 7352 76 7408
rect 20 7300 22 7352
rect 22 7300 74 7352
rect 74 7300 76 7352
rect 20 7244 76 7300
rect 20 7192 22 7244
rect 22 7192 74 7244
rect 74 7192 76 7244
rect 20 7136 76 7192
rect 20 7084 22 7136
rect 22 7084 74 7136
rect 74 7084 76 7136
rect 20 7028 76 7084
rect 20 6976 22 7028
rect 22 6976 74 7028
rect 74 6976 76 7028
rect 20 6920 76 6976
rect 20 6868 22 6920
rect 22 6868 74 6920
rect 74 6868 76 6920
rect 20 6812 76 6868
rect 20 6760 22 6812
rect 22 6760 74 6812
rect 74 6760 76 6812
rect 20 6704 76 6760
rect 20 6652 22 6704
rect 22 6652 74 6704
rect 74 6652 76 6704
rect 20 6596 76 6652
rect 20 6544 22 6596
rect 22 6544 74 6596
rect 74 6544 76 6596
rect 20 6488 76 6544
rect 20 6436 22 6488
rect 22 6436 74 6488
rect 74 6436 76 6488
rect 20 6380 76 6436
rect 20 6328 22 6380
rect 22 6328 74 6380
rect 74 6328 76 6380
rect 20 6272 76 6328
rect 20 6220 22 6272
rect 22 6220 74 6272
rect 74 6220 76 6272
rect 20 6164 76 6220
rect 20 6112 22 6164
rect 22 6112 74 6164
rect 74 6112 76 6164
rect 20 6056 76 6112
rect 20 6004 22 6056
rect 22 6004 74 6056
rect 74 6004 76 6056
rect 20 5948 76 6004
rect 20 5896 22 5948
rect 22 5896 74 5948
rect 74 5896 76 5948
rect 20 5840 76 5896
rect 20 5788 22 5840
rect 22 5788 74 5840
rect 74 5788 76 5840
rect 20 5732 76 5788
rect 20 5680 22 5732
rect 22 5680 74 5732
rect 74 5680 76 5732
rect 20 5624 76 5680
rect 20 5572 22 5624
rect 22 5572 74 5624
rect 74 5572 76 5624
rect 20 5516 76 5572
rect 20 5464 22 5516
rect 22 5464 74 5516
rect 74 5464 76 5516
rect 20 5408 76 5464
rect 20 5356 22 5408
rect 22 5356 74 5408
rect 74 5356 76 5408
rect 20 5300 76 5356
rect 20 5248 22 5300
rect 22 5248 74 5300
rect 74 5248 76 5300
rect 20 5192 76 5248
rect 20 5140 22 5192
rect 22 5140 74 5192
rect 74 5140 76 5192
rect 20 5084 76 5140
rect 20 5032 22 5084
rect 22 5032 74 5084
rect 74 5032 76 5084
rect 20 4976 76 5032
rect 20 4924 22 4976
rect 22 4924 74 4976
rect 74 4924 76 4976
rect 20 4868 76 4924
rect 20 4816 22 4868
rect 22 4816 74 4868
rect 74 4816 76 4868
rect 20 4814 76 4816
rect 315 7698 371 7754
rect 439 7698 495 7754
rect 563 7698 619 7754
rect 687 7698 743 7754
rect 811 7698 867 7754
rect 935 7698 991 7754
rect 1059 7698 1115 7754
rect 1183 7698 1239 7754
rect 1307 7698 1363 7754
rect 1431 7698 1487 7754
rect 1555 7698 1611 7754
rect 1679 7698 1735 7754
rect 1803 7698 1859 7754
rect 1927 7698 1983 7754
rect 2051 7698 2107 7754
rect 315 7574 371 7630
rect 439 7574 495 7630
rect 563 7574 619 7630
rect 687 7574 743 7630
rect 811 7574 867 7630
rect 935 7574 991 7630
rect 1059 7574 1115 7630
rect 1183 7574 1239 7630
rect 1307 7574 1363 7630
rect 1431 7574 1487 7630
rect 1555 7574 1611 7630
rect 1679 7574 1735 7630
rect 1803 7574 1859 7630
rect 1927 7574 1983 7630
rect 2051 7574 2107 7630
rect 315 7450 371 7506
rect 439 7450 495 7506
rect 563 7450 619 7506
rect 687 7450 743 7506
rect 811 7450 867 7506
rect 935 7450 991 7506
rect 1059 7450 1115 7506
rect 1183 7450 1239 7506
rect 1307 7450 1363 7506
rect 1431 7450 1487 7506
rect 1555 7450 1611 7506
rect 1679 7450 1735 7506
rect 1803 7450 1859 7506
rect 1927 7450 1983 7506
rect 2051 7450 2107 7506
rect 315 7326 371 7382
rect 439 7326 495 7382
rect 563 7326 619 7382
rect 687 7326 743 7382
rect 811 7326 867 7382
rect 935 7326 991 7382
rect 1059 7326 1115 7382
rect 1183 7326 1239 7382
rect 1307 7326 1363 7382
rect 1431 7326 1487 7382
rect 1555 7326 1611 7382
rect 1679 7326 1735 7382
rect 1803 7326 1859 7382
rect 1927 7326 1983 7382
rect 2051 7326 2107 7382
rect 315 7202 371 7258
rect 439 7202 495 7258
rect 563 7202 619 7258
rect 687 7202 743 7258
rect 811 7202 867 7258
rect 935 7202 991 7258
rect 1059 7202 1115 7258
rect 1183 7202 1239 7258
rect 1307 7202 1363 7258
rect 1431 7202 1487 7258
rect 1555 7202 1611 7258
rect 1679 7202 1735 7258
rect 1803 7202 1859 7258
rect 1927 7202 1983 7258
rect 2051 7202 2107 7258
rect 315 7078 371 7134
rect 439 7078 495 7134
rect 563 7078 619 7134
rect 687 7078 743 7134
rect 811 7078 867 7134
rect 935 7078 991 7134
rect 1059 7078 1115 7134
rect 1183 7078 1239 7134
rect 1307 7078 1363 7134
rect 1431 7078 1487 7134
rect 1555 7078 1611 7134
rect 1679 7078 1735 7134
rect 1803 7078 1859 7134
rect 1927 7078 1983 7134
rect 2051 7078 2107 7134
rect 315 6954 371 7010
rect 439 6954 495 7010
rect 563 6954 619 7010
rect 687 6954 743 7010
rect 811 6954 867 7010
rect 935 6954 991 7010
rect 1059 6954 1115 7010
rect 1183 6954 1239 7010
rect 1307 6954 1363 7010
rect 1431 6954 1487 7010
rect 1555 6954 1611 7010
rect 1679 6954 1735 7010
rect 1803 6954 1859 7010
rect 1927 6954 1983 7010
rect 2051 6954 2107 7010
rect 315 6830 371 6886
rect 439 6830 495 6886
rect 563 6830 619 6886
rect 687 6830 743 6886
rect 811 6830 867 6886
rect 935 6830 991 6886
rect 1059 6830 1115 6886
rect 1183 6830 1239 6886
rect 1307 6830 1363 6886
rect 1431 6830 1487 6886
rect 1555 6830 1611 6886
rect 1679 6830 1735 6886
rect 1803 6830 1859 6886
rect 1927 6830 1983 6886
rect 2051 6830 2107 6886
rect 315 6706 371 6762
rect 439 6706 495 6762
rect 563 6706 619 6762
rect 687 6706 743 6762
rect 811 6706 867 6762
rect 935 6706 991 6762
rect 1059 6706 1115 6762
rect 1183 6706 1239 6762
rect 1307 6706 1363 6762
rect 1431 6706 1487 6762
rect 1555 6706 1611 6762
rect 1679 6706 1735 6762
rect 1803 6706 1859 6762
rect 1927 6706 1983 6762
rect 2051 6706 2107 6762
rect 315 6582 371 6638
rect 439 6582 495 6638
rect 563 6582 619 6638
rect 687 6582 743 6638
rect 811 6582 867 6638
rect 935 6582 991 6638
rect 1059 6582 1115 6638
rect 1183 6582 1239 6638
rect 1307 6582 1363 6638
rect 1431 6582 1487 6638
rect 1555 6582 1611 6638
rect 1679 6582 1735 6638
rect 1803 6582 1859 6638
rect 1927 6582 1983 6638
rect 2051 6582 2107 6638
rect 315 6458 371 6514
rect 439 6458 495 6514
rect 563 6458 619 6514
rect 687 6458 743 6514
rect 811 6458 867 6514
rect 935 6458 991 6514
rect 1059 6458 1115 6514
rect 1183 6458 1239 6514
rect 1307 6458 1363 6514
rect 1431 6458 1487 6514
rect 1555 6458 1611 6514
rect 1679 6458 1735 6514
rect 1803 6458 1859 6514
rect 1927 6458 1983 6514
rect 2051 6458 2107 6514
rect 315 6334 371 6390
rect 439 6334 495 6390
rect 563 6334 619 6390
rect 687 6334 743 6390
rect 811 6334 867 6390
rect 935 6334 991 6390
rect 1059 6334 1115 6390
rect 1183 6334 1239 6390
rect 1307 6334 1363 6390
rect 1431 6334 1487 6390
rect 1555 6334 1611 6390
rect 1679 6334 1735 6390
rect 1803 6334 1859 6390
rect 1927 6334 1983 6390
rect 2051 6334 2107 6390
rect 315 6210 371 6266
rect 439 6210 495 6266
rect 563 6210 619 6266
rect 687 6210 743 6266
rect 811 6210 867 6266
rect 935 6210 991 6266
rect 1059 6210 1115 6266
rect 1183 6210 1239 6266
rect 1307 6210 1363 6266
rect 1431 6210 1487 6266
rect 1555 6210 1611 6266
rect 1679 6210 1735 6266
rect 1803 6210 1859 6266
rect 1927 6210 1983 6266
rect 2051 6210 2107 6266
rect 315 6086 371 6142
rect 439 6086 495 6142
rect 563 6086 619 6142
rect 687 6086 743 6142
rect 811 6086 867 6142
rect 935 6086 991 6142
rect 1059 6086 1115 6142
rect 1183 6086 1239 6142
rect 1307 6086 1363 6142
rect 1431 6086 1487 6142
rect 1555 6086 1611 6142
rect 1679 6086 1735 6142
rect 1803 6086 1859 6142
rect 1927 6086 1983 6142
rect 2051 6086 2107 6142
rect 315 5962 371 6018
rect 439 5962 495 6018
rect 563 5962 619 6018
rect 687 5962 743 6018
rect 811 5962 867 6018
rect 935 5962 991 6018
rect 1059 5962 1115 6018
rect 1183 5962 1239 6018
rect 1307 5962 1363 6018
rect 1431 5962 1487 6018
rect 1555 5962 1611 6018
rect 1679 5962 1735 6018
rect 1803 5962 1859 6018
rect 1927 5962 1983 6018
rect 2051 5962 2107 6018
rect 315 5838 371 5894
rect 439 5838 495 5894
rect 563 5838 619 5894
rect 687 5838 743 5894
rect 811 5838 867 5894
rect 935 5838 991 5894
rect 1059 5838 1115 5894
rect 1183 5838 1239 5894
rect 1307 5838 1363 5894
rect 1431 5838 1487 5894
rect 1555 5838 1611 5894
rect 1679 5838 1735 5894
rect 1803 5838 1859 5894
rect 1927 5838 1983 5894
rect 2051 5838 2107 5894
rect 315 5714 371 5770
rect 439 5714 495 5770
rect 563 5714 619 5770
rect 687 5714 743 5770
rect 811 5714 867 5770
rect 935 5714 991 5770
rect 1059 5714 1115 5770
rect 1183 5714 1239 5770
rect 1307 5714 1363 5770
rect 1431 5714 1487 5770
rect 1555 5714 1611 5770
rect 1679 5714 1735 5770
rect 1803 5714 1859 5770
rect 1927 5714 1983 5770
rect 2051 5714 2107 5770
rect 315 5590 371 5646
rect 439 5590 495 5646
rect 563 5590 619 5646
rect 687 5590 743 5646
rect 811 5590 867 5646
rect 935 5590 991 5646
rect 1059 5590 1115 5646
rect 1183 5590 1239 5646
rect 1307 5590 1363 5646
rect 1431 5590 1487 5646
rect 1555 5590 1611 5646
rect 1679 5590 1735 5646
rect 1803 5590 1859 5646
rect 1927 5590 1983 5646
rect 2051 5590 2107 5646
rect 315 5466 371 5522
rect 439 5466 495 5522
rect 563 5466 619 5522
rect 687 5466 743 5522
rect 811 5466 867 5522
rect 935 5466 991 5522
rect 1059 5466 1115 5522
rect 1183 5466 1239 5522
rect 1307 5466 1363 5522
rect 1431 5466 1487 5522
rect 1555 5466 1611 5522
rect 1679 5466 1735 5522
rect 1803 5466 1859 5522
rect 1927 5466 1983 5522
rect 2051 5466 2107 5522
rect 315 5342 371 5398
rect 439 5342 495 5398
rect 563 5342 619 5398
rect 687 5342 743 5398
rect 811 5342 867 5398
rect 935 5342 991 5398
rect 1059 5342 1115 5398
rect 1183 5342 1239 5398
rect 1307 5342 1363 5398
rect 1431 5342 1487 5398
rect 1555 5342 1611 5398
rect 1679 5342 1735 5398
rect 1803 5342 1859 5398
rect 1927 5342 1983 5398
rect 2051 5342 2107 5398
rect 315 5218 371 5274
rect 439 5218 495 5274
rect 563 5218 619 5274
rect 687 5218 743 5274
rect 811 5218 867 5274
rect 935 5218 991 5274
rect 1059 5218 1115 5274
rect 1183 5218 1239 5274
rect 1307 5218 1363 5274
rect 1431 5218 1487 5274
rect 1555 5218 1611 5274
rect 1679 5218 1735 5274
rect 1803 5218 1859 5274
rect 1927 5218 1983 5274
rect 2051 5218 2107 5274
rect 315 5094 371 5150
rect 439 5094 495 5150
rect 563 5094 619 5150
rect 687 5094 743 5150
rect 811 5094 867 5150
rect 935 5094 991 5150
rect 1059 5094 1115 5150
rect 1183 5094 1239 5150
rect 1307 5094 1363 5150
rect 1431 5094 1487 5150
rect 1555 5094 1611 5150
rect 1679 5094 1735 5150
rect 1803 5094 1859 5150
rect 1927 5094 1983 5150
rect 2051 5094 2107 5150
rect 315 4970 371 5026
rect 439 4970 495 5026
rect 563 4970 619 5026
rect 687 4970 743 5026
rect 811 4970 867 5026
rect 935 4970 991 5026
rect 1059 4970 1115 5026
rect 1183 4970 1239 5026
rect 1307 4970 1363 5026
rect 1431 4970 1487 5026
rect 1555 4970 1611 5026
rect 1679 4970 1735 5026
rect 1803 4970 1859 5026
rect 1927 4970 1983 5026
rect 2051 4970 2107 5026
rect 315 4846 371 4902
rect 439 4846 495 4902
rect 563 4846 619 4902
rect 687 4846 743 4902
rect 811 4846 867 4902
rect 935 4846 991 4902
rect 1059 4846 1115 4902
rect 1183 4846 1239 4902
rect 1307 4846 1363 4902
rect 1431 4846 1487 4902
rect 1555 4846 1611 4902
rect 1679 4846 1735 4902
rect 1803 4846 1859 4902
rect 1927 4846 1983 4902
rect 2051 4846 2107 4902
rect 2808 7698 2864 7754
rect 2932 7698 2988 7754
rect 3056 7698 3112 7754
rect 3180 7698 3236 7754
rect 3304 7698 3360 7754
rect 3428 7698 3484 7754
rect 3552 7698 3608 7754
rect 3676 7698 3732 7754
rect 3800 7698 3856 7754
rect 3924 7698 3980 7754
rect 4048 7698 4104 7754
rect 4172 7698 4228 7754
rect 4296 7698 4352 7754
rect 4420 7698 4476 7754
rect 4544 7698 4600 7754
rect 4668 7698 4724 7754
rect 2808 7574 2864 7630
rect 2932 7574 2988 7630
rect 3056 7574 3112 7630
rect 3180 7574 3236 7630
rect 3304 7574 3360 7630
rect 3428 7574 3484 7630
rect 3552 7574 3608 7630
rect 3676 7574 3732 7630
rect 3800 7574 3856 7630
rect 3924 7574 3980 7630
rect 4048 7574 4104 7630
rect 4172 7574 4228 7630
rect 4296 7574 4352 7630
rect 4420 7574 4476 7630
rect 4544 7574 4600 7630
rect 4668 7574 4724 7630
rect 2808 7450 2864 7506
rect 2932 7450 2988 7506
rect 3056 7450 3112 7506
rect 3180 7450 3236 7506
rect 3304 7450 3360 7506
rect 3428 7450 3484 7506
rect 3552 7450 3608 7506
rect 3676 7450 3732 7506
rect 3800 7450 3856 7506
rect 3924 7450 3980 7506
rect 4048 7450 4104 7506
rect 4172 7450 4228 7506
rect 4296 7450 4352 7506
rect 4420 7450 4476 7506
rect 4544 7450 4600 7506
rect 4668 7450 4724 7506
rect 2808 7326 2864 7382
rect 2932 7326 2988 7382
rect 3056 7326 3112 7382
rect 3180 7326 3236 7382
rect 3304 7326 3360 7382
rect 3428 7326 3484 7382
rect 3552 7326 3608 7382
rect 3676 7326 3732 7382
rect 3800 7326 3856 7382
rect 3924 7326 3980 7382
rect 4048 7326 4104 7382
rect 4172 7326 4228 7382
rect 4296 7326 4352 7382
rect 4420 7326 4476 7382
rect 4544 7326 4600 7382
rect 4668 7326 4724 7382
rect 2808 7202 2864 7258
rect 2932 7202 2988 7258
rect 3056 7202 3112 7258
rect 3180 7202 3236 7258
rect 3304 7202 3360 7258
rect 3428 7202 3484 7258
rect 3552 7202 3608 7258
rect 3676 7202 3732 7258
rect 3800 7202 3856 7258
rect 3924 7202 3980 7258
rect 4048 7202 4104 7258
rect 4172 7202 4228 7258
rect 4296 7202 4352 7258
rect 4420 7202 4476 7258
rect 4544 7202 4600 7258
rect 4668 7202 4724 7258
rect 2808 7078 2864 7134
rect 2932 7078 2988 7134
rect 3056 7078 3112 7134
rect 3180 7078 3236 7134
rect 3304 7078 3360 7134
rect 3428 7078 3484 7134
rect 3552 7078 3608 7134
rect 3676 7078 3732 7134
rect 3800 7078 3856 7134
rect 3924 7078 3980 7134
rect 4048 7078 4104 7134
rect 4172 7078 4228 7134
rect 4296 7078 4352 7134
rect 4420 7078 4476 7134
rect 4544 7078 4600 7134
rect 4668 7078 4724 7134
rect 2808 6954 2864 7010
rect 2932 6954 2988 7010
rect 3056 6954 3112 7010
rect 3180 6954 3236 7010
rect 3304 6954 3360 7010
rect 3428 6954 3484 7010
rect 3552 6954 3608 7010
rect 3676 6954 3732 7010
rect 3800 6954 3856 7010
rect 3924 6954 3980 7010
rect 4048 6954 4104 7010
rect 4172 6954 4228 7010
rect 4296 6954 4352 7010
rect 4420 6954 4476 7010
rect 4544 6954 4600 7010
rect 4668 6954 4724 7010
rect 2808 6830 2864 6886
rect 2932 6830 2988 6886
rect 3056 6830 3112 6886
rect 3180 6830 3236 6886
rect 3304 6830 3360 6886
rect 3428 6830 3484 6886
rect 3552 6830 3608 6886
rect 3676 6830 3732 6886
rect 3800 6830 3856 6886
rect 3924 6830 3980 6886
rect 4048 6830 4104 6886
rect 4172 6830 4228 6886
rect 4296 6830 4352 6886
rect 4420 6830 4476 6886
rect 4544 6830 4600 6886
rect 4668 6830 4724 6886
rect 2808 6706 2864 6762
rect 2932 6706 2988 6762
rect 3056 6706 3112 6762
rect 3180 6706 3236 6762
rect 3304 6706 3360 6762
rect 3428 6706 3484 6762
rect 3552 6706 3608 6762
rect 3676 6706 3732 6762
rect 3800 6706 3856 6762
rect 3924 6706 3980 6762
rect 4048 6706 4104 6762
rect 4172 6706 4228 6762
rect 4296 6706 4352 6762
rect 4420 6706 4476 6762
rect 4544 6706 4600 6762
rect 4668 6706 4724 6762
rect 2808 6582 2864 6638
rect 2932 6582 2988 6638
rect 3056 6582 3112 6638
rect 3180 6582 3236 6638
rect 3304 6582 3360 6638
rect 3428 6582 3484 6638
rect 3552 6582 3608 6638
rect 3676 6582 3732 6638
rect 3800 6582 3856 6638
rect 3924 6582 3980 6638
rect 4048 6582 4104 6638
rect 4172 6582 4228 6638
rect 4296 6582 4352 6638
rect 4420 6582 4476 6638
rect 4544 6582 4600 6638
rect 4668 6582 4724 6638
rect 2808 6458 2864 6514
rect 2932 6458 2988 6514
rect 3056 6458 3112 6514
rect 3180 6458 3236 6514
rect 3304 6458 3360 6514
rect 3428 6458 3484 6514
rect 3552 6458 3608 6514
rect 3676 6458 3732 6514
rect 3800 6458 3856 6514
rect 3924 6458 3980 6514
rect 4048 6458 4104 6514
rect 4172 6458 4228 6514
rect 4296 6458 4352 6514
rect 4420 6458 4476 6514
rect 4544 6458 4600 6514
rect 4668 6458 4724 6514
rect 2808 6334 2864 6390
rect 2932 6334 2988 6390
rect 3056 6334 3112 6390
rect 3180 6334 3236 6390
rect 3304 6334 3360 6390
rect 3428 6334 3484 6390
rect 3552 6334 3608 6390
rect 3676 6334 3732 6390
rect 3800 6334 3856 6390
rect 3924 6334 3980 6390
rect 4048 6334 4104 6390
rect 4172 6334 4228 6390
rect 4296 6334 4352 6390
rect 4420 6334 4476 6390
rect 4544 6334 4600 6390
rect 4668 6334 4724 6390
rect 2808 6210 2864 6266
rect 2932 6210 2988 6266
rect 3056 6210 3112 6266
rect 3180 6210 3236 6266
rect 3304 6210 3360 6266
rect 3428 6210 3484 6266
rect 3552 6210 3608 6266
rect 3676 6210 3732 6266
rect 3800 6210 3856 6266
rect 3924 6210 3980 6266
rect 4048 6210 4104 6266
rect 4172 6210 4228 6266
rect 4296 6210 4352 6266
rect 4420 6210 4476 6266
rect 4544 6210 4600 6266
rect 4668 6210 4724 6266
rect 2808 6086 2864 6142
rect 2932 6086 2988 6142
rect 3056 6086 3112 6142
rect 3180 6086 3236 6142
rect 3304 6086 3360 6142
rect 3428 6086 3484 6142
rect 3552 6086 3608 6142
rect 3676 6086 3732 6142
rect 3800 6086 3856 6142
rect 3924 6086 3980 6142
rect 4048 6086 4104 6142
rect 4172 6086 4228 6142
rect 4296 6086 4352 6142
rect 4420 6086 4476 6142
rect 4544 6086 4600 6142
rect 4668 6086 4724 6142
rect 2808 5962 2864 6018
rect 2932 5962 2988 6018
rect 3056 5962 3112 6018
rect 3180 5962 3236 6018
rect 3304 5962 3360 6018
rect 3428 5962 3484 6018
rect 3552 5962 3608 6018
rect 3676 5962 3732 6018
rect 3800 5962 3856 6018
rect 3924 5962 3980 6018
rect 4048 5962 4104 6018
rect 4172 5962 4228 6018
rect 4296 5962 4352 6018
rect 4420 5962 4476 6018
rect 4544 5962 4600 6018
rect 4668 5962 4724 6018
rect 2808 5838 2864 5894
rect 2932 5838 2988 5894
rect 3056 5838 3112 5894
rect 3180 5838 3236 5894
rect 3304 5838 3360 5894
rect 3428 5838 3484 5894
rect 3552 5838 3608 5894
rect 3676 5838 3732 5894
rect 3800 5838 3856 5894
rect 3924 5838 3980 5894
rect 4048 5838 4104 5894
rect 4172 5838 4228 5894
rect 4296 5838 4352 5894
rect 4420 5838 4476 5894
rect 4544 5838 4600 5894
rect 4668 5838 4724 5894
rect 2808 5714 2864 5770
rect 2932 5714 2988 5770
rect 3056 5714 3112 5770
rect 3180 5714 3236 5770
rect 3304 5714 3360 5770
rect 3428 5714 3484 5770
rect 3552 5714 3608 5770
rect 3676 5714 3732 5770
rect 3800 5714 3856 5770
rect 3924 5714 3980 5770
rect 4048 5714 4104 5770
rect 4172 5714 4228 5770
rect 4296 5714 4352 5770
rect 4420 5714 4476 5770
rect 4544 5714 4600 5770
rect 4668 5714 4724 5770
rect 2808 5590 2864 5646
rect 2932 5590 2988 5646
rect 3056 5590 3112 5646
rect 3180 5590 3236 5646
rect 3304 5590 3360 5646
rect 3428 5590 3484 5646
rect 3552 5590 3608 5646
rect 3676 5590 3732 5646
rect 3800 5590 3856 5646
rect 3924 5590 3980 5646
rect 4048 5590 4104 5646
rect 4172 5590 4228 5646
rect 4296 5590 4352 5646
rect 4420 5590 4476 5646
rect 4544 5590 4600 5646
rect 4668 5590 4724 5646
rect 2808 5466 2864 5522
rect 2932 5466 2988 5522
rect 3056 5466 3112 5522
rect 3180 5466 3236 5522
rect 3304 5466 3360 5522
rect 3428 5466 3484 5522
rect 3552 5466 3608 5522
rect 3676 5466 3732 5522
rect 3800 5466 3856 5522
rect 3924 5466 3980 5522
rect 4048 5466 4104 5522
rect 4172 5466 4228 5522
rect 4296 5466 4352 5522
rect 4420 5466 4476 5522
rect 4544 5466 4600 5522
rect 4668 5466 4724 5522
rect 2808 5342 2864 5398
rect 2932 5342 2988 5398
rect 3056 5342 3112 5398
rect 3180 5342 3236 5398
rect 3304 5342 3360 5398
rect 3428 5342 3484 5398
rect 3552 5342 3608 5398
rect 3676 5342 3732 5398
rect 3800 5342 3856 5398
rect 3924 5342 3980 5398
rect 4048 5342 4104 5398
rect 4172 5342 4228 5398
rect 4296 5342 4352 5398
rect 4420 5342 4476 5398
rect 4544 5342 4600 5398
rect 4668 5342 4724 5398
rect 2808 5218 2864 5274
rect 2932 5218 2988 5274
rect 3056 5218 3112 5274
rect 3180 5218 3236 5274
rect 3304 5218 3360 5274
rect 3428 5218 3484 5274
rect 3552 5218 3608 5274
rect 3676 5218 3732 5274
rect 3800 5218 3856 5274
rect 3924 5218 3980 5274
rect 4048 5218 4104 5274
rect 4172 5218 4228 5274
rect 4296 5218 4352 5274
rect 4420 5218 4476 5274
rect 4544 5218 4600 5274
rect 4668 5218 4724 5274
rect 2808 5094 2864 5150
rect 2932 5094 2988 5150
rect 3056 5094 3112 5150
rect 3180 5094 3236 5150
rect 3304 5094 3360 5150
rect 3428 5094 3484 5150
rect 3552 5094 3608 5150
rect 3676 5094 3732 5150
rect 3800 5094 3856 5150
rect 3924 5094 3980 5150
rect 4048 5094 4104 5150
rect 4172 5094 4228 5150
rect 4296 5094 4352 5150
rect 4420 5094 4476 5150
rect 4544 5094 4600 5150
rect 4668 5094 4724 5150
rect 2808 4970 2864 5026
rect 2932 4970 2988 5026
rect 3056 4970 3112 5026
rect 3180 4970 3236 5026
rect 3304 4970 3360 5026
rect 3428 4970 3484 5026
rect 3552 4970 3608 5026
rect 3676 4970 3732 5026
rect 3800 4970 3856 5026
rect 3924 4970 3980 5026
rect 4048 4970 4104 5026
rect 4172 4970 4228 5026
rect 4296 4970 4352 5026
rect 4420 4970 4476 5026
rect 4544 4970 4600 5026
rect 4668 4970 4724 5026
rect 2808 4846 2864 4902
rect 2932 4846 2988 4902
rect 3056 4846 3112 4902
rect 3180 4846 3236 4902
rect 3304 4846 3360 4902
rect 3428 4846 3484 4902
rect 3552 4846 3608 4902
rect 3676 4846 3732 4902
rect 3800 4846 3856 4902
rect 3924 4846 3980 4902
rect 4048 4846 4104 4902
rect 4172 4846 4228 4902
rect 4296 4846 4352 4902
rect 4420 4846 4476 4902
rect 4544 4846 4600 4902
rect 4668 4846 4724 4902
rect 5178 7698 5234 7754
rect 5302 7698 5358 7754
rect 5426 7698 5482 7754
rect 5550 7698 5606 7754
rect 5674 7698 5730 7754
rect 5798 7698 5854 7754
rect 5922 7698 5978 7754
rect 6046 7698 6102 7754
rect 6170 7698 6226 7754
rect 6294 7698 6350 7754
rect 6418 7698 6474 7754
rect 6542 7698 6598 7754
rect 6666 7698 6722 7754
rect 6790 7698 6846 7754
rect 6914 7698 6970 7754
rect 7038 7698 7094 7754
rect 5178 7574 5234 7630
rect 5302 7574 5358 7630
rect 5426 7574 5482 7630
rect 5550 7574 5606 7630
rect 5674 7574 5730 7630
rect 5798 7574 5854 7630
rect 5922 7574 5978 7630
rect 6046 7574 6102 7630
rect 6170 7574 6226 7630
rect 6294 7574 6350 7630
rect 6418 7574 6474 7630
rect 6542 7574 6598 7630
rect 6666 7574 6722 7630
rect 6790 7574 6846 7630
rect 6914 7574 6970 7630
rect 7038 7574 7094 7630
rect 5178 7450 5234 7506
rect 5302 7450 5358 7506
rect 5426 7450 5482 7506
rect 5550 7450 5606 7506
rect 5674 7450 5730 7506
rect 5798 7450 5854 7506
rect 5922 7450 5978 7506
rect 6046 7450 6102 7506
rect 6170 7450 6226 7506
rect 6294 7450 6350 7506
rect 6418 7450 6474 7506
rect 6542 7450 6598 7506
rect 6666 7450 6722 7506
rect 6790 7450 6846 7506
rect 6914 7450 6970 7506
rect 7038 7450 7094 7506
rect 5178 7326 5234 7382
rect 5302 7326 5358 7382
rect 5426 7326 5482 7382
rect 5550 7326 5606 7382
rect 5674 7326 5730 7382
rect 5798 7326 5854 7382
rect 5922 7326 5978 7382
rect 6046 7326 6102 7382
rect 6170 7326 6226 7382
rect 6294 7326 6350 7382
rect 6418 7326 6474 7382
rect 6542 7326 6598 7382
rect 6666 7326 6722 7382
rect 6790 7326 6846 7382
rect 6914 7326 6970 7382
rect 7038 7326 7094 7382
rect 5178 7202 5234 7258
rect 5302 7202 5358 7258
rect 5426 7202 5482 7258
rect 5550 7202 5606 7258
rect 5674 7202 5730 7258
rect 5798 7202 5854 7258
rect 5922 7202 5978 7258
rect 6046 7202 6102 7258
rect 6170 7202 6226 7258
rect 6294 7202 6350 7258
rect 6418 7202 6474 7258
rect 6542 7202 6598 7258
rect 6666 7202 6722 7258
rect 6790 7202 6846 7258
rect 6914 7202 6970 7258
rect 7038 7202 7094 7258
rect 5178 7078 5234 7134
rect 5302 7078 5358 7134
rect 5426 7078 5482 7134
rect 5550 7078 5606 7134
rect 5674 7078 5730 7134
rect 5798 7078 5854 7134
rect 5922 7078 5978 7134
rect 6046 7078 6102 7134
rect 6170 7078 6226 7134
rect 6294 7078 6350 7134
rect 6418 7078 6474 7134
rect 6542 7078 6598 7134
rect 6666 7078 6722 7134
rect 6790 7078 6846 7134
rect 6914 7078 6970 7134
rect 7038 7078 7094 7134
rect 5178 6954 5234 7010
rect 5302 6954 5358 7010
rect 5426 6954 5482 7010
rect 5550 6954 5606 7010
rect 5674 6954 5730 7010
rect 5798 6954 5854 7010
rect 5922 6954 5978 7010
rect 6046 6954 6102 7010
rect 6170 6954 6226 7010
rect 6294 6954 6350 7010
rect 6418 6954 6474 7010
rect 6542 6954 6598 7010
rect 6666 6954 6722 7010
rect 6790 6954 6846 7010
rect 6914 6954 6970 7010
rect 7038 6954 7094 7010
rect 5178 6830 5234 6886
rect 5302 6830 5358 6886
rect 5426 6830 5482 6886
rect 5550 6830 5606 6886
rect 5674 6830 5730 6886
rect 5798 6830 5854 6886
rect 5922 6830 5978 6886
rect 6046 6830 6102 6886
rect 6170 6830 6226 6886
rect 6294 6830 6350 6886
rect 6418 6830 6474 6886
rect 6542 6830 6598 6886
rect 6666 6830 6722 6886
rect 6790 6830 6846 6886
rect 6914 6830 6970 6886
rect 7038 6830 7094 6886
rect 5178 6706 5234 6762
rect 5302 6706 5358 6762
rect 5426 6706 5482 6762
rect 5550 6706 5606 6762
rect 5674 6706 5730 6762
rect 5798 6706 5854 6762
rect 5922 6706 5978 6762
rect 6046 6706 6102 6762
rect 6170 6706 6226 6762
rect 6294 6706 6350 6762
rect 6418 6706 6474 6762
rect 6542 6706 6598 6762
rect 6666 6706 6722 6762
rect 6790 6706 6846 6762
rect 6914 6706 6970 6762
rect 7038 6706 7094 6762
rect 5178 6582 5234 6638
rect 5302 6582 5358 6638
rect 5426 6582 5482 6638
rect 5550 6582 5606 6638
rect 5674 6582 5730 6638
rect 5798 6582 5854 6638
rect 5922 6582 5978 6638
rect 6046 6582 6102 6638
rect 6170 6582 6226 6638
rect 6294 6582 6350 6638
rect 6418 6582 6474 6638
rect 6542 6582 6598 6638
rect 6666 6582 6722 6638
rect 6790 6582 6846 6638
rect 6914 6582 6970 6638
rect 7038 6582 7094 6638
rect 5178 6458 5234 6514
rect 5302 6458 5358 6514
rect 5426 6458 5482 6514
rect 5550 6458 5606 6514
rect 5674 6458 5730 6514
rect 5798 6458 5854 6514
rect 5922 6458 5978 6514
rect 6046 6458 6102 6514
rect 6170 6458 6226 6514
rect 6294 6458 6350 6514
rect 6418 6458 6474 6514
rect 6542 6458 6598 6514
rect 6666 6458 6722 6514
rect 6790 6458 6846 6514
rect 6914 6458 6970 6514
rect 7038 6458 7094 6514
rect 5178 6334 5234 6390
rect 5302 6334 5358 6390
rect 5426 6334 5482 6390
rect 5550 6334 5606 6390
rect 5674 6334 5730 6390
rect 5798 6334 5854 6390
rect 5922 6334 5978 6390
rect 6046 6334 6102 6390
rect 6170 6334 6226 6390
rect 6294 6334 6350 6390
rect 6418 6334 6474 6390
rect 6542 6334 6598 6390
rect 6666 6334 6722 6390
rect 6790 6334 6846 6390
rect 6914 6334 6970 6390
rect 7038 6334 7094 6390
rect 5178 6210 5234 6266
rect 5302 6210 5358 6266
rect 5426 6210 5482 6266
rect 5550 6210 5606 6266
rect 5674 6210 5730 6266
rect 5798 6210 5854 6266
rect 5922 6210 5978 6266
rect 6046 6210 6102 6266
rect 6170 6210 6226 6266
rect 6294 6210 6350 6266
rect 6418 6210 6474 6266
rect 6542 6210 6598 6266
rect 6666 6210 6722 6266
rect 6790 6210 6846 6266
rect 6914 6210 6970 6266
rect 7038 6210 7094 6266
rect 5178 6086 5234 6142
rect 5302 6086 5358 6142
rect 5426 6086 5482 6142
rect 5550 6086 5606 6142
rect 5674 6086 5730 6142
rect 5798 6086 5854 6142
rect 5922 6086 5978 6142
rect 6046 6086 6102 6142
rect 6170 6086 6226 6142
rect 6294 6086 6350 6142
rect 6418 6086 6474 6142
rect 6542 6086 6598 6142
rect 6666 6086 6722 6142
rect 6790 6086 6846 6142
rect 6914 6086 6970 6142
rect 7038 6086 7094 6142
rect 5178 5962 5234 6018
rect 5302 5962 5358 6018
rect 5426 5962 5482 6018
rect 5550 5962 5606 6018
rect 5674 5962 5730 6018
rect 5798 5962 5854 6018
rect 5922 5962 5978 6018
rect 6046 5962 6102 6018
rect 6170 5962 6226 6018
rect 6294 5962 6350 6018
rect 6418 5962 6474 6018
rect 6542 5962 6598 6018
rect 6666 5962 6722 6018
rect 6790 5962 6846 6018
rect 6914 5962 6970 6018
rect 7038 5962 7094 6018
rect 5178 5838 5234 5894
rect 5302 5838 5358 5894
rect 5426 5838 5482 5894
rect 5550 5838 5606 5894
rect 5674 5838 5730 5894
rect 5798 5838 5854 5894
rect 5922 5838 5978 5894
rect 6046 5838 6102 5894
rect 6170 5838 6226 5894
rect 6294 5838 6350 5894
rect 6418 5838 6474 5894
rect 6542 5838 6598 5894
rect 6666 5838 6722 5894
rect 6790 5838 6846 5894
rect 6914 5838 6970 5894
rect 7038 5838 7094 5894
rect 5178 5714 5234 5770
rect 5302 5714 5358 5770
rect 5426 5714 5482 5770
rect 5550 5714 5606 5770
rect 5674 5714 5730 5770
rect 5798 5714 5854 5770
rect 5922 5714 5978 5770
rect 6046 5714 6102 5770
rect 6170 5714 6226 5770
rect 6294 5714 6350 5770
rect 6418 5714 6474 5770
rect 6542 5714 6598 5770
rect 6666 5714 6722 5770
rect 6790 5714 6846 5770
rect 6914 5714 6970 5770
rect 7038 5714 7094 5770
rect 5178 5590 5234 5646
rect 5302 5590 5358 5646
rect 5426 5590 5482 5646
rect 5550 5590 5606 5646
rect 5674 5590 5730 5646
rect 5798 5590 5854 5646
rect 5922 5590 5978 5646
rect 6046 5590 6102 5646
rect 6170 5590 6226 5646
rect 6294 5590 6350 5646
rect 6418 5590 6474 5646
rect 6542 5590 6598 5646
rect 6666 5590 6722 5646
rect 6790 5590 6846 5646
rect 6914 5590 6970 5646
rect 7038 5590 7094 5646
rect 5178 5466 5234 5522
rect 5302 5466 5358 5522
rect 5426 5466 5482 5522
rect 5550 5466 5606 5522
rect 5674 5466 5730 5522
rect 5798 5466 5854 5522
rect 5922 5466 5978 5522
rect 6046 5466 6102 5522
rect 6170 5466 6226 5522
rect 6294 5466 6350 5522
rect 6418 5466 6474 5522
rect 6542 5466 6598 5522
rect 6666 5466 6722 5522
rect 6790 5466 6846 5522
rect 6914 5466 6970 5522
rect 7038 5466 7094 5522
rect 5178 5342 5234 5398
rect 5302 5342 5358 5398
rect 5426 5342 5482 5398
rect 5550 5342 5606 5398
rect 5674 5342 5730 5398
rect 5798 5342 5854 5398
rect 5922 5342 5978 5398
rect 6046 5342 6102 5398
rect 6170 5342 6226 5398
rect 6294 5342 6350 5398
rect 6418 5342 6474 5398
rect 6542 5342 6598 5398
rect 6666 5342 6722 5398
rect 6790 5342 6846 5398
rect 6914 5342 6970 5398
rect 7038 5342 7094 5398
rect 5178 5218 5234 5274
rect 5302 5218 5358 5274
rect 5426 5218 5482 5274
rect 5550 5218 5606 5274
rect 5674 5218 5730 5274
rect 5798 5218 5854 5274
rect 5922 5218 5978 5274
rect 6046 5218 6102 5274
rect 6170 5218 6226 5274
rect 6294 5218 6350 5274
rect 6418 5218 6474 5274
rect 6542 5218 6598 5274
rect 6666 5218 6722 5274
rect 6790 5218 6846 5274
rect 6914 5218 6970 5274
rect 7038 5218 7094 5274
rect 5178 5094 5234 5150
rect 5302 5094 5358 5150
rect 5426 5094 5482 5150
rect 5550 5094 5606 5150
rect 5674 5094 5730 5150
rect 5798 5094 5854 5150
rect 5922 5094 5978 5150
rect 6046 5094 6102 5150
rect 6170 5094 6226 5150
rect 6294 5094 6350 5150
rect 6418 5094 6474 5150
rect 6542 5094 6598 5150
rect 6666 5094 6722 5150
rect 6790 5094 6846 5150
rect 6914 5094 6970 5150
rect 7038 5094 7094 5150
rect 5178 4970 5234 5026
rect 5302 4970 5358 5026
rect 5426 4970 5482 5026
rect 5550 4970 5606 5026
rect 5674 4970 5730 5026
rect 5798 4970 5854 5026
rect 5922 4970 5978 5026
rect 6046 4970 6102 5026
rect 6170 4970 6226 5026
rect 6294 4970 6350 5026
rect 6418 4970 6474 5026
rect 6542 4970 6598 5026
rect 6666 4970 6722 5026
rect 6790 4970 6846 5026
rect 6914 4970 6970 5026
rect 7038 4970 7094 5026
rect 5178 4846 5234 4902
rect 5302 4846 5358 4902
rect 5426 4846 5482 4902
rect 5550 4846 5606 4902
rect 5674 4846 5730 4902
rect 5798 4846 5854 4902
rect 5922 4846 5978 4902
rect 6046 4846 6102 4902
rect 6170 4846 6226 4902
rect 6294 4846 6350 4902
rect 6418 4846 6474 4902
rect 6542 4846 6598 4902
rect 6666 4846 6722 4902
rect 6790 4846 6846 4902
rect 6914 4846 6970 4902
rect 7038 4846 7094 4902
rect 7884 7698 7940 7754
rect 8008 7698 8064 7754
rect 8132 7698 8188 7754
rect 8256 7698 8312 7754
rect 8380 7698 8436 7754
rect 8504 7698 8560 7754
rect 8628 7698 8684 7754
rect 8752 7698 8808 7754
rect 8876 7698 8932 7754
rect 9000 7698 9056 7754
rect 9124 7698 9180 7754
rect 9248 7698 9304 7754
rect 9372 7698 9428 7754
rect 9496 7698 9552 7754
rect 9620 7698 9676 7754
rect 9744 7698 9800 7754
rect 7884 7574 7940 7630
rect 8008 7574 8064 7630
rect 8132 7574 8188 7630
rect 8256 7574 8312 7630
rect 8380 7574 8436 7630
rect 8504 7574 8560 7630
rect 8628 7574 8684 7630
rect 8752 7574 8808 7630
rect 8876 7574 8932 7630
rect 9000 7574 9056 7630
rect 9124 7574 9180 7630
rect 9248 7574 9304 7630
rect 9372 7574 9428 7630
rect 9496 7574 9552 7630
rect 9620 7574 9676 7630
rect 9744 7574 9800 7630
rect 7884 7450 7940 7506
rect 8008 7450 8064 7506
rect 8132 7450 8188 7506
rect 8256 7450 8312 7506
rect 8380 7450 8436 7506
rect 8504 7450 8560 7506
rect 8628 7450 8684 7506
rect 8752 7450 8808 7506
rect 8876 7450 8932 7506
rect 9000 7450 9056 7506
rect 9124 7450 9180 7506
rect 9248 7450 9304 7506
rect 9372 7450 9428 7506
rect 9496 7450 9552 7506
rect 9620 7450 9676 7506
rect 9744 7450 9800 7506
rect 7884 7326 7940 7382
rect 8008 7326 8064 7382
rect 8132 7326 8188 7382
rect 8256 7326 8312 7382
rect 8380 7326 8436 7382
rect 8504 7326 8560 7382
rect 8628 7326 8684 7382
rect 8752 7326 8808 7382
rect 8876 7326 8932 7382
rect 9000 7326 9056 7382
rect 9124 7326 9180 7382
rect 9248 7326 9304 7382
rect 9372 7326 9428 7382
rect 9496 7326 9552 7382
rect 9620 7326 9676 7382
rect 9744 7326 9800 7382
rect 7884 7202 7940 7258
rect 8008 7202 8064 7258
rect 8132 7202 8188 7258
rect 8256 7202 8312 7258
rect 8380 7202 8436 7258
rect 8504 7202 8560 7258
rect 8628 7202 8684 7258
rect 8752 7202 8808 7258
rect 8876 7202 8932 7258
rect 9000 7202 9056 7258
rect 9124 7202 9180 7258
rect 9248 7202 9304 7258
rect 9372 7202 9428 7258
rect 9496 7202 9552 7258
rect 9620 7202 9676 7258
rect 9744 7202 9800 7258
rect 7884 7078 7940 7134
rect 8008 7078 8064 7134
rect 8132 7078 8188 7134
rect 8256 7078 8312 7134
rect 8380 7078 8436 7134
rect 8504 7078 8560 7134
rect 8628 7078 8684 7134
rect 8752 7078 8808 7134
rect 8876 7078 8932 7134
rect 9000 7078 9056 7134
rect 9124 7078 9180 7134
rect 9248 7078 9304 7134
rect 9372 7078 9428 7134
rect 9496 7078 9552 7134
rect 9620 7078 9676 7134
rect 9744 7078 9800 7134
rect 7884 6954 7940 7010
rect 8008 6954 8064 7010
rect 8132 6954 8188 7010
rect 8256 6954 8312 7010
rect 8380 6954 8436 7010
rect 8504 6954 8560 7010
rect 8628 6954 8684 7010
rect 8752 6954 8808 7010
rect 8876 6954 8932 7010
rect 9000 6954 9056 7010
rect 9124 6954 9180 7010
rect 9248 6954 9304 7010
rect 9372 6954 9428 7010
rect 9496 6954 9552 7010
rect 9620 6954 9676 7010
rect 9744 6954 9800 7010
rect 7884 6830 7940 6886
rect 8008 6830 8064 6886
rect 8132 6830 8188 6886
rect 8256 6830 8312 6886
rect 8380 6830 8436 6886
rect 8504 6830 8560 6886
rect 8628 6830 8684 6886
rect 8752 6830 8808 6886
rect 8876 6830 8932 6886
rect 9000 6830 9056 6886
rect 9124 6830 9180 6886
rect 9248 6830 9304 6886
rect 9372 6830 9428 6886
rect 9496 6830 9552 6886
rect 9620 6830 9676 6886
rect 9744 6830 9800 6886
rect 7884 6706 7940 6762
rect 8008 6706 8064 6762
rect 8132 6706 8188 6762
rect 8256 6706 8312 6762
rect 8380 6706 8436 6762
rect 8504 6706 8560 6762
rect 8628 6706 8684 6762
rect 8752 6706 8808 6762
rect 8876 6706 8932 6762
rect 9000 6706 9056 6762
rect 9124 6706 9180 6762
rect 9248 6706 9304 6762
rect 9372 6706 9428 6762
rect 9496 6706 9552 6762
rect 9620 6706 9676 6762
rect 9744 6706 9800 6762
rect 7884 6582 7940 6638
rect 8008 6582 8064 6638
rect 8132 6582 8188 6638
rect 8256 6582 8312 6638
rect 8380 6582 8436 6638
rect 8504 6582 8560 6638
rect 8628 6582 8684 6638
rect 8752 6582 8808 6638
rect 8876 6582 8932 6638
rect 9000 6582 9056 6638
rect 9124 6582 9180 6638
rect 9248 6582 9304 6638
rect 9372 6582 9428 6638
rect 9496 6582 9552 6638
rect 9620 6582 9676 6638
rect 9744 6582 9800 6638
rect 7884 6458 7940 6514
rect 8008 6458 8064 6514
rect 8132 6458 8188 6514
rect 8256 6458 8312 6514
rect 8380 6458 8436 6514
rect 8504 6458 8560 6514
rect 8628 6458 8684 6514
rect 8752 6458 8808 6514
rect 8876 6458 8932 6514
rect 9000 6458 9056 6514
rect 9124 6458 9180 6514
rect 9248 6458 9304 6514
rect 9372 6458 9428 6514
rect 9496 6458 9552 6514
rect 9620 6458 9676 6514
rect 9744 6458 9800 6514
rect 7884 6334 7940 6390
rect 8008 6334 8064 6390
rect 8132 6334 8188 6390
rect 8256 6334 8312 6390
rect 8380 6334 8436 6390
rect 8504 6334 8560 6390
rect 8628 6334 8684 6390
rect 8752 6334 8808 6390
rect 8876 6334 8932 6390
rect 9000 6334 9056 6390
rect 9124 6334 9180 6390
rect 9248 6334 9304 6390
rect 9372 6334 9428 6390
rect 9496 6334 9552 6390
rect 9620 6334 9676 6390
rect 9744 6334 9800 6390
rect 7884 6210 7940 6266
rect 8008 6210 8064 6266
rect 8132 6210 8188 6266
rect 8256 6210 8312 6266
rect 8380 6210 8436 6266
rect 8504 6210 8560 6266
rect 8628 6210 8684 6266
rect 8752 6210 8808 6266
rect 8876 6210 8932 6266
rect 9000 6210 9056 6266
rect 9124 6210 9180 6266
rect 9248 6210 9304 6266
rect 9372 6210 9428 6266
rect 9496 6210 9552 6266
rect 9620 6210 9676 6266
rect 9744 6210 9800 6266
rect 7884 6086 7940 6142
rect 8008 6086 8064 6142
rect 8132 6086 8188 6142
rect 8256 6086 8312 6142
rect 8380 6086 8436 6142
rect 8504 6086 8560 6142
rect 8628 6086 8684 6142
rect 8752 6086 8808 6142
rect 8876 6086 8932 6142
rect 9000 6086 9056 6142
rect 9124 6086 9180 6142
rect 9248 6086 9304 6142
rect 9372 6086 9428 6142
rect 9496 6086 9552 6142
rect 9620 6086 9676 6142
rect 9744 6086 9800 6142
rect 7884 5962 7940 6018
rect 8008 5962 8064 6018
rect 8132 5962 8188 6018
rect 8256 5962 8312 6018
rect 8380 5962 8436 6018
rect 8504 5962 8560 6018
rect 8628 5962 8684 6018
rect 8752 5962 8808 6018
rect 8876 5962 8932 6018
rect 9000 5962 9056 6018
rect 9124 5962 9180 6018
rect 9248 5962 9304 6018
rect 9372 5962 9428 6018
rect 9496 5962 9552 6018
rect 9620 5962 9676 6018
rect 9744 5962 9800 6018
rect 7884 5838 7940 5894
rect 8008 5838 8064 5894
rect 8132 5838 8188 5894
rect 8256 5838 8312 5894
rect 8380 5838 8436 5894
rect 8504 5838 8560 5894
rect 8628 5838 8684 5894
rect 8752 5838 8808 5894
rect 8876 5838 8932 5894
rect 9000 5838 9056 5894
rect 9124 5838 9180 5894
rect 9248 5838 9304 5894
rect 9372 5838 9428 5894
rect 9496 5838 9552 5894
rect 9620 5838 9676 5894
rect 9744 5838 9800 5894
rect 7884 5714 7940 5770
rect 8008 5714 8064 5770
rect 8132 5714 8188 5770
rect 8256 5714 8312 5770
rect 8380 5714 8436 5770
rect 8504 5714 8560 5770
rect 8628 5714 8684 5770
rect 8752 5714 8808 5770
rect 8876 5714 8932 5770
rect 9000 5714 9056 5770
rect 9124 5714 9180 5770
rect 9248 5714 9304 5770
rect 9372 5714 9428 5770
rect 9496 5714 9552 5770
rect 9620 5714 9676 5770
rect 9744 5714 9800 5770
rect 7884 5590 7940 5646
rect 8008 5590 8064 5646
rect 8132 5590 8188 5646
rect 8256 5590 8312 5646
rect 8380 5590 8436 5646
rect 8504 5590 8560 5646
rect 8628 5590 8684 5646
rect 8752 5590 8808 5646
rect 8876 5590 8932 5646
rect 9000 5590 9056 5646
rect 9124 5590 9180 5646
rect 9248 5590 9304 5646
rect 9372 5590 9428 5646
rect 9496 5590 9552 5646
rect 9620 5590 9676 5646
rect 9744 5590 9800 5646
rect 7884 5466 7940 5522
rect 8008 5466 8064 5522
rect 8132 5466 8188 5522
rect 8256 5466 8312 5522
rect 8380 5466 8436 5522
rect 8504 5466 8560 5522
rect 8628 5466 8684 5522
rect 8752 5466 8808 5522
rect 8876 5466 8932 5522
rect 9000 5466 9056 5522
rect 9124 5466 9180 5522
rect 9248 5466 9304 5522
rect 9372 5466 9428 5522
rect 9496 5466 9552 5522
rect 9620 5466 9676 5522
rect 9744 5466 9800 5522
rect 7884 5342 7940 5398
rect 8008 5342 8064 5398
rect 8132 5342 8188 5398
rect 8256 5342 8312 5398
rect 8380 5342 8436 5398
rect 8504 5342 8560 5398
rect 8628 5342 8684 5398
rect 8752 5342 8808 5398
rect 8876 5342 8932 5398
rect 9000 5342 9056 5398
rect 9124 5342 9180 5398
rect 9248 5342 9304 5398
rect 9372 5342 9428 5398
rect 9496 5342 9552 5398
rect 9620 5342 9676 5398
rect 9744 5342 9800 5398
rect 7884 5218 7940 5274
rect 8008 5218 8064 5274
rect 8132 5218 8188 5274
rect 8256 5218 8312 5274
rect 8380 5218 8436 5274
rect 8504 5218 8560 5274
rect 8628 5218 8684 5274
rect 8752 5218 8808 5274
rect 8876 5218 8932 5274
rect 9000 5218 9056 5274
rect 9124 5218 9180 5274
rect 9248 5218 9304 5274
rect 9372 5218 9428 5274
rect 9496 5218 9552 5274
rect 9620 5218 9676 5274
rect 9744 5218 9800 5274
rect 7884 5094 7940 5150
rect 8008 5094 8064 5150
rect 8132 5094 8188 5150
rect 8256 5094 8312 5150
rect 8380 5094 8436 5150
rect 8504 5094 8560 5150
rect 8628 5094 8684 5150
rect 8752 5094 8808 5150
rect 8876 5094 8932 5150
rect 9000 5094 9056 5150
rect 9124 5094 9180 5150
rect 9248 5094 9304 5150
rect 9372 5094 9428 5150
rect 9496 5094 9552 5150
rect 9620 5094 9676 5150
rect 9744 5094 9800 5150
rect 7884 4970 7940 5026
rect 8008 4970 8064 5026
rect 8132 4970 8188 5026
rect 8256 4970 8312 5026
rect 8380 4970 8436 5026
rect 8504 4970 8560 5026
rect 8628 4970 8684 5026
rect 8752 4970 8808 5026
rect 8876 4970 8932 5026
rect 9000 4970 9056 5026
rect 9124 4970 9180 5026
rect 9248 4970 9304 5026
rect 9372 4970 9428 5026
rect 9496 4970 9552 5026
rect 9620 4970 9676 5026
rect 9744 4970 9800 5026
rect 7884 4846 7940 4902
rect 8008 4846 8064 4902
rect 8132 4846 8188 4902
rect 8256 4846 8312 4902
rect 8380 4846 8436 4902
rect 8504 4846 8560 4902
rect 8628 4846 8684 4902
rect 8752 4846 8808 4902
rect 8876 4846 8932 4902
rect 9000 4846 9056 4902
rect 9124 4846 9180 4902
rect 9248 4846 9304 4902
rect 9372 4846 9428 4902
rect 9496 4846 9552 4902
rect 9620 4846 9676 4902
rect 9744 4846 9800 4902
rect 10254 7698 10310 7754
rect 10378 7698 10434 7754
rect 10502 7698 10558 7754
rect 10626 7698 10682 7754
rect 10750 7698 10806 7754
rect 10874 7698 10930 7754
rect 10998 7698 11054 7754
rect 11122 7698 11178 7754
rect 11246 7698 11302 7754
rect 11370 7698 11426 7754
rect 11494 7698 11550 7754
rect 11618 7698 11674 7754
rect 11742 7698 11798 7754
rect 11866 7698 11922 7754
rect 11990 7698 12046 7754
rect 12114 7698 12170 7754
rect 10254 7574 10310 7630
rect 10378 7574 10434 7630
rect 10502 7574 10558 7630
rect 10626 7574 10682 7630
rect 10750 7574 10806 7630
rect 10874 7574 10930 7630
rect 10998 7574 11054 7630
rect 11122 7574 11178 7630
rect 11246 7574 11302 7630
rect 11370 7574 11426 7630
rect 11494 7574 11550 7630
rect 11618 7574 11674 7630
rect 11742 7574 11798 7630
rect 11866 7574 11922 7630
rect 11990 7574 12046 7630
rect 12114 7574 12170 7630
rect 10254 7450 10310 7506
rect 10378 7450 10434 7506
rect 10502 7450 10558 7506
rect 10626 7450 10682 7506
rect 10750 7450 10806 7506
rect 10874 7450 10930 7506
rect 10998 7450 11054 7506
rect 11122 7450 11178 7506
rect 11246 7450 11302 7506
rect 11370 7450 11426 7506
rect 11494 7450 11550 7506
rect 11618 7450 11674 7506
rect 11742 7450 11798 7506
rect 11866 7450 11922 7506
rect 11990 7450 12046 7506
rect 12114 7450 12170 7506
rect 10254 7326 10310 7382
rect 10378 7326 10434 7382
rect 10502 7326 10558 7382
rect 10626 7326 10682 7382
rect 10750 7326 10806 7382
rect 10874 7326 10930 7382
rect 10998 7326 11054 7382
rect 11122 7326 11178 7382
rect 11246 7326 11302 7382
rect 11370 7326 11426 7382
rect 11494 7326 11550 7382
rect 11618 7326 11674 7382
rect 11742 7326 11798 7382
rect 11866 7326 11922 7382
rect 11990 7326 12046 7382
rect 12114 7326 12170 7382
rect 10254 7202 10310 7258
rect 10378 7202 10434 7258
rect 10502 7202 10558 7258
rect 10626 7202 10682 7258
rect 10750 7202 10806 7258
rect 10874 7202 10930 7258
rect 10998 7202 11054 7258
rect 11122 7202 11178 7258
rect 11246 7202 11302 7258
rect 11370 7202 11426 7258
rect 11494 7202 11550 7258
rect 11618 7202 11674 7258
rect 11742 7202 11798 7258
rect 11866 7202 11922 7258
rect 11990 7202 12046 7258
rect 12114 7202 12170 7258
rect 10254 7078 10310 7134
rect 10378 7078 10434 7134
rect 10502 7078 10558 7134
rect 10626 7078 10682 7134
rect 10750 7078 10806 7134
rect 10874 7078 10930 7134
rect 10998 7078 11054 7134
rect 11122 7078 11178 7134
rect 11246 7078 11302 7134
rect 11370 7078 11426 7134
rect 11494 7078 11550 7134
rect 11618 7078 11674 7134
rect 11742 7078 11798 7134
rect 11866 7078 11922 7134
rect 11990 7078 12046 7134
rect 12114 7078 12170 7134
rect 10254 6954 10310 7010
rect 10378 6954 10434 7010
rect 10502 6954 10558 7010
rect 10626 6954 10682 7010
rect 10750 6954 10806 7010
rect 10874 6954 10930 7010
rect 10998 6954 11054 7010
rect 11122 6954 11178 7010
rect 11246 6954 11302 7010
rect 11370 6954 11426 7010
rect 11494 6954 11550 7010
rect 11618 6954 11674 7010
rect 11742 6954 11798 7010
rect 11866 6954 11922 7010
rect 11990 6954 12046 7010
rect 12114 6954 12170 7010
rect 10254 6830 10310 6886
rect 10378 6830 10434 6886
rect 10502 6830 10558 6886
rect 10626 6830 10682 6886
rect 10750 6830 10806 6886
rect 10874 6830 10930 6886
rect 10998 6830 11054 6886
rect 11122 6830 11178 6886
rect 11246 6830 11302 6886
rect 11370 6830 11426 6886
rect 11494 6830 11550 6886
rect 11618 6830 11674 6886
rect 11742 6830 11798 6886
rect 11866 6830 11922 6886
rect 11990 6830 12046 6886
rect 12114 6830 12170 6886
rect 10254 6706 10310 6762
rect 10378 6706 10434 6762
rect 10502 6706 10558 6762
rect 10626 6706 10682 6762
rect 10750 6706 10806 6762
rect 10874 6706 10930 6762
rect 10998 6706 11054 6762
rect 11122 6706 11178 6762
rect 11246 6706 11302 6762
rect 11370 6706 11426 6762
rect 11494 6706 11550 6762
rect 11618 6706 11674 6762
rect 11742 6706 11798 6762
rect 11866 6706 11922 6762
rect 11990 6706 12046 6762
rect 12114 6706 12170 6762
rect 10254 6582 10310 6638
rect 10378 6582 10434 6638
rect 10502 6582 10558 6638
rect 10626 6582 10682 6638
rect 10750 6582 10806 6638
rect 10874 6582 10930 6638
rect 10998 6582 11054 6638
rect 11122 6582 11178 6638
rect 11246 6582 11302 6638
rect 11370 6582 11426 6638
rect 11494 6582 11550 6638
rect 11618 6582 11674 6638
rect 11742 6582 11798 6638
rect 11866 6582 11922 6638
rect 11990 6582 12046 6638
rect 12114 6582 12170 6638
rect 10254 6458 10310 6514
rect 10378 6458 10434 6514
rect 10502 6458 10558 6514
rect 10626 6458 10682 6514
rect 10750 6458 10806 6514
rect 10874 6458 10930 6514
rect 10998 6458 11054 6514
rect 11122 6458 11178 6514
rect 11246 6458 11302 6514
rect 11370 6458 11426 6514
rect 11494 6458 11550 6514
rect 11618 6458 11674 6514
rect 11742 6458 11798 6514
rect 11866 6458 11922 6514
rect 11990 6458 12046 6514
rect 12114 6458 12170 6514
rect 10254 6334 10310 6390
rect 10378 6334 10434 6390
rect 10502 6334 10558 6390
rect 10626 6334 10682 6390
rect 10750 6334 10806 6390
rect 10874 6334 10930 6390
rect 10998 6334 11054 6390
rect 11122 6334 11178 6390
rect 11246 6334 11302 6390
rect 11370 6334 11426 6390
rect 11494 6334 11550 6390
rect 11618 6334 11674 6390
rect 11742 6334 11798 6390
rect 11866 6334 11922 6390
rect 11990 6334 12046 6390
rect 12114 6334 12170 6390
rect 10254 6210 10310 6266
rect 10378 6210 10434 6266
rect 10502 6210 10558 6266
rect 10626 6210 10682 6266
rect 10750 6210 10806 6266
rect 10874 6210 10930 6266
rect 10998 6210 11054 6266
rect 11122 6210 11178 6266
rect 11246 6210 11302 6266
rect 11370 6210 11426 6266
rect 11494 6210 11550 6266
rect 11618 6210 11674 6266
rect 11742 6210 11798 6266
rect 11866 6210 11922 6266
rect 11990 6210 12046 6266
rect 12114 6210 12170 6266
rect 10254 6086 10310 6142
rect 10378 6086 10434 6142
rect 10502 6086 10558 6142
rect 10626 6086 10682 6142
rect 10750 6086 10806 6142
rect 10874 6086 10930 6142
rect 10998 6086 11054 6142
rect 11122 6086 11178 6142
rect 11246 6086 11302 6142
rect 11370 6086 11426 6142
rect 11494 6086 11550 6142
rect 11618 6086 11674 6142
rect 11742 6086 11798 6142
rect 11866 6086 11922 6142
rect 11990 6086 12046 6142
rect 12114 6086 12170 6142
rect 10254 5962 10310 6018
rect 10378 5962 10434 6018
rect 10502 5962 10558 6018
rect 10626 5962 10682 6018
rect 10750 5962 10806 6018
rect 10874 5962 10930 6018
rect 10998 5962 11054 6018
rect 11122 5962 11178 6018
rect 11246 5962 11302 6018
rect 11370 5962 11426 6018
rect 11494 5962 11550 6018
rect 11618 5962 11674 6018
rect 11742 5962 11798 6018
rect 11866 5962 11922 6018
rect 11990 5962 12046 6018
rect 12114 5962 12170 6018
rect 10254 5838 10310 5894
rect 10378 5838 10434 5894
rect 10502 5838 10558 5894
rect 10626 5838 10682 5894
rect 10750 5838 10806 5894
rect 10874 5838 10930 5894
rect 10998 5838 11054 5894
rect 11122 5838 11178 5894
rect 11246 5838 11302 5894
rect 11370 5838 11426 5894
rect 11494 5838 11550 5894
rect 11618 5838 11674 5894
rect 11742 5838 11798 5894
rect 11866 5838 11922 5894
rect 11990 5838 12046 5894
rect 12114 5838 12170 5894
rect 10254 5714 10310 5770
rect 10378 5714 10434 5770
rect 10502 5714 10558 5770
rect 10626 5714 10682 5770
rect 10750 5714 10806 5770
rect 10874 5714 10930 5770
rect 10998 5714 11054 5770
rect 11122 5714 11178 5770
rect 11246 5714 11302 5770
rect 11370 5714 11426 5770
rect 11494 5714 11550 5770
rect 11618 5714 11674 5770
rect 11742 5714 11798 5770
rect 11866 5714 11922 5770
rect 11990 5714 12046 5770
rect 12114 5714 12170 5770
rect 10254 5590 10310 5646
rect 10378 5590 10434 5646
rect 10502 5590 10558 5646
rect 10626 5590 10682 5646
rect 10750 5590 10806 5646
rect 10874 5590 10930 5646
rect 10998 5590 11054 5646
rect 11122 5590 11178 5646
rect 11246 5590 11302 5646
rect 11370 5590 11426 5646
rect 11494 5590 11550 5646
rect 11618 5590 11674 5646
rect 11742 5590 11798 5646
rect 11866 5590 11922 5646
rect 11990 5590 12046 5646
rect 12114 5590 12170 5646
rect 10254 5466 10310 5522
rect 10378 5466 10434 5522
rect 10502 5466 10558 5522
rect 10626 5466 10682 5522
rect 10750 5466 10806 5522
rect 10874 5466 10930 5522
rect 10998 5466 11054 5522
rect 11122 5466 11178 5522
rect 11246 5466 11302 5522
rect 11370 5466 11426 5522
rect 11494 5466 11550 5522
rect 11618 5466 11674 5522
rect 11742 5466 11798 5522
rect 11866 5466 11922 5522
rect 11990 5466 12046 5522
rect 12114 5466 12170 5522
rect 10254 5342 10310 5398
rect 10378 5342 10434 5398
rect 10502 5342 10558 5398
rect 10626 5342 10682 5398
rect 10750 5342 10806 5398
rect 10874 5342 10930 5398
rect 10998 5342 11054 5398
rect 11122 5342 11178 5398
rect 11246 5342 11302 5398
rect 11370 5342 11426 5398
rect 11494 5342 11550 5398
rect 11618 5342 11674 5398
rect 11742 5342 11798 5398
rect 11866 5342 11922 5398
rect 11990 5342 12046 5398
rect 12114 5342 12170 5398
rect 10254 5218 10310 5274
rect 10378 5218 10434 5274
rect 10502 5218 10558 5274
rect 10626 5218 10682 5274
rect 10750 5218 10806 5274
rect 10874 5218 10930 5274
rect 10998 5218 11054 5274
rect 11122 5218 11178 5274
rect 11246 5218 11302 5274
rect 11370 5218 11426 5274
rect 11494 5218 11550 5274
rect 11618 5218 11674 5274
rect 11742 5218 11798 5274
rect 11866 5218 11922 5274
rect 11990 5218 12046 5274
rect 12114 5218 12170 5274
rect 10254 5094 10310 5150
rect 10378 5094 10434 5150
rect 10502 5094 10558 5150
rect 10626 5094 10682 5150
rect 10750 5094 10806 5150
rect 10874 5094 10930 5150
rect 10998 5094 11054 5150
rect 11122 5094 11178 5150
rect 11246 5094 11302 5150
rect 11370 5094 11426 5150
rect 11494 5094 11550 5150
rect 11618 5094 11674 5150
rect 11742 5094 11798 5150
rect 11866 5094 11922 5150
rect 11990 5094 12046 5150
rect 12114 5094 12170 5150
rect 10254 4970 10310 5026
rect 10378 4970 10434 5026
rect 10502 4970 10558 5026
rect 10626 4970 10682 5026
rect 10750 4970 10806 5026
rect 10874 4970 10930 5026
rect 10998 4970 11054 5026
rect 11122 4970 11178 5026
rect 11246 4970 11302 5026
rect 11370 4970 11426 5026
rect 11494 4970 11550 5026
rect 11618 4970 11674 5026
rect 11742 4970 11798 5026
rect 11866 4970 11922 5026
rect 11990 4970 12046 5026
rect 12114 4970 12170 5026
rect 10254 4846 10310 4902
rect 10378 4846 10434 4902
rect 10502 4846 10558 4902
rect 10626 4846 10682 4902
rect 10750 4846 10806 4902
rect 10874 4846 10930 4902
rect 10998 4846 11054 4902
rect 11122 4846 11178 4902
rect 11246 4846 11302 4902
rect 11370 4846 11426 4902
rect 11494 4846 11550 4902
rect 11618 4846 11674 4902
rect 11742 4846 11798 4902
rect 11866 4846 11922 4902
rect 11990 4846 12046 4902
rect 12114 4846 12170 4902
rect 12871 7698 12927 7754
rect 12995 7698 13051 7754
rect 13119 7698 13175 7754
rect 13243 7698 13299 7754
rect 13367 7698 13423 7754
rect 13491 7698 13547 7754
rect 13615 7698 13671 7754
rect 13739 7698 13795 7754
rect 13863 7698 13919 7754
rect 13987 7698 14043 7754
rect 14111 7698 14167 7754
rect 14235 7698 14291 7754
rect 14359 7698 14415 7754
rect 14483 7698 14539 7754
rect 14607 7698 14663 7754
rect 12871 7574 12927 7630
rect 12995 7574 13051 7630
rect 13119 7574 13175 7630
rect 13243 7574 13299 7630
rect 13367 7574 13423 7630
rect 13491 7574 13547 7630
rect 13615 7574 13671 7630
rect 13739 7574 13795 7630
rect 13863 7574 13919 7630
rect 13987 7574 14043 7630
rect 14111 7574 14167 7630
rect 14235 7574 14291 7630
rect 14359 7574 14415 7630
rect 14483 7574 14539 7630
rect 14607 7574 14663 7630
rect 12871 7450 12927 7506
rect 12995 7450 13051 7506
rect 13119 7450 13175 7506
rect 13243 7450 13299 7506
rect 13367 7450 13423 7506
rect 13491 7450 13547 7506
rect 13615 7450 13671 7506
rect 13739 7450 13795 7506
rect 13863 7450 13919 7506
rect 13987 7450 14043 7506
rect 14111 7450 14167 7506
rect 14235 7450 14291 7506
rect 14359 7450 14415 7506
rect 14483 7450 14539 7506
rect 14607 7450 14663 7506
rect 12871 7326 12927 7382
rect 12995 7326 13051 7382
rect 13119 7326 13175 7382
rect 13243 7326 13299 7382
rect 13367 7326 13423 7382
rect 13491 7326 13547 7382
rect 13615 7326 13671 7382
rect 13739 7326 13795 7382
rect 13863 7326 13919 7382
rect 13987 7326 14043 7382
rect 14111 7326 14167 7382
rect 14235 7326 14291 7382
rect 14359 7326 14415 7382
rect 14483 7326 14539 7382
rect 14607 7326 14663 7382
rect 12871 7202 12927 7258
rect 12995 7202 13051 7258
rect 13119 7202 13175 7258
rect 13243 7202 13299 7258
rect 13367 7202 13423 7258
rect 13491 7202 13547 7258
rect 13615 7202 13671 7258
rect 13739 7202 13795 7258
rect 13863 7202 13919 7258
rect 13987 7202 14043 7258
rect 14111 7202 14167 7258
rect 14235 7202 14291 7258
rect 14359 7202 14415 7258
rect 14483 7202 14539 7258
rect 14607 7202 14663 7258
rect 12871 7078 12927 7134
rect 12995 7078 13051 7134
rect 13119 7078 13175 7134
rect 13243 7078 13299 7134
rect 13367 7078 13423 7134
rect 13491 7078 13547 7134
rect 13615 7078 13671 7134
rect 13739 7078 13795 7134
rect 13863 7078 13919 7134
rect 13987 7078 14043 7134
rect 14111 7078 14167 7134
rect 14235 7078 14291 7134
rect 14359 7078 14415 7134
rect 14483 7078 14539 7134
rect 14607 7078 14663 7134
rect 12871 6954 12927 7010
rect 12995 6954 13051 7010
rect 13119 6954 13175 7010
rect 13243 6954 13299 7010
rect 13367 6954 13423 7010
rect 13491 6954 13547 7010
rect 13615 6954 13671 7010
rect 13739 6954 13795 7010
rect 13863 6954 13919 7010
rect 13987 6954 14043 7010
rect 14111 6954 14167 7010
rect 14235 6954 14291 7010
rect 14359 6954 14415 7010
rect 14483 6954 14539 7010
rect 14607 6954 14663 7010
rect 12871 6830 12927 6886
rect 12995 6830 13051 6886
rect 13119 6830 13175 6886
rect 13243 6830 13299 6886
rect 13367 6830 13423 6886
rect 13491 6830 13547 6886
rect 13615 6830 13671 6886
rect 13739 6830 13795 6886
rect 13863 6830 13919 6886
rect 13987 6830 14043 6886
rect 14111 6830 14167 6886
rect 14235 6830 14291 6886
rect 14359 6830 14415 6886
rect 14483 6830 14539 6886
rect 14607 6830 14663 6886
rect 12871 6706 12927 6762
rect 12995 6706 13051 6762
rect 13119 6706 13175 6762
rect 13243 6706 13299 6762
rect 13367 6706 13423 6762
rect 13491 6706 13547 6762
rect 13615 6706 13671 6762
rect 13739 6706 13795 6762
rect 13863 6706 13919 6762
rect 13987 6706 14043 6762
rect 14111 6706 14167 6762
rect 14235 6706 14291 6762
rect 14359 6706 14415 6762
rect 14483 6706 14539 6762
rect 14607 6706 14663 6762
rect 12871 6582 12927 6638
rect 12995 6582 13051 6638
rect 13119 6582 13175 6638
rect 13243 6582 13299 6638
rect 13367 6582 13423 6638
rect 13491 6582 13547 6638
rect 13615 6582 13671 6638
rect 13739 6582 13795 6638
rect 13863 6582 13919 6638
rect 13987 6582 14043 6638
rect 14111 6582 14167 6638
rect 14235 6582 14291 6638
rect 14359 6582 14415 6638
rect 14483 6582 14539 6638
rect 14607 6582 14663 6638
rect 12871 6458 12927 6514
rect 12995 6458 13051 6514
rect 13119 6458 13175 6514
rect 13243 6458 13299 6514
rect 13367 6458 13423 6514
rect 13491 6458 13547 6514
rect 13615 6458 13671 6514
rect 13739 6458 13795 6514
rect 13863 6458 13919 6514
rect 13987 6458 14043 6514
rect 14111 6458 14167 6514
rect 14235 6458 14291 6514
rect 14359 6458 14415 6514
rect 14483 6458 14539 6514
rect 14607 6458 14663 6514
rect 12871 6334 12927 6390
rect 12995 6334 13051 6390
rect 13119 6334 13175 6390
rect 13243 6334 13299 6390
rect 13367 6334 13423 6390
rect 13491 6334 13547 6390
rect 13615 6334 13671 6390
rect 13739 6334 13795 6390
rect 13863 6334 13919 6390
rect 13987 6334 14043 6390
rect 14111 6334 14167 6390
rect 14235 6334 14291 6390
rect 14359 6334 14415 6390
rect 14483 6334 14539 6390
rect 14607 6334 14663 6390
rect 12871 6210 12927 6266
rect 12995 6210 13051 6266
rect 13119 6210 13175 6266
rect 13243 6210 13299 6266
rect 13367 6210 13423 6266
rect 13491 6210 13547 6266
rect 13615 6210 13671 6266
rect 13739 6210 13795 6266
rect 13863 6210 13919 6266
rect 13987 6210 14043 6266
rect 14111 6210 14167 6266
rect 14235 6210 14291 6266
rect 14359 6210 14415 6266
rect 14483 6210 14539 6266
rect 14607 6210 14663 6266
rect 12871 6086 12927 6142
rect 12995 6086 13051 6142
rect 13119 6086 13175 6142
rect 13243 6086 13299 6142
rect 13367 6086 13423 6142
rect 13491 6086 13547 6142
rect 13615 6086 13671 6142
rect 13739 6086 13795 6142
rect 13863 6086 13919 6142
rect 13987 6086 14043 6142
rect 14111 6086 14167 6142
rect 14235 6086 14291 6142
rect 14359 6086 14415 6142
rect 14483 6086 14539 6142
rect 14607 6086 14663 6142
rect 12871 5962 12927 6018
rect 12995 5962 13051 6018
rect 13119 5962 13175 6018
rect 13243 5962 13299 6018
rect 13367 5962 13423 6018
rect 13491 5962 13547 6018
rect 13615 5962 13671 6018
rect 13739 5962 13795 6018
rect 13863 5962 13919 6018
rect 13987 5962 14043 6018
rect 14111 5962 14167 6018
rect 14235 5962 14291 6018
rect 14359 5962 14415 6018
rect 14483 5962 14539 6018
rect 14607 5962 14663 6018
rect 12871 5838 12927 5894
rect 12995 5838 13051 5894
rect 13119 5838 13175 5894
rect 13243 5838 13299 5894
rect 13367 5838 13423 5894
rect 13491 5838 13547 5894
rect 13615 5838 13671 5894
rect 13739 5838 13795 5894
rect 13863 5838 13919 5894
rect 13987 5838 14043 5894
rect 14111 5838 14167 5894
rect 14235 5838 14291 5894
rect 14359 5838 14415 5894
rect 14483 5838 14539 5894
rect 14607 5838 14663 5894
rect 12871 5714 12927 5770
rect 12995 5714 13051 5770
rect 13119 5714 13175 5770
rect 13243 5714 13299 5770
rect 13367 5714 13423 5770
rect 13491 5714 13547 5770
rect 13615 5714 13671 5770
rect 13739 5714 13795 5770
rect 13863 5714 13919 5770
rect 13987 5714 14043 5770
rect 14111 5714 14167 5770
rect 14235 5714 14291 5770
rect 14359 5714 14415 5770
rect 14483 5714 14539 5770
rect 14607 5714 14663 5770
rect 12871 5590 12927 5646
rect 12995 5590 13051 5646
rect 13119 5590 13175 5646
rect 13243 5590 13299 5646
rect 13367 5590 13423 5646
rect 13491 5590 13547 5646
rect 13615 5590 13671 5646
rect 13739 5590 13795 5646
rect 13863 5590 13919 5646
rect 13987 5590 14043 5646
rect 14111 5590 14167 5646
rect 14235 5590 14291 5646
rect 14359 5590 14415 5646
rect 14483 5590 14539 5646
rect 14607 5590 14663 5646
rect 12871 5466 12927 5522
rect 12995 5466 13051 5522
rect 13119 5466 13175 5522
rect 13243 5466 13299 5522
rect 13367 5466 13423 5522
rect 13491 5466 13547 5522
rect 13615 5466 13671 5522
rect 13739 5466 13795 5522
rect 13863 5466 13919 5522
rect 13987 5466 14043 5522
rect 14111 5466 14167 5522
rect 14235 5466 14291 5522
rect 14359 5466 14415 5522
rect 14483 5466 14539 5522
rect 14607 5466 14663 5522
rect 12871 5342 12927 5398
rect 12995 5342 13051 5398
rect 13119 5342 13175 5398
rect 13243 5342 13299 5398
rect 13367 5342 13423 5398
rect 13491 5342 13547 5398
rect 13615 5342 13671 5398
rect 13739 5342 13795 5398
rect 13863 5342 13919 5398
rect 13987 5342 14043 5398
rect 14111 5342 14167 5398
rect 14235 5342 14291 5398
rect 14359 5342 14415 5398
rect 14483 5342 14539 5398
rect 14607 5342 14663 5398
rect 12871 5218 12927 5274
rect 12995 5218 13051 5274
rect 13119 5218 13175 5274
rect 13243 5218 13299 5274
rect 13367 5218 13423 5274
rect 13491 5218 13547 5274
rect 13615 5218 13671 5274
rect 13739 5218 13795 5274
rect 13863 5218 13919 5274
rect 13987 5218 14043 5274
rect 14111 5218 14167 5274
rect 14235 5218 14291 5274
rect 14359 5218 14415 5274
rect 14483 5218 14539 5274
rect 14607 5218 14663 5274
rect 12871 5094 12927 5150
rect 12995 5094 13051 5150
rect 13119 5094 13175 5150
rect 13243 5094 13299 5150
rect 13367 5094 13423 5150
rect 13491 5094 13547 5150
rect 13615 5094 13671 5150
rect 13739 5094 13795 5150
rect 13863 5094 13919 5150
rect 13987 5094 14043 5150
rect 14111 5094 14167 5150
rect 14235 5094 14291 5150
rect 14359 5094 14415 5150
rect 14483 5094 14539 5150
rect 14607 5094 14663 5150
rect 12871 4970 12927 5026
rect 12995 4970 13051 5026
rect 13119 4970 13175 5026
rect 13243 4970 13299 5026
rect 13367 4970 13423 5026
rect 13491 4970 13547 5026
rect 13615 4970 13671 5026
rect 13739 4970 13795 5026
rect 13863 4970 13919 5026
rect 13987 4970 14043 5026
rect 14111 4970 14167 5026
rect 14235 4970 14291 5026
rect 14359 4970 14415 5026
rect 14483 4970 14539 5026
rect 14607 4970 14663 5026
rect 12871 4846 12927 4902
rect 12995 4846 13051 4902
rect 13119 4846 13175 4902
rect 13243 4846 13299 4902
rect 13367 4846 13423 4902
rect 13491 4846 13547 4902
rect 13615 4846 13671 4902
rect 13739 4846 13795 4902
rect 13863 4846 13919 4902
rect 13987 4846 14043 4902
rect 14111 4846 14167 4902
rect 14235 4846 14291 4902
rect 14359 4846 14415 4902
rect 14483 4846 14539 4902
rect 14607 4846 14663 4902
rect 14902 7784 14958 7786
rect 14902 7732 14904 7784
rect 14904 7732 14956 7784
rect 14956 7732 14958 7784
rect 14902 7676 14958 7732
rect 14902 7624 14904 7676
rect 14904 7624 14956 7676
rect 14956 7624 14958 7676
rect 14902 7568 14958 7624
rect 14902 7516 14904 7568
rect 14904 7516 14956 7568
rect 14956 7516 14958 7568
rect 14902 7460 14958 7516
rect 14902 7408 14904 7460
rect 14904 7408 14956 7460
rect 14956 7408 14958 7460
rect 14902 7352 14958 7408
rect 14902 7300 14904 7352
rect 14904 7300 14956 7352
rect 14956 7300 14958 7352
rect 14902 7244 14958 7300
rect 14902 7192 14904 7244
rect 14904 7192 14956 7244
rect 14956 7192 14958 7244
rect 14902 7136 14958 7192
rect 14902 7084 14904 7136
rect 14904 7084 14956 7136
rect 14956 7084 14958 7136
rect 14902 7028 14958 7084
rect 14902 6976 14904 7028
rect 14904 6976 14956 7028
rect 14956 6976 14958 7028
rect 14902 6920 14958 6976
rect 14902 6868 14904 6920
rect 14904 6868 14956 6920
rect 14956 6868 14958 6920
rect 14902 6812 14958 6868
rect 14902 6760 14904 6812
rect 14904 6760 14956 6812
rect 14956 6760 14958 6812
rect 14902 6704 14958 6760
rect 14902 6652 14904 6704
rect 14904 6652 14956 6704
rect 14956 6652 14958 6704
rect 14902 6596 14958 6652
rect 14902 6544 14904 6596
rect 14904 6544 14956 6596
rect 14956 6544 14958 6596
rect 14902 6488 14958 6544
rect 14902 6436 14904 6488
rect 14904 6436 14956 6488
rect 14956 6436 14958 6488
rect 14902 6380 14958 6436
rect 14902 6328 14904 6380
rect 14904 6328 14956 6380
rect 14956 6328 14958 6380
rect 14902 6272 14958 6328
rect 14902 6220 14904 6272
rect 14904 6220 14956 6272
rect 14956 6220 14958 6272
rect 14902 6164 14958 6220
rect 14902 6112 14904 6164
rect 14904 6112 14956 6164
rect 14956 6112 14958 6164
rect 14902 6056 14958 6112
rect 14902 6004 14904 6056
rect 14904 6004 14956 6056
rect 14956 6004 14958 6056
rect 14902 5948 14958 6004
rect 14902 5896 14904 5948
rect 14904 5896 14956 5948
rect 14956 5896 14958 5948
rect 14902 5840 14958 5896
rect 14902 5788 14904 5840
rect 14904 5788 14956 5840
rect 14956 5788 14958 5840
rect 14902 5732 14958 5788
rect 14902 5680 14904 5732
rect 14904 5680 14956 5732
rect 14956 5680 14958 5732
rect 14902 5624 14958 5680
rect 14902 5572 14904 5624
rect 14904 5572 14956 5624
rect 14956 5572 14958 5624
rect 14902 5516 14958 5572
rect 14902 5464 14904 5516
rect 14904 5464 14956 5516
rect 14956 5464 14958 5516
rect 14902 5408 14958 5464
rect 14902 5356 14904 5408
rect 14904 5356 14956 5408
rect 14956 5356 14958 5408
rect 14902 5300 14958 5356
rect 14902 5248 14904 5300
rect 14904 5248 14956 5300
rect 14956 5248 14958 5300
rect 14902 5192 14958 5248
rect 14902 5140 14904 5192
rect 14904 5140 14956 5192
rect 14956 5140 14958 5192
rect 14902 5084 14958 5140
rect 14902 5032 14904 5084
rect 14904 5032 14956 5084
rect 14956 5032 14958 5084
rect 14902 4976 14958 5032
rect 14902 4924 14904 4976
rect 14904 4924 14956 4976
rect 14956 4924 14958 4976
rect 14902 4868 14958 4924
rect 14902 4816 14904 4868
rect 14904 4816 14956 4868
rect 14956 4816 14958 4868
rect 14902 4814 14958 4816
rect 20 4584 76 4586
rect 20 4532 22 4584
rect 22 4532 74 4584
rect 74 4532 76 4584
rect 20 4476 76 4532
rect 20 4424 22 4476
rect 22 4424 74 4476
rect 74 4424 76 4476
rect 20 4368 76 4424
rect 20 4316 22 4368
rect 22 4316 74 4368
rect 74 4316 76 4368
rect 20 4260 76 4316
rect 20 4208 22 4260
rect 22 4208 74 4260
rect 74 4208 76 4260
rect 20 4152 76 4208
rect 20 4100 22 4152
rect 22 4100 74 4152
rect 74 4100 76 4152
rect 20 4044 76 4100
rect 20 3992 22 4044
rect 22 3992 74 4044
rect 74 3992 76 4044
rect 20 3936 76 3992
rect 20 3884 22 3936
rect 22 3884 74 3936
rect 74 3884 76 3936
rect 20 3828 76 3884
rect 20 3776 22 3828
rect 22 3776 74 3828
rect 74 3776 76 3828
rect 20 3720 76 3776
rect 20 3668 22 3720
rect 22 3668 74 3720
rect 74 3668 76 3720
rect 20 3612 76 3668
rect 20 3560 22 3612
rect 22 3560 74 3612
rect 74 3560 76 3612
rect 20 3504 76 3560
rect 20 3452 22 3504
rect 22 3452 74 3504
rect 74 3452 76 3504
rect 20 3396 76 3452
rect 20 3344 22 3396
rect 22 3344 74 3396
rect 74 3344 76 3396
rect 20 3288 76 3344
rect 20 3236 22 3288
rect 22 3236 74 3288
rect 74 3236 76 3288
rect 20 3180 76 3236
rect 20 3128 22 3180
rect 22 3128 74 3180
rect 74 3128 76 3180
rect 20 3072 76 3128
rect 20 3020 22 3072
rect 22 3020 74 3072
rect 74 3020 76 3072
rect 20 2964 76 3020
rect 20 2912 22 2964
rect 22 2912 74 2964
rect 74 2912 76 2964
rect 20 2856 76 2912
rect 20 2804 22 2856
rect 22 2804 74 2856
rect 74 2804 76 2856
rect 20 2748 76 2804
rect 20 2696 22 2748
rect 22 2696 74 2748
rect 74 2696 76 2748
rect 20 2640 76 2696
rect 20 2588 22 2640
rect 22 2588 74 2640
rect 74 2588 76 2640
rect 20 2532 76 2588
rect 20 2480 22 2532
rect 22 2480 74 2532
rect 74 2480 76 2532
rect 20 2424 76 2480
rect 20 2372 22 2424
rect 22 2372 74 2424
rect 74 2372 76 2424
rect 20 2316 76 2372
rect 20 2264 22 2316
rect 22 2264 74 2316
rect 74 2264 76 2316
rect 20 2208 76 2264
rect 20 2156 22 2208
rect 22 2156 74 2208
rect 74 2156 76 2208
rect 20 2100 76 2156
rect 20 2048 22 2100
rect 22 2048 74 2100
rect 74 2048 76 2100
rect 20 1992 76 2048
rect 20 1940 22 1992
rect 22 1940 74 1992
rect 74 1940 76 1992
rect 20 1884 76 1940
rect 20 1832 22 1884
rect 22 1832 74 1884
rect 74 1832 76 1884
rect 20 1776 76 1832
rect 20 1724 22 1776
rect 22 1724 74 1776
rect 74 1724 76 1776
rect 20 1668 76 1724
rect 20 1616 22 1668
rect 22 1616 74 1668
rect 74 1616 76 1668
rect 20 1614 76 1616
rect 315 4498 371 4554
rect 439 4498 495 4554
rect 563 4498 619 4554
rect 687 4498 743 4554
rect 811 4498 867 4554
rect 935 4498 991 4554
rect 1059 4498 1115 4554
rect 1183 4498 1239 4554
rect 1307 4498 1363 4554
rect 1431 4498 1487 4554
rect 1555 4498 1611 4554
rect 1679 4498 1735 4554
rect 1803 4498 1859 4554
rect 1927 4498 1983 4554
rect 2051 4498 2107 4554
rect 315 4374 371 4430
rect 439 4374 495 4430
rect 563 4374 619 4430
rect 687 4374 743 4430
rect 811 4374 867 4430
rect 935 4374 991 4430
rect 1059 4374 1115 4430
rect 1183 4374 1239 4430
rect 1307 4374 1363 4430
rect 1431 4374 1487 4430
rect 1555 4374 1611 4430
rect 1679 4374 1735 4430
rect 1803 4374 1859 4430
rect 1927 4374 1983 4430
rect 2051 4374 2107 4430
rect 315 4250 371 4306
rect 439 4250 495 4306
rect 563 4250 619 4306
rect 687 4250 743 4306
rect 811 4250 867 4306
rect 935 4250 991 4306
rect 1059 4250 1115 4306
rect 1183 4250 1239 4306
rect 1307 4250 1363 4306
rect 1431 4250 1487 4306
rect 1555 4250 1611 4306
rect 1679 4250 1735 4306
rect 1803 4250 1859 4306
rect 1927 4250 1983 4306
rect 2051 4250 2107 4306
rect 315 4126 371 4182
rect 439 4126 495 4182
rect 563 4126 619 4182
rect 687 4126 743 4182
rect 811 4126 867 4182
rect 935 4126 991 4182
rect 1059 4126 1115 4182
rect 1183 4126 1239 4182
rect 1307 4126 1363 4182
rect 1431 4126 1487 4182
rect 1555 4126 1611 4182
rect 1679 4126 1735 4182
rect 1803 4126 1859 4182
rect 1927 4126 1983 4182
rect 2051 4126 2107 4182
rect 315 4002 371 4058
rect 439 4002 495 4058
rect 563 4002 619 4058
rect 687 4002 743 4058
rect 811 4002 867 4058
rect 935 4002 991 4058
rect 1059 4002 1115 4058
rect 1183 4002 1239 4058
rect 1307 4002 1363 4058
rect 1431 4002 1487 4058
rect 1555 4002 1611 4058
rect 1679 4002 1735 4058
rect 1803 4002 1859 4058
rect 1927 4002 1983 4058
rect 2051 4002 2107 4058
rect 315 3878 371 3934
rect 439 3878 495 3934
rect 563 3878 619 3934
rect 687 3878 743 3934
rect 811 3878 867 3934
rect 935 3878 991 3934
rect 1059 3878 1115 3934
rect 1183 3878 1239 3934
rect 1307 3878 1363 3934
rect 1431 3878 1487 3934
rect 1555 3878 1611 3934
rect 1679 3878 1735 3934
rect 1803 3878 1859 3934
rect 1927 3878 1983 3934
rect 2051 3878 2107 3934
rect 315 3754 371 3810
rect 439 3754 495 3810
rect 563 3754 619 3810
rect 687 3754 743 3810
rect 811 3754 867 3810
rect 935 3754 991 3810
rect 1059 3754 1115 3810
rect 1183 3754 1239 3810
rect 1307 3754 1363 3810
rect 1431 3754 1487 3810
rect 1555 3754 1611 3810
rect 1679 3754 1735 3810
rect 1803 3754 1859 3810
rect 1927 3754 1983 3810
rect 2051 3754 2107 3810
rect 315 3630 371 3686
rect 439 3630 495 3686
rect 563 3630 619 3686
rect 687 3630 743 3686
rect 811 3630 867 3686
rect 935 3630 991 3686
rect 1059 3630 1115 3686
rect 1183 3630 1239 3686
rect 1307 3630 1363 3686
rect 1431 3630 1487 3686
rect 1555 3630 1611 3686
rect 1679 3630 1735 3686
rect 1803 3630 1859 3686
rect 1927 3630 1983 3686
rect 2051 3630 2107 3686
rect 315 3506 371 3562
rect 439 3506 495 3562
rect 563 3506 619 3562
rect 687 3506 743 3562
rect 811 3506 867 3562
rect 935 3506 991 3562
rect 1059 3506 1115 3562
rect 1183 3506 1239 3562
rect 1307 3506 1363 3562
rect 1431 3506 1487 3562
rect 1555 3506 1611 3562
rect 1679 3506 1735 3562
rect 1803 3506 1859 3562
rect 1927 3506 1983 3562
rect 2051 3506 2107 3562
rect 315 3382 371 3438
rect 439 3382 495 3438
rect 563 3382 619 3438
rect 687 3382 743 3438
rect 811 3382 867 3438
rect 935 3382 991 3438
rect 1059 3382 1115 3438
rect 1183 3382 1239 3438
rect 1307 3382 1363 3438
rect 1431 3382 1487 3438
rect 1555 3382 1611 3438
rect 1679 3382 1735 3438
rect 1803 3382 1859 3438
rect 1927 3382 1983 3438
rect 2051 3382 2107 3438
rect 315 3258 371 3314
rect 439 3258 495 3314
rect 563 3258 619 3314
rect 687 3258 743 3314
rect 811 3258 867 3314
rect 935 3258 991 3314
rect 1059 3258 1115 3314
rect 1183 3258 1239 3314
rect 1307 3258 1363 3314
rect 1431 3258 1487 3314
rect 1555 3258 1611 3314
rect 1679 3258 1735 3314
rect 1803 3258 1859 3314
rect 1927 3258 1983 3314
rect 2051 3258 2107 3314
rect 315 3134 371 3190
rect 439 3134 495 3190
rect 563 3134 619 3190
rect 687 3134 743 3190
rect 811 3134 867 3190
rect 935 3134 991 3190
rect 1059 3134 1115 3190
rect 1183 3134 1239 3190
rect 1307 3134 1363 3190
rect 1431 3134 1487 3190
rect 1555 3134 1611 3190
rect 1679 3134 1735 3190
rect 1803 3134 1859 3190
rect 1927 3134 1983 3190
rect 2051 3134 2107 3190
rect 315 3010 371 3066
rect 439 3010 495 3066
rect 563 3010 619 3066
rect 687 3010 743 3066
rect 811 3010 867 3066
rect 935 3010 991 3066
rect 1059 3010 1115 3066
rect 1183 3010 1239 3066
rect 1307 3010 1363 3066
rect 1431 3010 1487 3066
rect 1555 3010 1611 3066
rect 1679 3010 1735 3066
rect 1803 3010 1859 3066
rect 1927 3010 1983 3066
rect 2051 3010 2107 3066
rect 315 2886 371 2942
rect 439 2886 495 2942
rect 563 2886 619 2942
rect 687 2886 743 2942
rect 811 2886 867 2942
rect 935 2886 991 2942
rect 1059 2886 1115 2942
rect 1183 2886 1239 2942
rect 1307 2886 1363 2942
rect 1431 2886 1487 2942
rect 1555 2886 1611 2942
rect 1679 2886 1735 2942
rect 1803 2886 1859 2942
rect 1927 2886 1983 2942
rect 2051 2886 2107 2942
rect 315 2762 371 2818
rect 439 2762 495 2818
rect 563 2762 619 2818
rect 687 2762 743 2818
rect 811 2762 867 2818
rect 935 2762 991 2818
rect 1059 2762 1115 2818
rect 1183 2762 1239 2818
rect 1307 2762 1363 2818
rect 1431 2762 1487 2818
rect 1555 2762 1611 2818
rect 1679 2762 1735 2818
rect 1803 2762 1859 2818
rect 1927 2762 1983 2818
rect 2051 2762 2107 2818
rect 315 2638 371 2694
rect 439 2638 495 2694
rect 563 2638 619 2694
rect 687 2638 743 2694
rect 811 2638 867 2694
rect 935 2638 991 2694
rect 1059 2638 1115 2694
rect 1183 2638 1239 2694
rect 1307 2638 1363 2694
rect 1431 2638 1487 2694
rect 1555 2638 1611 2694
rect 1679 2638 1735 2694
rect 1803 2638 1859 2694
rect 1927 2638 1983 2694
rect 2051 2638 2107 2694
rect 315 2514 371 2570
rect 439 2514 495 2570
rect 563 2514 619 2570
rect 687 2514 743 2570
rect 811 2514 867 2570
rect 935 2514 991 2570
rect 1059 2514 1115 2570
rect 1183 2514 1239 2570
rect 1307 2514 1363 2570
rect 1431 2514 1487 2570
rect 1555 2514 1611 2570
rect 1679 2514 1735 2570
rect 1803 2514 1859 2570
rect 1927 2514 1983 2570
rect 2051 2514 2107 2570
rect 315 2390 371 2446
rect 439 2390 495 2446
rect 563 2390 619 2446
rect 687 2390 743 2446
rect 811 2390 867 2446
rect 935 2390 991 2446
rect 1059 2390 1115 2446
rect 1183 2390 1239 2446
rect 1307 2390 1363 2446
rect 1431 2390 1487 2446
rect 1555 2390 1611 2446
rect 1679 2390 1735 2446
rect 1803 2390 1859 2446
rect 1927 2390 1983 2446
rect 2051 2390 2107 2446
rect 315 2266 371 2322
rect 439 2266 495 2322
rect 563 2266 619 2322
rect 687 2266 743 2322
rect 811 2266 867 2322
rect 935 2266 991 2322
rect 1059 2266 1115 2322
rect 1183 2266 1239 2322
rect 1307 2266 1363 2322
rect 1431 2266 1487 2322
rect 1555 2266 1611 2322
rect 1679 2266 1735 2322
rect 1803 2266 1859 2322
rect 1927 2266 1983 2322
rect 2051 2266 2107 2322
rect 315 2142 371 2198
rect 439 2142 495 2198
rect 563 2142 619 2198
rect 687 2142 743 2198
rect 811 2142 867 2198
rect 935 2142 991 2198
rect 1059 2142 1115 2198
rect 1183 2142 1239 2198
rect 1307 2142 1363 2198
rect 1431 2142 1487 2198
rect 1555 2142 1611 2198
rect 1679 2142 1735 2198
rect 1803 2142 1859 2198
rect 1927 2142 1983 2198
rect 2051 2142 2107 2198
rect 315 2018 371 2074
rect 439 2018 495 2074
rect 563 2018 619 2074
rect 687 2018 743 2074
rect 811 2018 867 2074
rect 935 2018 991 2074
rect 1059 2018 1115 2074
rect 1183 2018 1239 2074
rect 1307 2018 1363 2074
rect 1431 2018 1487 2074
rect 1555 2018 1611 2074
rect 1679 2018 1735 2074
rect 1803 2018 1859 2074
rect 1927 2018 1983 2074
rect 2051 2018 2107 2074
rect 315 1894 371 1950
rect 439 1894 495 1950
rect 563 1894 619 1950
rect 687 1894 743 1950
rect 811 1894 867 1950
rect 935 1894 991 1950
rect 1059 1894 1115 1950
rect 1183 1894 1239 1950
rect 1307 1894 1363 1950
rect 1431 1894 1487 1950
rect 1555 1894 1611 1950
rect 1679 1894 1735 1950
rect 1803 1894 1859 1950
rect 1927 1894 1983 1950
rect 2051 1894 2107 1950
rect 315 1770 371 1826
rect 439 1770 495 1826
rect 563 1770 619 1826
rect 687 1770 743 1826
rect 811 1770 867 1826
rect 935 1770 991 1826
rect 1059 1770 1115 1826
rect 1183 1770 1239 1826
rect 1307 1770 1363 1826
rect 1431 1770 1487 1826
rect 1555 1770 1611 1826
rect 1679 1770 1735 1826
rect 1803 1770 1859 1826
rect 1927 1770 1983 1826
rect 2051 1770 2107 1826
rect 315 1646 371 1702
rect 439 1646 495 1702
rect 563 1646 619 1702
rect 687 1646 743 1702
rect 811 1646 867 1702
rect 935 1646 991 1702
rect 1059 1646 1115 1702
rect 1183 1646 1239 1702
rect 1307 1646 1363 1702
rect 1431 1646 1487 1702
rect 1555 1646 1611 1702
rect 1679 1646 1735 1702
rect 1803 1646 1859 1702
rect 1927 1646 1983 1702
rect 2051 1646 2107 1702
rect 2808 4498 2864 4554
rect 2932 4498 2988 4554
rect 3056 4498 3112 4554
rect 3180 4498 3236 4554
rect 3304 4498 3360 4554
rect 3428 4498 3484 4554
rect 3552 4498 3608 4554
rect 3676 4498 3732 4554
rect 3800 4498 3856 4554
rect 3924 4498 3980 4554
rect 4048 4498 4104 4554
rect 4172 4498 4228 4554
rect 4296 4498 4352 4554
rect 4420 4498 4476 4554
rect 4544 4498 4600 4554
rect 4668 4498 4724 4554
rect 2808 4374 2864 4430
rect 2932 4374 2988 4430
rect 3056 4374 3112 4430
rect 3180 4374 3236 4430
rect 3304 4374 3360 4430
rect 3428 4374 3484 4430
rect 3552 4374 3608 4430
rect 3676 4374 3732 4430
rect 3800 4374 3856 4430
rect 3924 4374 3980 4430
rect 4048 4374 4104 4430
rect 4172 4374 4228 4430
rect 4296 4374 4352 4430
rect 4420 4374 4476 4430
rect 4544 4374 4600 4430
rect 4668 4374 4724 4430
rect 2808 4250 2864 4306
rect 2932 4250 2988 4306
rect 3056 4250 3112 4306
rect 3180 4250 3236 4306
rect 3304 4250 3360 4306
rect 3428 4250 3484 4306
rect 3552 4250 3608 4306
rect 3676 4250 3732 4306
rect 3800 4250 3856 4306
rect 3924 4250 3980 4306
rect 4048 4250 4104 4306
rect 4172 4250 4228 4306
rect 4296 4250 4352 4306
rect 4420 4250 4476 4306
rect 4544 4250 4600 4306
rect 4668 4250 4724 4306
rect 2808 4126 2864 4182
rect 2932 4126 2988 4182
rect 3056 4126 3112 4182
rect 3180 4126 3236 4182
rect 3304 4126 3360 4182
rect 3428 4126 3484 4182
rect 3552 4126 3608 4182
rect 3676 4126 3732 4182
rect 3800 4126 3856 4182
rect 3924 4126 3980 4182
rect 4048 4126 4104 4182
rect 4172 4126 4228 4182
rect 4296 4126 4352 4182
rect 4420 4126 4476 4182
rect 4544 4126 4600 4182
rect 4668 4126 4724 4182
rect 2808 4002 2864 4058
rect 2932 4002 2988 4058
rect 3056 4002 3112 4058
rect 3180 4002 3236 4058
rect 3304 4002 3360 4058
rect 3428 4002 3484 4058
rect 3552 4002 3608 4058
rect 3676 4002 3732 4058
rect 3800 4002 3856 4058
rect 3924 4002 3980 4058
rect 4048 4002 4104 4058
rect 4172 4002 4228 4058
rect 4296 4002 4352 4058
rect 4420 4002 4476 4058
rect 4544 4002 4600 4058
rect 4668 4002 4724 4058
rect 2808 3878 2864 3934
rect 2932 3878 2988 3934
rect 3056 3878 3112 3934
rect 3180 3878 3236 3934
rect 3304 3878 3360 3934
rect 3428 3878 3484 3934
rect 3552 3878 3608 3934
rect 3676 3878 3732 3934
rect 3800 3878 3856 3934
rect 3924 3878 3980 3934
rect 4048 3878 4104 3934
rect 4172 3878 4228 3934
rect 4296 3878 4352 3934
rect 4420 3878 4476 3934
rect 4544 3878 4600 3934
rect 4668 3878 4724 3934
rect 2808 3754 2864 3810
rect 2932 3754 2988 3810
rect 3056 3754 3112 3810
rect 3180 3754 3236 3810
rect 3304 3754 3360 3810
rect 3428 3754 3484 3810
rect 3552 3754 3608 3810
rect 3676 3754 3732 3810
rect 3800 3754 3856 3810
rect 3924 3754 3980 3810
rect 4048 3754 4104 3810
rect 4172 3754 4228 3810
rect 4296 3754 4352 3810
rect 4420 3754 4476 3810
rect 4544 3754 4600 3810
rect 4668 3754 4724 3810
rect 2808 3630 2864 3686
rect 2932 3630 2988 3686
rect 3056 3630 3112 3686
rect 3180 3630 3236 3686
rect 3304 3630 3360 3686
rect 3428 3630 3484 3686
rect 3552 3630 3608 3686
rect 3676 3630 3732 3686
rect 3800 3630 3856 3686
rect 3924 3630 3980 3686
rect 4048 3630 4104 3686
rect 4172 3630 4228 3686
rect 4296 3630 4352 3686
rect 4420 3630 4476 3686
rect 4544 3630 4600 3686
rect 4668 3630 4724 3686
rect 2808 3506 2864 3562
rect 2932 3506 2988 3562
rect 3056 3506 3112 3562
rect 3180 3506 3236 3562
rect 3304 3506 3360 3562
rect 3428 3506 3484 3562
rect 3552 3506 3608 3562
rect 3676 3506 3732 3562
rect 3800 3506 3856 3562
rect 3924 3506 3980 3562
rect 4048 3506 4104 3562
rect 4172 3506 4228 3562
rect 4296 3506 4352 3562
rect 4420 3506 4476 3562
rect 4544 3506 4600 3562
rect 4668 3506 4724 3562
rect 2808 3382 2864 3438
rect 2932 3382 2988 3438
rect 3056 3382 3112 3438
rect 3180 3382 3236 3438
rect 3304 3382 3360 3438
rect 3428 3382 3484 3438
rect 3552 3382 3608 3438
rect 3676 3382 3732 3438
rect 3800 3382 3856 3438
rect 3924 3382 3980 3438
rect 4048 3382 4104 3438
rect 4172 3382 4228 3438
rect 4296 3382 4352 3438
rect 4420 3382 4476 3438
rect 4544 3382 4600 3438
rect 4668 3382 4724 3438
rect 2808 3258 2864 3314
rect 2932 3258 2988 3314
rect 3056 3258 3112 3314
rect 3180 3258 3236 3314
rect 3304 3258 3360 3314
rect 3428 3258 3484 3314
rect 3552 3258 3608 3314
rect 3676 3258 3732 3314
rect 3800 3258 3856 3314
rect 3924 3258 3980 3314
rect 4048 3258 4104 3314
rect 4172 3258 4228 3314
rect 4296 3258 4352 3314
rect 4420 3258 4476 3314
rect 4544 3258 4600 3314
rect 4668 3258 4724 3314
rect 2808 3134 2864 3190
rect 2932 3134 2988 3190
rect 3056 3134 3112 3190
rect 3180 3134 3236 3190
rect 3304 3134 3360 3190
rect 3428 3134 3484 3190
rect 3552 3134 3608 3190
rect 3676 3134 3732 3190
rect 3800 3134 3856 3190
rect 3924 3134 3980 3190
rect 4048 3134 4104 3190
rect 4172 3134 4228 3190
rect 4296 3134 4352 3190
rect 4420 3134 4476 3190
rect 4544 3134 4600 3190
rect 4668 3134 4724 3190
rect 2808 3010 2864 3066
rect 2932 3010 2988 3066
rect 3056 3010 3112 3066
rect 3180 3010 3236 3066
rect 3304 3010 3360 3066
rect 3428 3010 3484 3066
rect 3552 3010 3608 3066
rect 3676 3010 3732 3066
rect 3800 3010 3856 3066
rect 3924 3010 3980 3066
rect 4048 3010 4104 3066
rect 4172 3010 4228 3066
rect 4296 3010 4352 3066
rect 4420 3010 4476 3066
rect 4544 3010 4600 3066
rect 4668 3010 4724 3066
rect 2808 2886 2864 2942
rect 2932 2886 2988 2942
rect 3056 2886 3112 2942
rect 3180 2886 3236 2942
rect 3304 2886 3360 2942
rect 3428 2886 3484 2942
rect 3552 2886 3608 2942
rect 3676 2886 3732 2942
rect 3800 2886 3856 2942
rect 3924 2886 3980 2942
rect 4048 2886 4104 2942
rect 4172 2886 4228 2942
rect 4296 2886 4352 2942
rect 4420 2886 4476 2942
rect 4544 2886 4600 2942
rect 4668 2886 4724 2942
rect 2808 2762 2864 2818
rect 2932 2762 2988 2818
rect 3056 2762 3112 2818
rect 3180 2762 3236 2818
rect 3304 2762 3360 2818
rect 3428 2762 3484 2818
rect 3552 2762 3608 2818
rect 3676 2762 3732 2818
rect 3800 2762 3856 2818
rect 3924 2762 3980 2818
rect 4048 2762 4104 2818
rect 4172 2762 4228 2818
rect 4296 2762 4352 2818
rect 4420 2762 4476 2818
rect 4544 2762 4600 2818
rect 4668 2762 4724 2818
rect 2808 2638 2864 2694
rect 2932 2638 2988 2694
rect 3056 2638 3112 2694
rect 3180 2638 3236 2694
rect 3304 2638 3360 2694
rect 3428 2638 3484 2694
rect 3552 2638 3608 2694
rect 3676 2638 3732 2694
rect 3800 2638 3856 2694
rect 3924 2638 3980 2694
rect 4048 2638 4104 2694
rect 4172 2638 4228 2694
rect 4296 2638 4352 2694
rect 4420 2638 4476 2694
rect 4544 2638 4600 2694
rect 4668 2638 4724 2694
rect 2808 2514 2864 2570
rect 2932 2514 2988 2570
rect 3056 2514 3112 2570
rect 3180 2514 3236 2570
rect 3304 2514 3360 2570
rect 3428 2514 3484 2570
rect 3552 2514 3608 2570
rect 3676 2514 3732 2570
rect 3800 2514 3856 2570
rect 3924 2514 3980 2570
rect 4048 2514 4104 2570
rect 4172 2514 4228 2570
rect 4296 2514 4352 2570
rect 4420 2514 4476 2570
rect 4544 2514 4600 2570
rect 4668 2514 4724 2570
rect 2808 2390 2864 2446
rect 2932 2390 2988 2446
rect 3056 2390 3112 2446
rect 3180 2390 3236 2446
rect 3304 2390 3360 2446
rect 3428 2390 3484 2446
rect 3552 2390 3608 2446
rect 3676 2390 3732 2446
rect 3800 2390 3856 2446
rect 3924 2390 3980 2446
rect 4048 2390 4104 2446
rect 4172 2390 4228 2446
rect 4296 2390 4352 2446
rect 4420 2390 4476 2446
rect 4544 2390 4600 2446
rect 4668 2390 4724 2446
rect 2808 2266 2864 2322
rect 2932 2266 2988 2322
rect 3056 2266 3112 2322
rect 3180 2266 3236 2322
rect 3304 2266 3360 2322
rect 3428 2266 3484 2322
rect 3552 2266 3608 2322
rect 3676 2266 3732 2322
rect 3800 2266 3856 2322
rect 3924 2266 3980 2322
rect 4048 2266 4104 2322
rect 4172 2266 4228 2322
rect 4296 2266 4352 2322
rect 4420 2266 4476 2322
rect 4544 2266 4600 2322
rect 4668 2266 4724 2322
rect 2808 2142 2864 2198
rect 2932 2142 2988 2198
rect 3056 2142 3112 2198
rect 3180 2142 3236 2198
rect 3304 2142 3360 2198
rect 3428 2142 3484 2198
rect 3552 2142 3608 2198
rect 3676 2142 3732 2198
rect 3800 2142 3856 2198
rect 3924 2142 3980 2198
rect 4048 2142 4104 2198
rect 4172 2142 4228 2198
rect 4296 2142 4352 2198
rect 4420 2142 4476 2198
rect 4544 2142 4600 2198
rect 4668 2142 4724 2198
rect 2808 2018 2864 2074
rect 2932 2018 2988 2074
rect 3056 2018 3112 2074
rect 3180 2018 3236 2074
rect 3304 2018 3360 2074
rect 3428 2018 3484 2074
rect 3552 2018 3608 2074
rect 3676 2018 3732 2074
rect 3800 2018 3856 2074
rect 3924 2018 3980 2074
rect 4048 2018 4104 2074
rect 4172 2018 4228 2074
rect 4296 2018 4352 2074
rect 4420 2018 4476 2074
rect 4544 2018 4600 2074
rect 4668 2018 4724 2074
rect 2808 1894 2864 1950
rect 2932 1894 2988 1950
rect 3056 1894 3112 1950
rect 3180 1894 3236 1950
rect 3304 1894 3360 1950
rect 3428 1894 3484 1950
rect 3552 1894 3608 1950
rect 3676 1894 3732 1950
rect 3800 1894 3856 1950
rect 3924 1894 3980 1950
rect 4048 1894 4104 1950
rect 4172 1894 4228 1950
rect 4296 1894 4352 1950
rect 4420 1894 4476 1950
rect 4544 1894 4600 1950
rect 4668 1894 4724 1950
rect 2808 1770 2864 1826
rect 2932 1770 2988 1826
rect 3056 1770 3112 1826
rect 3180 1770 3236 1826
rect 3304 1770 3360 1826
rect 3428 1770 3484 1826
rect 3552 1770 3608 1826
rect 3676 1770 3732 1826
rect 3800 1770 3856 1826
rect 3924 1770 3980 1826
rect 4048 1770 4104 1826
rect 4172 1770 4228 1826
rect 4296 1770 4352 1826
rect 4420 1770 4476 1826
rect 4544 1770 4600 1826
rect 4668 1770 4724 1826
rect 2808 1646 2864 1702
rect 2932 1646 2988 1702
rect 3056 1646 3112 1702
rect 3180 1646 3236 1702
rect 3304 1646 3360 1702
rect 3428 1646 3484 1702
rect 3552 1646 3608 1702
rect 3676 1646 3732 1702
rect 3800 1646 3856 1702
rect 3924 1646 3980 1702
rect 4048 1646 4104 1702
rect 4172 1646 4228 1702
rect 4296 1646 4352 1702
rect 4420 1646 4476 1702
rect 4544 1646 4600 1702
rect 4668 1646 4724 1702
rect 5178 4498 5234 4554
rect 5302 4498 5358 4554
rect 5426 4498 5482 4554
rect 5550 4498 5606 4554
rect 5674 4498 5730 4554
rect 5798 4498 5854 4554
rect 5922 4498 5978 4554
rect 6046 4498 6102 4554
rect 6170 4498 6226 4554
rect 6294 4498 6350 4554
rect 6418 4498 6474 4554
rect 6542 4498 6598 4554
rect 6666 4498 6722 4554
rect 6790 4498 6846 4554
rect 6914 4498 6970 4554
rect 7038 4498 7094 4554
rect 5178 4374 5234 4430
rect 5302 4374 5358 4430
rect 5426 4374 5482 4430
rect 5550 4374 5606 4430
rect 5674 4374 5730 4430
rect 5798 4374 5854 4430
rect 5922 4374 5978 4430
rect 6046 4374 6102 4430
rect 6170 4374 6226 4430
rect 6294 4374 6350 4430
rect 6418 4374 6474 4430
rect 6542 4374 6598 4430
rect 6666 4374 6722 4430
rect 6790 4374 6846 4430
rect 6914 4374 6970 4430
rect 7038 4374 7094 4430
rect 5178 4250 5234 4306
rect 5302 4250 5358 4306
rect 5426 4250 5482 4306
rect 5550 4250 5606 4306
rect 5674 4250 5730 4306
rect 5798 4250 5854 4306
rect 5922 4250 5978 4306
rect 6046 4250 6102 4306
rect 6170 4250 6226 4306
rect 6294 4250 6350 4306
rect 6418 4250 6474 4306
rect 6542 4250 6598 4306
rect 6666 4250 6722 4306
rect 6790 4250 6846 4306
rect 6914 4250 6970 4306
rect 7038 4250 7094 4306
rect 5178 4126 5234 4182
rect 5302 4126 5358 4182
rect 5426 4126 5482 4182
rect 5550 4126 5606 4182
rect 5674 4126 5730 4182
rect 5798 4126 5854 4182
rect 5922 4126 5978 4182
rect 6046 4126 6102 4182
rect 6170 4126 6226 4182
rect 6294 4126 6350 4182
rect 6418 4126 6474 4182
rect 6542 4126 6598 4182
rect 6666 4126 6722 4182
rect 6790 4126 6846 4182
rect 6914 4126 6970 4182
rect 7038 4126 7094 4182
rect 5178 4002 5234 4058
rect 5302 4002 5358 4058
rect 5426 4002 5482 4058
rect 5550 4002 5606 4058
rect 5674 4002 5730 4058
rect 5798 4002 5854 4058
rect 5922 4002 5978 4058
rect 6046 4002 6102 4058
rect 6170 4002 6226 4058
rect 6294 4002 6350 4058
rect 6418 4002 6474 4058
rect 6542 4002 6598 4058
rect 6666 4002 6722 4058
rect 6790 4002 6846 4058
rect 6914 4002 6970 4058
rect 7038 4002 7094 4058
rect 5178 3878 5234 3934
rect 5302 3878 5358 3934
rect 5426 3878 5482 3934
rect 5550 3878 5606 3934
rect 5674 3878 5730 3934
rect 5798 3878 5854 3934
rect 5922 3878 5978 3934
rect 6046 3878 6102 3934
rect 6170 3878 6226 3934
rect 6294 3878 6350 3934
rect 6418 3878 6474 3934
rect 6542 3878 6598 3934
rect 6666 3878 6722 3934
rect 6790 3878 6846 3934
rect 6914 3878 6970 3934
rect 7038 3878 7094 3934
rect 5178 3754 5234 3810
rect 5302 3754 5358 3810
rect 5426 3754 5482 3810
rect 5550 3754 5606 3810
rect 5674 3754 5730 3810
rect 5798 3754 5854 3810
rect 5922 3754 5978 3810
rect 6046 3754 6102 3810
rect 6170 3754 6226 3810
rect 6294 3754 6350 3810
rect 6418 3754 6474 3810
rect 6542 3754 6598 3810
rect 6666 3754 6722 3810
rect 6790 3754 6846 3810
rect 6914 3754 6970 3810
rect 7038 3754 7094 3810
rect 5178 3630 5234 3686
rect 5302 3630 5358 3686
rect 5426 3630 5482 3686
rect 5550 3630 5606 3686
rect 5674 3630 5730 3686
rect 5798 3630 5854 3686
rect 5922 3630 5978 3686
rect 6046 3630 6102 3686
rect 6170 3630 6226 3686
rect 6294 3630 6350 3686
rect 6418 3630 6474 3686
rect 6542 3630 6598 3686
rect 6666 3630 6722 3686
rect 6790 3630 6846 3686
rect 6914 3630 6970 3686
rect 7038 3630 7094 3686
rect 5178 3506 5234 3562
rect 5302 3506 5358 3562
rect 5426 3506 5482 3562
rect 5550 3506 5606 3562
rect 5674 3506 5730 3562
rect 5798 3506 5854 3562
rect 5922 3506 5978 3562
rect 6046 3506 6102 3562
rect 6170 3506 6226 3562
rect 6294 3506 6350 3562
rect 6418 3506 6474 3562
rect 6542 3506 6598 3562
rect 6666 3506 6722 3562
rect 6790 3506 6846 3562
rect 6914 3506 6970 3562
rect 7038 3506 7094 3562
rect 5178 3382 5234 3438
rect 5302 3382 5358 3438
rect 5426 3382 5482 3438
rect 5550 3382 5606 3438
rect 5674 3382 5730 3438
rect 5798 3382 5854 3438
rect 5922 3382 5978 3438
rect 6046 3382 6102 3438
rect 6170 3382 6226 3438
rect 6294 3382 6350 3438
rect 6418 3382 6474 3438
rect 6542 3382 6598 3438
rect 6666 3382 6722 3438
rect 6790 3382 6846 3438
rect 6914 3382 6970 3438
rect 7038 3382 7094 3438
rect 5178 3258 5234 3314
rect 5302 3258 5358 3314
rect 5426 3258 5482 3314
rect 5550 3258 5606 3314
rect 5674 3258 5730 3314
rect 5798 3258 5854 3314
rect 5922 3258 5978 3314
rect 6046 3258 6102 3314
rect 6170 3258 6226 3314
rect 6294 3258 6350 3314
rect 6418 3258 6474 3314
rect 6542 3258 6598 3314
rect 6666 3258 6722 3314
rect 6790 3258 6846 3314
rect 6914 3258 6970 3314
rect 7038 3258 7094 3314
rect 5178 3134 5234 3190
rect 5302 3134 5358 3190
rect 5426 3134 5482 3190
rect 5550 3134 5606 3190
rect 5674 3134 5730 3190
rect 5798 3134 5854 3190
rect 5922 3134 5978 3190
rect 6046 3134 6102 3190
rect 6170 3134 6226 3190
rect 6294 3134 6350 3190
rect 6418 3134 6474 3190
rect 6542 3134 6598 3190
rect 6666 3134 6722 3190
rect 6790 3134 6846 3190
rect 6914 3134 6970 3190
rect 7038 3134 7094 3190
rect 5178 3010 5234 3066
rect 5302 3010 5358 3066
rect 5426 3010 5482 3066
rect 5550 3010 5606 3066
rect 5674 3010 5730 3066
rect 5798 3010 5854 3066
rect 5922 3010 5978 3066
rect 6046 3010 6102 3066
rect 6170 3010 6226 3066
rect 6294 3010 6350 3066
rect 6418 3010 6474 3066
rect 6542 3010 6598 3066
rect 6666 3010 6722 3066
rect 6790 3010 6846 3066
rect 6914 3010 6970 3066
rect 7038 3010 7094 3066
rect 5178 2886 5234 2942
rect 5302 2886 5358 2942
rect 5426 2886 5482 2942
rect 5550 2886 5606 2942
rect 5674 2886 5730 2942
rect 5798 2886 5854 2942
rect 5922 2886 5978 2942
rect 6046 2886 6102 2942
rect 6170 2886 6226 2942
rect 6294 2886 6350 2942
rect 6418 2886 6474 2942
rect 6542 2886 6598 2942
rect 6666 2886 6722 2942
rect 6790 2886 6846 2942
rect 6914 2886 6970 2942
rect 7038 2886 7094 2942
rect 5178 2762 5234 2818
rect 5302 2762 5358 2818
rect 5426 2762 5482 2818
rect 5550 2762 5606 2818
rect 5674 2762 5730 2818
rect 5798 2762 5854 2818
rect 5922 2762 5978 2818
rect 6046 2762 6102 2818
rect 6170 2762 6226 2818
rect 6294 2762 6350 2818
rect 6418 2762 6474 2818
rect 6542 2762 6598 2818
rect 6666 2762 6722 2818
rect 6790 2762 6846 2818
rect 6914 2762 6970 2818
rect 7038 2762 7094 2818
rect 5178 2638 5234 2694
rect 5302 2638 5358 2694
rect 5426 2638 5482 2694
rect 5550 2638 5606 2694
rect 5674 2638 5730 2694
rect 5798 2638 5854 2694
rect 5922 2638 5978 2694
rect 6046 2638 6102 2694
rect 6170 2638 6226 2694
rect 6294 2638 6350 2694
rect 6418 2638 6474 2694
rect 6542 2638 6598 2694
rect 6666 2638 6722 2694
rect 6790 2638 6846 2694
rect 6914 2638 6970 2694
rect 7038 2638 7094 2694
rect 5178 2514 5234 2570
rect 5302 2514 5358 2570
rect 5426 2514 5482 2570
rect 5550 2514 5606 2570
rect 5674 2514 5730 2570
rect 5798 2514 5854 2570
rect 5922 2514 5978 2570
rect 6046 2514 6102 2570
rect 6170 2514 6226 2570
rect 6294 2514 6350 2570
rect 6418 2514 6474 2570
rect 6542 2514 6598 2570
rect 6666 2514 6722 2570
rect 6790 2514 6846 2570
rect 6914 2514 6970 2570
rect 7038 2514 7094 2570
rect 5178 2390 5234 2446
rect 5302 2390 5358 2446
rect 5426 2390 5482 2446
rect 5550 2390 5606 2446
rect 5674 2390 5730 2446
rect 5798 2390 5854 2446
rect 5922 2390 5978 2446
rect 6046 2390 6102 2446
rect 6170 2390 6226 2446
rect 6294 2390 6350 2446
rect 6418 2390 6474 2446
rect 6542 2390 6598 2446
rect 6666 2390 6722 2446
rect 6790 2390 6846 2446
rect 6914 2390 6970 2446
rect 7038 2390 7094 2446
rect 5178 2266 5234 2322
rect 5302 2266 5358 2322
rect 5426 2266 5482 2322
rect 5550 2266 5606 2322
rect 5674 2266 5730 2322
rect 5798 2266 5854 2322
rect 5922 2266 5978 2322
rect 6046 2266 6102 2322
rect 6170 2266 6226 2322
rect 6294 2266 6350 2322
rect 6418 2266 6474 2322
rect 6542 2266 6598 2322
rect 6666 2266 6722 2322
rect 6790 2266 6846 2322
rect 6914 2266 6970 2322
rect 7038 2266 7094 2322
rect 5178 2142 5234 2198
rect 5302 2142 5358 2198
rect 5426 2142 5482 2198
rect 5550 2142 5606 2198
rect 5674 2142 5730 2198
rect 5798 2142 5854 2198
rect 5922 2142 5978 2198
rect 6046 2142 6102 2198
rect 6170 2142 6226 2198
rect 6294 2142 6350 2198
rect 6418 2142 6474 2198
rect 6542 2142 6598 2198
rect 6666 2142 6722 2198
rect 6790 2142 6846 2198
rect 6914 2142 6970 2198
rect 7038 2142 7094 2198
rect 5178 2018 5234 2074
rect 5302 2018 5358 2074
rect 5426 2018 5482 2074
rect 5550 2018 5606 2074
rect 5674 2018 5730 2074
rect 5798 2018 5854 2074
rect 5922 2018 5978 2074
rect 6046 2018 6102 2074
rect 6170 2018 6226 2074
rect 6294 2018 6350 2074
rect 6418 2018 6474 2074
rect 6542 2018 6598 2074
rect 6666 2018 6722 2074
rect 6790 2018 6846 2074
rect 6914 2018 6970 2074
rect 7038 2018 7094 2074
rect 5178 1894 5234 1950
rect 5302 1894 5358 1950
rect 5426 1894 5482 1950
rect 5550 1894 5606 1950
rect 5674 1894 5730 1950
rect 5798 1894 5854 1950
rect 5922 1894 5978 1950
rect 6046 1894 6102 1950
rect 6170 1894 6226 1950
rect 6294 1894 6350 1950
rect 6418 1894 6474 1950
rect 6542 1894 6598 1950
rect 6666 1894 6722 1950
rect 6790 1894 6846 1950
rect 6914 1894 6970 1950
rect 7038 1894 7094 1950
rect 5178 1770 5234 1826
rect 5302 1770 5358 1826
rect 5426 1770 5482 1826
rect 5550 1770 5606 1826
rect 5674 1770 5730 1826
rect 5798 1770 5854 1826
rect 5922 1770 5978 1826
rect 6046 1770 6102 1826
rect 6170 1770 6226 1826
rect 6294 1770 6350 1826
rect 6418 1770 6474 1826
rect 6542 1770 6598 1826
rect 6666 1770 6722 1826
rect 6790 1770 6846 1826
rect 6914 1770 6970 1826
rect 7038 1770 7094 1826
rect 5178 1646 5234 1702
rect 5302 1646 5358 1702
rect 5426 1646 5482 1702
rect 5550 1646 5606 1702
rect 5674 1646 5730 1702
rect 5798 1646 5854 1702
rect 5922 1646 5978 1702
rect 6046 1646 6102 1702
rect 6170 1646 6226 1702
rect 6294 1646 6350 1702
rect 6418 1646 6474 1702
rect 6542 1646 6598 1702
rect 6666 1646 6722 1702
rect 6790 1646 6846 1702
rect 6914 1646 6970 1702
rect 7038 1646 7094 1702
rect 7884 4498 7940 4554
rect 8008 4498 8064 4554
rect 8132 4498 8188 4554
rect 8256 4498 8312 4554
rect 8380 4498 8436 4554
rect 8504 4498 8560 4554
rect 8628 4498 8684 4554
rect 8752 4498 8808 4554
rect 8876 4498 8932 4554
rect 9000 4498 9056 4554
rect 9124 4498 9180 4554
rect 9248 4498 9304 4554
rect 9372 4498 9428 4554
rect 9496 4498 9552 4554
rect 9620 4498 9676 4554
rect 9744 4498 9800 4554
rect 7884 4374 7940 4430
rect 8008 4374 8064 4430
rect 8132 4374 8188 4430
rect 8256 4374 8312 4430
rect 8380 4374 8436 4430
rect 8504 4374 8560 4430
rect 8628 4374 8684 4430
rect 8752 4374 8808 4430
rect 8876 4374 8932 4430
rect 9000 4374 9056 4430
rect 9124 4374 9180 4430
rect 9248 4374 9304 4430
rect 9372 4374 9428 4430
rect 9496 4374 9552 4430
rect 9620 4374 9676 4430
rect 9744 4374 9800 4430
rect 7884 4250 7940 4306
rect 8008 4250 8064 4306
rect 8132 4250 8188 4306
rect 8256 4250 8312 4306
rect 8380 4250 8436 4306
rect 8504 4250 8560 4306
rect 8628 4250 8684 4306
rect 8752 4250 8808 4306
rect 8876 4250 8932 4306
rect 9000 4250 9056 4306
rect 9124 4250 9180 4306
rect 9248 4250 9304 4306
rect 9372 4250 9428 4306
rect 9496 4250 9552 4306
rect 9620 4250 9676 4306
rect 9744 4250 9800 4306
rect 7884 4126 7940 4182
rect 8008 4126 8064 4182
rect 8132 4126 8188 4182
rect 8256 4126 8312 4182
rect 8380 4126 8436 4182
rect 8504 4126 8560 4182
rect 8628 4126 8684 4182
rect 8752 4126 8808 4182
rect 8876 4126 8932 4182
rect 9000 4126 9056 4182
rect 9124 4126 9180 4182
rect 9248 4126 9304 4182
rect 9372 4126 9428 4182
rect 9496 4126 9552 4182
rect 9620 4126 9676 4182
rect 9744 4126 9800 4182
rect 7884 4002 7940 4058
rect 8008 4002 8064 4058
rect 8132 4002 8188 4058
rect 8256 4002 8312 4058
rect 8380 4002 8436 4058
rect 8504 4002 8560 4058
rect 8628 4002 8684 4058
rect 8752 4002 8808 4058
rect 8876 4002 8932 4058
rect 9000 4002 9056 4058
rect 9124 4002 9180 4058
rect 9248 4002 9304 4058
rect 9372 4002 9428 4058
rect 9496 4002 9552 4058
rect 9620 4002 9676 4058
rect 9744 4002 9800 4058
rect 7884 3878 7940 3934
rect 8008 3878 8064 3934
rect 8132 3878 8188 3934
rect 8256 3878 8312 3934
rect 8380 3878 8436 3934
rect 8504 3878 8560 3934
rect 8628 3878 8684 3934
rect 8752 3878 8808 3934
rect 8876 3878 8932 3934
rect 9000 3878 9056 3934
rect 9124 3878 9180 3934
rect 9248 3878 9304 3934
rect 9372 3878 9428 3934
rect 9496 3878 9552 3934
rect 9620 3878 9676 3934
rect 9744 3878 9800 3934
rect 7884 3754 7940 3810
rect 8008 3754 8064 3810
rect 8132 3754 8188 3810
rect 8256 3754 8312 3810
rect 8380 3754 8436 3810
rect 8504 3754 8560 3810
rect 8628 3754 8684 3810
rect 8752 3754 8808 3810
rect 8876 3754 8932 3810
rect 9000 3754 9056 3810
rect 9124 3754 9180 3810
rect 9248 3754 9304 3810
rect 9372 3754 9428 3810
rect 9496 3754 9552 3810
rect 9620 3754 9676 3810
rect 9744 3754 9800 3810
rect 7884 3630 7940 3686
rect 8008 3630 8064 3686
rect 8132 3630 8188 3686
rect 8256 3630 8312 3686
rect 8380 3630 8436 3686
rect 8504 3630 8560 3686
rect 8628 3630 8684 3686
rect 8752 3630 8808 3686
rect 8876 3630 8932 3686
rect 9000 3630 9056 3686
rect 9124 3630 9180 3686
rect 9248 3630 9304 3686
rect 9372 3630 9428 3686
rect 9496 3630 9552 3686
rect 9620 3630 9676 3686
rect 9744 3630 9800 3686
rect 7884 3506 7940 3562
rect 8008 3506 8064 3562
rect 8132 3506 8188 3562
rect 8256 3506 8312 3562
rect 8380 3506 8436 3562
rect 8504 3506 8560 3562
rect 8628 3506 8684 3562
rect 8752 3506 8808 3562
rect 8876 3506 8932 3562
rect 9000 3506 9056 3562
rect 9124 3506 9180 3562
rect 9248 3506 9304 3562
rect 9372 3506 9428 3562
rect 9496 3506 9552 3562
rect 9620 3506 9676 3562
rect 9744 3506 9800 3562
rect 7884 3382 7940 3438
rect 8008 3382 8064 3438
rect 8132 3382 8188 3438
rect 8256 3382 8312 3438
rect 8380 3382 8436 3438
rect 8504 3382 8560 3438
rect 8628 3382 8684 3438
rect 8752 3382 8808 3438
rect 8876 3382 8932 3438
rect 9000 3382 9056 3438
rect 9124 3382 9180 3438
rect 9248 3382 9304 3438
rect 9372 3382 9428 3438
rect 9496 3382 9552 3438
rect 9620 3382 9676 3438
rect 9744 3382 9800 3438
rect 7884 3258 7940 3314
rect 8008 3258 8064 3314
rect 8132 3258 8188 3314
rect 8256 3258 8312 3314
rect 8380 3258 8436 3314
rect 8504 3258 8560 3314
rect 8628 3258 8684 3314
rect 8752 3258 8808 3314
rect 8876 3258 8932 3314
rect 9000 3258 9056 3314
rect 9124 3258 9180 3314
rect 9248 3258 9304 3314
rect 9372 3258 9428 3314
rect 9496 3258 9552 3314
rect 9620 3258 9676 3314
rect 9744 3258 9800 3314
rect 7884 3134 7940 3190
rect 8008 3134 8064 3190
rect 8132 3134 8188 3190
rect 8256 3134 8312 3190
rect 8380 3134 8436 3190
rect 8504 3134 8560 3190
rect 8628 3134 8684 3190
rect 8752 3134 8808 3190
rect 8876 3134 8932 3190
rect 9000 3134 9056 3190
rect 9124 3134 9180 3190
rect 9248 3134 9304 3190
rect 9372 3134 9428 3190
rect 9496 3134 9552 3190
rect 9620 3134 9676 3190
rect 9744 3134 9800 3190
rect 7884 3010 7940 3066
rect 8008 3010 8064 3066
rect 8132 3010 8188 3066
rect 8256 3010 8312 3066
rect 8380 3010 8436 3066
rect 8504 3010 8560 3066
rect 8628 3010 8684 3066
rect 8752 3010 8808 3066
rect 8876 3010 8932 3066
rect 9000 3010 9056 3066
rect 9124 3010 9180 3066
rect 9248 3010 9304 3066
rect 9372 3010 9428 3066
rect 9496 3010 9552 3066
rect 9620 3010 9676 3066
rect 9744 3010 9800 3066
rect 7884 2886 7940 2942
rect 8008 2886 8064 2942
rect 8132 2886 8188 2942
rect 8256 2886 8312 2942
rect 8380 2886 8436 2942
rect 8504 2886 8560 2942
rect 8628 2886 8684 2942
rect 8752 2886 8808 2942
rect 8876 2886 8932 2942
rect 9000 2886 9056 2942
rect 9124 2886 9180 2942
rect 9248 2886 9304 2942
rect 9372 2886 9428 2942
rect 9496 2886 9552 2942
rect 9620 2886 9676 2942
rect 9744 2886 9800 2942
rect 7884 2762 7940 2818
rect 8008 2762 8064 2818
rect 8132 2762 8188 2818
rect 8256 2762 8312 2818
rect 8380 2762 8436 2818
rect 8504 2762 8560 2818
rect 8628 2762 8684 2818
rect 8752 2762 8808 2818
rect 8876 2762 8932 2818
rect 9000 2762 9056 2818
rect 9124 2762 9180 2818
rect 9248 2762 9304 2818
rect 9372 2762 9428 2818
rect 9496 2762 9552 2818
rect 9620 2762 9676 2818
rect 9744 2762 9800 2818
rect 7884 2638 7940 2694
rect 8008 2638 8064 2694
rect 8132 2638 8188 2694
rect 8256 2638 8312 2694
rect 8380 2638 8436 2694
rect 8504 2638 8560 2694
rect 8628 2638 8684 2694
rect 8752 2638 8808 2694
rect 8876 2638 8932 2694
rect 9000 2638 9056 2694
rect 9124 2638 9180 2694
rect 9248 2638 9304 2694
rect 9372 2638 9428 2694
rect 9496 2638 9552 2694
rect 9620 2638 9676 2694
rect 9744 2638 9800 2694
rect 7884 2514 7940 2570
rect 8008 2514 8064 2570
rect 8132 2514 8188 2570
rect 8256 2514 8312 2570
rect 8380 2514 8436 2570
rect 8504 2514 8560 2570
rect 8628 2514 8684 2570
rect 8752 2514 8808 2570
rect 8876 2514 8932 2570
rect 9000 2514 9056 2570
rect 9124 2514 9180 2570
rect 9248 2514 9304 2570
rect 9372 2514 9428 2570
rect 9496 2514 9552 2570
rect 9620 2514 9676 2570
rect 9744 2514 9800 2570
rect 7884 2390 7940 2446
rect 8008 2390 8064 2446
rect 8132 2390 8188 2446
rect 8256 2390 8312 2446
rect 8380 2390 8436 2446
rect 8504 2390 8560 2446
rect 8628 2390 8684 2446
rect 8752 2390 8808 2446
rect 8876 2390 8932 2446
rect 9000 2390 9056 2446
rect 9124 2390 9180 2446
rect 9248 2390 9304 2446
rect 9372 2390 9428 2446
rect 9496 2390 9552 2446
rect 9620 2390 9676 2446
rect 9744 2390 9800 2446
rect 7884 2266 7940 2322
rect 8008 2266 8064 2322
rect 8132 2266 8188 2322
rect 8256 2266 8312 2322
rect 8380 2266 8436 2322
rect 8504 2266 8560 2322
rect 8628 2266 8684 2322
rect 8752 2266 8808 2322
rect 8876 2266 8932 2322
rect 9000 2266 9056 2322
rect 9124 2266 9180 2322
rect 9248 2266 9304 2322
rect 9372 2266 9428 2322
rect 9496 2266 9552 2322
rect 9620 2266 9676 2322
rect 9744 2266 9800 2322
rect 7884 2142 7940 2198
rect 8008 2142 8064 2198
rect 8132 2142 8188 2198
rect 8256 2142 8312 2198
rect 8380 2142 8436 2198
rect 8504 2142 8560 2198
rect 8628 2142 8684 2198
rect 8752 2142 8808 2198
rect 8876 2142 8932 2198
rect 9000 2142 9056 2198
rect 9124 2142 9180 2198
rect 9248 2142 9304 2198
rect 9372 2142 9428 2198
rect 9496 2142 9552 2198
rect 9620 2142 9676 2198
rect 9744 2142 9800 2198
rect 7884 2018 7940 2074
rect 8008 2018 8064 2074
rect 8132 2018 8188 2074
rect 8256 2018 8312 2074
rect 8380 2018 8436 2074
rect 8504 2018 8560 2074
rect 8628 2018 8684 2074
rect 8752 2018 8808 2074
rect 8876 2018 8932 2074
rect 9000 2018 9056 2074
rect 9124 2018 9180 2074
rect 9248 2018 9304 2074
rect 9372 2018 9428 2074
rect 9496 2018 9552 2074
rect 9620 2018 9676 2074
rect 9744 2018 9800 2074
rect 7884 1894 7940 1950
rect 8008 1894 8064 1950
rect 8132 1894 8188 1950
rect 8256 1894 8312 1950
rect 8380 1894 8436 1950
rect 8504 1894 8560 1950
rect 8628 1894 8684 1950
rect 8752 1894 8808 1950
rect 8876 1894 8932 1950
rect 9000 1894 9056 1950
rect 9124 1894 9180 1950
rect 9248 1894 9304 1950
rect 9372 1894 9428 1950
rect 9496 1894 9552 1950
rect 9620 1894 9676 1950
rect 9744 1894 9800 1950
rect 7884 1770 7940 1826
rect 8008 1770 8064 1826
rect 8132 1770 8188 1826
rect 8256 1770 8312 1826
rect 8380 1770 8436 1826
rect 8504 1770 8560 1826
rect 8628 1770 8684 1826
rect 8752 1770 8808 1826
rect 8876 1770 8932 1826
rect 9000 1770 9056 1826
rect 9124 1770 9180 1826
rect 9248 1770 9304 1826
rect 9372 1770 9428 1826
rect 9496 1770 9552 1826
rect 9620 1770 9676 1826
rect 9744 1770 9800 1826
rect 7884 1646 7940 1702
rect 8008 1646 8064 1702
rect 8132 1646 8188 1702
rect 8256 1646 8312 1702
rect 8380 1646 8436 1702
rect 8504 1646 8560 1702
rect 8628 1646 8684 1702
rect 8752 1646 8808 1702
rect 8876 1646 8932 1702
rect 9000 1646 9056 1702
rect 9124 1646 9180 1702
rect 9248 1646 9304 1702
rect 9372 1646 9428 1702
rect 9496 1646 9552 1702
rect 9620 1646 9676 1702
rect 9744 1646 9800 1702
rect 10254 4498 10310 4554
rect 10378 4498 10434 4554
rect 10502 4498 10558 4554
rect 10626 4498 10682 4554
rect 10750 4498 10806 4554
rect 10874 4498 10930 4554
rect 10998 4498 11054 4554
rect 11122 4498 11178 4554
rect 11246 4498 11302 4554
rect 11370 4498 11426 4554
rect 11494 4498 11550 4554
rect 11618 4498 11674 4554
rect 11742 4498 11798 4554
rect 11866 4498 11922 4554
rect 11990 4498 12046 4554
rect 12114 4498 12170 4554
rect 10254 4374 10310 4430
rect 10378 4374 10434 4430
rect 10502 4374 10558 4430
rect 10626 4374 10682 4430
rect 10750 4374 10806 4430
rect 10874 4374 10930 4430
rect 10998 4374 11054 4430
rect 11122 4374 11178 4430
rect 11246 4374 11302 4430
rect 11370 4374 11426 4430
rect 11494 4374 11550 4430
rect 11618 4374 11674 4430
rect 11742 4374 11798 4430
rect 11866 4374 11922 4430
rect 11990 4374 12046 4430
rect 12114 4374 12170 4430
rect 10254 4250 10310 4306
rect 10378 4250 10434 4306
rect 10502 4250 10558 4306
rect 10626 4250 10682 4306
rect 10750 4250 10806 4306
rect 10874 4250 10930 4306
rect 10998 4250 11054 4306
rect 11122 4250 11178 4306
rect 11246 4250 11302 4306
rect 11370 4250 11426 4306
rect 11494 4250 11550 4306
rect 11618 4250 11674 4306
rect 11742 4250 11798 4306
rect 11866 4250 11922 4306
rect 11990 4250 12046 4306
rect 12114 4250 12170 4306
rect 10254 4126 10310 4182
rect 10378 4126 10434 4182
rect 10502 4126 10558 4182
rect 10626 4126 10682 4182
rect 10750 4126 10806 4182
rect 10874 4126 10930 4182
rect 10998 4126 11054 4182
rect 11122 4126 11178 4182
rect 11246 4126 11302 4182
rect 11370 4126 11426 4182
rect 11494 4126 11550 4182
rect 11618 4126 11674 4182
rect 11742 4126 11798 4182
rect 11866 4126 11922 4182
rect 11990 4126 12046 4182
rect 12114 4126 12170 4182
rect 10254 4002 10310 4058
rect 10378 4002 10434 4058
rect 10502 4002 10558 4058
rect 10626 4002 10682 4058
rect 10750 4002 10806 4058
rect 10874 4002 10930 4058
rect 10998 4002 11054 4058
rect 11122 4002 11178 4058
rect 11246 4002 11302 4058
rect 11370 4002 11426 4058
rect 11494 4002 11550 4058
rect 11618 4002 11674 4058
rect 11742 4002 11798 4058
rect 11866 4002 11922 4058
rect 11990 4002 12046 4058
rect 12114 4002 12170 4058
rect 10254 3878 10310 3934
rect 10378 3878 10434 3934
rect 10502 3878 10558 3934
rect 10626 3878 10682 3934
rect 10750 3878 10806 3934
rect 10874 3878 10930 3934
rect 10998 3878 11054 3934
rect 11122 3878 11178 3934
rect 11246 3878 11302 3934
rect 11370 3878 11426 3934
rect 11494 3878 11550 3934
rect 11618 3878 11674 3934
rect 11742 3878 11798 3934
rect 11866 3878 11922 3934
rect 11990 3878 12046 3934
rect 12114 3878 12170 3934
rect 10254 3754 10310 3810
rect 10378 3754 10434 3810
rect 10502 3754 10558 3810
rect 10626 3754 10682 3810
rect 10750 3754 10806 3810
rect 10874 3754 10930 3810
rect 10998 3754 11054 3810
rect 11122 3754 11178 3810
rect 11246 3754 11302 3810
rect 11370 3754 11426 3810
rect 11494 3754 11550 3810
rect 11618 3754 11674 3810
rect 11742 3754 11798 3810
rect 11866 3754 11922 3810
rect 11990 3754 12046 3810
rect 12114 3754 12170 3810
rect 10254 3630 10310 3686
rect 10378 3630 10434 3686
rect 10502 3630 10558 3686
rect 10626 3630 10682 3686
rect 10750 3630 10806 3686
rect 10874 3630 10930 3686
rect 10998 3630 11054 3686
rect 11122 3630 11178 3686
rect 11246 3630 11302 3686
rect 11370 3630 11426 3686
rect 11494 3630 11550 3686
rect 11618 3630 11674 3686
rect 11742 3630 11798 3686
rect 11866 3630 11922 3686
rect 11990 3630 12046 3686
rect 12114 3630 12170 3686
rect 10254 3506 10310 3562
rect 10378 3506 10434 3562
rect 10502 3506 10558 3562
rect 10626 3506 10682 3562
rect 10750 3506 10806 3562
rect 10874 3506 10930 3562
rect 10998 3506 11054 3562
rect 11122 3506 11178 3562
rect 11246 3506 11302 3562
rect 11370 3506 11426 3562
rect 11494 3506 11550 3562
rect 11618 3506 11674 3562
rect 11742 3506 11798 3562
rect 11866 3506 11922 3562
rect 11990 3506 12046 3562
rect 12114 3506 12170 3562
rect 10254 3382 10310 3438
rect 10378 3382 10434 3438
rect 10502 3382 10558 3438
rect 10626 3382 10682 3438
rect 10750 3382 10806 3438
rect 10874 3382 10930 3438
rect 10998 3382 11054 3438
rect 11122 3382 11178 3438
rect 11246 3382 11302 3438
rect 11370 3382 11426 3438
rect 11494 3382 11550 3438
rect 11618 3382 11674 3438
rect 11742 3382 11798 3438
rect 11866 3382 11922 3438
rect 11990 3382 12046 3438
rect 12114 3382 12170 3438
rect 10254 3258 10310 3314
rect 10378 3258 10434 3314
rect 10502 3258 10558 3314
rect 10626 3258 10682 3314
rect 10750 3258 10806 3314
rect 10874 3258 10930 3314
rect 10998 3258 11054 3314
rect 11122 3258 11178 3314
rect 11246 3258 11302 3314
rect 11370 3258 11426 3314
rect 11494 3258 11550 3314
rect 11618 3258 11674 3314
rect 11742 3258 11798 3314
rect 11866 3258 11922 3314
rect 11990 3258 12046 3314
rect 12114 3258 12170 3314
rect 10254 3134 10310 3190
rect 10378 3134 10434 3190
rect 10502 3134 10558 3190
rect 10626 3134 10682 3190
rect 10750 3134 10806 3190
rect 10874 3134 10930 3190
rect 10998 3134 11054 3190
rect 11122 3134 11178 3190
rect 11246 3134 11302 3190
rect 11370 3134 11426 3190
rect 11494 3134 11550 3190
rect 11618 3134 11674 3190
rect 11742 3134 11798 3190
rect 11866 3134 11922 3190
rect 11990 3134 12046 3190
rect 12114 3134 12170 3190
rect 10254 3010 10310 3066
rect 10378 3010 10434 3066
rect 10502 3010 10558 3066
rect 10626 3010 10682 3066
rect 10750 3010 10806 3066
rect 10874 3010 10930 3066
rect 10998 3010 11054 3066
rect 11122 3010 11178 3066
rect 11246 3010 11302 3066
rect 11370 3010 11426 3066
rect 11494 3010 11550 3066
rect 11618 3010 11674 3066
rect 11742 3010 11798 3066
rect 11866 3010 11922 3066
rect 11990 3010 12046 3066
rect 12114 3010 12170 3066
rect 10254 2886 10310 2942
rect 10378 2886 10434 2942
rect 10502 2886 10558 2942
rect 10626 2886 10682 2942
rect 10750 2886 10806 2942
rect 10874 2886 10930 2942
rect 10998 2886 11054 2942
rect 11122 2886 11178 2942
rect 11246 2886 11302 2942
rect 11370 2886 11426 2942
rect 11494 2886 11550 2942
rect 11618 2886 11674 2942
rect 11742 2886 11798 2942
rect 11866 2886 11922 2942
rect 11990 2886 12046 2942
rect 12114 2886 12170 2942
rect 10254 2762 10310 2818
rect 10378 2762 10434 2818
rect 10502 2762 10558 2818
rect 10626 2762 10682 2818
rect 10750 2762 10806 2818
rect 10874 2762 10930 2818
rect 10998 2762 11054 2818
rect 11122 2762 11178 2818
rect 11246 2762 11302 2818
rect 11370 2762 11426 2818
rect 11494 2762 11550 2818
rect 11618 2762 11674 2818
rect 11742 2762 11798 2818
rect 11866 2762 11922 2818
rect 11990 2762 12046 2818
rect 12114 2762 12170 2818
rect 10254 2638 10310 2694
rect 10378 2638 10434 2694
rect 10502 2638 10558 2694
rect 10626 2638 10682 2694
rect 10750 2638 10806 2694
rect 10874 2638 10930 2694
rect 10998 2638 11054 2694
rect 11122 2638 11178 2694
rect 11246 2638 11302 2694
rect 11370 2638 11426 2694
rect 11494 2638 11550 2694
rect 11618 2638 11674 2694
rect 11742 2638 11798 2694
rect 11866 2638 11922 2694
rect 11990 2638 12046 2694
rect 12114 2638 12170 2694
rect 10254 2514 10310 2570
rect 10378 2514 10434 2570
rect 10502 2514 10558 2570
rect 10626 2514 10682 2570
rect 10750 2514 10806 2570
rect 10874 2514 10930 2570
rect 10998 2514 11054 2570
rect 11122 2514 11178 2570
rect 11246 2514 11302 2570
rect 11370 2514 11426 2570
rect 11494 2514 11550 2570
rect 11618 2514 11674 2570
rect 11742 2514 11798 2570
rect 11866 2514 11922 2570
rect 11990 2514 12046 2570
rect 12114 2514 12170 2570
rect 10254 2390 10310 2446
rect 10378 2390 10434 2446
rect 10502 2390 10558 2446
rect 10626 2390 10682 2446
rect 10750 2390 10806 2446
rect 10874 2390 10930 2446
rect 10998 2390 11054 2446
rect 11122 2390 11178 2446
rect 11246 2390 11302 2446
rect 11370 2390 11426 2446
rect 11494 2390 11550 2446
rect 11618 2390 11674 2446
rect 11742 2390 11798 2446
rect 11866 2390 11922 2446
rect 11990 2390 12046 2446
rect 12114 2390 12170 2446
rect 10254 2266 10310 2322
rect 10378 2266 10434 2322
rect 10502 2266 10558 2322
rect 10626 2266 10682 2322
rect 10750 2266 10806 2322
rect 10874 2266 10930 2322
rect 10998 2266 11054 2322
rect 11122 2266 11178 2322
rect 11246 2266 11302 2322
rect 11370 2266 11426 2322
rect 11494 2266 11550 2322
rect 11618 2266 11674 2322
rect 11742 2266 11798 2322
rect 11866 2266 11922 2322
rect 11990 2266 12046 2322
rect 12114 2266 12170 2322
rect 10254 2142 10310 2198
rect 10378 2142 10434 2198
rect 10502 2142 10558 2198
rect 10626 2142 10682 2198
rect 10750 2142 10806 2198
rect 10874 2142 10930 2198
rect 10998 2142 11054 2198
rect 11122 2142 11178 2198
rect 11246 2142 11302 2198
rect 11370 2142 11426 2198
rect 11494 2142 11550 2198
rect 11618 2142 11674 2198
rect 11742 2142 11798 2198
rect 11866 2142 11922 2198
rect 11990 2142 12046 2198
rect 12114 2142 12170 2198
rect 10254 2018 10310 2074
rect 10378 2018 10434 2074
rect 10502 2018 10558 2074
rect 10626 2018 10682 2074
rect 10750 2018 10806 2074
rect 10874 2018 10930 2074
rect 10998 2018 11054 2074
rect 11122 2018 11178 2074
rect 11246 2018 11302 2074
rect 11370 2018 11426 2074
rect 11494 2018 11550 2074
rect 11618 2018 11674 2074
rect 11742 2018 11798 2074
rect 11866 2018 11922 2074
rect 11990 2018 12046 2074
rect 12114 2018 12170 2074
rect 10254 1894 10310 1950
rect 10378 1894 10434 1950
rect 10502 1894 10558 1950
rect 10626 1894 10682 1950
rect 10750 1894 10806 1950
rect 10874 1894 10930 1950
rect 10998 1894 11054 1950
rect 11122 1894 11178 1950
rect 11246 1894 11302 1950
rect 11370 1894 11426 1950
rect 11494 1894 11550 1950
rect 11618 1894 11674 1950
rect 11742 1894 11798 1950
rect 11866 1894 11922 1950
rect 11990 1894 12046 1950
rect 12114 1894 12170 1950
rect 10254 1770 10310 1826
rect 10378 1770 10434 1826
rect 10502 1770 10558 1826
rect 10626 1770 10682 1826
rect 10750 1770 10806 1826
rect 10874 1770 10930 1826
rect 10998 1770 11054 1826
rect 11122 1770 11178 1826
rect 11246 1770 11302 1826
rect 11370 1770 11426 1826
rect 11494 1770 11550 1826
rect 11618 1770 11674 1826
rect 11742 1770 11798 1826
rect 11866 1770 11922 1826
rect 11990 1770 12046 1826
rect 12114 1770 12170 1826
rect 10254 1646 10310 1702
rect 10378 1646 10434 1702
rect 10502 1646 10558 1702
rect 10626 1646 10682 1702
rect 10750 1646 10806 1702
rect 10874 1646 10930 1702
rect 10998 1646 11054 1702
rect 11122 1646 11178 1702
rect 11246 1646 11302 1702
rect 11370 1646 11426 1702
rect 11494 1646 11550 1702
rect 11618 1646 11674 1702
rect 11742 1646 11798 1702
rect 11866 1646 11922 1702
rect 11990 1646 12046 1702
rect 12114 1646 12170 1702
rect 12871 4498 12927 4554
rect 12995 4498 13051 4554
rect 13119 4498 13175 4554
rect 13243 4498 13299 4554
rect 13367 4498 13423 4554
rect 13491 4498 13547 4554
rect 13615 4498 13671 4554
rect 13739 4498 13795 4554
rect 13863 4498 13919 4554
rect 13987 4498 14043 4554
rect 14111 4498 14167 4554
rect 14235 4498 14291 4554
rect 14359 4498 14415 4554
rect 14483 4498 14539 4554
rect 14607 4498 14663 4554
rect 12871 4374 12927 4430
rect 12995 4374 13051 4430
rect 13119 4374 13175 4430
rect 13243 4374 13299 4430
rect 13367 4374 13423 4430
rect 13491 4374 13547 4430
rect 13615 4374 13671 4430
rect 13739 4374 13795 4430
rect 13863 4374 13919 4430
rect 13987 4374 14043 4430
rect 14111 4374 14167 4430
rect 14235 4374 14291 4430
rect 14359 4374 14415 4430
rect 14483 4374 14539 4430
rect 14607 4374 14663 4430
rect 12871 4250 12927 4306
rect 12995 4250 13051 4306
rect 13119 4250 13175 4306
rect 13243 4250 13299 4306
rect 13367 4250 13423 4306
rect 13491 4250 13547 4306
rect 13615 4250 13671 4306
rect 13739 4250 13795 4306
rect 13863 4250 13919 4306
rect 13987 4250 14043 4306
rect 14111 4250 14167 4306
rect 14235 4250 14291 4306
rect 14359 4250 14415 4306
rect 14483 4250 14539 4306
rect 14607 4250 14663 4306
rect 12871 4126 12927 4182
rect 12995 4126 13051 4182
rect 13119 4126 13175 4182
rect 13243 4126 13299 4182
rect 13367 4126 13423 4182
rect 13491 4126 13547 4182
rect 13615 4126 13671 4182
rect 13739 4126 13795 4182
rect 13863 4126 13919 4182
rect 13987 4126 14043 4182
rect 14111 4126 14167 4182
rect 14235 4126 14291 4182
rect 14359 4126 14415 4182
rect 14483 4126 14539 4182
rect 14607 4126 14663 4182
rect 12871 4002 12927 4058
rect 12995 4002 13051 4058
rect 13119 4002 13175 4058
rect 13243 4002 13299 4058
rect 13367 4002 13423 4058
rect 13491 4002 13547 4058
rect 13615 4002 13671 4058
rect 13739 4002 13795 4058
rect 13863 4002 13919 4058
rect 13987 4002 14043 4058
rect 14111 4002 14167 4058
rect 14235 4002 14291 4058
rect 14359 4002 14415 4058
rect 14483 4002 14539 4058
rect 14607 4002 14663 4058
rect 12871 3878 12927 3934
rect 12995 3878 13051 3934
rect 13119 3878 13175 3934
rect 13243 3878 13299 3934
rect 13367 3878 13423 3934
rect 13491 3878 13547 3934
rect 13615 3878 13671 3934
rect 13739 3878 13795 3934
rect 13863 3878 13919 3934
rect 13987 3878 14043 3934
rect 14111 3878 14167 3934
rect 14235 3878 14291 3934
rect 14359 3878 14415 3934
rect 14483 3878 14539 3934
rect 14607 3878 14663 3934
rect 12871 3754 12927 3810
rect 12995 3754 13051 3810
rect 13119 3754 13175 3810
rect 13243 3754 13299 3810
rect 13367 3754 13423 3810
rect 13491 3754 13547 3810
rect 13615 3754 13671 3810
rect 13739 3754 13795 3810
rect 13863 3754 13919 3810
rect 13987 3754 14043 3810
rect 14111 3754 14167 3810
rect 14235 3754 14291 3810
rect 14359 3754 14415 3810
rect 14483 3754 14539 3810
rect 14607 3754 14663 3810
rect 12871 3630 12927 3686
rect 12995 3630 13051 3686
rect 13119 3630 13175 3686
rect 13243 3630 13299 3686
rect 13367 3630 13423 3686
rect 13491 3630 13547 3686
rect 13615 3630 13671 3686
rect 13739 3630 13795 3686
rect 13863 3630 13919 3686
rect 13987 3630 14043 3686
rect 14111 3630 14167 3686
rect 14235 3630 14291 3686
rect 14359 3630 14415 3686
rect 14483 3630 14539 3686
rect 14607 3630 14663 3686
rect 12871 3506 12927 3562
rect 12995 3506 13051 3562
rect 13119 3506 13175 3562
rect 13243 3506 13299 3562
rect 13367 3506 13423 3562
rect 13491 3506 13547 3562
rect 13615 3506 13671 3562
rect 13739 3506 13795 3562
rect 13863 3506 13919 3562
rect 13987 3506 14043 3562
rect 14111 3506 14167 3562
rect 14235 3506 14291 3562
rect 14359 3506 14415 3562
rect 14483 3506 14539 3562
rect 14607 3506 14663 3562
rect 12871 3382 12927 3438
rect 12995 3382 13051 3438
rect 13119 3382 13175 3438
rect 13243 3382 13299 3438
rect 13367 3382 13423 3438
rect 13491 3382 13547 3438
rect 13615 3382 13671 3438
rect 13739 3382 13795 3438
rect 13863 3382 13919 3438
rect 13987 3382 14043 3438
rect 14111 3382 14167 3438
rect 14235 3382 14291 3438
rect 14359 3382 14415 3438
rect 14483 3382 14539 3438
rect 14607 3382 14663 3438
rect 12871 3258 12927 3314
rect 12995 3258 13051 3314
rect 13119 3258 13175 3314
rect 13243 3258 13299 3314
rect 13367 3258 13423 3314
rect 13491 3258 13547 3314
rect 13615 3258 13671 3314
rect 13739 3258 13795 3314
rect 13863 3258 13919 3314
rect 13987 3258 14043 3314
rect 14111 3258 14167 3314
rect 14235 3258 14291 3314
rect 14359 3258 14415 3314
rect 14483 3258 14539 3314
rect 14607 3258 14663 3314
rect 12871 3134 12927 3190
rect 12995 3134 13051 3190
rect 13119 3134 13175 3190
rect 13243 3134 13299 3190
rect 13367 3134 13423 3190
rect 13491 3134 13547 3190
rect 13615 3134 13671 3190
rect 13739 3134 13795 3190
rect 13863 3134 13919 3190
rect 13987 3134 14043 3190
rect 14111 3134 14167 3190
rect 14235 3134 14291 3190
rect 14359 3134 14415 3190
rect 14483 3134 14539 3190
rect 14607 3134 14663 3190
rect 12871 3010 12927 3066
rect 12995 3010 13051 3066
rect 13119 3010 13175 3066
rect 13243 3010 13299 3066
rect 13367 3010 13423 3066
rect 13491 3010 13547 3066
rect 13615 3010 13671 3066
rect 13739 3010 13795 3066
rect 13863 3010 13919 3066
rect 13987 3010 14043 3066
rect 14111 3010 14167 3066
rect 14235 3010 14291 3066
rect 14359 3010 14415 3066
rect 14483 3010 14539 3066
rect 14607 3010 14663 3066
rect 12871 2886 12927 2942
rect 12995 2886 13051 2942
rect 13119 2886 13175 2942
rect 13243 2886 13299 2942
rect 13367 2886 13423 2942
rect 13491 2886 13547 2942
rect 13615 2886 13671 2942
rect 13739 2886 13795 2942
rect 13863 2886 13919 2942
rect 13987 2886 14043 2942
rect 14111 2886 14167 2942
rect 14235 2886 14291 2942
rect 14359 2886 14415 2942
rect 14483 2886 14539 2942
rect 14607 2886 14663 2942
rect 12871 2762 12927 2818
rect 12995 2762 13051 2818
rect 13119 2762 13175 2818
rect 13243 2762 13299 2818
rect 13367 2762 13423 2818
rect 13491 2762 13547 2818
rect 13615 2762 13671 2818
rect 13739 2762 13795 2818
rect 13863 2762 13919 2818
rect 13987 2762 14043 2818
rect 14111 2762 14167 2818
rect 14235 2762 14291 2818
rect 14359 2762 14415 2818
rect 14483 2762 14539 2818
rect 14607 2762 14663 2818
rect 12871 2638 12927 2694
rect 12995 2638 13051 2694
rect 13119 2638 13175 2694
rect 13243 2638 13299 2694
rect 13367 2638 13423 2694
rect 13491 2638 13547 2694
rect 13615 2638 13671 2694
rect 13739 2638 13795 2694
rect 13863 2638 13919 2694
rect 13987 2638 14043 2694
rect 14111 2638 14167 2694
rect 14235 2638 14291 2694
rect 14359 2638 14415 2694
rect 14483 2638 14539 2694
rect 14607 2638 14663 2694
rect 12871 2514 12927 2570
rect 12995 2514 13051 2570
rect 13119 2514 13175 2570
rect 13243 2514 13299 2570
rect 13367 2514 13423 2570
rect 13491 2514 13547 2570
rect 13615 2514 13671 2570
rect 13739 2514 13795 2570
rect 13863 2514 13919 2570
rect 13987 2514 14043 2570
rect 14111 2514 14167 2570
rect 14235 2514 14291 2570
rect 14359 2514 14415 2570
rect 14483 2514 14539 2570
rect 14607 2514 14663 2570
rect 12871 2390 12927 2446
rect 12995 2390 13051 2446
rect 13119 2390 13175 2446
rect 13243 2390 13299 2446
rect 13367 2390 13423 2446
rect 13491 2390 13547 2446
rect 13615 2390 13671 2446
rect 13739 2390 13795 2446
rect 13863 2390 13919 2446
rect 13987 2390 14043 2446
rect 14111 2390 14167 2446
rect 14235 2390 14291 2446
rect 14359 2390 14415 2446
rect 14483 2390 14539 2446
rect 14607 2390 14663 2446
rect 12871 2266 12927 2322
rect 12995 2266 13051 2322
rect 13119 2266 13175 2322
rect 13243 2266 13299 2322
rect 13367 2266 13423 2322
rect 13491 2266 13547 2322
rect 13615 2266 13671 2322
rect 13739 2266 13795 2322
rect 13863 2266 13919 2322
rect 13987 2266 14043 2322
rect 14111 2266 14167 2322
rect 14235 2266 14291 2322
rect 14359 2266 14415 2322
rect 14483 2266 14539 2322
rect 14607 2266 14663 2322
rect 12871 2142 12927 2198
rect 12995 2142 13051 2198
rect 13119 2142 13175 2198
rect 13243 2142 13299 2198
rect 13367 2142 13423 2198
rect 13491 2142 13547 2198
rect 13615 2142 13671 2198
rect 13739 2142 13795 2198
rect 13863 2142 13919 2198
rect 13987 2142 14043 2198
rect 14111 2142 14167 2198
rect 14235 2142 14291 2198
rect 14359 2142 14415 2198
rect 14483 2142 14539 2198
rect 14607 2142 14663 2198
rect 12871 2018 12927 2074
rect 12995 2018 13051 2074
rect 13119 2018 13175 2074
rect 13243 2018 13299 2074
rect 13367 2018 13423 2074
rect 13491 2018 13547 2074
rect 13615 2018 13671 2074
rect 13739 2018 13795 2074
rect 13863 2018 13919 2074
rect 13987 2018 14043 2074
rect 14111 2018 14167 2074
rect 14235 2018 14291 2074
rect 14359 2018 14415 2074
rect 14483 2018 14539 2074
rect 14607 2018 14663 2074
rect 12871 1894 12927 1950
rect 12995 1894 13051 1950
rect 13119 1894 13175 1950
rect 13243 1894 13299 1950
rect 13367 1894 13423 1950
rect 13491 1894 13547 1950
rect 13615 1894 13671 1950
rect 13739 1894 13795 1950
rect 13863 1894 13919 1950
rect 13987 1894 14043 1950
rect 14111 1894 14167 1950
rect 14235 1894 14291 1950
rect 14359 1894 14415 1950
rect 14483 1894 14539 1950
rect 14607 1894 14663 1950
rect 12871 1770 12927 1826
rect 12995 1770 13051 1826
rect 13119 1770 13175 1826
rect 13243 1770 13299 1826
rect 13367 1770 13423 1826
rect 13491 1770 13547 1826
rect 13615 1770 13671 1826
rect 13739 1770 13795 1826
rect 13863 1770 13919 1826
rect 13987 1770 14043 1826
rect 14111 1770 14167 1826
rect 14235 1770 14291 1826
rect 14359 1770 14415 1826
rect 14483 1770 14539 1826
rect 14607 1770 14663 1826
rect 12871 1646 12927 1702
rect 12995 1646 13051 1702
rect 13119 1646 13175 1702
rect 13243 1646 13299 1702
rect 13367 1646 13423 1702
rect 13491 1646 13547 1702
rect 13615 1646 13671 1702
rect 13739 1646 13795 1702
rect 13863 1646 13919 1702
rect 13987 1646 14043 1702
rect 14111 1646 14167 1702
rect 14235 1646 14291 1702
rect 14359 1646 14415 1702
rect 14483 1646 14539 1702
rect 14607 1646 14663 1702
rect 14902 4584 14958 4586
rect 14902 4532 14904 4584
rect 14904 4532 14956 4584
rect 14956 4532 14958 4584
rect 14902 4476 14958 4532
rect 14902 4424 14904 4476
rect 14904 4424 14956 4476
rect 14956 4424 14958 4476
rect 14902 4368 14958 4424
rect 14902 4316 14904 4368
rect 14904 4316 14956 4368
rect 14956 4316 14958 4368
rect 14902 4260 14958 4316
rect 14902 4208 14904 4260
rect 14904 4208 14956 4260
rect 14956 4208 14958 4260
rect 14902 4152 14958 4208
rect 14902 4100 14904 4152
rect 14904 4100 14956 4152
rect 14956 4100 14958 4152
rect 14902 4044 14958 4100
rect 14902 3992 14904 4044
rect 14904 3992 14956 4044
rect 14956 3992 14958 4044
rect 14902 3936 14958 3992
rect 14902 3884 14904 3936
rect 14904 3884 14956 3936
rect 14956 3884 14958 3936
rect 14902 3828 14958 3884
rect 14902 3776 14904 3828
rect 14904 3776 14956 3828
rect 14956 3776 14958 3828
rect 14902 3720 14958 3776
rect 14902 3668 14904 3720
rect 14904 3668 14956 3720
rect 14956 3668 14958 3720
rect 14902 3612 14958 3668
rect 14902 3560 14904 3612
rect 14904 3560 14956 3612
rect 14956 3560 14958 3612
rect 14902 3504 14958 3560
rect 14902 3452 14904 3504
rect 14904 3452 14956 3504
rect 14956 3452 14958 3504
rect 14902 3396 14958 3452
rect 14902 3344 14904 3396
rect 14904 3344 14956 3396
rect 14956 3344 14958 3396
rect 14902 3288 14958 3344
rect 14902 3236 14904 3288
rect 14904 3236 14956 3288
rect 14956 3236 14958 3288
rect 14902 3180 14958 3236
rect 14902 3128 14904 3180
rect 14904 3128 14956 3180
rect 14956 3128 14958 3180
rect 14902 3072 14958 3128
rect 14902 3020 14904 3072
rect 14904 3020 14956 3072
rect 14956 3020 14958 3072
rect 14902 2964 14958 3020
rect 14902 2912 14904 2964
rect 14904 2912 14956 2964
rect 14956 2912 14958 2964
rect 14902 2856 14958 2912
rect 14902 2804 14904 2856
rect 14904 2804 14956 2856
rect 14956 2804 14958 2856
rect 14902 2748 14958 2804
rect 14902 2696 14904 2748
rect 14904 2696 14956 2748
rect 14956 2696 14958 2748
rect 14902 2640 14958 2696
rect 14902 2588 14904 2640
rect 14904 2588 14956 2640
rect 14956 2588 14958 2640
rect 14902 2532 14958 2588
rect 14902 2480 14904 2532
rect 14904 2480 14956 2532
rect 14956 2480 14958 2532
rect 14902 2424 14958 2480
rect 14902 2372 14904 2424
rect 14904 2372 14956 2424
rect 14956 2372 14958 2424
rect 14902 2316 14958 2372
rect 14902 2264 14904 2316
rect 14904 2264 14956 2316
rect 14956 2264 14958 2316
rect 14902 2208 14958 2264
rect 14902 2156 14904 2208
rect 14904 2156 14956 2208
rect 14956 2156 14958 2208
rect 14902 2100 14958 2156
rect 14902 2048 14904 2100
rect 14904 2048 14956 2100
rect 14956 2048 14958 2100
rect 14902 1992 14958 2048
rect 14902 1940 14904 1992
rect 14904 1940 14956 1992
rect 14956 1940 14958 1992
rect 14902 1884 14958 1940
rect 14902 1832 14904 1884
rect 14904 1832 14956 1884
rect 14956 1832 14958 1884
rect 14902 1776 14958 1832
rect 14902 1724 14904 1776
rect 14904 1724 14956 1776
rect 14956 1724 14958 1776
rect 14902 1668 14958 1724
rect 14902 1616 14904 1668
rect 14904 1616 14956 1668
rect 14956 1616 14958 1668
rect 14902 1614 14958 1616
<< metal3 >>
rect 10 57261 86 57271
rect 10 56017 20 57261
rect 76 56017 86 57261
rect 14892 57261 14968 57271
rect 305 57225 2117 57235
rect 305 57169 315 57225
rect 371 57169 439 57225
rect 495 57169 563 57225
rect 619 57169 687 57225
rect 743 57169 811 57225
rect 867 57169 935 57225
rect 991 57169 1059 57225
rect 1115 57169 1183 57225
rect 1239 57169 1307 57225
rect 1363 57169 1431 57225
rect 1487 57169 1555 57225
rect 1611 57169 1679 57225
rect 1735 57169 1803 57225
rect 1859 57169 1927 57225
rect 1983 57169 2051 57225
rect 2107 57169 2117 57225
rect 305 57101 2117 57169
rect 305 57045 315 57101
rect 371 57045 439 57101
rect 495 57045 563 57101
rect 619 57045 687 57101
rect 743 57045 811 57101
rect 867 57045 935 57101
rect 991 57045 1059 57101
rect 1115 57045 1183 57101
rect 1239 57045 1307 57101
rect 1363 57045 1431 57101
rect 1487 57045 1555 57101
rect 1611 57045 1679 57101
rect 1735 57045 1803 57101
rect 1859 57045 1927 57101
rect 1983 57045 2051 57101
rect 2107 57045 2117 57101
rect 305 56977 2117 57045
rect 305 56921 315 56977
rect 371 56921 439 56977
rect 495 56921 563 56977
rect 619 56921 687 56977
rect 743 56921 811 56977
rect 867 56921 935 56977
rect 991 56921 1059 56977
rect 1115 56921 1183 56977
rect 1239 56921 1307 56977
rect 1363 56921 1431 56977
rect 1487 56921 1555 56977
rect 1611 56921 1679 56977
rect 1735 56921 1803 56977
rect 1859 56921 1927 56977
rect 1983 56921 2051 56977
rect 2107 56921 2117 56977
rect 305 56853 2117 56921
rect 305 56797 315 56853
rect 371 56797 439 56853
rect 495 56797 563 56853
rect 619 56797 687 56853
rect 743 56797 811 56853
rect 867 56797 935 56853
rect 991 56797 1059 56853
rect 1115 56797 1183 56853
rect 1239 56797 1307 56853
rect 1363 56797 1431 56853
rect 1487 56797 1555 56853
rect 1611 56797 1679 56853
rect 1735 56797 1803 56853
rect 1859 56797 1927 56853
rect 1983 56797 2051 56853
rect 2107 56797 2117 56853
rect 305 56729 2117 56797
rect 305 56673 315 56729
rect 371 56673 439 56729
rect 495 56673 563 56729
rect 619 56673 687 56729
rect 743 56673 811 56729
rect 867 56673 935 56729
rect 991 56673 1059 56729
rect 1115 56673 1183 56729
rect 1239 56673 1307 56729
rect 1363 56673 1431 56729
rect 1487 56673 1555 56729
rect 1611 56673 1679 56729
rect 1735 56673 1803 56729
rect 1859 56673 1927 56729
rect 1983 56673 2051 56729
rect 2107 56673 2117 56729
rect 305 56605 2117 56673
rect 305 56549 315 56605
rect 371 56549 439 56605
rect 495 56549 563 56605
rect 619 56549 687 56605
rect 743 56549 811 56605
rect 867 56549 935 56605
rect 991 56549 1059 56605
rect 1115 56549 1183 56605
rect 1239 56549 1307 56605
rect 1363 56549 1431 56605
rect 1487 56549 1555 56605
rect 1611 56549 1679 56605
rect 1735 56549 1803 56605
rect 1859 56549 1927 56605
rect 1983 56549 2051 56605
rect 2107 56549 2117 56605
rect 305 56481 2117 56549
rect 305 56425 315 56481
rect 371 56425 439 56481
rect 495 56425 563 56481
rect 619 56425 687 56481
rect 743 56425 811 56481
rect 867 56425 935 56481
rect 991 56425 1059 56481
rect 1115 56425 1183 56481
rect 1239 56425 1307 56481
rect 1363 56425 1431 56481
rect 1487 56425 1555 56481
rect 1611 56425 1679 56481
rect 1735 56425 1803 56481
rect 1859 56425 1927 56481
rect 1983 56425 2051 56481
rect 2107 56425 2117 56481
rect 305 56357 2117 56425
rect 305 56301 315 56357
rect 371 56301 439 56357
rect 495 56301 563 56357
rect 619 56301 687 56357
rect 743 56301 811 56357
rect 867 56301 935 56357
rect 991 56301 1059 56357
rect 1115 56301 1183 56357
rect 1239 56301 1307 56357
rect 1363 56301 1431 56357
rect 1487 56301 1555 56357
rect 1611 56301 1679 56357
rect 1735 56301 1803 56357
rect 1859 56301 1927 56357
rect 1983 56301 2051 56357
rect 2107 56301 2117 56357
rect 305 56233 2117 56301
rect 305 56177 315 56233
rect 371 56177 439 56233
rect 495 56177 563 56233
rect 619 56177 687 56233
rect 743 56177 811 56233
rect 867 56177 935 56233
rect 991 56177 1059 56233
rect 1115 56177 1183 56233
rect 1239 56177 1307 56233
rect 1363 56177 1431 56233
rect 1487 56177 1555 56233
rect 1611 56177 1679 56233
rect 1735 56177 1803 56233
rect 1859 56177 1927 56233
rect 1983 56177 2051 56233
rect 2107 56177 2117 56233
rect 305 56109 2117 56177
rect 305 56053 315 56109
rect 371 56053 439 56109
rect 495 56053 563 56109
rect 619 56053 687 56109
rect 743 56053 811 56109
rect 867 56053 935 56109
rect 991 56053 1059 56109
rect 1115 56053 1183 56109
rect 1239 56053 1307 56109
rect 1363 56053 1431 56109
rect 1487 56053 1555 56109
rect 1611 56053 1679 56109
rect 1735 56053 1803 56109
rect 1859 56053 1927 56109
rect 1983 56053 2051 56109
rect 2107 56053 2117 56109
rect 305 56043 2117 56053
rect 2798 57225 4734 57235
rect 2798 57169 2808 57225
rect 2864 57169 2932 57225
rect 2988 57169 3056 57225
rect 3112 57169 3180 57225
rect 3236 57169 3304 57225
rect 3360 57169 3428 57225
rect 3484 57169 3552 57225
rect 3608 57169 3676 57225
rect 3732 57169 3800 57225
rect 3856 57169 3924 57225
rect 3980 57169 4048 57225
rect 4104 57169 4172 57225
rect 4228 57169 4296 57225
rect 4352 57169 4420 57225
rect 4476 57169 4544 57225
rect 4600 57169 4668 57225
rect 4724 57169 4734 57225
rect 2798 57101 4734 57169
rect 2798 57045 2808 57101
rect 2864 57045 2932 57101
rect 2988 57045 3056 57101
rect 3112 57045 3180 57101
rect 3236 57045 3304 57101
rect 3360 57045 3428 57101
rect 3484 57045 3552 57101
rect 3608 57045 3676 57101
rect 3732 57045 3800 57101
rect 3856 57045 3924 57101
rect 3980 57045 4048 57101
rect 4104 57045 4172 57101
rect 4228 57045 4296 57101
rect 4352 57045 4420 57101
rect 4476 57045 4544 57101
rect 4600 57045 4668 57101
rect 4724 57045 4734 57101
rect 2798 56977 4734 57045
rect 2798 56921 2808 56977
rect 2864 56921 2932 56977
rect 2988 56921 3056 56977
rect 3112 56921 3180 56977
rect 3236 56921 3304 56977
rect 3360 56921 3428 56977
rect 3484 56921 3552 56977
rect 3608 56921 3676 56977
rect 3732 56921 3800 56977
rect 3856 56921 3924 56977
rect 3980 56921 4048 56977
rect 4104 56921 4172 56977
rect 4228 56921 4296 56977
rect 4352 56921 4420 56977
rect 4476 56921 4544 56977
rect 4600 56921 4668 56977
rect 4724 56921 4734 56977
rect 2798 56853 4734 56921
rect 2798 56797 2808 56853
rect 2864 56797 2932 56853
rect 2988 56797 3056 56853
rect 3112 56797 3180 56853
rect 3236 56797 3304 56853
rect 3360 56797 3428 56853
rect 3484 56797 3552 56853
rect 3608 56797 3676 56853
rect 3732 56797 3800 56853
rect 3856 56797 3924 56853
rect 3980 56797 4048 56853
rect 4104 56797 4172 56853
rect 4228 56797 4296 56853
rect 4352 56797 4420 56853
rect 4476 56797 4544 56853
rect 4600 56797 4668 56853
rect 4724 56797 4734 56853
rect 2798 56729 4734 56797
rect 2798 56673 2808 56729
rect 2864 56673 2932 56729
rect 2988 56673 3056 56729
rect 3112 56673 3180 56729
rect 3236 56673 3304 56729
rect 3360 56673 3428 56729
rect 3484 56673 3552 56729
rect 3608 56673 3676 56729
rect 3732 56673 3800 56729
rect 3856 56673 3924 56729
rect 3980 56673 4048 56729
rect 4104 56673 4172 56729
rect 4228 56673 4296 56729
rect 4352 56673 4420 56729
rect 4476 56673 4544 56729
rect 4600 56673 4668 56729
rect 4724 56673 4734 56729
rect 2798 56605 4734 56673
rect 2798 56549 2808 56605
rect 2864 56549 2932 56605
rect 2988 56549 3056 56605
rect 3112 56549 3180 56605
rect 3236 56549 3304 56605
rect 3360 56549 3428 56605
rect 3484 56549 3552 56605
rect 3608 56549 3676 56605
rect 3732 56549 3800 56605
rect 3856 56549 3924 56605
rect 3980 56549 4048 56605
rect 4104 56549 4172 56605
rect 4228 56549 4296 56605
rect 4352 56549 4420 56605
rect 4476 56549 4544 56605
rect 4600 56549 4668 56605
rect 4724 56549 4734 56605
rect 2798 56481 4734 56549
rect 2798 56425 2808 56481
rect 2864 56425 2932 56481
rect 2988 56425 3056 56481
rect 3112 56425 3180 56481
rect 3236 56425 3304 56481
rect 3360 56425 3428 56481
rect 3484 56425 3552 56481
rect 3608 56425 3676 56481
rect 3732 56425 3800 56481
rect 3856 56425 3924 56481
rect 3980 56425 4048 56481
rect 4104 56425 4172 56481
rect 4228 56425 4296 56481
rect 4352 56425 4420 56481
rect 4476 56425 4544 56481
rect 4600 56425 4668 56481
rect 4724 56425 4734 56481
rect 2798 56357 4734 56425
rect 2798 56301 2808 56357
rect 2864 56301 2932 56357
rect 2988 56301 3056 56357
rect 3112 56301 3180 56357
rect 3236 56301 3304 56357
rect 3360 56301 3428 56357
rect 3484 56301 3552 56357
rect 3608 56301 3676 56357
rect 3732 56301 3800 56357
rect 3856 56301 3924 56357
rect 3980 56301 4048 56357
rect 4104 56301 4172 56357
rect 4228 56301 4296 56357
rect 4352 56301 4420 56357
rect 4476 56301 4544 56357
rect 4600 56301 4668 56357
rect 4724 56301 4734 56357
rect 2798 56233 4734 56301
rect 2798 56177 2808 56233
rect 2864 56177 2932 56233
rect 2988 56177 3056 56233
rect 3112 56177 3180 56233
rect 3236 56177 3304 56233
rect 3360 56177 3428 56233
rect 3484 56177 3552 56233
rect 3608 56177 3676 56233
rect 3732 56177 3800 56233
rect 3856 56177 3924 56233
rect 3980 56177 4048 56233
rect 4104 56177 4172 56233
rect 4228 56177 4296 56233
rect 4352 56177 4420 56233
rect 4476 56177 4544 56233
rect 4600 56177 4668 56233
rect 4724 56177 4734 56233
rect 2798 56109 4734 56177
rect 2798 56053 2808 56109
rect 2864 56053 2932 56109
rect 2988 56053 3056 56109
rect 3112 56053 3180 56109
rect 3236 56053 3304 56109
rect 3360 56053 3428 56109
rect 3484 56053 3552 56109
rect 3608 56053 3676 56109
rect 3732 56053 3800 56109
rect 3856 56053 3924 56109
rect 3980 56053 4048 56109
rect 4104 56053 4172 56109
rect 4228 56053 4296 56109
rect 4352 56053 4420 56109
rect 4476 56053 4544 56109
rect 4600 56053 4668 56109
rect 4724 56053 4734 56109
rect 2798 56043 4734 56053
rect 5168 57225 7104 57235
rect 5168 57169 5178 57225
rect 5234 57169 5302 57225
rect 5358 57169 5426 57225
rect 5482 57169 5550 57225
rect 5606 57169 5674 57225
rect 5730 57169 5798 57225
rect 5854 57169 5922 57225
rect 5978 57169 6046 57225
rect 6102 57169 6170 57225
rect 6226 57169 6294 57225
rect 6350 57169 6418 57225
rect 6474 57169 6542 57225
rect 6598 57169 6666 57225
rect 6722 57169 6790 57225
rect 6846 57169 6914 57225
rect 6970 57169 7038 57225
rect 7094 57169 7104 57225
rect 5168 57101 7104 57169
rect 5168 57045 5178 57101
rect 5234 57045 5302 57101
rect 5358 57045 5426 57101
rect 5482 57045 5550 57101
rect 5606 57045 5674 57101
rect 5730 57045 5798 57101
rect 5854 57045 5922 57101
rect 5978 57045 6046 57101
rect 6102 57045 6170 57101
rect 6226 57045 6294 57101
rect 6350 57045 6418 57101
rect 6474 57045 6542 57101
rect 6598 57045 6666 57101
rect 6722 57045 6790 57101
rect 6846 57045 6914 57101
rect 6970 57045 7038 57101
rect 7094 57045 7104 57101
rect 5168 56977 7104 57045
rect 5168 56921 5178 56977
rect 5234 56921 5302 56977
rect 5358 56921 5426 56977
rect 5482 56921 5550 56977
rect 5606 56921 5674 56977
rect 5730 56921 5798 56977
rect 5854 56921 5922 56977
rect 5978 56921 6046 56977
rect 6102 56921 6170 56977
rect 6226 56921 6294 56977
rect 6350 56921 6418 56977
rect 6474 56921 6542 56977
rect 6598 56921 6666 56977
rect 6722 56921 6790 56977
rect 6846 56921 6914 56977
rect 6970 56921 7038 56977
rect 7094 56921 7104 56977
rect 5168 56853 7104 56921
rect 5168 56797 5178 56853
rect 5234 56797 5302 56853
rect 5358 56797 5426 56853
rect 5482 56797 5550 56853
rect 5606 56797 5674 56853
rect 5730 56797 5798 56853
rect 5854 56797 5922 56853
rect 5978 56797 6046 56853
rect 6102 56797 6170 56853
rect 6226 56797 6294 56853
rect 6350 56797 6418 56853
rect 6474 56797 6542 56853
rect 6598 56797 6666 56853
rect 6722 56797 6790 56853
rect 6846 56797 6914 56853
rect 6970 56797 7038 56853
rect 7094 56797 7104 56853
rect 5168 56729 7104 56797
rect 5168 56673 5178 56729
rect 5234 56673 5302 56729
rect 5358 56673 5426 56729
rect 5482 56673 5550 56729
rect 5606 56673 5674 56729
rect 5730 56673 5798 56729
rect 5854 56673 5922 56729
rect 5978 56673 6046 56729
rect 6102 56673 6170 56729
rect 6226 56673 6294 56729
rect 6350 56673 6418 56729
rect 6474 56673 6542 56729
rect 6598 56673 6666 56729
rect 6722 56673 6790 56729
rect 6846 56673 6914 56729
rect 6970 56673 7038 56729
rect 7094 56673 7104 56729
rect 5168 56605 7104 56673
rect 5168 56549 5178 56605
rect 5234 56549 5302 56605
rect 5358 56549 5426 56605
rect 5482 56549 5550 56605
rect 5606 56549 5674 56605
rect 5730 56549 5798 56605
rect 5854 56549 5922 56605
rect 5978 56549 6046 56605
rect 6102 56549 6170 56605
rect 6226 56549 6294 56605
rect 6350 56549 6418 56605
rect 6474 56549 6542 56605
rect 6598 56549 6666 56605
rect 6722 56549 6790 56605
rect 6846 56549 6914 56605
rect 6970 56549 7038 56605
rect 7094 56549 7104 56605
rect 5168 56481 7104 56549
rect 5168 56425 5178 56481
rect 5234 56425 5302 56481
rect 5358 56425 5426 56481
rect 5482 56425 5550 56481
rect 5606 56425 5674 56481
rect 5730 56425 5798 56481
rect 5854 56425 5922 56481
rect 5978 56425 6046 56481
rect 6102 56425 6170 56481
rect 6226 56425 6294 56481
rect 6350 56425 6418 56481
rect 6474 56425 6542 56481
rect 6598 56425 6666 56481
rect 6722 56425 6790 56481
rect 6846 56425 6914 56481
rect 6970 56425 7038 56481
rect 7094 56425 7104 56481
rect 5168 56357 7104 56425
rect 5168 56301 5178 56357
rect 5234 56301 5302 56357
rect 5358 56301 5426 56357
rect 5482 56301 5550 56357
rect 5606 56301 5674 56357
rect 5730 56301 5798 56357
rect 5854 56301 5922 56357
rect 5978 56301 6046 56357
rect 6102 56301 6170 56357
rect 6226 56301 6294 56357
rect 6350 56301 6418 56357
rect 6474 56301 6542 56357
rect 6598 56301 6666 56357
rect 6722 56301 6790 56357
rect 6846 56301 6914 56357
rect 6970 56301 7038 56357
rect 7094 56301 7104 56357
rect 5168 56233 7104 56301
rect 5168 56177 5178 56233
rect 5234 56177 5302 56233
rect 5358 56177 5426 56233
rect 5482 56177 5550 56233
rect 5606 56177 5674 56233
rect 5730 56177 5798 56233
rect 5854 56177 5922 56233
rect 5978 56177 6046 56233
rect 6102 56177 6170 56233
rect 6226 56177 6294 56233
rect 6350 56177 6418 56233
rect 6474 56177 6542 56233
rect 6598 56177 6666 56233
rect 6722 56177 6790 56233
rect 6846 56177 6914 56233
rect 6970 56177 7038 56233
rect 7094 56177 7104 56233
rect 5168 56109 7104 56177
rect 5168 56053 5178 56109
rect 5234 56053 5302 56109
rect 5358 56053 5426 56109
rect 5482 56053 5550 56109
rect 5606 56053 5674 56109
rect 5730 56053 5798 56109
rect 5854 56053 5922 56109
rect 5978 56053 6046 56109
rect 6102 56053 6170 56109
rect 6226 56053 6294 56109
rect 6350 56053 6418 56109
rect 6474 56053 6542 56109
rect 6598 56053 6666 56109
rect 6722 56053 6790 56109
rect 6846 56053 6914 56109
rect 6970 56053 7038 56109
rect 7094 56053 7104 56109
rect 5168 56043 7104 56053
rect 7874 57225 9810 57235
rect 7874 57169 7884 57225
rect 7940 57169 8008 57225
rect 8064 57169 8132 57225
rect 8188 57169 8256 57225
rect 8312 57169 8380 57225
rect 8436 57169 8504 57225
rect 8560 57169 8628 57225
rect 8684 57169 8752 57225
rect 8808 57169 8876 57225
rect 8932 57169 9000 57225
rect 9056 57169 9124 57225
rect 9180 57169 9248 57225
rect 9304 57169 9372 57225
rect 9428 57169 9496 57225
rect 9552 57169 9620 57225
rect 9676 57169 9744 57225
rect 9800 57169 9810 57225
rect 7874 57101 9810 57169
rect 7874 57045 7884 57101
rect 7940 57045 8008 57101
rect 8064 57045 8132 57101
rect 8188 57045 8256 57101
rect 8312 57045 8380 57101
rect 8436 57045 8504 57101
rect 8560 57045 8628 57101
rect 8684 57045 8752 57101
rect 8808 57045 8876 57101
rect 8932 57045 9000 57101
rect 9056 57045 9124 57101
rect 9180 57045 9248 57101
rect 9304 57045 9372 57101
rect 9428 57045 9496 57101
rect 9552 57045 9620 57101
rect 9676 57045 9744 57101
rect 9800 57045 9810 57101
rect 7874 56977 9810 57045
rect 7874 56921 7884 56977
rect 7940 56921 8008 56977
rect 8064 56921 8132 56977
rect 8188 56921 8256 56977
rect 8312 56921 8380 56977
rect 8436 56921 8504 56977
rect 8560 56921 8628 56977
rect 8684 56921 8752 56977
rect 8808 56921 8876 56977
rect 8932 56921 9000 56977
rect 9056 56921 9124 56977
rect 9180 56921 9248 56977
rect 9304 56921 9372 56977
rect 9428 56921 9496 56977
rect 9552 56921 9620 56977
rect 9676 56921 9744 56977
rect 9800 56921 9810 56977
rect 7874 56853 9810 56921
rect 7874 56797 7884 56853
rect 7940 56797 8008 56853
rect 8064 56797 8132 56853
rect 8188 56797 8256 56853
rect 8312 56797 8380 56853
rect 8436 56797 8504 56853
rect 8560 56797 8628 56853
rect 8684 56797 8752 56853
rect 8808 56797 8876 56853
rect 8932 56797 9000 56853
rect 9056 56797 9124 56853
rect 9180 56797 9248 56853
rect 9304 56797 9372 56853
rect 9428 56797 9496 56853
rect 9552 56797 9620 56853
rect 9676 56797 9744 56853
rect 9800 56797 9810 56853
rect 7874 56729 9810 56797
rect 7874 56673 7884 56729
rect 7940 56673 8008 56729
rect 8064 56673 8132 56729
rect 8188 56673 8256 56729
rect 8312 56673 8380 56729
rect 8436 56673 8504 56729
rect 8560 56673 8628 56729
rect 8684 56673 8752 56729
rect 8808 56673 8876 56729
rect 8932 56673 9000 56729
rect 9056 56673 9124 56729
rect 9180 56673 9248 56729
rect 9304 56673 9372 56729
rect 9428 56673 9496 56729
rect 9552 56673 9620 56729
rect 9676 56673 9744 56729
rect 9800 56673 9810 56729
rect 7874 56605 9810 56673
rect 7874 56549 7884 56605
rect 7940 56549 8008 56605
rect 8064 56549 8132 56605
rect 8188 56549 8256 56605
rect 8312 56549 8380 56605
rect 8436 56549 8504 56605
rect 8560 56549 8628 56605
rect 8684 56549 8752 56605
rect 8808 56549 8876 56605
rect 8932 56549 9000 56605
rect 9056 56549 9124 56605
rect 9180 56549 9248 56605
rect 9304 56549 9372 56605
rect 9428 56549 9496 56605
rect 9552 56549 9620 56605
rect 9676 56549 9744 56605
rect 9800 56549 9810 56605
rect 7874 56481 9810 56549
rect 7874 56425 7884 56481
rect 7940 56425 8008 56481
rect 8064 56425 8132 56481
rect 8188 56425 8256 56481
rect 8312 56425 8380 56481
rect 8436 56425 8504 56481
rect 8560 56425 8628 56481
rect 8684 56425 8752 56481
rect 8808 56425 8876 56481
rect 8932 56425 9000 56481
rect 9056 56425 9124 56481
rect 9180 56425 9248 56481
rect 9304 56425 9372 56481
rect 9428 56425 9496 56481
rect 9552 56425 9620 56481
rect 9676 56425 9744 56481
rect 9800 56425 9810 56481
rect 7874 56357 9810 56425
rect 7874 56301 7884 56357
rect 7940 56301 8008 56357
rect 8064 56301 8132 56357
rect 8188 56301 8256 56357
rect 8312 56301 8380 56357
rect 8436 56301 8504 56357
rect 8560 56301 8628 56357
rect 8684 56301 8752 56357
rect 8808 56301 8876 56357
rect 8932 56301 9000 56357
rect 9056 56301 9124 56357
rect 9180 56301 9248 56357
rect 9304 56301 9372 56357
rect 9428 56301 9496 56357
rect 9552 56301 9620 56357
rect 9676 56301 9744 56357
rect 9800 56301 9810 56357
rect 7874 56233 9810 56301
rect 7874 56177 7884 56233
rect 7940 56177 8008 56233
rect 8064 56177 8132 56233
rect 8188 56177 8256 56233
rect 8312 56177 8380 56233
rect 8436 56177 8504 56233
rect 8560 56177 8628 56233
rect 8684 56177 8752 56233
rect 8808 56177 8876 56233
rect 8932 56177 9000 56233
rect 9056 56177 9124 56233
rect 9180 56177 9248 56233
rect 9304 56177 9372 56233
rect 9428 56177 9496 56233
rect 9552 56177 9620 56233
rect 9676 56177 9744 56233
rect 9800 56177 9810 56233
rect 7874 56109 9810 56177
rect 7874 56053 7884 56109
rect 7940 56053 8008 56109
rect 8064 56053 8132 56109
rect 8188 56053 8256 56109
rect 8312 56053 8380 56109
rect 8436 56053 8504 56109
rect 8560 56053 8628 56109
rect 8684 56053 8752 56109
rect 8808 56053 8876 56109
rect 8932 56053 9000 56109
rect 9056 56053 9124 56109
rect 9180 56053 9248 56109
rect 9304 56053 9372 56109
rect 9428 56053 9496 56109
rect 9552 56053 9620 56109
rect 9676 56053 9744 56109
rect 9800 56053 9810 56109
rect 7874 56043 9810 56053
rect 10244 57225 12180 57235
rect 10244 57169 10254 57225
rect 10310 57169 10378 57225
rect 10434 57169 10502 57225
rect 10558 57169 10626 57225
rect 10682 57169 10750 57225
rect 10806 57169 10874 57225
rect 10930 57169 10998 57225
rect 11054 57169 11122 57225
rect 11178 57169 11246 57225
rect 11302 57169 11370 57225
rect 11426 57169 11494 57225
rect 11550 57169 11618 57225
rect 11674 57169 11742 57225
rect 11798 57169 11866 57225
rect 11922 57169 11990 57225
rect 12046 57169 12114 57225
rect 12170 57169 12180 57225
rect 10244 57101 12180 57169
rect 10244 57045 10254 57101
rect 10310 57045 10378 57101
rect 10434 57045 10502 57101
rect 10558 57045 10626 57101
rect 10682 57045 10750 57101
rect 10806 57045 10874 57101
rect 10930 57045 10998 57101
rect 11054 57045 11122 57101
rect 11178 57045 11246 57101
rect 11302 57045 11370 57101
rect 11426 57045 11494 57101
rect 11550 57045 11618 57101
rect 11674 57045 11742 57101
rect 11798 57045 11866 57101
rect 11922 57045 11990 57101
rect 12046 57045 12114 57101
rect 12170 57045 12180 57101
rect 10244 56977 12180 57045
rect 10244 56921 10254 56977
rect 10310 56921 10378 56977
rect 10434 56921 10502 56977
rect 10558 56921 10626 56977
rect 10682 56921 10750 56977
rect 10806 56921 10874 56977
rect 10930 56921 10998 56977
rect 11054 56921 11122 56977
rect 11178 56921 11246 56977
rect 11302 56921 11370 56977
rect 11426 56921 11494 56977
rect 11550 56921 11618 56977
rect 11674 56921 11742 56977
rect 11798 56921 11866 56977
rect 11922 56921 11990 56977
rect 12046 56921 12114 56977
rect 12170 56921 12180 56977
rect 10244 56853 12180 56921
rect 10244 56797 10254 56853
rect 10310 56797 10378 56853
rect 10434 56797 10502 56853
rect 10558 56797 10626 56853
rect 10682 56797 10750 56853
rect 10806 56797 10874 56853
rect 10930 56797 10998 56853
rect 11054 56797 11122 56853
rect 11178 56797 11246 56853
rect 11302 56797 11370 56853
rect 11426 56797 11494 56853
rect 11550 56797 11618 56853
rect 11674 56797 11742 56853
rect 11798 56797 11866 56853
rect 11922 56797 11990 56853
rect 12046 56797 12114 56853
rect 12170 56797 12180 56853
rect 10244 56729 12180 56797
rect 10244 56673 10254 56729
rect 10310 56673 10378 56729
rect 10434 56673 10502 56729
rect 10558 56673 10626 56729
rect 10682 56673 10750 56729
rect 10806 56673 10874 56729
rect 10930 56673 10998 56729
rect 11054 56673 11122 56729
rect 11178 56673 11246 56729
rect 11302 56673 11370 56729
rect 11426 56673 11494 56729
rect 11550 56673 11618 56729
rect 11674 56673 11742 56729
rect 11798 56673 11866 56729
rect 11922 56673 11990 56729
rect 12046 56673 12114 56729
rect 12170 56673 12180 56729
rect 10244 56605 12180 56673
rect 10244 56549 10254 56605
rect 10310 56549 10378 56605
rect 10434 56549 10502 56605
rect 10558 56549 10626 56605
rect 10682 56549 10750 56605
rect 10806 56549 10874 56605
rect 10930 56549 10998 56605
rect 11054 56549 11122 56605
rect 11178 56549 11246 56605
rect 11302 56549 11370 56605
rect 11426 56549 11494 56605
rect 11550 56549 11618 56605
rect 11674 56549 11742 56605
rect 11798 56549 11866 56605
rect 11922 56549 11990 56605
rect 12046 56549 12114 56605
rect 12170 56549 12180 56605
rect 10244 56481 12180 56549
rect 10244 56425 10254 56481
rect 10310 56425 10378 56481
rect 10434 56425 10502 56481
rect 10558 56425 10626 56481
rect 10682 56425 10750 56481
rect 10806 56425 10874 56481
rect 10930 56425 10998 56481
rect 11054 56425 11122 56481
rect 11178 56425 11246 56481
rect 11302 56425 11370 56481
rect 11426 56425 11494 56481
rect 11550 56425 11618 56481
rect 11674 56425 11742 56481
rect 11798 56425 11866 56481
rect 11922 56425 11990 56481
rect 12046 56425 12114 56481
rect 12170 56425 12180 56481
rect 10244 56357 12180 56425
rect 10244 56301 10254 56357
rect 10310 56301 10378 56357
rect 10434 56301 10502 56357
rect 10558 56301 10626 56357
rect 10682 56301 10750 56357
rect 10806 56301 10874 56357
rect 10930 56301 10998 56357
rect 11054 56301 11122 56357
rect 11178 56301 11246 56357
rect 11302 56301 11370 56357
rect 11426 56301 11494 56357
rect 11550 56301 11618 56357
rect 11674 56301 11742 56357
rect 11798 56301 11866 56357
rect 11922 56301 11990 56357
rect 12046 56301 12114 56357
rect 12170 56301 12180 56357
rect 10244 56233 12180 56301
rect 10244 56177 10254 56233
rect 10310 56177 10378 56233
rect 10434 56177 10502 56233
rect 10558 56177 10626 56233
rect 10682 56177 10750 56233
rect 10806 56177 10874 56233
rect 10930 56177 10998 56233
rect 11054 56177 11122 56233
rect 11178 56177 11246 56233
rect 11302 56177 11370 56233
rect 11426 56177 11494 56233
rect 11550 56177 11618 56233
rect 11674 56177 11742 56233
rect 11798 56177 11866 56233
rect 11922 56177 11990 56233
rect 12046 56177 12114 56233
rect 12170 56177 12180 56233
rect 10244 56109 12180 56177
rect 10244 56053 10254 56109
rect 10310 56053 10378 56109
rect 10434 56053 10502 56109
rect 10558 56053 10626 56109
rect 10682 56053 10750 56109
rect 10806 56053 10874 56109
rect 10930 56053 10998 56109
rect 11054 56053 11122 56109
rect 11178 56053 11246 56109
rect 11302 56053 11370 56109
rect 11426 56053 11494 56109
rect 11550 56053 11618 56109
rect 11674 56053 11742 56109
rect 11798 56053 11866 56109
rect 11922 56053 11990 56109
rect 12046 56053 12114 56109
rect 12170 56053 12180 56109
rect 10244 56043 12180 56053
rect 12861 57225 14673 57235
rect 12861 57169 12871 57225
rect 12927 57169 12995 57225
rect 13051 57169 13119 57225
rect 13175 57169 13243 57225
rect 13299 57169 13367 57225
rect 13423 57169 13491 57225
rect 13547 57169 13615 57225
rect 13671 57169 13739 57225
rect 13795 57169 13863 57225
rect 13919 57169 13987 57225
rect 14043 57169 14111 57225
rect 14167 57169 14235 57225
rect 14291 57169 14359 57225
rect 14415 57169 14483 57225
rect 14539 57169 14607 57225
rect 14663 57169 14673 57225
rect 12861 57101 14673 57169
rect 12861 57045 12871 57101
rect 12927 57045 12995 57101
rect 13051 57045 13119 57101
rect 13175 57045 13243 57101
rect 13299 57045 13367 57101
rect 13423 57045 13491 57101
rect 13547 57045 13615 57101
rect 13671 57045 13739 57101
rect 13795 57045 13863 57101
rect 13919 57045 13987 57101
rect 14043 57045 14111 57101
rect 14167 57045 14235 57101
rect 14291 57045 14359 57101
rect 14415 57045 14483 57101
rect 14539 57045 14607 57101
rect 14663 57045 14673 57101
rect 12861 56977 14673 57045
rect 12861 56921 12871 56977
rect 12927 56921 12995 56977
rect 13051 56921 13119 56977
rect 13175 56921 13243 56977
rect 13299 56921 13367 56977
rect 13423 56921 13491 56977
rect 13547 56921 13615 56977
rect 13671 56921 13739 56977
rect 13795 56921 13863 56977
rect 13919 56921 13987 56977
rect 14043 56921 14111 56977
rect 14167 56921 14235 56977
rect 14291 56921 14359 56977
rect 14415 56921 14483 56977
rect 14539 56921 14607 56977
rect 14663 56921 14673 56977
rect 12861 56853 14673 56921
rect 12861 56797 12871 56853
rect 12927 56797 12995 56853
rect 13051 56797 13119 56853
rect 13175 56797 13243 56853
rect 13299 56797 13367 56853
rect 13423 56797 13491 56853
rect 13547 56797 13615 56853
rect 13671 56797 13739 56853
rect 13795 56797 13863 56853
rect 13919 56797 13987 56853
rect 14043 56797 14111 56853
rect 14167 56797 14235 56853
rect 14291 56797 14359 56853
rect 14415 56797 14483 56853
rect 14539 56797 14607 56853
rect 14663 56797 14673 56853
rect 12861 56729 14673 56797
rect 12861 56673 12871 56729
rect 12927 56673 12995 56729
rect 13051 56673 13119 56729
rect 13175 56673 13243 56729
rect 13299 56673 13367 56729
rect 13423 56673 13491 56729
rect 13547 56673 13615 56729
rect 13671 56673 13739 56729
rect 13795 56673 13863 56729
rect 13919 56673 13987 56729
rect 14043 56673 14111 56729
rect 14167 56673 14235 56729
rect 14291 56673 14359 56729
rect 14415 56673 14483 56729
rect 14539 56673 14607 56729
rect 14663 56673 14673 56729
rect 12861 56605 14673 56673
rect 12861 56549 12871 56605
rect 12927 56549 12995 56605
rect 13051 56549 13119 56605
rect 13175 56549 13243 56605
rect 13299 56549 13367 56605
rect 13423 56549 13491 56605
rect 13547 56549 13615 56605
rect 13671 56549 13739 56605
rect 13795 56549 13863 56605
rect 13919 56549 13987 56605
rect 14043 56549 14111 56605
rect 14167 56549 14235 56605
rect 14291 56549 14359 56605
rect 14415 56549 14483 56605
rect 14539 56549 14607 56605
rect 14663 56549 14673 56605
rect 12861 56481 14673 56549
rect 12861 56425 12871 56481
rect 12927 56425 12995 56481
rect 13051 56425 13119 56481
rect 13175 56425 13243 56481
rect 13299 56425 13367 56481
rect 13423 56425 13491 56481
rect 13547 56425 13615 56481
rect 13671 56425 13739 56481
rect 13795 56425 13863 56481
rect 13919 56425 13987 56481
rect 14043 56425 14111 56481
rect 14167 56425 14235 56481
rect 14291 56425 14359 56481
rect 14415 56425 14483 56481
rect 14539 56425 14607 56481
rect 14663 56425 14673 56481
rect 12861 56357 14673 56425
rect 12861 56301 12871 56357
rect 12927 56301 12995 56357
rect 13051 56301 13119 56357
rect 13175 56301 13243 56357
rect 13299 56301 13367 56357
rect 13423 56301 13491 56357
rect 13547 56301 13615 56357
rect 13671 56301 13739 56357
rect 13795 56301 13863 56357
rect 13919 56301 13987 56357
rect 14043 56301 14111 56357
rect 14167 56301 14235 56357
rect 14291 56301 14359 56357
rect 14415 56301 14483 56357
rect 14539 56301 14607 56357
rect 14663 56301 14673 56357
rect 12861 56233 14673 56301
rect 12861 56177 12871 56233
rect 12927 56177 12995 56233
rect 13051 56177 13119 56233
rect 13175 56177 13243 56233
rect 13299 56177 13367 56233
rect 13423 56177 13491 56233
rect 13547 56177 13615 56233
rect 13671 56177 13739 56233
rect 13795 56177 13863 56233
rect 13919 56177 13987 56233
rect 14043 56177 14111 56233
rect 14167 56177 14235 56233
rect 14291 56177 14359 56233
rect 14415 56177 14483 56233
rect 14539 56177 14607 56233
rect 14663 56177 14673 56233
rect 12861 56109 14673 56177
rect 12861 56053 12871 56109
rect 12927 56053 12995 56109
rect 13051 56053 13119 56109
rect 13175 56053 13243 56109
rect 13299 56053 13367 56109
rect 13423 56053 13491 56109
rect 13547 56053 13615 56109
rect 13671 56053 13739 56109
rect 13795 56053 13863 56109
rect 13919 56053 13987 56109
rect 14043 56053 14111 56109
rect 14167 56053 14235 56109
rect 14291 56053 14359 56109
rect 14415 56053 14483 56109
rect 14539 56053 14607 56109
rect 14663 56053 14673 56109
rect 12861 56043 14673 56053
rect 10 56007 86 56017
rect 14892 56017 14902 57261
rect 14958 56017 14968 57261
rect 14892 56007 14968 56017
rect 2481 55748 2681 55758
rect 2481 55692 2491 55748
rect 2547 55692 2615 55748
rect 2671 55692 2681 55748
rect 2481 55624 2681 55692
rect 2481 55568 2491 55624
rect 2547 55568 2615 55624
rect 2671 55568 2681 55624
rect 2481 55500 2681 55568
rect 2481 55444 2491 55500
rect 2547 55444 2615 55500
rect 2671 55444 2681 55500
rect 2481 55376 2681 55444
rect 2481 55320 2491 55376
rect 2547 55320 2615 55376
rect 2671 55320 2681 55376
rect 2481 55252 2681 55320
rect 2481 55196 2491 55252
rect 2547 55196 2615 55252
rect 2671 55196 2681 55252
rect 2481 55128 2681 55196
rect 2481 55072 2491 55128
rect 2547 55072 2615 55128
rect 2671 55072 2681 55128
rect 2481 55004 2681 55072
rect 2481 54948 2491 55004
rect 2547 54948 2615 55004
rect 2671 54948 2681 55004
rect 2481 54880 2681 54948
rect 2481 54824 2491 54880
rect 2547 54824 2615 54880
rect 2671 54824 2681 54880
rect 2481 54756 2681 54824
rect 2481 54700 2491 54756
rect 2547 54700 2615 54756
rect 2671 54700 2681 54756
rect 2481 54632 2681 54700
rect 2481 54576 2491 54632
rect 2547 54576 2615 54632
rect 2671 54576 2681 54632
rect 2481 54508 2681 54576
rect 2481 54452 2491 54508
rect 2547 54452 2615 54508
rect 2671 54452 2681 54508
rect 2481 54442 2681 54452
rect 4851 55748 5051 55758
rect 4851 55692 4861 55748
rect 4917 55692 4985 55748
rect 5041 55692 5051 55748
rect 4851 55624 5051 55692
rect 4851 55568 4861 55624
rect 4917 55568 4985 55624
rect 5041 55568 5051 55624
rect 4851 55500 5051 55568
rect 4851 55444 4861 55500
rect 4917 55444 4985 55500
rect 5041 55444 5051 55500
rect 4851 55376 5051 55444
rect 4851 55320 4861 55376
rect 4917 55320 4985 55376
rect 5041 55320 5051 55376
rect 4851 55252 5051 55320
rect 4851 55196 4861 55252
rect 4917 55196 4985 55252
rect 5041 55196 5051 55252
rect 4851 55128 5051 55196
rect 4851 55072 4861 55128
rect 4917 55072 4985 55128
rect 5041 55072 5051 55128
rect 4851 55004 5051 55072
rect 4851 54948 4861 55004
rect 4917 54948 4985 55004
rect 5041 54948 5051 55004
rect 4851 54880 5051 54948
rect 4851 54824 4861 54880
rect 4917 54824 4985 54880
rect 5041 54824 5051 54880
rect 4851 54756 5051 54824
rect 4851 54700 4861 54756
rect 4917 54700 4985 54756
rect 5041 54700 5051 54756
rect 4851 54632 5051 54700
rect 4851 54576 4861 54632
rect 4917 54576 4985 54632
rect 5041 54576 5051 54632
rect 4851 54508 5051 54576
rect 4851 54452 4861 54508
rect 4917 54452 4985 54508
rect 5041 54452 5051 54508
rect 4851 54442 5051 54452
rect 7265 55748 7713 55758
rect 7265 55692 7275 55748
rect 7331 55692 7399 55748
rect 7455 55692 7523 55748
rect 7579 55692 7647 55748
rect 7703 55692 7713 55748
rect 7265 55624 7713 55692
rect 7265 55568 7275 55624
rect 7331 55568 7399 55624
rect 7455 55568 7523 55624
rect 7579 55568 7647 55624
rect 7703 55568 7713 55624
rect 7265 55500 7713 55568
rect 7265 55444 7275 55500
rect 7331 55444 7399 55500
rect 7455 55444 7523 55500
rect 7579 55444 7647 55500
rect 7703 55444 7713 55500
rect 7265 55376 7713 55444
rect 7265 55320 7275 55376
rect 7331 55320 7399 55376
rect 7455 55320 7523 55376
rect 7579 55320 7647 55376
rect 7703 55320 7713 55376
rect 7265 55252 7713 55320
rect 7265 55196 7275 55252
rect 7331 55196 7399 55252
rect 7455 55196 7523 55252
rect 7579 55196 7647 55252
rect 7703 55196 7713 55252
rect 7265 55128 7713 55196
rect 7265 55072 7275 55128
rect 7331 55072 7399 55128
rect 7455 55072 7523 55128
rect 7579 55072 7647 55128
rect 7703 55072 7713 55128
rect 7265 55004 7713 55072
rect 7265 54948 7275 55004
rect 7331 54948 7399 55004
rect 7455 54948 7523 55004
rect 7579 54948 7647 55004
rect 7703 54948 7713 55004
rect 7265 54880 7713 54948
rect 7265 54824 7275 54880
rect 7331 54824 7399 54880
rect 7455 54824 7523 54880
rect 7579 54824 7647 54880
rect 7703 54824 7713 54880
rect 7265 54756 7713 54824
rect 7265 54700 7275 54756
rect 7331 54700 7399 54756
rect 7455 54700 7523 54756
rect 7579 54700 7647 54756
rect 7703 54700 7713 54756
rect 7265 54632 7713 54700
rect 7265 54576 7275 54632
rect 7331 54576 7399 54632
rect 7455 54576 7523 54632
rect 7579 54576 7647 54632
rect 7703 54576 7713 54632
rect 7265 54508 7713 54576
rect 7265 54452 7275 54508
rect 7331 54452 7399 54508
rect 7455 54452 7523 54508
rect 7579 54452 7647 54508
rect 7703 54452 7713 54508
rect 7265 54442 7713 54452
rect 9927 55748 10127 55758
rect 9927 55692 9937 55748
rect 9993 55692 10061 55748
rect 10117 55692 10127 55748
rect 9927 55624 10127 55692
rect 9927 55568 9937 55624
rect 9993 55568 10061 55624
rect 10117 55568 10127 55624
rect 9927 55500 10127 55568
rect 9927 55444 9937 55500
rect 9993 55444 10061 55500
rect 10117 55444 10127 55500
rect 9927 55376 10127 55444
rect 9927 55320 9937 55376
rect 9993 55320 10061 55376
rect 10117 55320 10127 55376
rect 9927 55252 10127 55320
rect 9927 55196 9937 55252
rect 9993 55196 10061 55252
rect 10117 55196 10127 55252
rect 9927 55128 10127 55196
rect 9927 55072 9937 55128
rect 9993 55072 10061 55128
rect 10117 55072 10127 55128
rect 9927 55004 10127 55072
rect 9927 54948 9937 55004
rect 9993 54948 10061 55004
rect 10117 54948 10127 55004
rect 9927 54880 10127 54948
rect 9927 54824 9937 54880
rect 9993 54824 10061 54880
rect 10117 54824 10127 54880
rect 9927 54756 10127 54824
rect 9927 54700 9937 54756
rect 9993 54700 10061 54756
rect 10117 54700 10127 54756
rect 9927 54632 10127 54700
rect 9927 54576 9937 54632
rect 9993 54576 10061 54632
rect 10117 54576 10127 54632
rect 9927 54508 10127 54576
rect 9927 54452 9937 54508
rect 9993 54452 10061 54508
rect 10117 54452 10127 54508
rect 9927 54442 10127 54452
rect 12297 55748 12497 55758
rect 12297 55692 12307 55748
rect 12363 55692 12431 55748
rect 12487 55692 12497 55748
rect 12297 55624 12497 55692
rect 12297 55568 12307 55624
rect 12363 55568 12431 55624
rect 12487 55568 12497 55624
rect 12297 55500 12497 55568
rect 12297 55444 12307 55500
rect 12363 55444 12431 55500
rect 12487 55444 12497 55500
rect 12297 55376 12497 55444
rect 12297 55320 12307 55376
rect 12363 55320 12431 55376
rect 12487 55320 12497 55376
rect 12297 55252 12497 55320
rect 12297 55196 12307 55252
rect 12363 55196 12431 55252
rect 12487 55196 12497 55252
rect 12297 55128 12497 55196
rect 12297 55072 12307 55128
rect 12363 55072 12431 55128
rect 12487 55072 12497 55128
rect 12297 55004 12497 55072
rect 12297 54948 12307 55004
rect 12363 54948 12431 55004
rect 12487 54948 12497 55004
rect 12297 54880 12497 54948
rect 12297 54824 12307 54880
rect 12363 54824 12431 54880
rect 12487 54824 12497 54880
rect 12297 54756 12497 54824
rect 12297 54700 12307 54756
rect 12363 54700 12431 54756
rect 12487 54700 12497 54756
rect 12297 54632 12497 54700
rect 12297 54576 12307 54632
rect 12363 54576 12431 54632
rect 12487 54576 12497 54632
rect 12297 54508 12497 54576
rect 12297 54452 12307 54508
rect 12363 54452 12431 54508
rect 12487 54452 12497 54508
rect 12297 54442 12497 54452
rect 10 54176 86 54186
rect 10 52824 20 54176
rect 76 52824 86 54176
rect 14892 54176 14968 54186
rect 305 54148 2117 54158
rect 305 54092 315 54148
rect 371 54092 439 54148
rect 495 54092 563 54148
rect 619 54092 687 54148
rect 743 54092 811 54148
rect 867 54092 935 54148
rect 991 54092 1059 54148
rect 1115 54092 1183 54148
rect 1239 54092 1307 54148
rect 1363 54092 1431 54148
rect 1487 54092 1555 54148
rect 1611 54092 1679 54148
rect 1735 54092 1803 54148
rect 1859 54092 1927 54148
rect 1983 54092 2051 54148
rect 2107 54092 2117 54148
rect 305 54024 2117 54092
rect 305 53968 315 54024
rect 371 53968 439 54024
rect 495 53968 563 54024
rect 619 53968 687 54024
rect 743 53968 811 54024
rect 867 53968 935 54024
rect 991 53968 1059 54024
rect 1115 53968 1183 54024
rect 1239 53968 1307 54024
rect 1363 53968 1431 54024
rect 1487 53968 1555 54024
rect 1611 53968 1679 54024
rect 1735 53968 1803 54024
rect 1859 53968 1927 54024
rect 1983 53968 2051 54024
rect 2107 53968 2117 54024
rect 305 53900 2117 53968
rect 305 53844 315 53900
rect 371 53844 439 53900
rect 495 53844 563 53900
rect 619 53844 687 53900
rect 743 53844 811 53900
rect 867 53844 935 53900
rect 991 53844 1059 53900
rect 1115 53844 1183 53900
rect 1239 53844 1307 53900
rect 1363 53844 1431 53900
rect 1487 53844 1555 53900
rect 1611 53844 1679 53900
rect 1735 53844 1803 53900
rect 1859 53844 1927 53900
rect 1983 53844 2051 53900
rect 2107 53844 2117 53900
rect 305 53776 2117 53844
rect 305 53720 315 53776
rect 371 53720 439 53776
rect 495 53720 563 53776
rect 619 53720 687 53776
rect 743 53720 811 53776
rect 867 53720 935 53776
rect 991 53720 1059 53776
rect 1115 53720 1183 53776
rect 1239 53720 1307 53776
rect 1363 53720 1431 53776
rect 1487 53720 1555 53776
rect 1611 53720 1679 53776
rect 1735 53720 1803 53776
rect 1859 53720 1927 53776
rect 1983 53720 2051 53776
rect 2107 53720 2117 53776
rect 305 53652 2117 53720
rect 305 53596 315 53652
rect 371 53596 439 53652
rect 495 53596 563 53652
rect 619 53596 687 53652
rect 743 53596 811 53652
rect 867 53596 935 53652
rect 991 53596 1059 53652
rect 1115 53596 1183 53652
rect 1239 53596 1307 53652
rect 1363 53596 1431 53652
rect 1487 53596 1555 53652
rect 1611 53596 1679 53652
rect 1735 53596 1803 53652
rect 1859 53596 1927 53652
rect 1983 53596 2051 53652
rect 2107 53596 2117 53652
rect 305 53528 2117 53596
rect 305 53472 315 53528
rect 371 53472 439 53528
rect 495 53472 563 53528
rect 619 53472 687 53528
rect 743 53472 811 53528
rect 867 53472 935 53528
rect 991 53472 1059 53528
rect 1115 53472 1183 53528
rect 1239 53472 1307 53528
rect 1363 53472 1431 53528
rect 1487 53472 1555 53528
rect 1611 53472 1679 53528
rect 1735 53472 1803 53528
rect 1859 53472 1927 53528
rect 1983 53472 2051 53528
rect 2107 53472 2117 53528
rect 305 53404 2117 53472
rect 305 53348 315 53404
rect 371 53348 439 53404
rect 495 53348 563 53404
rect 619 53348 687 53404
rect 743 53348 811 53404
rect 867 53348 935 53404
rect 991 53348 1059 53404
rect 1115 53348 1183 53404
rect 1239 53348 1307 53404
rect 1363 53348 1431 53404
rect 1487 53348 1555 53404
rect 1611 53348 1679 53404
rect 1735 53348 1803 53404
rect 1859 53348 1927 53404
rect 1983 53348 2051 53404
rect 2107 53348 2117 53404
rect 305 53280 2117 53348
rect 305 53224 315 53280
rect 371 53224 439 53280
rect 495 53224 563 53280
rect 619 53224 687 53280
rect 743 53224 811 53280
rect 867 53224 935 53280
rect 991 53224 1059 53280
rect 1115 53224 1183 53280
rect 1239 53224 1307 53280
rect 1363 53224 1431 53280
rect 1487 53224 1555 53280
rect 1611 53224 1679 53280
rect 1735 53224 1803 53280
rect 1859 53224 1927 53280
rect 1983 53224 2051 53280
rect 2107 53224 2117 53280
rect 305 53156 2117 53224
rect 305 53100 315 53156
rect 371 53100 439 53156
rect 495 53100 563 53156
rect 619 53100 687 53156
rect 743 53100 811 53156
rect 867 53100 935 53156
rect 991 53100 1059 53156
rect 1115 53100 1183 53156
rect 1239 53100 1307 53156
rect 1363 53100 1431 53156
rect 1487 53100 1555 53156
rect 1611 53100 1679 53156
rect 1735 53100 1803 53156
rect 1859 53100 1927 53156
rect 1983 53100 2051 53156
rect 2107 53100 2117 53156
rect 305 53032 2117 53100
rect 305 52976 315 53032
rect 371 52976 439 53032
rect 495 52976 563 53032
rect 619 52976 687 53032
rect 743 52976 811 53032
rect 867 52976 935 53032
rect 991 52976 1059 53032
rect 1115 52976 1183 53032
rect 1239 52976 1307 53032
rect 1363 52976 1431 53032
rect 1487 52976 1555 53032
rect 1611 52976 1679 53032
rect 1735 52976 1803 53032
rect 1859 52976 1927 53032
rect 1983 52976 2051 53032
rect 2107 52976 2117 53032
rect 305 52908 2117 52976
rect 305 52852 315 52908
rect 371 52852 439 52908
rect 495 52852 563 52908
rect 619 52852 687 52908
rect 743 52852 811 52908
rect 867 52852 935 52908
rect 991 52852 1059 52908
rect 1115 52852 1183 52908
rect 1239 52852 1307 52908
rect 1363 52852 1431 52908
rect 1487 52852 1555 52908
rect 1611 52852 1679 52908
rect 1735 52852 1803 52908
rect 1859 52852 1927 52908
rect 1983 52852 2051 52908
rect 2107 52852 2117 52908
rect 305 52842 2117 52852
rect 2798 54148 4734 54158
rect 2798 54092 2808 54148
rect 2864 54092 2932 54148
rect 2988 54092 3056 54148
rect 3112 54092 3180 54148
rect 3236 54092 3304 54148
rect 3360 54092 3428 54148
rect 3484 54092 3552 54148
rect 3608 54092 3676 54148
rect 3732 54092 3800 54148
rect 3856 54092 3924 54148
rect 3980 54092 4048 54148
rect 4104 54092 4172 54148
rect 4228 54092 4296 54148
rect 4352 54092 4420 54148
rect 4476 54092 4544 54148
rect 4600 54092 4668 54148
rect 4724 54092 4734 54148
rect 2798 54024 4734 54092
rect 2798 53968 2808 54024
rect 2864 53968 2932 54024
rect 2988 53968 3056 54024
rect 3112 53968 3180 54024
rect 3236 53968 3304 54024
rect 3360 53968 3428 54024
rect 3484 53968 3552 54024
rect 3608 53968 3676 54024
rect 3732 53968 3800 54024
rect 3856 53968 3924 54024
rect 3980 53968 4048 54024
rect 4104 53968 4172 54024
rect 4228 53968 4296 54024
rect 4352 53968 4420 54024
rect 4476 53968 4544 54024
rect 4600 53968 4668 54024
rect 4724 53968 4734 54024
rect 2798 53900 4734 53968
rect 2798 53844 2808 53900
rect 2864 53844 2932 53900
rect 2988 53844 3056 53900
rect 3112 53844 3180 53900
rect 3236 53844 3304 53900
rect 3360 53844 3428 53900
rect 3484 53844 3552 53900
rect 3608 53844 3676 53900
rect 3732 53844 3800 53900
rect 3856 53844 3924 53900
rect 3980 53844 4048 53900
rect 4104 53844 4172 53900
rect 4228 53844 4296 53900
rect 4352 53844 4420 53900
rect 4476 53844 4544 53900
rect 4600 53844 4668 53900
rect 4724 53844 4734 53900
rect 2798 53776 4734 53844
rect 2798 53720 2808 53776
rect 2864 53720 2932 53776
rect 2988 53720 3056 53776
rect 3112 53720 3180 53776
rect 3236 53720 3304 53776
rect 3360 53720 3428 53776
rect 3484 53720 3552 53776
rect 3608 53720 3676 53776
rect 3732 53720 3800 53776
rect 3856 53720 3924 53776
rect 3980 53720 4048 53776
rect 4104 53720 4172 53776
rect 4228 53720 4296 53776
rect 4352 53720 4420 53776
rect 4476 53720 4544 53776
rect 4600 53720 4668 53776
rect 4724 53720 4734 53776
rect 2798 53652 4734 53720
rect 2798 53596 2808 53652
rect 2864 53596 2932 53652
rect 2988 53596 3056 53652
rect 3112 53596 3180 53652
rect 3236 53596 3304 53652
rect 3360 53596 3428 53652
rect 3484 53596 3552 53652
rect 3608 53596 3676 53652
rect 3732 53596 3800 53652
rect 3856 53596 3924 53652
rect 3980 53596 4048 53652
rect 4104 53596 4172 53652
rect 4228 53596 4296 53652
rect 4352 53596 4420 53652
rect 4476 53596 4544 53652
rect 4600 53596 4668 53652
rect 4724 53596 4734 53652
rect 2798 53528 4734 53596
rect 2798 53472 2808 53528
rect 2864 53472 2932 53528
rect 2988 53472 3056 53528
rect 3112 53472 3180 53528
rect 3236 53472 3304 53528
rect 3360 53472 3428 53528
rect 3484 53472 3552 53528
rect 3608 53472 3676 53528
rect 3732 53472 3800 53528
rect 3856 53472 3924 53528
rect 3980 53472 4048 53528
rect 4104 53472 4172 53528
rect 4228 53472 4296 53528
rect 4352 53472 4420 53528
rect 4476 53472 4544 53528
rect 4600 53472 4668 53528
rect 4724 53472 4734 53528
rect 2798 53404 4734 53472
rect 2798 53348 2808 53404
rect 2864 53348 2932 53404
rect 2988 53348 3056 53404
rect 3112 53348 3180 53404
rect 3236 53348 3304 53404
rect 3360 53348 3428 53404
rect 3484 53348 3552 53404
rect 3608 53348 3676 53404
rect 3732 53348 3800 53404
rect 3856 53348 3924 53404
rect 3980 53348 4048 53404
rect 4104 53348 4172 53404
rect 4228 53348 4296 53404
rect 4352 53348 4420 53404
rect 4476 53348 4544 53404
rect 4600 53348 4668 53404
rect 4724 53348 4734 53404
rect 2798 53280 4734 53348
rect 2798 53224 2808 53280
rect 2864 53224 2932 53280
rect 2988 53224 3056 53280
rect 3112 53224 3180 53280
rect 3236 53224 3304 53280
rect 3360 53224 3428 53280
rect 3484 53224 3552 53280
rect 3608 53224 3676 53280
rect 3732 53224 3800 53280
rect 3856 53224 3924 53280
rect 3980 53224 4048 53280
rect 4104 53224 4172 53280
rect 4228 53224 4296 53280
rect 4352 53224 4420 53280
rect 4476 53224 4544 53280
rect 4600 53224 4668 53280
rect 4724 53224 4734 53280
rect 2798 53156 4734 53224
rect 2798 53100 2808 53156
rect 2864 53100 2932 53156
rect 2988 53100 3056 53156
rect 3112 53100 3180 53156
rect 3236 53100 3304 53156
rect 3360 53100 3428 53156
rect 3484 53100 3552 53156
rect 3608 53100 3676 53156
rect 3732 53100 3800 53156
rect 3856 53100 3924 53156
rect 3980 53100 4048 53156
rect 4104 53100 4172 53156
rect 4228 53100 4296 53156
rect 4352 53100 4420 53156
rect 4476 53100 4544 53156
rect 4600 53100 4668 53156
rect 4724 53100 4734 53156
rect 2798 53032 4734 53100
rect 2798 52976 2808 53032
rect 2864 52976 2932 53032
rect 2988 52976 3056 53032
rect 3112 52976 3180 53032
rect 3236 52976 3304 53032
rect 3360 52976 3428 53032
rect 3484 52976 3552 53032
rect 3608 52976 3676 53032
rect 3732 52976 3800 53032
rect 3856 52976 3924 53032
rect 3980 52976 4048 53032
rect 4104 52976 4172 53032
rect 4228 52976 4296 53032
rect 4352 52976 4420 53032
rect 4476 52976 4544 53032
rect 4600 52976 4668 53032
rect 4724 52976 4734 53032
rect 2798 52908 4734 52976
rect 2798 52852 2808 52908
rect 2864 52852 2932 52908
rect 2988 52852 3056 52908
rect 3112 52852 3180 52908
rect 3236 52852 3304 52908
rect 3360 52852 3428 52908
rect 3484 52852 3552 52908
rect 3608 52852 3676 52908
rect 3732 52852 3800 52908
rect 3856 52852 3924 52908
rect 3980 52852 4048 52908
rect 4104 52852 4172 52908
rect 4228 52852 4296 52908
rect 4352 52852 4420 52908
rect 4476 52852 4544 52908
rect 4600 52852 4668 52908
rect 4724 52852 4734 52908
rect 2798 52842 4734 52852
rect 5168 54148 7104 54158
rect 5168 54092 5178 54148
rect 5234 54092 5302 54148
rect 5358 54092 5426 54148
rect 5482 54092 5550 54148
rect 5606 54092 5674 54148
rect 5730 54092 5798 54148
rect 5854 54092 5922 54148
rect 5978 54092 6046 54148
rect 6102 54092 6170 54148
rect 6226 54092 6294 54148
rect 6350 54092 6418 54148
rect 6474 54092 6542 54148
rect 6598 54092 6666 54148
rect 6722 54092 6790 54148
rect 6846 54092 6914 54148
rect 6970 54092 7038 54148
rect 7094 54092 7104 54148
rect 5168 54024 7104 54092
rect 5168 53968 5178 54024
rect 5234 53968 5302 54024
rect 5358 53968 5426 54024
rect 5482 53968 5550 54024
rect 5606 53968 5674 54024
rect 5730 53968 5798 54024
rect 5854 53968 5922 54024
rect 5978 53968 6046 54024
rect 6102 53968 6170 54024
rect 6226 53968 6294 54024
rect 6350 53968 6418 54024
rect 6474 53968 6542 54024
rect 6598 53968 6666 54024
rect 6722 53968 6790 54024
rect 6846 53968 6914 54024
rect 6970 53968 7038 54024
rect 7094 53968 7104 54024
rect 5168 53900 7104 53968
rect 5168 53844 5178 53900
rect 5234 53844 5302 53900
rect 5358 53844 5426 53900
rect 5482 53844 5550 53900
rect 5606 53844 5674 53900
rect 5730 53844 5798 53900
rect 5854 53844 5922 53900
rect 5978 53844 6046 53900
rect 6102 53844 6170 53900
rect 6226 53844 6294 53900
rect 6350 53844 6418 53900
rect 6474 53844 6542 53900
rect 6598 53844 6666 53900
rect 6722 53844 6790 53900
rect 6846 53844 6914 53900
rect 6970 53844 7038 53900
rect 7094 53844 7104 53900
rect 5168 53776 7104 53844
rect 5168 53720 5178 53776
rect 5234 53720 5302 53776
rect 5358 53720 5426 53776
rect 5482 53720 5550 53776
rect 5606 53720 5674 53776
rect 5730 53720 5798 53776
rect 5854 53720 5922 53776
rect 5978 53720 6046 53776
rect 6102 53720 6170 53776
rect 6226 53720 6294 53776
rect 6350 53720 6418 53776
rect 6474 53720 6542 53776
rect 6598 53720 6666 53776
rect 6722 53720 6790 53776
rect 6846 53720 6914 53776
rect 6970 53720 7038 53776
rect 7094 53720 7104 53776
rect 5168 53652 7104 53720
rect 5168 53596 5178 53652
rect 5234 53596 5302 53652
rect 5358 53596 5426 53652
rect 5482 53596 5550 53652
rect 5606 53596 5674 53652
rect 5730 53596 5798 53652
rect 5854 53596 5922 53652
rect 5978 53596 6046 53652
rect 6102 53596 6170 53652
rect 6226 53596 6294 53652
rect 6350 53596 6418 53652
rect 6474 53596 6542 53652
rect 6598 53596 6666 53652
rect 6722 53596 6790 53652
rect 6846 53596 6914 53652
rect 6970 53596 7038 53652
rect 7094 53596 7104 53652
rect 5168 53528 7104 53596
rect 5168 53472 5178 53528
rect 5234 53472 5302 53528
rect 5358 53472 5426 53528
rect 5482 53472 5550 53528
rect 5606 53472 5674 53528
rect 5730 53472 5798 53528
rect 5854 53472 5922 53528
rect 5978 53472 6046 53528
rect 6102 53472 6170 53528
rect 6226 53472 6294 53528
rect 6350 53472 6418 53528
rect 6474 53472 6542 53528
rect 6598 53472 6666 53528
rect 6722 53472 6790 53528
rect 6846 53472 6914 53528
rect 6970 53472 7038 53528
rect 7094 53472 7104 53528
rect 5168 53404 7104 53472
rect 5168 53348 5178 53404
rect 5234 53348 5302 53404
rect 5358 53348 5426 53404
rect 5482 53348 5550 53404
rect 5606 53348 5674 53404
rect 5730 53348 5798 53404
rect 5854 53348 5922 53404
rect 5978 53348 6046 53404
rect 6102 53348 6170 53404
rect 6226 53348 6294 53404
rect 6350 53348 6418 53404
rect 6474 53348 6542 53404
rect 6598 53348 6666 53404
rect 6722 53348 6790 53404
rect 6846 53348 6914 53404
rect 6970 53348 7038 53404
rect 7094 53348 7104 53404
rect 5168 53280 7104 53348
rect 5168 53224 5178 53280
rect 5234 53224 5302 53280
rect 5358 53224 5426 53280
rect 5482 53224 5550 53280
rect 5606 53224 5674 53280
rect 5730 53224 5798 53280
rect 5854 53224 5922 53280
rect 5978 53224 6046 53280
rect 6102 53224 6170 53280
rect 6226 53224 6294 53280
rect 6350 53224 6418 53280
rect 6474 53224 6542 53280
rect 6598 53224 6666 53280
rect 6722 53224 6790 53280
rect 6846 53224 6914 53280
rect 6970 53224 7038 53280
rect 7094 53224 7104 53280
rect 5168 53156 7104 53224
rect 5168 53100 5178 53156
rect 5234 53100 5302 53156
rect 5358 53100 5426 53156
rect 5482 53100 5550 53156
rect 5606 53100 5674 53156
rect 5730 53100 5798 53156
rect 5854 53100 5922 53156
rect 5978 53100 6046 53156
rect 6102 53100 6170 53156
rect 6226 53100 6294 53156
rect 6350 53100 6418 53156
rect 6474 53100 6542 53156
rect 6598 53100 6666 53156
rect 6722 53100 6790 53156
rect 6846 53100 6914 53156
rect 6970 53100 7038 53156
rect 7094 53100 7104 53156
rect 5168 53032 7104 53100
rect 5168 52976 5178 53032
rect 5234 52976 5302 53032
rect 5358 52976 5426 53032
rect 5482 52976 5550 53032
rect 5606 52976 5674 53032
rect 5730 52976 5798 53032
rect 5854 52976 5922 53032
rect 5978 52976 6046 53032
rect 6102 52976 6170 53032
rect 6226 52976 6294 53032
rect 6350 52976 6418 53032
rect 6474 52976 6542 53032
rect 6598 52976 6666 53032
rect 6722 52976 6790 53032
rect 6846 52976 6914 53032
rect 6970 52976 7038 53032
rect 7094 52976 7104 53032
rect 5168 52908 7104 52976
rect 5168 52852 5178 52908
rect 5234 52852 5302 52908
rect 5358 52852 5426 52908
rect 5482 52852 5550 52908
rect 5606 52852 5674 52908
rect 5730 52852 5798 52908
rect 5854 52852 5922 52908
rect 5978 52852 6046 52908
rect 6102 52852 6170 52908
rect 6226 52852 6294 52908
rect 6350 52852 6418 52908
rect 6474 52852 6542 52908
rect 6598 52852 6666 52908
rect 6722 52852 6790 52908
rect 6846 52852 6914 52908
rect 6970 52852 7038 52908
rect 7094 52852 7104 52908
rect 5168 52842 7104 52852
rect 7874 54148 9810 54158
rect 7874 54092 7884 54148
rect 7940 54092 8008 54148
rect 8064 54092 8132 54148
rect 8188 54092 8256 54148
rect 8312 54092 8380 54148
rect 8436 54092 8504 54148
rect 8560 54092 8628 54148
rect 8684 54092 8752 54148
rect 8808 54092 8876 54148
rect 8932 54092 9000 54148
rect 9056 54092 9124 54148
rect 9180 54092 9248 54148
rect 9304 54092 9372 54148
rect 9428 54092 9496 54148
rect 9552 54092 9620 54148
rect 9676 54092 9744 54148
rect 9800 54092 9810 54148
rect 7874 54024 9810 54092
rect 7874 53968 7884 54024
rect 7940 53968 8008 54024
rect 8064 53968 8132 54024
rect 8188 53968 8256 54024
rect 8312 53968 8380 54024
rect 8436 53968 8504 54024
rect 8560 53968 8628 54024
rect 8684 53968 8752 54024
rect 8808 53968 8876 54024
rect 8932 53968 9000 54024
rect 9056 53968 9124 54024
rect 9180 53968 9248 54024
rect 9304 53968 9372 54024
rect 9428 53968 9496 54024
rect 9552 53968 9620 54024
rect 9676 53968 9744 54024
rect 9800 53968 9810 54024
rect 7874 53900 9810 53968
rect 7874 53844 7884 53900
rect 7940 53844 8008 53900
rect 8064 53844 8132 53900
rect 8188 53844 8256 53900
rect 8312 53844 8380 53900
rect 8436 53844 8504 53900
rect 8560 53844 8628 53900
rect 8684 53844 8752 53900
rect 8808 53844 8876 53900
rect 8932 53844 9000 53900
rect 9056 53844 9124 53900
rect 9180 53844 9248 53900
rect 9304 53844 9372 53900
rect 9428 53844 9496 53900
rect 9552 53844 9620 53900
rect 9676 53844 9744 53900
rect 9800 53844 9810 53900
rect 7874 53776 9810 53844
rect 7874 53720 7884 53776
rect 7940 53720 8008 53776
rect 8064 53720 8132 53776
rect 8188 53720 8256 53776
rect 8312 53720 8380 53776
rect 8436 53720 8504 53776
rect 8560 53720 8628 53776
rect 8684 53720 8752 53776
rect 8808 53720 8876 53776
rect 8932 53720 9000 53776
rect 9056 53720 9124 53776
rect 9180 53720 9248 53776
rect 9304 53720 9372 53776
rect 9428 53720 9496 53776
rect 9552 53720 9620 53776
rect 9676 53720 9744 53776
rect 9800 53720 9810 53776
rect 7874 53652 9810 53720
rect 7874 53596 7884 53652
rect 7940 53596 8008 53652
rect 8064 53596 8132 53652
rect 8188 53596 8256 53652
rect 8312 53596 8380 53652
rect 8436 53596 8504 53652
rect 8560 53596 8628 53652
rect 8684 53596 8752 53652
rect 8808 53596 8876 53652
rect 8932 53596 9000 53652
rect 9056 53596 9124 53652
rect 9180 53596 9248 53652
rect 9304 53596 9372 53652
rect 9428 53596 9496 53652
rect 9552 53596 9620 53652
rect 9676 53596 9744 53652
rect 9800 53596 9810 53652
rect 7874 53528 9810 53596
rect 7874 53472 7884 53528
rect 7940 53472 8008 53528
rect 8064 53472 8132 53528
rect 8188 53472 8256 53528
rect 8312 53472 8380 53528
rect 8436 53472 8504 53528
rect 8560 53472 8628 53528
rect 8684 53472 8752 53528
rect 8808 53472 8876 53528
rect 8932 53472 9000 53528
rect 9056 53472 9124 53528
rect 9180 53472 9248 53528
rect 9304 53472 9372 53528
rect 9428 53472 9496 53528
rect 9552 53472 9620 53528
rect 9676 53472 9744 53528
rect 9800 53472 9810 53528
rect 7874 53404 9810 53472
rect 7874 53348 7884 53404
rect 7940 53348 8008 53404
rect 8064 53348 8132 53404
rect 8188 53348 8256 53404
rect 8312 53348 8380 53404
rect 8436 53348 8504 53404
rect 8560 53348 8628 53404
rect 8684 53348 8752 53404
rect 8808 53348 8876 53404
rect 8932 53348 9000 53404
rect 9056 53348 9124 53404
rect 9180 53348 9248 53404
rect 9304 53348 9372 53404
rect 9428 53348 9496 53404
rect 9552 53348 9620 53404
rect 9676 53348 9744 53404
rect 9800 53348 9810 53404
rect 7874 53280 9810 53348
rect 7874 53224 7884 53280
rect 7940 53224 8008 53280
rect 8064 53224 8132 53280
rect 8188 53224 8256 53280
rect 8312 53224 8380 53280
rect 8436 53224 8504 53280
rect 8560 53224 8628 53280
rect 8684 53224 8752 53280
rect 8808 53224 8876 53280
rect 8932 53224 9000 53280
rect 9056 53224 9124 53280
rect 9180 53224 9248 53280
rect 9304 53224 9372 53280
rect 9428 53224 9496 53280
rect 9552 53224 9620 53280
rect 9676 53224 9744 53280
rect 9800 53224 9810 53280
rect 7874 53156 9810 53224
rect 7874 53100 7884 53156
rect 7940 53100 8008 53156
rect 8064 53100 8132 53156
rect 8188 53100 8256 53156
rect 8312 53100 8380 53156
rect 8436 53100 8504 53156
rect 8560 53100 8628 53156
rect 8684 53100 8752 53156
rect 8808 53100 8876 53156
rect 8932 53100 9000 53156
rect 9056 53100 9124 53156
rect 9180 53100 9248 53156
rect 9304 53100 9372 53156
rect 9428 53100 9496 53156
rect 9552 53100 9620 53156
rect 9676 53100 9744 53156
rect 9800 53100 9810 53156
rect 7874 53032 9810 53100
rect 7874 52976 7884 53032
rect 7940 52976 8008 53032
rect 8064 52976 8132 53032
rect 8188 52976 8256 53032
rect 8312 52976 8380 53032
rect 8436 52976 8504 53032
rect 8560 52976 8628 53032
rect 8684 52976 8752 53032
rect 8808 52976 8876 53032
rect 8932 52976 9000 53032
rect 9056 52976 9124 53032
rect 9180 52976 9248 53032
rect 9304 52976 9372 53032
rect 9428 52976 9496 53032
rect 9552 52976 9620 53032
rect 9676 52976 9744 53032
rect 9800 52976 9810 53032
rect 7874 52908 9810 52976
rect 7874 52852 7884 52908
rect 7940 52852 8008 52908
rect 8064 52852 8132 52908
rect 8188 52852 8256 52908
rect 8312 52852 8380 52908
rect 8436 52852 8504 52908
rect 8560 52852 8628 52908
rect 8684 52852 8752 52908
rect 8808 52852 8876 52908
rect 8932 52852 9000 52908
rect 9056 52852 9124 52908
rect 9180 52852 9248 52908
rect 9304 52852 9372 52908
rect 9428 52852 9496 52908
rect 9552 52852 9620 52908
rect 9676 52852 9744 52908
rect 9800 52852 9810 52908
rect 7874 52842 9810 52852
rect 10244 54148 12180 54158
rect 10244 54092 10254 54148
rect 10310 54092 10378 54148
rect 10434 54092 10502 54148
rect 10558 54092 10626 54148
rect 10682 54092 10750 54148
rect 10806 54092 10874 54148
rect 10930 54092 10998 54148
rect 11054 54092 11122 54148
rect 11178 54092 11246 54148
rect 11302 54092 11370 54148
rect 11426 54092 11494 54148
rect 11550 54092 11618 54148
rect 11674 54092 11742 54148
rect 11798 54092 11866 54148
rect 11922 54092 11990 54148
rect 12046 54092 12114 54148
rect 12170 54092 12180 54148
rect 10244 54024 12180 54092
rect 10244 53968 10254 54024
rect 10310 53968 10378 54024
rect 10434 53968 10502 54024
rect 10558 53968 10626 54024
rect 10682 53968 10750 54024
rect 10806 53968 10874 54024
rect 10930 53968 10998 54024
rect 11054 53968 11122 54024
rect 11178 53968 11246 54024
rect 11302 53968 11370 54024
rect 11426 53968 11494 54024
rect 11550 53968 11618 54024
rect 11674 53968 11742 54024
rect 11798 53968 11866 54024
rect 11922 53968 11990 54024
rect 12046 53968 12114 54024
rect 12170 53968 12180 54024
rect 10244 53900 12180 53968
rect 10244 53844 10254 53900
rect 10310 53844 10378 53900
rect 10434 53844 10502 53900
rect 10558 53844 10626 53900
rect 10682 53844 10750 53900
rect 10806 53844 10874 53900
rect 10930 53844 10998 53900
rect 11054 53844 11122 53900
rect 11178 53844 11246 53900
rect 11302 53844 11370 53900
rect 11426 53844 11494 53900
rect 11550 53844 11618 53900
rect 11674 53844 11742 53900
rect 11798 53844 11866 53900
rect 11922 53844 11990 53900
rect 12046 53844 12114 53900
rect 12170 53844 12180 53900
rect 10244 53776 12180 53844
rect 10244 53720 10254 53776
rect 10310 53720 10378 53776
rect 10434 53720 10502 53776
rect 10558 53720 10626 53776
rect 10682 53720 10750 53776
rect 10806 53720 10874 53776
rect 10930 53720 10998 53776
rect 11054 53720 11122 53776
rect 11178 53720 11246 53776
rect 11302 53720 11370 53776
rect 11426 53720 11494 53776
rect 11550 53720 11618 53776
rect 11674 53720 11742 53776
rect 11798 53720 11866 53776
rect 11922 53720 11990 53776
rect 12046 53720 12114 53776
rect 12170 53720 12180 53776
rect 10244 53652 12180 53720
rect 10244 53596 10254 53652
rect 10310 53596 10378 53652
rect 10434 53596 10502 53652
rect 10558 53596 10626 53652
rect 10682 53596 10750 53652
rect 10806 53596 10874 53652
rect 10930 53596 10998 53652
rect 11054 53596 11122 53652
rect 11178 53596 11246 53652
rect 11302 53596 11370 53652
rect 11426 53596 11494 53652
rect 11550 53596 11618 53652
rect 11674 53596 11742 53652
rect 11798 53596 11866 53652
rect 11922 53596 11990 53652
rect 12046 53596 12114 53652
rect 12170 53596 12180 53652
rect 10244 53528 12180 53596
rect 10244 53472 10254 53528
rect 10310 53472 10378 53528
rect 10434 53472 10502 53528
rect 10558 53472 10626 53528
rect 10682 53472 10750 53528
rect 10806 53472 10874 53528
rect 10930 53472 10998 53528
rect 11054 53472 11122 53528
rect 11178 53472 11246 53528
rect 11302 53472 11370 53528
rect 11426 53472 11494 53528
rect 11550 53472 11618 53528
rect 11674 53472 11742 53528
rect 11798 53472 11866 53528
rect 11922 53472 11990 53528
rect 12046 53472 12114 53528
rect 12170 53472 12180 53528
rect 10244 53404 12180 53472
rect 10244 53348 10254 53404
rect 10310 53348 10378 53404
rect 10434 53348 10502 53404
rect 10558 53348 10626 53404
rect 10682 53348 10750 53404
rect 10806 53348 10874 53404
rect 10930 53348 10998 53404
rect 11054 53348 11122 53404
rect 11178 53348 11246 53404
rect 11302 53348 11370 53404
rect 11426 53348 11494 53404
rect 11550 53348 11618 53404
rect 11674 53348 11742 53404
rect 11798 53348 11866 53404
rect 11922 53348 11990 53404
rect 12046 53348 12114 53404
rect 12170 53348 12180 53404
rect 10244 53280 12180 53348
rect 10244 53224 10254 53280
rect 10310 53224 10378 53280
rect 10434 53224 10502 53280
rect 10558 53224 10626 53280
rect 10682 53224 10750 53280
rect 10806 53224 10874 53280
rect 10930 53224 10998 53280
rect 11054 53224 11122 53280
rect 11178 53224 11246 53280
rect 11302 53224 11370 53280
rect 11426 53224 11494 53280
rect 11550 53224 11618 53280
rect 11674 53224 11742 53280
rect 11798 53224 11866 53280
rect 11922 53224 11990 53280
rect 12046 53224 12114 53280
rect 12170 53224 12180 53280
rect 10244 53156 12180 53224
rect 10244 53100 10254 53156
rect 10310 53100 10378 53156
rect 10434 53100 10502 53156
rect 10558 53100 10626 53156
rect 10682 53100 10750 53156
rect 10806 53100 10874 53156
rect 10930 53100 10998 53156
rect 11054 53100 11122 53156
rect 11178 53100 11246 53156
rect 11302 53100 11370 53156
rect 11426 53100 11494 53156
rect 11550 53100 11618 53156
rect 11674 53100 11742 53156
rect 11798 53100 11866 53156
rect 11922 53100 11990 53156
rect 12046 53100 12114 53156
rect 12170 53100 12180 53156
rect 10244 53032 12180 53100
rect 10244 52976 10254 53032
rect 10310 52976 10378 53032
rect 10434 52976 10502 53032
rect 10558 52976 10626 53032
rect 10682 52976 10750 53032
rect 10806 52976 10874 53032
rect 10930 52976 10998 53032
rect 11054 52976 11122 53032
rect 11178 52976 11246 53032
rect 11302 52976 11370 53032
rect 11426 52976 11494 53032
rect 11550 52976 11618 53032
rect 11674 52976 11742 53032
rect 11798 52976 11866 53032
rect 11922 52976 11990 53032
rect 12046 52976 12114 53032
rect 12170 52976 12180 53032
rect 10244 52908 12180 52976
rect 10244 52852 10254 52908
rect 10310 52852 10378 52908
rect 10434 52852 10502 52908
rect 10558 52852 10626 52908
rect 10682 52852 10750 52908
rect 10806 52852 10874 52908
rect 10930 52852 10998 52908
rect 11054 52852 11122 52908
rect 11178 52852 11246 52908
rect 11302 52852 11370 52908
rect 11426 52852 11494 52908
rect 11550 52852 11618 52908
rect 11674 52852 11742 52908
rect 11798 52852 11866 52908
rect 11922 52852 11990 52908
rect 12046 52852 12114 52908
rect 12170 52852 12180 52908
rect 10244 52842 12180 52852
rect 12861 54148 14673 54158
rect 12861 54092 12871 54148
rect 12927 54092 12995 54148
rect 13051 54092 13119 54148
rect 13175 54092 13243 54148
rect 13299 54092 13367 54148
rect 13423 54092 13491 54148
rect 13547 54092 13615 54148
rect 13671 54092 13739 54148
rect 13795 54092 13863 54148
rect 13919 54092 13987 54148
rect 14043 54092 14111 54148
rect 14167 54092 14235 54148
rect 14291 54092 14359 54148
rect 14415 54092 14483 54148
rect 14539 54092 14607 54148
rect 14663 54092 14673 54148
rect 12861 54024 14673 54092
rect 12861 53968 12871 54024
rect 12927 53968 12995 54024
rect 13051 53968 13119 54024
rect 13175 53968 13243 54024
rect 13299 53968 13367 54024
rect 13423 53968 13491 54024
rect 13547 53968 13615 54024
rect 13671 53968 13739 54024
rect 13795 53968 13863 54024
rect 13919 53968 13987 54024
rect 14043 53968 14111 54024
rect 14167 53968 14235 54024
rect 14291 53968 14359 54024
rect 14415 53968 14483 54024
rect 14539 53968 14607 54024
rect 14663 53968 14673 54024
rect 12861 53900 14673 53968
rect 12861 53844 12871 53900
rect 12927 53844 12995 53900
rect 13051 53844 13119 53900
rect 13175 53844 13243 53900
rect 13299 53844 13367 53900
rect 13423 53844 13491 53900
rect 13547 53844 13615 53900
rect 13671 53844 13739 53900
rect 13795 53844 13863 53900
rect 13919 53844 13987 53900
rect 14043 53844 14111 53900
rect 14167 53844 14235 53900
rect 14291 53844 14359 53900
rect 14415 53844 14483 53900
rect 14539 53844 14607 53900
rect 14663 53844 14673 53900
rect 12861 53776 14673 53844
rect 12861 53720 12871 53776
rect 12927 53720 12995 53776
rect 13051 53720 13119 53776
rect 13175 53720 13243 53776
rect 13299 53720 13367 53776
rect 13423 53720 13491 53776
rect 13547 53720 13615 53776
rect 13671 53720 13739 53776
rect 13795 53720 13863 53776
rect 13919 53720 13987 53776
rect 14043 53720 14111 53776
rect 14167 53720 14235 53776
rect 14291 53720 14359 53776
rect 14415 53720 14483 53776
rect 14539 53720 14607 53776
rect 14663 53720 14673 53776
rect 12861 53652 14673 53720
rect 12861 53596 12871 53652
rect 12927 53596 12995 53652
rect 13051 53596 13119 53652
rect 13175 53596 13243 53652
rect 13299 53596 13367 53652
rect 13423 53596 13491 53652
rect 13547 53596 13615 53652
rect 13671 53596 13739 53652
rect 13795 53596 13863 53652
rect 13919 53596 13987 53652
rect 14043 53596 14111 53652
rect 14167 53596 14235 53652
rect 14291 53596 14359 53652
rect 14415 53596 14483 53652
rect 14539 53596 14607 53652
rect 14663 53596 14673 53652
rect 12861 53528 14673 53596
rect 12861 53472 12871 53528
rect 12927 53472 12995 53528
rect 13051 53472 13119 53528
rect 13175 53472 13243 53528
rect 13299 53472 13367 53528
rect 13423 53472 13491 53528
rect 13547 53472 13615 53528
rect 13671 53472 13739 53528
rect 13795 53472 13863 53528
rect 13919 53472 13987 53528
rect 14043 53472 14111 53528
rect 14167 53472 14235 53528
rect 14291 53472 14359 53528
rect 14415 53472 14483 53528
rect 14539 53472 14607 53528
rect 14663 53472 14673 53528
rect 12861 53404 14673 53472
rect 12861 53348 12871 53404
rect 12927 53348 12995 53404
rect 13051 53348 13119 53404
rect 13175 53348 13243 53404
rect 13299 53348 13367 53404
rect 13423 53348 13491 53404
rect 13547 53348 13615 53404
rect 13671 53348 13739 53404
rect 13795 53348 13863 53404
rect 13919 53348 13987 53404
rect 14043 53348 14111 53404
rect 14167 53348 14235 53404
rect 14291 53348 14359 53404
rect 14415 53348 14483 53404
rect 14539 53348 14607 53404
rect 14663 53348 14673 53404
rect 12861 53280 14673 53348
rect 12861 53224 12871 53280
rect 12927 53224 12995 53280
rect 13051 53224 13119 53280
rect 13175 53224 13243 53280
rect 13299 53224 13367 53280
rect 13423 53224 13491 53280
rect 13547 53224 13615 53280
rect 13671 53224 13739 53280
rect 13795 53224 13863 53280
rect 13919 53224 13987 53280
rect 14043 53224 14111 53280
rect 14167 53224 14235 53280
rect 14291 53224 14359 53280
rect 14415 53224 14483 53280
rect 14539 53224 14607 53280
rect 14663 53224 14673 53280
rect 12861 53156 14673 53224
rect 12861 53100 12871 53156
rect 12927 53100 12995 53156
rect 13051 53100 13119 53156
rect 13175 53100 13243 53156
rect 13299 53100 13367 53156
rect 13423 53100 13491 53156
rect 13547 53100 13615 53156
rect 13671 53100 13739 53156
rect 13795 53100 13863 53156
rect 13919 53100 13987 53156
rect 14043 53100 14111 53156
rect 14167 53100 14235 53156
rect 14291 53100 14359 53156
rect 14415 53100 14483 53156
rect 14539 53100 14607 53156
rect 14663 53100 14673 53156
rect 12861 53032 14673 53100
rect 12861 52976 12871 53032
rect 12927 52976 12995 53032
rect 13051 52976 13119 53032
rect 13175 52976 13243 53032
rect 13299 52976 13367 53032
rect 13423 52976 13491 53032
rect 13547 52976 13615 53032
rect 13671 52976 13739 53032
rect 13795 52976 13863 53032
rect 13919 52976 13987 53032
rect 14043 52976 14111 53032
rect 14167 52976 14235 53032
rect 14291 52976 14359 53032
rect 14415 52976 14483 53032
rect 14539 52976 14607 53032
rect 14663 52976 14673 53032
rect 12861 52908 14673 52976
rect 12861 52852 12871 52908
rect 12927 52852 12995 52908
rect 13051 52852 13119 52908
rect 13175 52852 13243 52908
rect 13299 52852 13367 52908
rect 13423 52852 13491 52908
rect 13547 52852 13615 52908
rect 13671 52852 13739 52908
rect 13795 52852 13863 52908
rect 13919 52852 13987 52908
rect 14043 52852 14111 52908
rect 14167 52852 14235 52908
rect 14291 52852 14359 52908
rect 14415 52852 14483 52908
rect 14539 52852 14607 52908
rect 14663 52852 14673 52908
rect 12861 52842 14673 52852
rect 10 52814 86 52824
rect 14892 52824 14902 54176
rect 14958 52824 14968 54176
rect 14892 52814 14968 52824
rect 10 52576 86 52586
rect 10 51224 20 52576
rect 76 51224 86 52576
rect 14892 52576 14968 52586
rect 305 52548 2117 52558
rect 305 52492 315 52548
rect 371 52492 439 52548
rect 495 52492 563 52548
rect 619 52492 687 52548
rect 743 52492 811 52548
rect 867 52492 935 52548
rect 991 52492 1059 52548
rect 1115 52492 1183 52548
rect 1239 52492 1307 52548
rect 1363 52492 1431 52548
rect 1487 52492 1555 52548
rect 1611 52492 1679 52548
rect 1735 52492 1803 52548
rect 1859 52492 1927 52548
rect 1983 52492 2051 52548
rect 2107 52492 2117 52548
rect 305 52424 2117 52492
rect 305 52368 315 52424
rect 371 52368 439 52424
rect 495 52368 563 52424
rect 619 52368 687 52424
rect 743 52368 811 52424
rect 867 52368 935 52424
rect 991 52368 1059 52424
rect 1115 52368 1183 52424
rect 1239 52368 1307 52424
rect 1363 52368 1431 52424
rect 1487 52368 1555 52424
rect 1611 52368 1679 52424
rect 1735 52368 1803 52424
rect 1859 52368 1927 52424
rect 1983 52368 2051 52424
rect 2107 52368 2117 52424
rect 305 52300 2117 52368
rect 305 52244 315 52300
rect 371 52244 439 52300
rect 495 52244 563 52300
rect 619 52244 687 52300
rect 743 52244 811 52300
rect 867 52244 935 52300
rect 991 52244 1059 52300
rect 1115 52244 1183 52300
rect 1239 52244 1307 52300
rect 1363 52244 1431 52300
rect 1487 52244 1555 52300
rect 1611 52244 1679 52300
rect 1735 52244 1803 52300
rect 1859 52244 1927 52300
rect 1983 52244 2051 52300
rect 2107 52244 2117 52300
rect 305 52176 2117 52244
rect 305 52120 315 52176
rect 371 52120 439 52176
rect 495 52120 563 52176
rect 619 52120 687 52176
rect 743 52120 811 52176
rect 867 52120 935 52176
rect 991 52120 1059 52176
rect 1115 52120 1183 52176
rect 1239 52120 1307 52176
rect 1363 52120 1431 52176
rect 1487 52120 1555 52176
rect 1611 52120 1679 52176
rect 1735 52120 1803 52176
rect 1859 52120 1927 52176
rect 1983 52120 2051 52176
rect 2107 52120 2117 52176
rect 305 52052 2117 52120
rect 305 51996 315 52052
rect 371 51996 439 52052
rect 495 51996 563 52052
rect 619 51996 687 52052
rect 743 51996 811 52052
rect 867 51996 935 52052
rect 991 51996 1059 52052
rect 1115 51996 1183 52052
rect 1239 51996 1307 52052
rect 1363 51996 1431 52052
rect 1487 51996 1555 52052
rect 1611 51996 1679 52052
rect 1735 51996 1803 52052
rect 1859 51996 1927 52052
rect 1983 51996 2051 52052
rect 2107 51996 2117 52052
rect 305 51928 2117 51996
rect 305 51872 315 51928
rect 371 51872 439 51928
rect 495 51872 563 51928
rect 619 51872 687 51928
rect 743 51872 811 51928
rect 867 51872 935 51928
rect 991 51872 1059 51928
rect 1115 51872 1183 51928
rect 1239 51872 1307 51928
rect 1363 51872 1431 51928
rect 1487 51872 1555 51928
rect 1611 51872 1679 51928
rect 1735 51872 1803 51928
rect 1859 51872 1927 51928
rect 1983 51872 2051 51928
rect 2107 51872 2117 51928
rect 305 51804 2117 51872
rect 305 51748 315 51804
rect 371 51748 439 51804
rect 495 51748 563 51804
rect 619 51748 687 51804
rect 743 51748 811 51804
rect 867 51748 935 51804
rect 991 51748 1059 51804
rect 1115 51748 1183 51804
rect 1239 51748 1307 51804
rect 1363 51748 1431 51804
rect 1487 51748 1555 51804
rect 1611 51748 1679 51804
rect 1735 51748 1803 51804
rect 1859 51748 1927 51804
rect 1983 51748 2051 51804
rect 2107 51748 2117 51804
rect 305 51680 2117 51748
rect 305 51624 315 51680
rect 371 51624 439 51680
rect 495 51624 563 51680
rect 619 51624 687 51680
rect 743 51624 811 51680
rect 867 51624 935 51680
rect 991 51624 1059 51680
rect 1115 51624 1183 51680
rect 1239 51624 1307 51680
rect 1363 51624 1431 51680
rect 1487 51624 1555 51680
rect 1611 51624 1679 51680
rect 1735 51624 1803 51680
rect 1859 51624 1927 51680
rect 1983 51624 2051 51680
rect 2107 51624 2117 51680
rect 305 51556 2117 51624
rect 305 51500 315 51556
rect 371 51500 439 51556
rect 495 51500 563 51556
rect 619 51500 687 51556
rect 743 51500 811 51556
rect 867 51500 935 51556
rect 991 51500 1059 51556
rect 1115 51500 1183 51556
rect 1239 51500 1307 51556
rect 1363 51500 1431 51556
rect 1487 51500 1555 51556
rect 1611 51500 1679 51556
rect 1735 51500 1803 51556
rect 1859 51500 1927 51556
rect 1983 51500 2051 51556
rect 2107 51500 2117 51556
rect 305 51432 2117 51500
rect 305 51376 315 51432
rect 371 51376 439 51432
rect 495 51376 563 51432
rect 619 51376 687 51432
rect 743 51376 811 51432
rect 867 51376 935 51432
rect 991 51376 1059 51432
rect 1115 51376 1183 51432
rect 1239 51376 1307 51432
rect 1363 51376 1431 51432
rect 1487 51376 1555 51432
rect 1611 51376 1679 51432
rect 1735 51376 1803 51432
rect 1859 51376 1927 51432
rect 1983 51376 2051 51432
rect 2107 51376 2117 51432
rect 305 51308 2117 51376
rect 305 51252 315 51308
rect 371 51252 439 51308
rect 495 51252 563 51308
rect 619 51252 687 51308
rect 743 51252 811 51308
rect 867 51252 935 51308
rect 991 51252 1059 51308
rect 1115 51252 1183 51308
rect 1239 51252 1307 51308
rect 1363 51252 1431 51308
rect 1487 51252 1555 51308
rect 1611 51252 1679 51308
rect 1735 51252 1803 51308
rect 1859 51252 1927 51308
rect 1983 51252 2051 51308
rect 2107 51252 2117 51308
rect 305 51242 2117 51252
rect 2798 52548 4734 52558
rect 2798 52492 2808 52548
rect 2864 52492 2932 52548
rect 2988 52492 3056 52548
rect 3112 52492 3180 52548
rect 3236 52492 3304 52548
rect 3360 52492 3428 52548
rect 3484 52492 3552 52548
rect 3608 52492 3676 52548
rect 3732 52492 3800 52548
rect 3856 52492 3924 52548
rect 3980 52492 4048 52548
rect 4104 52492 4172 52548
rect 4228 52492 4296 52548
rect 4352 52492 4420 52548
rect 4476 52492 4544 52548
rect 4600 52492 4668 52548
rect 4724 52492 4734 52548
rect 2798 52424 4734 52492
rect 2798 52368 2808 52424
rect 2864 52368 2932 52424
rect 2988 52368 3056 52424
rect 3112 52368 3180 52424
rect 3236 52368 3304 52424
rect 3360 52368 3428 52424
rect 3484 52368 3552 52424
rect 3608 52368 3676 52424
rect 3732 52368 3800 52424
rect 3856 52368 3924 52424
rect 3980 52368 4048 52424
rect 4104 52368 4172 52424
rect 4228 52368 4296 52424
rect 4352 52368 4420 52424
rect 4476 52368 4544 52424
rect 4600 52368 4668 52424
rect 4724 52368 4734 52424
rect 2798 52300 4734 52368
rect 2798 52244 2808 52300
rect 2864 52244 2932 52300
rect 2988 52244 3056 52300
rect 3112 52244 3180 52300
rect 3236 52244 3304 52300
rect 3360 52244 3428 52300
rect 3484 52244 3552 52300
rect 3608 52244 3676 52300
rect 3732 52244 3800 52300
rect 3856 52244 3924 52300
rect 3980 52244 4048 52300
rect 4104 52244 4172 52300
rect 4228 52244 4296 52300
rect 4352 52244 4420 52300
rect 4476 52244 4544 52300
rect 4600 52244 4668 52300
rect 4724 52244 4734 52300
rect 2798 52176 4734 52244
rect 2798 52120 2808 52176
rect 2864 52120 2932 52176
rect 2988 52120 3056 52176
rect 3112 52120 3180 52176
rect 3236 52120 3304 52176
rect 3360 52120 3428 52176
rect 3484 52120 3552 52176
rect 3608 52120 3676 52176
rect 3732 52120 3800 52176
rect 3856 52120 3924 52176
rect 3980 52120 4048 52176
rect 4104 52120 4172 52176
rect 4228 52120 4296 52176
rect 4352 52120 4420 52176
rect 4476 52120 4544 52176
rect 4600 52120 4668 52176
rect 4724 52120 4734 52176
rect 2798 52052 4734 52120
rect 2798 51996 2808 52052
rect 2864 51996 2932 52052
rect 2988 51996 3056 52052
rect 3112 51996 3180 52052
rect 3236 51996 3304 52052
rect 3360 51996 3428 52052
rect 3484 51996 3552 52052
rect 3608 51996 3676 52052
rect 3732 51996 3800 52052
rect 3856 51996 3924 52052
rect 3980 51996 4048 52052
rect 4104 51996 4172 52052
rect 4228 51996 4296 52052
rect 4352 51996 4420 52052
rect 4476 51996 4544 52052
rect 4600 51996 4668 52052
rect 4724 51996 4734 52052
rect 2798 51928 4734 51996
rect 2798 51872 2808 51928
rect 2864 51872 2932 51928
rect 2988 51872 3056 51928
rect 3112 51872 3180 51928
rect 3236 51872 3304 51928
rect 3360 51872 3428 51928
rect 3484 51872 3552 51928
rect 3608 51872 3676 51928
rect 3732 51872 3800 51928
rect 3856 51872 3924 51928
rect 3980 51872 4048 51928
rect 4104 51872 4172 51928
rect 4228 51872 4296 51928
rect 4352 51872 4420 51928
rect 4476 51872 4544 51928
rect 4600 51872 4668 51928
rect 4724 51872 4734 51928
rect 2798 51804 4734 51872
rect 2798 51748 2808 51804
rect 2864 51748 2932 51804
rect 2988 51748 3056 51804
rect 3112 51748 3180 51804
rect 3236 51748 3304 51804
rect 3360 51748 3428 51804
rect 3484 51748 3552 51804
rect 3608 51748 3676 51804
rect 3732 51748 3800 51804
rect 3856 51748 3924 51804
rect 3980 51748 4048 51804
rect 4104 51748 4172 51804
rect 4228 51748 4296 51804
rect 4352 51748 4420 51804
rect 4476 51748 4544 51804
rect 4600 51748 4668 51804
rect 4724 51748 4734 51804
rect 2798 51680 4734 51748
rect 2798 51624 2808 51680
rect 2864 51624 2932 51680
rect 2988 51624 3056 51680
rect 3112 51624 3180 51680
rect 3236 51624 3304 51680
rect 3360 51624 3428 51680
rect 3484 51624 3552 51680
rect 3608 51624 3676 51680
rect 3732 51624 3800 51680
rect 3856 51624 3924 51680
rect 3980 51624 4048 51680
rect 4104 51624 4172 51680
rect 4228 51624 4296 51680
rect 4352 51624 4420 51680
rect 4476 51624 4544 51680
rect 4600 51624 4668 51680
rect 4724 51624 4734 51680
rect 2798 51556 4734 51624
rect 2798 51500 2808 51556
rect 2864 51500 2932 51556
rect 2988 51500 3056 51556
rect 3112 51500 3180 51556
rect 3236 51500 3304 51556
rect 3360 51500 3428 51556
rect 3484 51500 3552 51556
rect 3608 51500 3676 51556
rect 3732 51500 3800 51556
rect 3856 51500 3924 51556
rect 3980 51500 4048 51556
rect 4104 51500 4172 51556
rect 4228 51500 4296 51556
rect 4352 51500 4420 51556
rect 4476 51500 4544 51556
rect 4600 51500 4668 51556
rect 4724 51500 4734 51556
rect 2798 51432 4734 51500
rect 2798 51376 2808 51432
rect 2864 51376 2932 51432
rect 2988 51376 3056 51432
rect 3112 51376 3180 51432
rect 3236 51376 3304 51432
rect 3360 51376 3428 51432
rect 3484 51376 3552 51432
rect 3608 51376 3676 51432
rect 3732 51376 3800 51432
rect 3856 51376 3924 51432
rect 3980 51376 4048 51432
rect 4104 51376 4172 51432
rect 4228 51376 4296 51432
rect 4352 51376 4420 51432
rect 4476 51376 4544 51432
rect 4600 51376 4668 51432
rect 4724 51376 4734 51432
rect 2798 51308 4734 51376
rect 2798 51252 2808 51308
rect 2864 51252 2932 51308
rect 2988 51252 3056 51308
rect 3112 51252 3180 51308
rect 3236 51252 3304 51308
rect 3360 51252 3428 51308
rect 3484 51252 3552 51308
rect 3608 51252 3676 51308
rect 3732 51252 3800 51308
rect 3856 51252 3924 51308
rect 3980 51252 4048 51308
rect 4104 51252 4172 51308
rect 4228 51252 4296 51308
rect 4352 51252 4420 51308
rect 4476 51252 4544 51308
rect 4600 51252 4668 51308
rect 4724 51252 4734 51308
rect 2798 51242 4734 51252
rect 5168 52548 7104 52558
rect 5168 52492 5178 52548
rect 5234 52492 5302 52548
rect 5358 52492 5426 52548
rect 5482 52492 5550 52548
rect 5606 52492 5674 52548
rect 5730 52492 5798 52548
rect 5854 52492 5922 52548
rect 5978 52492 6046 52548
rect 6102 52492 6170 52548
rect 6226 52492 6294 52548
rect 6350 52492 6418 52548
rect 6474 52492 6542 52548
rect 6598 52492 6666 52548
rect 6722 52492 6790 52548
rect 6846 52492 6914 52548
rect 6970 52492 7038 52548
rect 7094 52492 7104 52548
rect 5168 52424 7104 52492
rect 5168 52368 5178 52424
rect 5234 52368 5302 52424
rect 5358 52368 5426 52424
rect 5482 52368 5550 52424
rect 5606 52368 5674 52424
rect 5730 52368 5798 52424
rect 5854 52368 5922 52424
rect 5978 52368 6046 52424
rect 6102 52368 6170 52424
rect 6226 52368 6294 52424
rect 6350 52368 6418 52424
rect 6474 52368 6542 52424
rect 6598 52368 6666 52424
rect 6722 52368 6790 52424
rect 6846 52368 6914 52424
rect 6970 52368 7038 52424
rect 7094 52368 7104 52424
rect 5168 52300 7104 52368
rect 5168 52244 5178 52300
rect 5234 52244 5302 52300
rect 5358 52244 5426 52300
rect 5482 52244 5550 52300
rect 5606 52244 5674 52300
rect 5730 52244 5798 52300
rect 5854 52244 5922 52300
rect 5978 52244 6046 52300
rect 6102 52244 6170 52300
rect 6226 52244 6294 52300
rect 6350 52244 6418 52300
rect 6474 52244 6542 52300
rect 6598 52244 6666 52300
rect 6722 52244 6790 52300
rect 6846 52244 6914 52300
rect 6970 52244 7038 52300
rect 7094 52244 7104 52300
rect 5168 52176 7104 52244
rect 5168 52120 5178 52176
rect 5234 52120 5302 52176
rect 5358 52120 5426 52176
rect 5482 52120 5550 52176
rect 5606 52120 5674 52176
rect 5730 52120 5798 52176
rect 5854 52120 5922 52176
rect 5978 52120 6046 52176
rect 6102 52120 6170 52176
rect 6226 52120 6294 52176
rect 6350 52120 6418 52176
rect 6474 52120 6542 52176
rect 6598 52120 6666 52176
rect 6722 52120 6790 52176
rect 6846 52120 6914 52176
rect 6970 52120 7038 52176
rect 7094 52120 7104 52176
rect 5168 52052 7104 52120
rect 5168 51996 5178 52052
rect 5234 51996 5302 52052
rect 5358 51996 5426 52052
rect 5482 51996 5550 52052
rect 5606 51996 5674 52052
rect 5730 51996 5798 52052
rect 5854 51996 5922 52052
rect 5978 51996 6046 52052
rect 6102 51996 6170 52052
rect 6226 51996 6294 52052
rect 6350 51996 6418 52052
rect 6474 51996 6542 52052
rect 6598 51996 6666 52052
rect 6722 51996 6790 52052
rect 6846 51996 6914 52052
rect 6970 51996 7038 52052
rect 7094 51996 7104 52052
rect 5168 51928 7104 51996
rect 5168 51872 5178 51928
rect 5234 51872 5302 51928
rect 5358 51872 5426 51928
rect 5482 51872 5550 51928
rect 5606 51872 5674 51928
rect 5730 51872 5798 51928
rect 5854 51872 5922 51928
rect 5978 51872 6046 51928
rect 6102 51872 6170 51928
rect 6226 51872 6294 51928
rect 6350 51872 6418 51928
rect 6474 51872 6542 51928
rect 6598 51872 6666 51928
rect 6722 51872 6790 51928
rect 6846 51872 6914 51928
rect 6970 51872 7038 51928
rect 7094 51872 7104 51928
rect 5168 51804 7104 51872
rect 5168 51748 5178 51804
rect 5234 51748 5302 51804
rect 5358 51748 5426 51804
rect 5482 51748 5550 51804
rect 5606 51748 5674 51804
rect 5730 51748 5798 51804
rect 5854 51748 5922 51804
rect 5978 51748 6046 51804
rect 6102 51748 6170 51804
rect 6226 51748 6294 51804
rect 6350 51748 6418 51804
rect 6474 51748 6542 51804
rect 6598 51748 6666 51804
rect 6722 51748 6790 51804
rect 6846 51748 6914 51804
rect 6970 51748 7038 51804
rect 7094 51748 7104 51804
rect 5168 51680 7104 51748
rect 5168 51624 5178 51680
rect 5234 51624 5302 51680
rect 5358 51624 5426 51680
rect 5482 51624 5550 51680
rect 5606 51624 5674 51680
rect 5730 51624 5798 51680
rect 5854 51624 5922 51680
rect 5978 51624 6046 51680
rect 6102 51624 6170 51680
rect 6226 51624 6294 51680
rect 6350 51624 6418 51680
rect 6474 51624 6542 51680
rect 6598 51624 6666 51680
rect 6722 51624 6790 51680
rect 6846 51624 6914 51680
rect 6970 51624 7038 51680
rect 7094 51624 7104 51680
rect 5168 51556 7104 51624
rect 5168 51500 5178 51556
rect 5234 51500 5302 51556
rect 5358 51500 5426 51556
rect 5482 51500 5550 51556
rect 5606 51500 5674 51556
rect 5730 51500 5798 51556
rect 5854 51500 5922 51556
rect 5978 51500 6046 51556
rect 6102 51500 6170 51556
rect 6226 51500 6294 51556
rect 6350 51500 6418 51556
rect 6474 51500 6542 51556
rect 6598 51500 6666 51556
rect 6722 51500 6790 51556
rect 6846 51500 6914 51556
rect 6970 51500 7038 51556
rect 7094 51500 7104 51556
rect 5168 51432 7104 51500
rect 5168 51376 5178 51432
rect 5234 51376 5302 51432
rect 5358 51376 5426 51432
rect 5482 51376 5550 51432
rect 5606 51376 5674 51432
rect 5730 51376 5798 51432
rect 5854 51376 5922 51432
rect 5978 51376 6046 51432
rect 6102 51376 6170 51432
rect 6226 51376 6294 51432
rect 6350 51376 6418 51432
rect 6474 51376 6542 51432
rect 6598 51376 6666 51432
rect 6722 51376 6790 51432
rect 6846 51376 6914 51432
rect 6970 51376 7038 51432
rect 7094 51376 7104 51432
rect 5168 51308 7104 51376
rect 5168 51252 5178 51308
rect 5234 51252 5302 51308
rect 5358 51252 5426 51308
rect 5482 51252 5550 51308
rect 5606 51252 5674 51308
rect 5730 51252 5798 51308
rect 5854 51252 5922 51308
rect 5978 51252 6046 51308
rect 6102 51252 6170 51308
rect 6226 51252 6294 51308
rect 6350 51252 6418 51308
rect 6474 51252 6542 51308
rect 6598 51252 6666 51308
rect 6722 51252 6790 51308
rect 6846 51252 6914 51308
rect 6970 51252 7038 51308
rect 7094 51252 7104 51308
rect 5168 51242 7104 51252
rect 7874 52548 9810 52558
rect 7874 52492 7884 52548
rect 7940 52492 8008 52548
rect 8064 52492 8132 52548
rect 8188 52492 8256 52548
rect 8312 52492 8380 52548
rect 8436 52492 8504 52548
rect 8560 52492 8628 52548
rect 8684 52492 8752 52548
rect 8808 52492 8876 52548
rect 8932 52492 9000 52548
rect 9056 52492 9124 52548
rect 9180 52492 9248 52548
rect 9304 52492 9372 52548
rect 9428 52492 9496 52548
rect 9552 52492 9620 52548
rect 9676 52492 9744 52548
rect 9800 52492 9810 52548
rect 7874 52424 9810 52492
rect 7874 52368 7884 52424
rect 7940 52368 8008 52424
rect 8064 52368 8132 52424
rect 8188 52368 8256 52424
rect 8312 52368 8380 52424
rect 8436 52368 8504 52424
rect 8560 52368 8628 52424
rect 8684 52368 8752 52424
rect 8808 52368 8876 52424
rect 8932 52368 9000 52424
rect 9056 52368 9124 52424
rect 9180 52368 9248 52424
rect 9304 52368 9372 52424
rect 9428 52368 9496 52424
rect 9552 52368 9620 52424
rect 9676 52368 9744 52424
rect 9800 52368 9810 52424
rect 7874 52300 9810 52368
rect 7874 52244 7884 52300
rect 7940 52244 8008 52300
rect 8064 52244 8132 52300
rect 8188 52244 8256 52300
rect 8312 52244 8380 52300
rect 8436 52244 8504 52300
rect 8560 52244 8628 52300
rect 8684 52244 8752 52300
rect 8808 52244 8876 52300
rect 8932 52244 9000 52300
rect 9056 52244 9124 52300
rect 9180 52244 9248 52300
rect 9304 52244 9372 52300
rect 9428 52244 9496 52300
rect 9552 52244 9620 52300
rect 9676 52244 9744 52300
rect 9800 52244 9810 52300
rect 7874 52176 9810 52244
rect 7874 52120 7884 52176
rect 7940 52120 8008 52176
rect 8064 52120 8132 52176
rect 8188 52120 8256 52176
rect 8312 52120 8380 52176
rect 8436 52120 8504 52176
rect 8560 52120 8628 52176
rect 8684 52120 8752 52176
rect 8808 52120 8876 52176
rect 8932 52120 9000 52176
rect 9056 52120 9124 52176
rect 9180 52120 9248 52176
rect 9304 52120 9372 52176
rect 9428 52120 9496 52176
rect 9552 52120 9620 52176
rect 9676 52120 9744 52176
rect 9800 52120 9810 52176
rect 7874 52052 9810 52120
rect 7874 51996 7884 52052
rect 7940 51996 8008 52052
rect 8064 51996 8132 52052
rect 8188 51996 8256 52052
rect 8312 51996 8380 52052
rect 8436 51996 8504 52052
rect 8560 51996 8628 52052
rect 8684 51996 8752 52052
rect 8808 51996 8876 52052
rect 8932 51996 9000 52052
rect 9056 51996 9124 52052
rect 9180 51996 9248 52052
rect 9304 51996 9372 52052
rect 9428 51996 9496 52052
rect 9552 51996 9620 52052
rect 9676 51996 9744 52052
rect 9800 51996 9810 52052
rect 7874 51928 9810 51996
rect 7874 51872 7884 51928
rect 7940 51872 8008 51928
rect 8064 51872 8132 51928
rect 8188 51872 8256 51928
rect 8312 51872 8380 51928
rect 8436 51872 8504 51928
rect 8560 51872 8628 51928
rect 8684 51872 8752 51928
rect 8808 51872 8876 51928
rect 8932 51872 9000 51928
rect 9056 51872 9124 51928
rect 9180 51872 9248 51928
rect 9304 51872 9372 51928
rect 9428 51872 9496 51928
rect 9552 51872 9620 51928
rect 9676 51872 9744 51928
rect 9800 51872 9810 51928
rect 7874 51804 9810 51872
rect 7874 51748 7884 51804
rect 7940 51748 8008 51804
rect 8064 51748 8132 51804
rect 8188 51748 8256 51804
rect 8312 51748 8380 51804
rect 8436 51748 8504 51804
rect 8560 51748 8628 51804
rect 8684 51748 8752 51804
rect 8808 51748 8876 51804
rect 8932 51748 9000 51804
rect 9056 51748 9124 51804
rect 9180 51748 9248 51804
rect 9304 51748 9372 51804
rect 9428 51748 9496 51804
rect 9552 51748 9620 51804
rect 9676 51748 9744 51804
rect 9800 51748 9810 51804
rect 7874 51680 9810 51748
rect 7874 51624 7884 51680
rect 7940 51624 8008 51680
rect 8064 51624 8132 51680
rect 8188 51624 8256 51680
rect 8312 51624 8380 51680
rect 8436 51624 8504 51680
rect 8560 51624 8628 51680
rect 8684 51624 8752 51680
rect 8808 51624 8876 51680
rect 8932 51624 9000 51680
rect 9056 51624 9124 51680
rect 9180 51624 9248 51680
rect 9304 51624 9372 51680
rect 9428 51624 9496 51680
rect 9552 51624 9620 51680
rect 9676 51624 9744 51680
rect 9800 51624 9810 51680
rect 7874 51556 9810 51624
rect 7874 51500 7884 51556
rect 7940 51500 8008 51556
rect 8064 51500 8132 51556
rect 8188 51500 8256 51556
rect 8312 51500 8380 51556
rect 8436 51500 8504 51556
rect 8560 51500 8628 51556
rect 8684 51500 8752 51556
rect 8808 51500 8876 51556
rect 8932 51500 9000 51556
rect 9056 51500 9124 51556
rect 9180 51500 9248 51556
rect 9304 51500 9372 51556
rect 9428 51500 9496 51556
rect 9552 51500 9620 51556
rect 9676 51500 9744 51556
rect 9800 51500 9810 51556
rect 7874 51432 9810 51500
rect 7874 51376 7884 51432
rect 7940 51376 8008 51432
rect 8064 51376 8132 51432
rect 8188 51376 8256 51432
rect 8312 51376 8380 51432
rect 8436 51376 8504 51432
rect 8560 51376 8628 51432
rect 8684 51376 8752 51432
rect 8808 51376 8876 51432
rect 8932 51376 9000 51432
rect 9056 51376 9124 51432
rect 9180 51376 9248 51432
rect 9304 51376 9372 51432
rect 9428 51376 9496 51432
rect 9552 51376 9620 51432
rect 9676 51376 9744 51432
rect 9800 51376 9810 51432
rect 7874 51308 9810 51376
rect 7874 51252 7884 51308
rect 7940 51252 8008 51308
rect 8064 51252 8132 51308
rect 8188 51252 8256 51308
rect 8312 51252 8380 51308
rect 8436 51252 8504 51308
rect 8560 51252 8628 51308
rect 8684 51252 8752 51308
rect 8808 51252 8876 51308
rect 8932 51252 9000 51308
rect 9056 51252 9124 51308
rect 9180 51252 9248 51308
rect 9304 51252 9372 51308
rect 9428 51252 9496 51308
rect 9552 51252 9620 51308
rect 9676 51252 9744 51308
rect 9800 51252 9810 51308
rect 7874 51242 9810 51252
rect 10244 52548 12180 52558
rect 10244 52492 10254 52548
rect 10310 52492 10378 52548
rect 10434 52492 10502 52548
rect 10558 52492 10626 52548
rect 10682 52492 10750 52548
rect 10806 52492 10874 52548
rect 10930 52492 10998 52548
rect 11054 52492 11122 52548
rect 11178 52492 11246 52548
rect 11302 52492 11370 52548
rect 11426 52492 11494 52548
rect 11550 52492 11618 52548
rect 11674 52492 11742 52548
rect 11798 52492 11866 52548
rect 11922 52492 11990 52548
rect 12046 52492 12114 52548
rect 12170 52492 12180 52548
rect 10244 52424 12180 52492
rect 10244 52368 10254 52424
rect 10310 52368 10378 52424
rect 10434 52368 10502 52424
rect 10558 52368 10626 52424
rect 10682 52368 10750 52424
rect 10806 52368 10874 52424
rect 10930 52368 10998 52424
rect 11054 52368 11122 52424
rect 11178 52368 11246 52424
rect 11302 52368 11370 52424
rect 11426 52368 11494 52424
rect 11550 52368 11618 52424
rect 11674 52368 11742 52424
rect 11798 52368 11866 52424
rect 11922 52368 11990 52424
rect 12046 52368 12114 52424
rect 12170 52368 12180 52424
rect 10244 52300 12180 52368
rect 10244 52244 10254 52300
rect 10310 52244 10378 52300
rect 10434 52244 10502 52300
rect 10558 52244 10626 52300
rect 10682 52244 10750 52300
rect 10806 52244 10874 52300
rect 10930 52244 10998 52300
rect 11054 52244 11122 52300
rect 11178 52244 11246 52300
rect 11302 52244 11370 52300
rect 11426 52244 11494 52300
rect 11550 52244 11618 52300
rect 11674 52244 11742 52300
rect 11798 52244 11866 52300
rect 11922 52244 11990 52300
rect 12046 52244 12114 52300
rect 12170 52244 12180 52300
rect 10244 52176 12180 52244
rect 10244 52120 10254 52176
rect 10310 52120 10378 52176
rect 10434 52120 10502 52176
rect 10558 52120 10626 52176
rect 10682 52120 10750 52176
rect 10806 52120 10874 52176
rect 10930 52120 10998 52176
rect 11054 52120 11122 52176
rect 11178 52120 11246 52176
rect 11302 52120 11370 52176
rect 11426 52120 11494 52176
rect 11550 52120 11618 52176
rect 11674 52120 11742 52176
rect 11798 52120 11866 52176
rect 11922 52120 11990 52176
rect 12046 52120 12114 52176
rect 12170 52120 12180 52176
rect 10244 52052 12180 52120
rect 10244 51996 10254 52052
rect 10310 51996 10378 52052
rect 10434 51996 10502 52052
rect 10558 51996 10626 52052
rect 10682 51996 10750 52052
rect 10806 51996 10874 52052
rect 10930 51996 10998 52052
rect 11054 51996 11122 52052
rect 11178 51996 11246 52052
rect 11302 51996 11370 52052
rect 11426 51996 11494 52052
rect 11550 51996 11618 52052
rect 11674 51996 11742 52052
rect 11798 51996 11866 52052
rect 11922 51996 11990 52052
rect 12046 51996 12114 52052
rect 12170 51996 12180 52052
rect 10244 51928 12180 51996
rect 10244 51872 10254 51928
rect 10310 51872 10378 51928
rect 10434 51872 10502 51928
rect 10558 51872 10626 51928
rect 10682 51872 10750 51928
rect 10806 51872 10874 51928
rect 10930 51872 10998 51928
rect 11054 51872 11122 51928
rect 11178 51872 11246 51928
rect 11302 51872 11370 51928
rect 11426 51872 11494 51928
rect 11550 51872 11618 51928
rect 11674 51872 11742 51928
rect 11798 51872 11866 51928
rect 11922 51872 11990 51928
rect 12046 51872 12114 51928
rect 12170 51872 12180 51928
rect 10244 51804 12180 51872
rect 10244 51748 10254 51804
rect 10310 51748 10378 51804
rect 10434 51748 10502 51804
rect 10558 51748 10626 51804
rect 10682 51748 10750 51804
rect 10806 51748 10874 51804
rect 10930 51748 10998 51804
rect 11054 51748 11122 51804
rect 11178 51748 11246 51804
rect 11302 51748 11370 51804
rect 11426 51748 11494 51804
rect 11550 51748 11618 51804
rect 11674 51748 11742 51804
rect 11798 51748 11866 51804
rect 11922 51748 11990 51804
rect 12046 51748 12114 51804
rect 12170 51748 12180 51804
rect 10244 51680 12180 51748
rect 10244 51624 10254 51680
rect 10310 51624 10378 51680
rect 10434 51624 10502 51680
rect 10558 51624 10626 51680
rect 10682 51624 10750 51680
rect 10806 51624 10874 51680
rect 10930 51624 10998 51680
rect 11054 51624 11122 51680
rect 11178 51624 11246 51680
rect 11302 51624 11370 51680
rect 11426 51624 11494 51680
rect 11550 51624 11618 51680
rect 11674 51624 11742 51680
rect 11798 51624 11866 51680
rect 11922 51624 11990 51680
rect 12046 51624 12114 51680
rect 12170 51624 12180 51680
rect 10244 51556 12180 51624
rect 10244 51500 10254 51556
rect 10310 51500 10378 51556
rect 10434 51500 10502 51556
rect 10558 51500 10626 51556
rect 10682 51500 10750 51556
rect 10806 51500 10874 51556
rect 10930 51500 10998 51556
rect 11054 51500 11122 51556
rect 11178 51500 11246 51556
rect 11302 51500 11370 51556
rect 11426 51500 11494 51556
rect 11550 51500 11618 51556
rect 11674 51500 11742 51556
rect 11798 51500 11866 51556
rect 11922 51500 11990 51556
rect 12046 51500 12114 51556
rect 12170 51500 12180 51556
rect 10244 51432 12180 51500
rect 10244 51376 10254 51432
rect 10310 51376 10378 51432
rect 10434 51376 10502 51432
rect 10558 51376 10626 51432
rect 10682 51376 10750 51432
rect 10806 51376 10874 51432
rect 10930 51376 10998 51432
rect 11054 51376 11122 51432
rect 11178 51376 11246 51432
rect 11302 51376 11370 51432
rect 11426 51376 11494 51432
rect 11550 51376 11618 51432
rect 11674 51376 11742 51432
rect 11798 51376 11866 51432
rect 11922 51376 11990 51432
rect 12046 51376 12114 51432
rect 12170 51376 12180 51432
rect 10244 51308 12180 51376
rect 10244 51252 10254 51308
rect 10310 51252 10378 51308
rect 10434 51252 10502 51308
rect 10558 51252 10626 51308
rect 10682 51252 10750 51308
rect 10806 51252 10874 51308
rect 10930 51252 10998 51308
rect 11054 51252 11122 51308
rect 11178 51252 11246 51308
rect 11302 51252 11370 51308
rect 11426 51252 11494 51308
rect 11550 51252 11618 51308
rect 11674 51252 11742 51308
rect 11798 51252 11866 51308
rect 11922 51252 11990 51308
rect 12046 51252 12114 51308
rect 12170 51252 12180 51308
rect 10244 51242 12180 51252
rect 12861 52548 14673 52558
rect 12861 52492 12871 52548
rect 12927 52492 12995 52548
rect 13051 52492 13119 52548
rect 13175 52492 13243 52548
rect 13299 52492 13367 52548
rect 13423 52492 13491 52548
rect 13547 52492 13615 52548
rect 13671 52492 13739 52548
rect 13795 52492 13863 52548
rect 13919 52492 13987 52548
rect 14043 52492 14111 52548
rect 14167 52492 14235 52548
rect 14291 52492 14359 52548
rect 14415 52492 14483 52548
rect 14539 52492 14607 52548
rect 14663 52492 14673 52548
rect 12861 52424 14673 52492
rect 12861 52368 12871 52424
rect 12927 52368 12995 52424
rect 13051 52368 13119 52424
rect 13175 52368 13243 52424
rect 13299 52368 13367 52424
rect 13423 52368 13491 52424
rect 13547 52368 13615 52424
rect 13671 52368 13739 52424
rect 13795 52368 13863 52424
rect 13919 52368 13987 52424
rect 14043 52368 14111 52424
rect 14167 52368 14235 52424
rect 14291 52368 14359 52424
rect 14415 52368 14483 52424
rect 14539 52368 14607 52424
rect 14663 52368 14673 52424
rect 12861 52300 14673 52368
rect 12861 52244 12871 52300
rect 12927 52244 12995 52300
rect 13051 52244 13119 52300
rect 13175 52244 13243 52300
rect 13299 52244 13367 52300
rect 13423 52244 13491 52300
rect 13547 52244 13615 52300
rect 13671 52244 13739 52300
rect 13795 52244 13863 52300
rect 13919 52244 13987 52300
rect 14043 52244 14111 52300
rect 14167 52244 14235 52300
rect 14291 52244 14359 52300
rect 14415 52244 14483 52300
rect 14539 52244 14607 52300
rect 14663 52244 14673 52300
rect 12861 52176 14673 52244
rect 12861 52120 12871 52176
rect 12927 52120 12995 52176
rect 13051 52120 13119 52176
rect 13175 52120 13243 52176
rect 13299 52120 13367 52176
rect 13423 52120 13491 52176
rect 13547 52120 13615 52176
rect 13671 52120 13739 52176
rect 13795 52120 13863 52176
rect 13919 52120 13987 52176
rect 14043 52120 14111 52176
rect 14167 52120 14235 52176
rect 14291 52120 14359 52176
rect 14415 52120 14483 52176
rect 14539 52120 14607 52176
rect 14663 52120 14673 52176
rect 12861 52052 14673 52120
rect 12861 51996 12871 52052
rect 12927 51996 12995 52052
rect 13051 51996 13119 52052
rect 13175 51996 13243 52052
rect 13299 51996 13367 52052
rect 13423 51996 13491 52052
rect 13547 51996 13615 52052
rect 13671 51996 13739 52052
rect 13795 51996 13863 52052
rect 13919 51996 13987 52052
rect 14043 51996 14111 52052
rect 14167 51996 14235 52052
rect 14291 51996 14359 52052
rect 14415 51996 14483 52052
rect 14539 51996 14607 52052
rect 14663 51996 14673 52052
rect 12861 51928 14673 51996
rect 12861 51872 12871 51928
rect 12927 51872 12995 51928
rect 13051 51872 13119 51928
rect 13175 51872 13243 51928
rect 13299 51872 13367 51928
rect 13423 51872 13491 51928
rect 13547 51872 13615 51928
rect 13671 51872 13739 51928
rect 13795 51872 13863 51928
rect 13919 51872 13987 51928
rect 14043 51872 14111 51928
rect 14167 51872 14235 51928
rect 14291 51872 14359 51928
rect 14415 51872 14483 51928
rect 14539 51872 14607 51928
rect 14663 51872 14673 51928
rect 12861 51804 14673 51872
rect 12861 51748 12871 51804
rect 12927 51748 12995 51804
rect 13051 51748 13119 51804
rect 13175 51748 13243 51804
rect 13299 51748 13367 51804
rect 13423 51748 13491 51804
rect 13547 51748 13615 51804
rect 13671 51748 13739 51804
rect 13795 51748 13863 51804
rect 13919 51748 13987 51804
rect 14043 51748 14111 51804
rect 14167 51748 14235 51804
rect 14291 51748 14359 51804
rect 14415 51748 14483 51804
rect 14539 51748 14607 51804
rect 14663 51748 14673 51804
rect 12861 51680 14673 51748
rect 12861 51624 12871 51680
rect 12927 51624 12995 51680
rect 13051 51624 13119 51680
rect 13175 51624 13243 51680
rect 13299 51624 13367 51680
rect 13423 51624 13491 51680
rect 13547 51624 13615 51680
rect 13671 51624 13739 51680
rect 13795 51624 13863 51680
rect 13919 51624 13987 51680
rect 14043 51624 14111 51680
rect 14167 51624 14235 51680
rect 14291 51624 14359 51680
rect 14415 51624 14483 51680
rect 14539 51624 14607 51680
rect 14663 51624 14673 51680
rect 12861 51556 14673 51624
rect 12861 51500 12871 51556
rect 12927 51500 12995 51556
rect 13051 51500 13119 51556
rect 13175 51500 13243 51556
rect 13299 51500 13367 51556
rect 13423 51500 13491 51556
rect 13547 51500 13615 51556
rect 13671 51500 13739 51556
rect 13795 51500 13863 51556
rect 13919 51500 13987 51556
rect 14043 51500 14111 51556
rect 14167 51500 14235 51556
rect 14291 51500 14359 51556
rect 14415 51500 14483 51556
rect 14539 51500 14607 51556
rect 14663 51500 14673 51556
rect 12861 51432 14673 51500
rect 12861 51376 12871 51432
rect 12927 51376 12995 51432
rect 13051 51376 13119 51432
rect 13175 51376 13243 51432
rect 13299 51376 13367 51432
rect 13423 51376 13491 51432
rect 13547 51376 13615 51432
rect 13671 51376 13739 51432
rect 13795 51376 13863 51432
rect 13919 51376 13987 51432
rect 14043 51376 14111 51432
rect 14167 51376 14235 51432
rect 14291 51376 14359 51432
rect 14415 51376 14483 51432
rect 14539 51376 14607 51432
rect 14663 51376 14673 51432
rect 12861 51308 14673 51376
rect 12861 51252 12871 51308
rect 12927 51252 12995 51308
rect 13051 51252 13119 51308
rect 13175 51252 13243 51308
rect 13299 51252 13367 51308
rect 13423 51252 13491 51308
rect 13547 51252 13615 51308
rect 13671 51252 13739 51308
rect 13795 51252 13863 51308
rect 13919 51252 13987 51308
rect 14043 51252 14111 51308
rect 14167 51252 14235 51308
rect 14291 51252 14359 51308
rect 14415 51252 14483 51308
rect 14539 51252 14607 51308
rect 14663 51252 14673 51308
rect 12861 51242 14673 51252
rect 10 51214 86 51224
rect 14892 51224 14902 52576
rect 14958 51224 14968 52576
rect 14892 51214 14968 51224
rect 2292 50926 2368 50936
rect 2292 50870 2302 50926
rect 2358 50870 2368 50926
rect 2292 50794 2368 50870
rect 2292 50738 2302 50794
rect 2358 50738 2368 50794
rect 2292 50662 2368 50738
rect 2292 50606 2302 50662
rect 2358 50606 2368 50662
rect 2292 50530 2368 50606
rect 2292 50474 2302 50530
rect 2358 50474 2368 50530
rect 2292 50398 2368 50474
rect 2292 50342 2302 50398
rect 2358 50342 2368 50398
rect 2292 50266 2368 50342
rect 2292 50210 2302 50266
rect 2358 50210 2368 50266
rect 2292 50134 2368 50210
rect 2292 50078 2302 50134
rect 2358 50078 2368 50134
rect 2292 50002 2368 50078
rect 2292 49946 2302 50002
rect 2358 49946 2368 50002
rect 2292 49870 2368 49946
rect 2292 49814 2302 49870
rect 2358 49814 2368 49870
rect 2292 49738 2368 49814
rect 2292 49682 2302 49738
rect 2358 49682 2368 49738
rect 2292 49672 2368 49682
rect 10 49376 86 49386
rect 10 48024 20 49376
rect 76 48024 86 49376
rect 14892 49376 14968 49386
rect 305 49348 2117 49358
rect 305 49292 315 49348
rect 371 49292 439 49348
rect 495 49292 563 49348
rect 619 49292 687 49348
rect 743 49292 811 49348
rect 867 49292 935 49348
rect 991 49292 1059 49348
rect 1115 49292 1183 49348
rect 1239 49292 1307 49348
rect 1363 49292 1431 49348
rect 1487 49292 1555 49348
rect 1611 49292 1679 49348
rect 1735 49292 1803 49348
rect 1859 49292 1927 49348
rect 1983 49292 2051 49348
rect 2107 49292 2117 49348
rect 305 49224 2117 49292
rect 305 49168 315 49224
rect 371 49168 439 49224
rect 495 49168 563 49224
rect 619 49168 687 49224
rect 743 49168 811 49224
rect 867 49168 935 49224
rect 991 49168 1059 49224
rect 1115 49168 1183 49224
rect 1239 49168 1307 49224
rect 1363 49168 1431 49224
rect 1487 49168 1555 49224
rect 1611 49168 1679 49224
rect 1735 49168 1803 49224
rect 1859 49168 1927 49224
rect 1983 49168 2051 49224
rect 2107 49168 2117 49224
rect 305 49100 2117 49168
rect 305 49044 315 49100
rect 371 49044 439 49100
rect 495 49044 563 49100
rect 619 49044 687 49100
rect 743 49044 811 49100
rect 867 49044 935 49100
rect 991 49044 1059 49100
rect 1115 49044 1183 49100
rect 1239 49044 1307 49100
rect 1363 49044 1431 49100
rect 1487 49044 1555 49100
rect 1611 49044 1679 49100
rect 1735 49044 1803 49100
rect 1859 49044 1927 49100
rect 1983 49044 2051 49100
rect 2107 49044 2117 49100
rect 305 48976 2117 49044
rect 305 48920 315 48976
rect 371 48920 439 48976
rect 495 48920 563 48976
rect 619 48920 687 48976
rect 743 48920 811 48976
rect 867 48920 935 48976
rect 991 48920 1059 48976
rect 1115 48920 1183 48976
rect 1239 48920 1307 48976
rect 1363 48920 1431 48976
rect 1487 48920 1555 48976
rect 1611 48920 1679 48976
rect 1735 48920 1803 48976
rect 1859 48920 1927 48976
rect 1983 48920 2051 48976
rect 2107 48920 2117 48976
rect 305 48852 2117 48920
rect 305 48796 315 48852
rect 371 48796 439 48852
rect 495 48796 563 48852
rect 619 48796 687 48852
rect 743 48796 811 48852
rect 867 48796 935 48852
rect 991 48796 1059 48852
rect 1115 48796 1183 48852
rect 1239 48796 1307 48852
rect 1363 48796 1431 48852
rect 1487 48796 1555 48852
rect 1611 48796 1679 48852
rect 1735 48796 1803 48852
rect 1859 48796 1927 48852
rect 1983 48796 2051 48852
rect 2107 48796 2117 48852
rect 305 48728 2117 48796
rect 305 48672 315 48728
rect 371 48672 439 48728
rect 495 48672 563 48728
rect 619 48672 687 48728
rect 743 48672 811 48728
rect 867 48672 935 48728
rect 991 48672 1059 48728
rect 1115 48672 1183 48728
rect 1239 48672 1307 48728
rect 1363 48672 1431 48728
rect 1487 48672 1555 48728
rect 1611 48672 1679 48728
rect 1735 48672 1803 48728
rect 1859 48672 1927 48728
rect 1983 48672 2051 48728
rect 2107 48672 2117 48728
rect 305 48604 2117 48672
rect 305 48548 315 48604
rect 371 48548 439 48604
rect 495 48548 563 48604
rect 619 48548 687 48604
rect 743 48548 811 48604
rect 867 48548 935 48604
rect 991 48548 1059 48604
rect 1115 48548 1183 48604
rect 1239 48548 1307 48604
rect 1363 48548 1431 48604
rect 1487 48548 1555 48604
rect 1611 48548 1679 48604
rect 1735 48548 1803 48604
rect 1859 48548 1927 48604
rect 1983 48548 2051 48604
rect 2107 48548 2117 48604
rect 305 48480 2117 48548
rect 305 48424 315 48480
rect 371 48424 439 48480
rect 495 48424 563 48480
rect 619 48424 687 48480
rect 743 48424 811 48480
rect 867 48424 935 48480
rect 991 48424 1059 48480
rect 1115 48424 1183 48480
rect 1239 48424 1307 48480
rect 1363 48424 1431 48480
rect 1487 48424 1555 48480
rect 1611 48424 1679 48480
rect 1735 48424 1803 48480
rect 1859 48424 1927 48480
rect 1983 48424 2051 48480
rect 2107 48424 2117 48480
rect 305 48356 2117 48424
rect 305 48300 315 48356
rect 371 48300 439 48356
rect 495 48300 563 48356
rect 619 48300 687 48356
rect 743 48300 811 48356
rect 867 48300 935 48356
rect 991 48300 1059 48356
rect 1115 48300 1183 48356
rect 1239 48300 1307 48356
rect 1363 48300 1431 48356
rect 1487 48300 1555 48356
rect 1611 48300 1679 48356
rect 1735 48300 1803 48356
rect 1859 48300 1927 48356
rect 1983 48300 2051 48356
rect 2107 48300 2117 48356
rect 305 48232 2117 48300
rect 305 48176 315 48232
rect 371 48176 439 48232
rect 495 48176 563 48232
rect 619 48176 687 48232
rect 743 48176 811 48232
rect 867 48176 935 48232
rect 991 48176 1059 48232
rect 1115 48176 1183 48232
rect 1239 48176 1307 48232
rect 1363 48176 1431 48232
rect 1487 48176 1555 48232
rect 1611 48176 1679 48232
rect 1735 48176 1803 48232
rect 1859 48176 1927 48232
rect 1983 48176 2051 48232
rect 2107 48176 2117 48232
rect 305 48108 2117 48176
rect 305 48052 315 48108
rect 371 48052 439 48108
rect 495 48052 563 48108
rect 619 48052 687 48108
rect 743 48052 811 48108
rect 867 48052 935 48108
rect 991 48052 1059 48108
rect 1115 48052 1183 48108
rect 1239 48052 1307 48108
rect 1363 48052 1431 48108
rect 1487 48052 1555 48108
rect 1611 48052 1679 48108
rect 1735 48052 1803 48108
rect 1859 48052 1927 48108
rect 1983 48052 2051 48108
rect 2107 48052 2117 48108
rect 305 48042 2117 48052
rect 2798 49348 4734 49358
rect 2798 49292 2808 49348
rect 2864 49292 2932 49348
rect 2988 49292 3056 49348
rect 3112 49292 3180 49348
rect 3236 49292 3304 49348
rect 3360 49292 3428 49348
rect 3484 49292 3552 49348
rect 3608 49292 3676 49348
rect 3732 49292 3800 49348
rect 3856 49292 3924 49348
rect 3980 49292 4048 49348
rect 4104 49292 4172 49348
rect 4228 49292 4296 49348
rect 4352 49292 4420 49348
rect 4476 49292 4544 49348
rect 4600 49292 4668 49348
rect 4724 49292 4734 49348
rect 2798 49224 4734 49292
rect 2798 49168 2808 49224
rect 2864 49168 2932 49224
rect 2988 49168 3056 49224
rect 3112 49168 3180 49224
rect 3236 49168 3304 49224
rect 3360 49168 3428 49224
rect 3484 49168 3552 49224
rect 3608 49168 3676 49224
rect 3732 49168 3800 49224
rect 3856 49168 3924 49224
rect 3980 49168 4048 49224
rect 4104 49168 4172 49224
rect 4228 49168 4296 49224
rect 4352 49168 4420 49224
rect 4476 49168 4544 49224
rect 4600 49168 4668 49224
rect 4724 49168 4734 49224
rect 2798 49100 4734 49168
rect 2798 49044 2808 49100
rect 2864 49044 2932 49100
rect 2988 49044 3056 49100
rect 3112 49044 3180 49100
rect 3236 49044 3304 49100
rect 3360 49044 3428 49100
rect 3484 49044 3552 49100
rect 3608 49044 3676 49100
rect 3732 49044 3800 49100
rect 3856 49044 3924 49100
rect 3980 49044 4048 49100
rect 4104 49044 4172 49100
rect 4228 49044 4296 49100
rect 4352 49044 4420 49100
rect 4476 49044 4544 49100
rect 4600 49044 4668 49100
rect 4724 49044 4734 49100
rect 2798 48976 4734 49044
rect 2798 48920 2808 48976
rect 2864 48920 2932 48976
rect 2988 48920 3056 48976
rect 3112 48920 3180 48976
rect 3236 48920 3304 48976
rect 3360 48920 3428 48976
rect 3484 48920 3552 48976
rect 3608 48920 3676 48976
rect 3732 48920 3800 48976
rect 3856 48920 3924 48976
rect 3980 48920 4048 48976
rect 4104 48920 4172 48976
rect 4228 48920 4296 48976
rect 4352 48920 4420 48976
rect 4476 48920 4544 48976
rect 4600 48920 4668 48976
rect 4724 48920 4734 48976
rect 2798 48852 4734 48920
rect 2798 48796 2808 48852
rect 2864 48796 2932 48852
rect 2988 48796 3056 48852
rect 3112 48796 3180 48852
rect 3236 48796 3304 48852
rect 3360 48796 3428 48852
rect 3484 48796 3552 48852
rect 3608 48796 3676 48852
rect 3732 48796 3800 48852
rect 3856 48796 3924 48852
rect 3980 48796 4048 48852
rect 4104 48796 4172 48852
rect 4228 48796 4296 48852
rect 4352 48796 4420 48852
rect 4476 48796 4544 48852
rect 4600 48796 4668 48852
rect 4724 48796 4734 48852
rect 2798 48728 4734 48796
rect 2798 48672 2808 48728
rect 2864 48672 2932 48728
rect 2988 48672 3056 48728
rect 3112 48672 3180 48728
rect 3236 48672 3304 48728
rect 3360 48672 3428 48728
rect 3484 48672 3552 48728
rect 3608 48672 3676 48728
rect 3732 48672 3800 48728
rect 3856 48672 3924 48728
rect 3980 48672 4048 48728
rect 4104 48672 4172 48728
rect 4228 48672 4296 48728
rect 4352 48672 4420 48728
rect 4476 48672 4544 48728
rect 4600 48672 4668 48728
rect 4724 48672 4734 48728
rect 2798 48604 4734 48672
rect 2798 48548 2808 48604
rect 2864 48548 2932 48604
rect 2988 48548 3056 48604
rect 3112 48548 3180 48604
rect 3236 48548 3304 48604
rect 3360 48548 3428 48604
rect 3484 48548 3552 48604
rect 3608 48548 3676 48604
rect 3732 48548 3800 48604
rect 3856 48548 3924 48604
rect 3980 48548 4048 48604
rect 4104 48548 4172 48604
rect 4228 48548 4296 48604
rect 4352 48548 4420 48604
rect 4476 48548 4544 48604
rect 4600 48548 4668 48604
rect 4724 48548 4734 48604
rect 2798 48480 4734 48548
rect 2798 48424 2808 48480
rect 2864 48424 2932 48480
rect 2988 48424 3056 48480
rect 3112 48424 3180 48480
rect 3236 48424 3304 48480
rect 3360 48424 3428 48480
rect 3484 48424 3552 48480
rect 3608 48424 3676 48480
rect 3732 48424 3800 48480
rect 3856 48424 3924 48480
rect 3980 48424 4048 48480
rect 4104 48424 4172 48480
rect 4228 48424 4296 48480
rect 4352 48424 4420 48480
rect 4476 48424 4544 48480
rect 4600 48424 4668 48480
rect 4724 48424 4734 48480
rect 2798 48356 4734 48424
rect 2798 48300 2808 48356
rect 2864 48300 2932 48356
rect 2988 48300 3056 48356
rect 3112 48300 3180 48356
rect 3236 48300 3304 48356
rect 3360 48300 3428 48356
rect 3484 48300 3552 48356
rect 3608 48300 3676 48356
rect 3732 48300 3800 48356
rect 3856 48300 3924 48356
rect 3980 48300 4048 48356
rect 4104 48300 4172 48356
rect 4228 48300 4296 48356
rect 4352 48300 4420 48356
rect 4476 48300 4544 48356
rect 4600 48300 4668 48356
rect 4724 48300 4734 48356
rect 2798 48232 4734 48300
rect 2798 48176 2808 48232
rect 2864 48176 2932 48232
rect 2988 48176 3056 48232
rect 3112 48176 3180 48232
rect 3236 48176 3304 48232
rect 3360 48176 3428 48232
rect 3484 48176 3552 48232
rect 3608 48176 3676 48232
rect 3732 48176 3800 48232
rect 3856 48176 3924 48232
rect 3980 48176 4048 48232
rect 4104 48176 4172 48232
rect 4228 48176 4296 48232
rect 4352 48176 4420 48232
rect 4476 48176 4544 48232
rect 4600 48176 4668 48232
rect 4724 48176 4734 48232
rect 2798 48108 4734 48176
rect 2798 48052 2808 48108
rect 2864 48052 2932 48108
rect 2988 48052 3056 48108
rect 3112 48052 3180 48108
rect 3236 48052 3304 48108
rect 3360 48052 3428 48108
rect 3484 48052 3552 48108
rect 3608 48052 3676 48108
rect 3732 48052 3800 48108
rect 3856 48052 3924 48108
rect 3980 48052 4048 48108
rect 4104 48052 4172 48108
rect 4228 48052 4296 48108
rect 4352 48052 4420 48108
rect 4476 48052 4544 48108
rect 4600 48052 4668 48108
rect 4724 48052 4734 48108
rect 2798 48042 4734 48052
rect 5168 49348 7104 49358
rect 5168 49292 5178 49348
rect 5234 49292 5302 49348
rect 5358 49292 5426 49348
rect 5482 49292 5550 49348
rect 5606 49292 5674 49348
rect 5730 49292 5798 49348
rect 5854 49292 5922 49348
rect 5978 49292 6046 49348
rect 6102 49292 6170 49348
rect 6226 49292 6294 49348
rect 6350 49292 6418 49348
rect 6474 49292 6542 49348
rect 6598 49292 6666 49348
rect 6722 49292 6790 49348
rect 6846 49292 6914 49348
rect 6970 49292 7038 49348
rect 7094 49292 7104 49348
rect 5168 49224 7104 49292
rect 5168 49168 5178 49224
rect 5234 49168 5302 49224
rect 5358 49168 5426 49224
rect 5482 49168 5550 49224
rect 5606 49168 5674 49224
rect 5730 49168 5798 49224
rect 5854 49168 5922 49224
rect 5978 49168 6046 49224
rect 6102 49168 6170 49224
rect 6226 49168 6294 49224
rect 6350 49168 6418 49224
rect 6474 49168 6542 49224
rect 6598 49168 6666 49224
rect 6722 49168 6790 49224
rect 6846 49168 6914 49224
rect 6970 49168 7038 49224
rect 7094 49168 7104 49224
rect 5168 49100 7104 49168
rect 5168 49044 5178 49100
rect 5234 49044 5302 49100
rect 5358 49044 5426 49100
rect 5482 49044 5550 49100
rect 5606 49044 5674 49100
rect 5730 49044 5798 49100
rect 5854 49044 5922 49100
rect 5978 49044 6046 49100
rect 6102 49044 6170 49100
rect 6226 49044 6294 49100
rect 6350 49044 6418 49100
rect 6474 49044 6542 49100
rect 6598 49044 6666 49100
rect 6722 49044 6790 49100
rect 6846 49044 6914 49100
rect 6970 49044 7038 49100
rect 7094 49044 7104 49100
rect 5168 48976 7104 49044
rect 5168 48920 5178 48976
rect 5234 48920 5302 48976
rect 5358 48920 5426 48976
rect 5482 48920 5550 48976
rect 5606 48920 5674 48976
rect 5730 48920 5798 48976
rect 5854 48920 5922 48976
rect 5978 48920 6046 48976
rect 6102 48920 6170 48976
rect 6226 48920 6294 48976
rect 6350 48920 6418 48976
rect 6474 48920 6542 48976
rect 6598 48920 6666 48976
rect 6722 48920 6790 48976
rect 6846 48920 6914 48976
rect 6970 48920 7038 48976
rect 7094 48920 7104 48976
rect 5168 48852 7104 48920
rect 5168 48796 5178 48852
rect 5234 48796 5302 48852
rect 5358 48796 5426 48852
rect 5482 48796 5550 48852
rect 5606 48796 5674 48852
rect 5730 48796 5798 48852
rect 5854 48796 5922 48852
rect 5978 48796 6046 48852
rect 6102 48796 6170 48852
rect 6226 48796 6294 48852
rect 6350 48796 6418 48852
rect 6474 48796 6542 48852
rect 6598 48796 6666 48852
rect 6722 48796 6790 48852
rect 6846 48796 6914 48852
rect 6970 48796 7038 48852
rect 7094 48796 7104 48852
rect 5168 48728 7104 48796
rect 5168 48672 5178 48728
rect 5234 48672 5302 48728
rect 5358 48672 5426 48728
rect 5482 48672 5550 48728
rect 5606 48672 5674 48728
rect 5730 48672 5798 48728
rect 5854 48672 5922 48728
rect 5978 48672 6046 48728
rect 6102 48672 6170 48728
rect 6226 48672 6294 48728
rect 6350 48672 6418 48728
rect 6474 48672 6542 48728
rect 6598 48672 6666 48728
rect 6722 48672 6790 48728
rect 6846 48672 6914 48728
rect 6970 48672 7038 48728
rect 7094 48672 7104 48728
rect 5168 48604 7104 48672
rect 5168 48548 5178 48604
rect 5234 48548 5302 48604
rect 5358 48548 5426 48604
rect 5482 48548 5550 48604
rect 5606 48548 5674 48604
rect 5730 48548 5798 48604
rect 5854 48548 5922 48604
rect 5978 48548 6046 48604
rect 6102 48548 6170 48604
rect 6226 48548 6294 48604
rect 6350 48548 6418 48604
rect 6474 48548 6542 48604
rect 6598 48548 6666 48604
rect 6722 48548 6790 48604
rect 6846 48548 6914 48604
rect 6970 48548 7038 48604
rect 7094 48548 7104 48604
rect 5168 48480 7104 48548
rect 5168 48424 5178 48480
rect 5234 48424 5302 48480
rect 5358 48424 5426 48480
rect 5482 48424 5550 48480
rect 5606 48424 5674 48480
rect 5730 48424 5798 48480
rect 5854 48424 5922 48480
rect 5978 48424 6046 48480
rect 6102 48424 6170 48480
rect 6226 48424 6294 48480
rect 6350 48424 6418 48480
rect 6474 48424 6542 48480
rect 6598 48424 6666 48480
rect 6722 48424 6790 48480
rect 6846 48424 6914 48480
rect 6970 48424 7038 48480
rect 7094 48424 7104 48480
rect 5168 48356 7104 48424
rect 5168 48300 5178 48356
rect 5234 48300 5302 48356
rect 5358 48300 5426 48356
rect 5482 48300 5550 48356
rect 5606 48300 5674 48356
rect 5730 48300 5798 48356
rect 5854 48300 5922 48356
rect 5978 48300 6046 48356
rect 6102 48300 6170 48356
rect 6226 48300 6294 48356
rect 6350 48300 6418 48356
rect 6474 48300 6542 48356
rect 6598 48300 6666 48356
rect 6722 48300 6790 48356
rect 6846 48300 6914 48356
rect 6970 48300 7038 48356
rect 7094 48300 7104 48356
rect 5168 48232 7104 48300
rect 5168 48176 5178 48232
rect 5234 48176 5302 48232
rect 5358 48176 5426 48232
rect 5482 48176 5550 48232
rect 5606 48176 5674 48232
rect 5730 48176 5798 48232
rect 5854 48176 5922 48232
rect 5978 48176 6046 48232
rect 6102 48176 6170 48232
rect 6226 48176 6294 48232
rect 6350 48176 6418 48232
rect 6474 48176 6542 48232
rect 6598 48176 6666 48232
rect 6722 48176 6790 48232
rect 6846 48176 6914 48232
rect 6970 48176 7038 48232
rect 7094 48176 7104 48232
rect 5168 48108 7104 48176
rect 5168 48052 5178 48108
rect 5234 48052 5302 48108
rect 5358 48052 5426 48108
rect 5482 48052 5550 48108
rect 5606 48052 5674 48108
rect 5730 48052 5798 48108
rect 5854 48052 5922 48108
rect 5978 48052 6046 48108
rect 6102 48052 6170 48108
rect 6226 48052 6294 48108
rect 6350 48052 6418 48108
rect 6474 48052 6542 48108
rect 6598 48052 6666 48108
rect 6722 48052 6790 48108
rect 6846 48052 6914 48108
rect 6970 48052 7038 48108
rect 7094 48052 7104 48108
rect 5168 48042 7104 48052
rect 7874 49348 9810 49358
rect 7874 49292 7884 49348
rect 7940 49292 8008 49348
rect 8064 49292 8132 49348
rect 8188 49292 8256 49348
rect 8312 49292 8380 49348
rect 8436 49292 8504 49348
rect 8560 49292 8628 49348
rect 8684 49292 8752 49348
rect 8808 49292 8876 49348
rect 8932 49292 9000 49348
rect 9056 49292 9124 49348
rect 9180 49292 9248 49348
rect 9304 49292 9372 49348
rect 9428 49292 9496 49348
rect 9552 49292 9620 49348
rect 9676 49292 9744 49348
rect 9800 49292 9810 49348
rect 7874 49224 9810 49292
rect 7874 49168 7884 49224
rect 7940 49168 8008 49224
rect 8064 49168 8132 49224
rect 8188 49168 8256 49224
rect 8312 49168 8380 49224
rect 8436 49168 8504 49224
rect 8560 49168 8628 49224
rect 8684 49168 8752 49224
rect 8808 49168 8876 49224
rect 8932 49168 9000 49224
rect 9056 49168 9124 49224
rect 9180 49168 9248 49224
rect 9304 49168 9372 49224
rect 9428 49168 9496 49224
rect 9552 49168 9620 49224
rect 9676 49168 9744 49224
rect 9800 49168 9810 49224
rect 7874 49100 9810 49168
rect 7874 49044 7884 49100
rect 7940 49044 8008 49100
rect 8064 49044 8132 49100
rect 8188 49044 8256 49100
rect 8312 49044 8380 49100
rect 8436 49044 8504 49100
rect 8560 49044 8628 49100
rect 8684 49044 8752 49100
rect 8808 49044 8876 49100
rect 8932 49044 9000 49100
rect 9056 49044 9124 49100
rect 9180 49044 9248 49100
rect 9304 49044 9372 49100
rect 9428 49044 9496 49100
rect 9552 49044 9620 49100
rect 9676 49044 9744 49100
rect 9800 49044 9810 49100
rect 7874 48976 9810 49044
rect 7874 48920 7884 48976
rect 7940 48920 8008 48976
rect 8064 48920 8132 48976
rect 8188 48920 8256 48976
rect 8312 48920 8380 48976
rect 8436 48920 8504 48976
rect 8560 48920 8628 48976
rect 8684 48920 8752 48976
rect 8808 48920 8876 48976
rect 8932 48920 9000 48976
rect 9056 48920 9124 48976
rect 9180 48920 9248 48976
rect 9304 48920 9372 48976
rect 9428 48920 9496 48976
rect 9552 48920 9620 48976
rect 9676 48920 9744 48976
rect 9800 48920 9810 48976
rect 7874 48852 9810 48920
rect 7874 48796 7884 48852
rect 7940 48796 8008 48852
rect 8064 48796 8132 48852
rect 8188 48796 8256 48852
rect 8312 48796 8380 48852
rect 8436 48796 8504 48852
rect 8560 48796 8628 48852
rect 8684 48796 8752 48852
rect 8808 48796 8876 48852
rect 8932 48796 9000 48852
rect 9056 48796 9124 48852
rect 9180 48796 9248 48852
rect 9304 48796 9372 48852
rect 9428 48796 9496 48852
rect 9552 48796 9620 48852
rect 9676 48796 9744 48852
rect 9800 48796 9810 48852
rect 7874 48728 9810 48796
rect 7874 48672 7884 48728
rect 7940 48672 8008 48728
rect 8064 48672 8132 48728
rect 8188 48672 8256 48728
rect 8312 48672 8380 48728
rect 8436 48672 8504 48728
rect 8560 48672 8628 48728
rect 8684 48672 8752 48728
rect 8808 48672 8876 48728
rect 8932 48672 9000 48728
rect 9056 48672 9124 48728
rect 9180 48672 9248 48728
rect 9304 48672 9372 48728
rect 9428 48672 9496 48728
rect 9552 48672 9620 48728
rect 9676 48672 9744 48728
rect 9800 48672 9810 48728
rect 7874 48604 9810 48672
rect 7874 48548 7884 48604
rect 7940 48548 8008 48604
rect 8064 48548 8132 48604
rect 8188 48548 8256 48604
rect 8312 48548 8380 48604
rect 8436 48548 8504 48604
rect 8560 48548 8628 48604
rect 8684 48548 8752 48604
rect 8808 48548 8876 48604
rect 8932 48548 9000 48604
rect 9056 48548 9124 48604
rect 9180 48548 9248 48604
rect 9304 48548 9372 48604
rect 9428 48548 9496 48604
rect 9552 48548 9620 48604
rect 9676 48548 9744 48604
rect 9800 48548 9810 48604
rect 7874 48480 9810 48548
rect 7874 48424 7884 48480
rect 7940 48424 8008 48480
rect 8064 48424 8132 48480
rect 8188 48424 8256 48480
rect 8312 48424 8380 48480
rect 8436 48424 8504 48480
rect 8560 48424 8628 48480
rect 8684 48424 8752 48480
rect 8808 48424 8876 48480
rect 8932 48424 9000 48480
rect 9056 48424 9124 48480
rect 9180 48424 9248 48480
rect 9304 48424 9372 48480
rect 9428 48424 9496 48480
rect 9552 48424 9620 48480
rect 9676 48424 9744 48480
rect 9800 48424 9810 48480
rect 7874 48356 9810 48424
rect 7874 48300 7884 48356
rect 7940 48300 8008 48356
rect 8064 48300 8132 48356
rect 8188 48300 8256 48356
rect 8312 48300 8380 48356
rect 8436 48300 8504 48356
rect 8560 48300 8628 48356
rect 8684 48300 8752 48356
rect 8808 48300 8876 48356
rect 8932 48300 9000 48356
rect 9056 48300 9124 48356
rect 9180 48300 9248 48356
rect 9304 48300 9372 48356
rect 9428 48300 9496 48356
rect 9552 48300 9620 48356
rect 9676 48300 9744 48356
rect 9800 48300 9810 48356
rect 7874 48232 9810 48300
rect 7874 48176 7884 48232
rect 7940 48176 8008 48232
rect 8064 48176 8132 48232
rect 8188 48176 8256 48232
rect 8312 48176 8380 48232
rect 8436 48176 8504 48232
rect 8560 48176 8628 48232
rect 8684 48176 8752 48232
rect 8808 48176 8876 48232
rect 8932 48176 9000 48232
rect 9056 48176 9124 48232
rect 9180 48176 9248 48232
rect 9304 48176 9372 48232
rect 9428 48176 9496 48232
rect 9552 48176 9620 48232
rect 9676 48176 9744 48232
rect 9800 48176 9810 48232
rect 7874 48108 9810 48176
rect 7874 48052 7884 48108
rect 7940 48052 8008 48108
rect 8064 48052 8132 48108
rect 8188 48052 8256 48108
rect 8312 48052 8380 48108
rect 8436 48052 8504 48108
rect 8560 48052 8628 48108
rect 8684 48052 8752 48108
rect 8808 48052 8876 48108
rect 8932 48052 9000 48108
rect 9056 48052 9124 48108
rect 9180 48052 9248 48108
rect 9304 48052 9372 48108
rect 9428 48052 9496 48108
rect 9552 48052 9620 48108
rect 9676 48052 9744 48108
rect 9800 48052 9810 48108
rect 7874 48042 9810 48052
rect 10244 49348 12180 49358
rect 10244 49292 10254 49348
rect 10310 49292 10378 49348
rect 10434 49292 10502 49348
rect 10558 49292 10626 49348
rect 10682 49292 10750 49348
rect 10806 49292 10874 49348
rect 10930 49292 10998 49348
rect 11054 49292 11122 49348
rect 11178 49292 11246 49348
rect 11302 49292 11370 49348
rect 11426 49292 11494 49348
rect 11550 49292 11618 49348
rect 11674 49292 11742 49348
rect 11798 49292 11866 49348
rect 11922 49292 11990 49348
rect 12046 49292 12114 49348
rect 12170 49292 12180 49348
rect 10244 49224 12180 49292
rect 10244 49168 10254 49224
rect 10310 49168 10378 49224
rect 10434 49168 10502 49224
rect 10558 49168 10626 49224
rect 10682 49168 10750 49224
rect 10806 49168 10874 49224
rect 10930 49168 10998 49224
rect 11054 49168 11122 49224
rect 11178 49168 11246 49224
rect 11302 49168 11370 49224
rect 11426 49168 11494 49224
rect 11550 49168 11618 49224
rect 11674 49168 11742 49224
rect 11798 49168 11866 49224
rect 11922 49168 11990 49224
rect 12046 49168 12114 49224
rect 12170 49168 12180 49224
rect 10244 49100 12180 49168
rect 10244 49044 10254 49100
rect 10310 49044 10378 49100
rect 10434 49044 10502 49100
rect 10558 49044 10626 49100
rect 10682 49044 10750 49100
rect 10806 49044 10874 49100
rect 10930 49044 10998 49100
rect 11054 49044 11122 49100
rect 11178 49044 11246 49100
rect 11302 49044 11370 49100
rect 11426 49044 11494 49100
rect 11550 49044 11618 49100
rect 11674 49044 11742 49100
rect 11798 49044 11866 49100
rect 11922 49044 11990 49100
rect 12046 49044 12114 49100
rect 12170 49044 12180 49100
rect 10244 48976 12180 49044
rect 10244 48920 10254 48976
rect 10310 48920 10378 48976
rect 10434 48920 10502 48976
rect 10558 48920 10626 48976
rect 10682 48920 10750 48976
rect 10806 48920 10874 48976
rect 10930 48920 10998 48976
rect 11054 48920 11122 48976
rect 11178 48920 11246 48976
rect 11302 48920 11370 48976
rect 11426 48920 11494 48976
rect 11550 48920 11618 48976
rect 11674 48920 11742 48976
rect 11798 48920 11866 48976
rect 11922 48920 11990 48976
rect 12046 48920 12114 48976
rect 12170 48920 12180 48976
rect 10244 48852 12180 48920
rect 10244 48796 10254 48852
rect 10310 48796 10378 48852
rect 10434 48796 10502 48852
rect 10558 48796 10626 48852
rect 10682 48796 10750 48852
rect 10806 48796 10874 48852
rect 10930 48796 10998 48852
rect 11054 48796 11122 48852
rect 11178 48796 11246 48852
rect 11302 48796 11370 48852
rect 11426 48796 11494 48852
rect 11550 48796 11618 48852
rect 11674 48796 11742 48852
rect 11798 48796 11866 48852
rect 11922 48796 11990 48852
rect 12046 48796 12114 48852
rect 12170 48796 12180 48852
rect 10244 48728 12180 48796
rect 10244 48672 10254 48728
rect 10310 48672 10378 48728
rect 10434 48672 10502 48728
rect 10558 48672 10626 48728
rect 10682 48672 10750 48728
rect 10806 48672 10874 48728
rect 10930 48672 10998 48728
rect 11054 48672 11122 48728
rect 11178 48672 11246 48728
rect 11302 48672 11370 48728
rect 11426 48672 11494 48728
rect 11550 48672 11618 48728
rect 11674 48672 11742 48728
rect 11798 48672 11866 48728
rect 11922 48672 11990 48728
rect 12046 48672 12114 48728
rect 12170 48672 12180 48728
rect 10244 48604 12180 48672
rect 10244 48548 10254 48604
rect 10310 48548 10378 48604
rect 10434 48548 10502 48604
rect 10558 48548 10626 48604
rect 10682 48548 10750 48604
rect 10806 48548 10874 48604
rect 10930 48548 10998 48604
rect 11054 48548 11122 48604
rect 11178 48548 11246 48604
rect 11302 48548 11370 48604
rect 11426 48548 11494 48604
rect 11550 48548 11618 48604
rect 11674 48548 11742 48604
rect 11798 48548 11866 48604
rect 11922 48548 11990 48604
rect 12046 48548 12114 48604
rect 12170 48548 12180 48604
rect 10244 48480 12180 48548
rect 10244 48424 10254 48480
rect 10310 48424 10378 48480
rect 10434 48424 10502 48480
rect 10558 48424 10626 48480
rect 10682 48424 10750 48480
rect 10806 48424 10874 48480
rect 10930 48424 10998 48480
rect 11054 48424 11122 48480
rect 11178 48424 11246 48480
rect 11302 48424 11370 48480
rect 11426 48424 11494 48480
rect 11550 48424 11618 48480
rect 11674 48424 11742 48480
rect 11798 48424 11866 48480
rect 11922 48424 11990 48480
rect 12046 48424 12114 48480
rect 12170 48424 12180 48480
rect 10244 48356 12180 48424
rect 10244 48300 10254 48356
rect 10310 48300 10378 48356
rect 10434 48300 10502 48356
rect 10558 48300 10626 48356
rect 10682 48300 10750 48356
rect 10806 48300 10874 48356
rect 10930 48300 10998 48356
rect 11054 48300 11122 48356
rect 11178 48300 11246 48356
rect 11302 48300 11370 48356
rect 11426 48300 11494 48356
rect 11550 48300 11618 48356
rect 11674 48300 11742 48356
rect 11798 48300 11866 48356
rect 11922 48300 11990 48356
rect 12046 48300 12114 48356
rect 12170 48300 12180 48356
rect 10244 48232 12180 48300
rect 10244 48176 10254 48232
rect 10310 48176 10378 48232
rect 10434 48176 10502 48232
rect 10558 48176 10626 48232
rect 10682 48176 10750 48232
rect 10806 48176 10874 48232
rect 10930 48176 10998 48232
rect 11054 48176 11122 48232
rect 11178 48176 11246 48232
rect 11302 48176 11370 48232
rect 11426 48176 11494 48232
rect 11550 48176 11618 48232
rect 11674 48176 11742 48232
rect 11798 48176 11866 48232
rect 11922 48176 11990 48232
rect 12046 48176 12114 48232
rect 12170 48176 12180 48232
rect 10244 48108 12180 48176
rect 10244 48052 10254 48108
rect 10310 48052 10378 48108
rect 10434 48052 10502 48108
rect 10558 48052 10626 48108
rect 10682 48052 10750 48108
rect 10806 48052 10874 48108
rect 10930 48052 10998 48108
rect 11054 48052 11122 48108
rect 11178 48052 11246 48108
rect 11302 48052 11370 48108
rect 11426 48052 11494 48108
rect 11550 48052 11618 48108
rect 11674 48052 11742 48108
rect 11798 48052 11866 48108
rect 11922 48052 11990 48108
rect 12046 48052 12114 48108
rect 12170 48052 12180 48108
rect 10244 48042 12180 48052
rect 12861 49348 14673 49358
rect 12861 49292 12871 49348
rect 12927 49292 12995 49348
rect 13051 49292 13119 49348
rect 13175 49292 13243 49348
rect 13299 49292 13367 49348
rect 13423 49292 13491 49348
rect 13547 49292 13615 49348
rect 13671 49292 13739 49348
rect 13795 49292 13863 49348
rect 13919 49292 13987 49348
rect 14043 49292 14111 49348
rect 14167 49292 14235 49348
rect 14291 49292 14359 49348
rect 14415 49292 14483 49348
rect 14539 49292 14607 49348
rect 14663 49292 14673 49348
rect 12861 49224 14673 49292
rect 12861 49168 12871 49224
rect 12927 49168 12995 49224
rect 13051 49168 13119 49224
rect 13175 49168 13243 49224
rect 13299 49168 13367 49224
rect 13423 49168 13491 49224
rect 13547 49168 13615 49224
rect 13671 49168 13739 49224
rect 13795 49168 13863 49224
rect 13919 49168 13987 49224
rect 14043 49168 14111 49224
rect 14167 49168 14235 49224
rect 14291 49168 14359 49224
rect 14415 49168 14483 49224
rect 14539 49168 14607 49224
rect 14663 49168 14673 49224
rect 12861 49100 14673 49168
rect 12861 49044 12871 49100
rect 12927 49044 12995 49100
rect 13051 49044 13119 49100
rect 13175 49044 13243 49100
rect 13299 49044 13367 49100
rect 13423 49044 13491 49100
rect 13547 49044 13615 49100
rect 13671 49044 13739 49100
rect 13795 49044 13863 49100
rect 13919 49044 13987 49100
rect 14043 49044 14111 49100
rect 14167 49044 14235 49100
rect 14291 49044 14359 49100
rect 14415 49044 14483 49100
rect 14539 49044 14607 49100
rect 14663 49044 14673 49100
rect 12861 48976 14673 49044
rect 12861 48920 12871 48976
rect 12927 48920 12995 48976
rect 13051 48920 13119 48976
rect 13175 48920 13243 48976
rect 13299 48920 13367 48976
rect 13423 48920 13491 48976
rect 13547 48920 13615 48976
rect 13671 48920 13739 48976
rect 13795 48920 13863 48976
rect 13919 48920 13987 48976
rect 14043 48920 14111 48976
rect 14167 48920 14235 48976
rect 14291 48920 14359 48976
rect 14415 48920 14483 48976
rect 14539 48920 14607 48976
rect 14663 48920 14673 48976
rect 12861 48852 14673 48920
rect 12861 48796 12871 48852
rect 12927 48796 12995 48852
rect 13051 48796 13119 48852
rect 13175 48796 13243 48852
rect 13299 48796 13367 48852
rect 13423 48796 13491 48852
rect 13547 48796 13615 48852
rect 13671 48796 13739 48852
rect 13795 48796 13863 48852
rect 13919 48796 13987 48852
rect 14043 48796 14111 48852
rect 14167 48796 14235 48852
rect 14291 48796 14359 48852
rect 14415 48796 14483 48852
rect 14539 48796 14607 48852
rect 14663 48796 14673 48852
rect 12861 48728 14673 48796
rect 12861 48672 12871 48728
rect 12927 48672 12995 48728
rect 13051 48672 13119 48728
rect 13175 48672 13243 48728
rect 13299 48672 13367 48728
rect 13423 48672 13491 48728
rect 13547 48672 13615 48728
rect 13671 48672 13739 48728
rect 13795 48672 13863 48728
rect 13919 48672 13987 48728
rect 14043 48672 14111 48728
rect 14167 48672 14235 48728
rect 14291 48672 14359 48728
rect 14415 48672 14483 48728
rect 14539 48672 14607 48728
rect 14663 48672 14673 48728
rect 12861 48604 14673 48672
rect 12861 48548 12871 48604
rect 12927 48548 12995 48604
rect 13051 48548 13119 48604
rect 13175 48548 13243 48604
rect 13299 48548 13367 48604
rect 13423 48548 13491 48604
rect 13547 48548 13615 48604
rect 13671 48548 13739 48604
rect 13795 48548 13863 48604
rect 13919 48548 13987 48604
rect 14043 48548 14111 48604
rect 14167 48548 14235 48604
rect 14291 48548 14359 48604
rect 14415 48548 14483 48604
rect 14539 48548 14607 48604
rect 14663 48548 14673 48604
rect 12861 48480 14673 48548
rect 12861 48424 12871 48480
rect 12927 48424 12995 48480
rect 13051 48424 13119 48480
rect 13175 48424 13243 48480
rect 13299 48424 13367 48480
rect 13423 48424 13491 48480
rect 13547 48424 13615 48480
rect 13671 48424 13739 48480
rect 13795 48424 13863 48480
rect 13919 48424 13987 48480
rect 14043 48424 14111 48480
rect 14167 48424 14235 48480
rect 14291 48424 14359 48480
rect 14415 48424 14483 48480
rect 14539 48424 14607 48480
rect 14663 48424 14673 48480
rect 12861 48356 14673 48424
rect 12861 48300 12871 48356
rect 12927 48300 12995 48356
rect 13051 48300 13119 48356
rect 13175 48300 13243 48356
rect 13299 48300 13367 48356
rect 13423 48300 13491 48356
rect 13547 48300 13615 48356
rect 13671 48300 13739 48356
rect 13795 48300 13863 48356
rect 13919 48300 13987 48356
rect 14043 48300 14111 48356
rect 14167 48300 14235 48356
rect 14291 48300 14359 48356
rect 14415 48300 14483 48356
rect 14539 48300 14607 48356
rect 14663 48300 14673 48356
rect 12861 48232 14673 48300
rect 12861 48176 12871 48232
rect 12927 48176 12995 48232
rect 13051 48176 13119 48232
rect 13175 48176 13243 48232
rect 13299 48176 13367 48232
rect 13423 48176 13491 48232
rect 13547 48176 13615 48232
rect 13671 48176 13739 48232
rect 13795 48176 13863 48232
rect 13919 48176 13987 48232
rect 14043 48176 14111 48232
rect 14167 48176 14235 48232
rect 14291 48176 14359 48232
rect 14415 48176 14483 48232
rect 14539 48176 14607 48232
rect 14663 48176 14673 48232
rect 12861 48108 14673 48176
rect 12861 48052 12871 48108
rect 12927 48052 12995 48108
rect 13051 48052 13119 48108
rect 13175 48052 13243 48108
rect 13299 48052 13367 48108
rect 13423 48052 13491 48108
rect 13547 48052 13615 48108
rect 13671 48052 13739 48108
rect 13795 48052 13863 48108
rect 13919 48052 13987 48108
rect 14043 48052 14111 48108
rect 14167 48052 14235 48108
rect 14291 48052 14359 48108
rect 14415 48052 14483 48108
rect 14539 48052 14607 48108
rect 14663 48052 14673 48108
rect 12861 48042 14673 48052
rect 10 48014 86 48024
rect 14892 48024 14902 49376
rect 14958 48024 14968 49376
rect 14892 48014 14968 48024
rect 2481 47748 2681 47758
rect 2481 47692 2491 47748
rect 2547 47692 2615 47748
rect 2671 47692 2681 47748
rect 2481 47624 2681 47692
rect 2481 47568 2491 47624
rect 2547 47568 2615 47624
rect 2671 47568 2681 47624
rect 2481 47500 2681 47568
rect 2481 47444 2491 47500
rect 2547 47444 2615 47500
rect 2671 47444 2681 47500
rect 2481 47376 2681 47444
rect 2481 47320 2491 47376
rect 2547 47320 2615 47376
rect 2671 47320 2681 47376
rect 2481 47252 2681 47320
rect 2481 47196 2491 47252
rect 2547 47196 2615 47252
rect 2671 47196 2681 47252
rect 2481 47128 2681 47196
rect 2481 47072 2491 47128
rect 2547 47072 2615 47128
rect 2671 47072 2681 47128
rect 2481 47004 2681 47072
rect 2481 46948 2491 47004
rect 2547 46948 2615 47004
rect 2671 46948 2681 47004
rect 2481 46880 2681 46948
rect 2481 46824 2491 46880
rect 2547 46824 2615 46880
rect 2671 46824 2681 46880
rect 2481 46756 2681 46824
rect 2481 46700 2491 46756
rect 2547 46700 2615 46756
rect 2671 46700 2681 46756
rect 2481 46632 2681 46700
rect 2481 46576 2491 46632
rect 2547 46576 2615 46632
rect 2671 46576 2681 46632
rect 2481 46508 2681 46576
rect 2481 46452 2491 46508
rect 2547 46452 2615 46508
rect 2671 46452 2681 46508
rect 2481 46442 2681 46452
rect 4851 47748 5051 47758
rect 4851 47692 4861 47748
rect 4917 47692 4985 47748
rect 5041 47692 5051 47748
rect 4851 47624 5051 47692
rect 4851 47568 4861 47624
rect 4917 47568 4985 47624
rect 5041 47568 5051 47624
rect 4851 47500 5051 47568
rect 4851 47444 4861 47500
rect 4917 47444 4985 47500
rect 5041 47444 5051 47500
rect 4851 47376 5051 47444
rect 4851 47320 4861 47376
rect 4917 47320 4985 47376
rect 5041 47320 5051 47376
rect 4851 47252 5051 47320
rect 4851 47196 4861 47252
rect 4917 47196 4985 47252
rect 5041 47196 5051 47252
rect 4851 47128 5051 47196
rect 4851 47072 4861 47128
rect 4917 47072 4985 47128
rect 5041 47072 5051 47128
rect 4851 47004 5051 47072
rect 4851 46948 4861 47004
rect 4917 46948 4985 47004
rect 5041 46948 5051 47004
rect 4851 46880 5051 46948
rect 4851 46824 4861 46880
rect 4917 46824 4985 46880
rect 5041 46824 5051 46880
rect 4851 46756 5051 46824
rect 4851 46700 4861 46756
rect 4917 46700 4985 46756
rect 5041 46700 5051 46756
rect 4851 46632 5051 46700
rect 4851 46576 4861 46632
rect 4917 46576 4985 46632
rect 5041 46576 5051 46632
rect 4851 46508 5051 46576
rect 4851 46452 4861 46508
rect 4917 46452 4985 46508
rect 5041 46452 5051 46508
rect 4851 46442 5051 46452
rect 7265 47748 7713 47758
rect 7265 47692 7275 47748
rect 7331 47692 7399 47748
rect 7455 47692 7523 47748
rect 7579 47692 7647 47748
rect 7703 47692 7713 47748
rect 7265 47624 7713 47692
rect 7265 47568 7275 47624
rect 7331 47568 7399 47624
rect 7455 47568 7523 47624
rect 7579 47568 7647 47624
rect 7703 47568 7713 47624
rect 7265 47500 7713 47568
rect 7265 47444 7275 47500
rect 7331 47444 7399 47500
rect 7455 47444 7523 47500
rect 7579 47444 7647 47500
rect 7703 47444 7713 47500
rect 7265 47376 7713 47444
rect 7265 47320 7275 47376
rect 7331 47320 7399 47376
rect 7455 47320 7523 47376
rect 7579 47320 7647 47376
rect 7703 47320 7713 47376
rect 7265 47252 7713 47320
rect 7265 47196 7275 47252
rect 7331 47196 7399 47252
rect 7455 47196 7523 47252
rect 7579 47196 7647 47252
rect 7703 47196 7713 47252
rect 7265 47128 7713 47196
rect 7265 47072 7275 47128
rect 7331 47072 7399 47128
rect 7455 47072 7523 47128
rect 7579 47072 7647 47128
rect 7703 47072 7713 47128
rect 7265 47004 7713 47072
rect 7265 46948 7275 47004
rect 7331 46948 7399 47004
rect 7455 46948 7523 47004
rect 7579 46948 7647 47004
rect 7703 46948 7713 47004
rect 7265 46880 7713 46948
rect 7265 46824 7275 46880
rect 7331 46824 7399 46880
rect 7455 46824 7523 46880
rect 7579 46824 7647 46880
rect 7703 46824 7713 46880
rect 7265 46756 7713 46824
rect 7265 46700 7275 46756
rect 7331 46700 7399 46756
rect 7455 46700 7523 46756
rect 7579 46700 7647 46756
rect 7703 46700 7713 46756
rect 7265 46632 7713 46700
rect 7265 46576 7275 46632
rect 7331 46576 7399 46632
rect 7455 46576 7523 46632
rect 7579 46576 7647 46632
rect 7703 46576 7713 46632
rect 7265 46508 7713 46576
rect 7265 46452 7275 46508
rect 7331 46452 7399 46508
rect 7455 46452 7523 46508
rect 7579 46452 7647 46508
rect 7703 46452 7713 46508
rect 7265 46442 7713 46452
rect 9927 47748 10127 47758
rect 9927 47692 9937 47748
rect 9993 47692 10061 47748
rect 10117 47692 10127 47748
rect 9927 47624 10127 47692
rect 9927 47568 9937 47624
rect 9993 47568 10061 47624
rect 10117 47568 10127 47624
rect 9927 47500 10127 47568
rect 9927 47444 9937 47500
rect 9993 47444 10061 47500
rect 10117 47444 10127 47500
rect 9927 47376 10127 47444
rect 9927 47320 9937 47376
rect 9993 47320 10061 47376
rect 10117 47320 10127 47376
rect 9927 47252 10127 47320
rect 9927 47196 9937 47252
rect 9993 47196 10061 47252
rect 10117 47196 10127 47252
rect 9927 47128 10127 47196
rect 9927 47072 9937 47128
rect 9993 47072 10061 47128
rect 10117 47072 10127 47128
rect 9927 47004 10127 47072
rect 9927 46948 9937 47004
rect 9993 46948 10061 47004
rect 10117 46948 10127 47004
rect 9927 46880 10127 46948
rect 9927 46824 9937 46880
rect 9993 46824 10061 46880
rect 10117 46824 10127 46880
rect 9927 46756 10127 46824
rect 9927 46700 9937 46756
rect 9993 46700 10061 46756
rect 10117 46700 10127 46756
rect 9927 46632 10127 46700
rect 9927 46576 9937 46632
rect 9993 46576 10061 46632
rect 10117 46576 10127 46632
rect 9927 46508 10127 46576
rect 9927 46452 9937 46508
rect 9993 46452 10061 46508
rect 10117 46452 10127 46508
rect 9927 46442 10127 46452
rect 12297 47748 12497 47758
rect 12297 47692 12307 47748
rect 12363 47692 12431 47748
rect 12487 47692 12497 47748
rect 12297 47624 12497 47692
rect 12297 47568 12307 47624
rect 12363 47568 12431 47624
rect 12487 47568 12497 47624
rect 12297 47500 12497 47568
rect 12297 47444 12307 47500
rect 12363 47444 12431 47500
rect 12487 47444 12497 47500
rect 12297 47376 12497 47444
rect 12297 47320 12307 47376
rect 12363 47320 12431 47376
rect 12487 47320 12497 47376
rect 12297 47252 12497 47320
rect 12297 47196 12307 47252
rect 12363 47196 12431 47252
rect 12487 47196 12497 47252
rect 12297 47128 12497 47196
rect 12297 47072 12307 47128
rect 12363 47072 12431 47128
rect 12487 47072 12497 47128
rect 12297 47004 12497 47072
rect 12297 46948 12307 47004
rect 12363 46948 12431 47004
rect 12487 46948 12497 47004
rect 12297 46880 12497 46948
rect 12297 46824 12307 46880
rect 12363 46824 12431 46880
rect 12487 46824 12497 46880
rect 12297 46756 12497 46824
rect 12297 46700 12307 46756
rect 12363 46700 12431 46756
rect 12487 46700 12497 46756
rect 12297 46632 12497 46700
rect 12297 46576 12307 46632
rect 12363 46576 12431 46632
rect 12487 46576 12497 46632
rect 12297 46508 12497 46576
rect 12297 46452 12307 46508
rect 12363 46452 12431 46508
rect 12487 46452 12497 46508
rect 12297 46442 12497 46452
rect 10 46176 86 46186
rect 10 44824 20 46176
rect 76 44824 86 46176
rect 14892 46176 14968 46186
rect 305 46148 2117 46158
rect 305 46092 315 46148
rect 371 46092 439 46148
rect 495 46092 563 46148
rect 619 46092 687 46148
rect 743 46092 811 46148
rect 867 46092 935 46148
rect 991 46092 1059 46148
rect 1115 46092 1183 46148
rect 1239 46092 1307 46148
rect 1363 46092 1431 46148
rect 1487 46092 1555 46148
rect 1611 46092 1679 46148
rect 1735 46092 1803 46148
rect 1859 46092 1927 46148
rect 1983 46092 2051 46148
rect 2107 46092 2117 46148
rect 305 46024 2117 46092
rect 305 45968 315 46024
rect 371 45968 439 46024
rect 495 45968 563 46024
rect 619 45968 687 46024
rect 743 45968 811 46024
rect 867 45968 935 46024
rect 991 45968 1059 46024
rect 1115 45968 1183 46024
rect 1239 45968 1307 46024
rect 1363 45968 1431 46024
rect 1487 45968 1555 46024
rect 1611 45968 1679 46024
rect 1735 45968 1803 46024
rect 1859 45968 1927 46024
rect 1983 45968 2051 46024
rect 2107 45968 2117 46024
rect 305 45900 2117 45968
rect 305 45844 315 45900
rect 371 45844 439 45900
rect 495 45844 563 45900
rect 619 45844 687 45900
rect 743 45844 811 45900
rect 867 45844 935 45900
rect 991 45844 1059 45900
rect 1115 45844 1183 45900
rect 1239 45844 1307 45900
rect 1363 45844 1431 45900
rect 1487 45844 1555 45900
rect 1611 45844 1679 45900
rect 1735 45844 1803 45900
rect 1859 45844 1927 45900
rect 1983 45844 2051 45900
rect 2107 45844 2117 45900
rect 305 45776 2117 45844
rect 305 45720 315 45776
rect 371 45720 439 45776
rect 495 45720 563 45776
rect 619 45720 687 45776
rect 743 45720 811 45776
rect 867 45720 935 45776
rect 991 45720 1059 45776
rect 1115 45720 1183 45776
rect 1239 45720 1307 45776
rect 1363 45720 1431 45776
rect 1487 45720 1555 45776
rect 1611 45720 1679 45776
rect 1735 45720 1803 45776
rect 1859 45720 1927 45776
rect 1983 45720 2051 45776
rect 2107 45720 2117 45776
rect 305 45652 2117 45720
rect 305 45596 315 45652
rect 371 45596 439 45652
rect 495 45596 563 45652
rect 619 45596 687 45652
rect 743 45596 811 45652
rect 867 45596 935 45652
rect 991 45596 1059 45652
rect 1115 45596 1183 45652
rect 1239 45596 1307 45652
rect 1363 45596 1431 45652
rect 1487 45596 1555 45652
rect 1611 45596 1679 45652
rect 1735 45596 1803 45652
rect 1859 45596 1927 45652
rect 1983 45596 2051 45652
rect 2107 45596 2117 45652
rect 305 45528 2117 45596
rect 305 45472 315 45528
rect 371 45472 439 45528
rect 495 45472 563 45528
rect 619 45472 687 45528
rect 743 45472 811 45528
rect 867 45472 935 45528
rect 991 45472 1059 45528
rect 1115 45472 1183 45528
rect 1239 45472 1307 45528
rect 1363 45472 1431 45528
rect 1487 45472 1555 45528
rect 1611 45472 1679 45528
rect 1735 45472 1803 45528
rect 1859 45472 1927 45528
rect 1983 45472 2051 45528
rect 2107 45472 2117 45528
rect 305 45404 2117 45472
rect 305 45348 315 45404
rect 371 45348 439 45404
rect 495 45348 563 45404
rect 619 45348 687 45404
rect 743 45348 811 45404
rect 867 45348 935 45404
rect 991 45348 1059 45404
rect 1115 45348 1183 45404
rect 1239 45348 1307 45404
rect 1363 45348 1431 45404
rect 1487 45348 1555 45404
rect 1611 45348 1679 45404
rect 1735 45348 1803 45404
rect 1859 45348 1927 45404
rect 1983 45348 2051 45404
rect 2107 45348 2117 45404
rect 305 45280 2117 45348
rect 305 45224 315 45280
rect 371 45224 439 45280
rect 495 45224 563 45280
rect 619 45224 687 45280
rect 743 45224 811 45280
rect 867 45224 935 45280
rect 991 45224 1059 45280
rect 1115 45224 1183 45280
rect 1239 45224 1307 45280
rect 1363 45224 1431 45280
rect 1487 45224 1555 45280
rect 1611 45224 1679 45280
rect 1735 45224 1803 45280
rect 1859 45224 1927 45280
rect 1983 45224 2051 45280
rect 2107 45224 2117 45280
rect 305 45156 2117 45224
rect 305 45100 315 45156
rect 371 45100 439 45156
rect 495 45100 563 45156
rect 619 45100 687 45156
rect 743 45100 811 45156
rect 867 45100 935 45156
rect 991 45100 1059 45156
rect 1115 45100 1183 45156
rect 1239 45100 1307 45156
rect 1363 45100 1431 45156
rect 1487 45100 1555 45156
rect 1611 45100 1679 45156
rect 1735 45100 1803 45156
rect 1859 45100 1927 45156
rect 1983 45100 2051 45156
rect 2107 45100 2117 45156
rect 305 45032 2117 45100
rect 305 44976 315 45032
rect 371 44976 439 45032
rect 495 44976 563 45032
rect 619 44976 687 45032
rect 743 44976 811 45032
rect 867 44976 935 45032
rect 991 44976 1059 45032
rect 1115 44976 1183 45032
rect 1239 44976 1307 45032
rect 1363 44976 1431 45032
rect 1487 44976 1555 45032
rect 1611 44976 1679 45032
rect 1735 44976 1803 45032
rect 1859 44976 1927 45032
rect 1983 44976 2051 45032
rect 2107 44976 2117 45032
rect 305 44908 2117 44976
rect 305 44852 315 44908
rect 371 44852 439 44908
rect 495 44852 563 44908
rect 619 44852 687 44908
rect 743 44852 811 44908
rect 867 44852 935 44908
rect 991 44852 1059 44908
rect 1115 44852 1183 44908
rect 1239 44852 1307 44908
rect 1363 44852 1431 44908
rect 1487 44852 1555 44908
rect 1611 44852 1679 44908
rect 1735 44852 1803 44908
rect 1859 44852 1927 44908
rect 1983 44852 2051 44908
rect 2107 44852 2117 44908
rect 305 44842 2117 44852
rect 2798 46148 4734 46158
rect 2798 46092 2808 46148
rect 2864 46092 2932 46148
rect 2988 46092 3056 46148
rect 3112 46092 3180 46148
rect 3236 46092 3304 46148
rect 3360 46092 3428 46148
rect 3484 46092 3552 46148
rect 3608 46092 3676 46148
rect 3732 46092 3800 46148
rect 3856 46092 3924 46148
rect 3980 46092 4048 46148
rect 4104 46092 4172 46148
rect 4228 46092 4296 46148
rect 4352 46092 4420 46148
rect 4476 46092 4544 46148
rect 4600 46092 4668 46148
rect 4724 46092 4734 46148
rect 2798 46024 4734 46092
rect 2798 45968 2808 46024
rect 2864 45968 2932 46024
rect 2988 45968 3056 46024
rect 3112 45968 3180 46024
rect 3236 45968 3304 46024
rect 3360 45968 3428 46024
rect 3484 45968 3552 46024
rect 3608 45968 3676 46024
rect 3732 45968 3800 46024
rect 3856 45968 3924 46024
rect 3980 45968 4048 46024
rect 4104 45968 4172 46024
rect 4228 45968 4296 46024
rect 4352 45968 4420 46024
rect 4476 45968 4544 46024
rect 4600 45968 4668 46024
rect 4724 45968 4734 46024
rect 2798 45900 4734 45968
rect 2798 45844 2808 45900
rect 2864 45844 2932 45900
rect 2988 45844 3056 45900
rect 3112 45844 3180 45900
rect 3236 45844 3304 45900
rect 3360 45844 3428 45900
rect 3484 45844 3552 45900
rect 3608 45844 3676 45900
rect 3732 45844 3800 45900
rect 3856 45844 3924 45900
rect 3980 45844 4048 45900
rect 4104 45844 4172 45900
rect 4228 45844 4296 45900
rect 4352 45844 4420 45900
rect 4476 45844 4544 45900
rect 4600 45844 4668 45900
rect 4724 45844 4734 45900
rect 2798 45776 4734 45844
rect 2798 45720 2808 45776
rect 2864 45720 2932 45776
rect 2988 45720 3056 45776
rect 3112 45720 3180 45776
rect 3236 45720 3304 45776
rect 3360 45720 3428 45776
rect 3484 45720 3552 45776
rect 3608 45720 3676 45776
rect 3732 45720 3800 45776
rect 3856 45720 3924 45776
rect 3980 45720 4048 45776
rect 4104 45720 4172 45776
rect 4228 45720 4296 45776
rect 4352 45720 4420 45776
rect 4476 45720 4544 45776
rect 4600 45720 4668 45776
rect 4724 45720 4734 45776
rect 2798 45652 4734 45720
rect 2798 45596 2808 45652
rect 2864 45596 2932 45652
rect 2988 45596 3056 45652
rect 3112 45596 3180 45652
rect 3236 45596 3304 45652
rect 3360 45596 3428 45652
rect 3484 45596 3552 45652
rect 3608 45596 3676 45652
rect 3732 45596 3800 45652
rect 3856 45596 3924 45652
rect 3980 45596 4048 45652
rect 4104 45596 4172 45652
rect 4228 45596 4296 45652
rect 4352 45596 4420 45652
rect 4476 45596 4544 45652
rect 4600 45596 4668 45652
rect 4724 45596 4734 45652
rect 2798 45528 4734 45596
rect 2798 45472 2808 45528
rect 2864 45472 2932 45528
rect 2988 45472 3056 45528
rect 3112 45472 3180 45528
rect 3236 45472 3304 45528
rect 3360 45472 3428 45528
rect 3484 45472 3552 45528
rect 3608 45472 3676 45528
rect 3732 45472 3800 45528
rect 3856 45472 3924 45528
rect 3980 45472 4048 45528
rect 4104 45472 4172 45528
rect 4228 45472 4296 45528
rect 4352 45472 4420 45528
rect 4476 45472 4544 45528
rect 4600 45472 4668 45528
rect 4724 45472 4734 45528
rect 2798 45404 4734 45472
rect 2798 45348 2808 45404
rect 2864 45348 2932 45404
rect 2988 45348 3056 45404
rect 3112 45348 3180 45404
rect 3236 45348 3304 45404
rect 3360 45348 3428 45404
rect 3484 45348 3552 45404
rect 3608 45348 3676 45404
rect 3732 45348 3800 45404
rect 3856 45348 3924 45404
rect 3980 45348 4048 45404
rect 4104 45348 4172 45404
rect 4228 45348 4296 45404
rect 4352 45348 4420 45404
rect 4476 45348 4544 45404
rect 4600 45348 4668 45404
rect 4724 45348 4734 45404
rect 2798 45280 4734 45348
rect 2798 45224 2808 45280
rect 2864 45224 2932 45280
rect 2988 45224 3056 45280
rect 3112 45224 3180 45280
rect 3236 45224 3304 45280
rect 3360 45224 3428 45280
rect 3484 45224 3552 45280
rect 3608 45224 3676 45280
rect 3732 45224 3800 45280
rect 3856 45224 3924 45280
rect 3980 45224 4048 45280
rect 4104 45224 4172 45280
rect 4228 45224 4296 45280
rect 4352 45224 4420 45280
rect 4476 45224 4544 45280
rect 4600 45224 4668 45280
rect 4724 45224 4734 45280
rect 2798 45156 4734 45224
rect 2798 45100 2808 45156
rect 2864 45100 2932 45156
rect 2988 45100 3056 45156
rect 3112 45100 3180 45156
rect 3236 45100 3304 45156
rect 3360 45100 3428 45156
rect 3484 45100 3552 45156
rect 3608 45100 3676 45156
rect 3732 45100 3800 45156
rect 3856 45100 3924 45156
rect 3980 45100 4048 45156
rect 4104 45100 4172 45156
rect 4228 45100 4296 45156
rect 4352 45100 4420 45156
rect 4476 45100 4544 45156
rect 4600 45100 4668 45156
rect 4724 45100 4734 45156
rect 2798 45032 4734 45100
rect 2798 44976 2808 45032
rect 2864 44976 2932 45032
rect 2988 44976 3056 45032
rect 3112 44976 3180 45032
rect 3236 44976 3304 45032
rect 3360 44976 3428 45032
rect 3484 44976 3552 45032
rect 3608 44976 3676 45032
rect 3732 44976 3800 45032
rect 3856 44976 3924 45032
rect 3980 44976 4048 45032
rect 4104 44976 4172 45032
rect 4228 44976 4296 45032
rect 4352 44976 4420 45032
rect 4476 44976 4544 45032
rect 4600 44976 4668 45032
rect 4724 44976 4734 45032
rect 2798 44908 4734 44976
rect 2798 44852 2808 44908
rect 2864 44852 2932 44908
rect 2988 44852 3056 44908
rect 3112 44852 3180 44908
rect 3236 44852 3304 44908
rect 3360 44852 3428 44908
rect 3484 44852 3552 44908
rect 3608 44852 3676 44908
rect 3732 44852 3800 44908
rect 3856 44852 3924 44908
rect 3980 44852 4048 44908
rect 4104 44852 4172 44908
rect 4228 44852 4296 44908
rect 4352 44852 4420 44908
rect 4476 44852 4544 44908
rect 4600 44852 4668 44908
rect 4724 44852 4734 44908
rect 2798 44842 4734 44852
rect 5168 46148 7104 46158
rect 5168 46092 5178 46148
rect 5234 46092 5302 46148
rect 5358 46092 5426 46148
rect 5482 46092 5550 46148
rect 5606 46092 5674 46148
rect 5730 46092 5798 46148
rect 5854 46092 5922 46148
rect 5978 46092 6046 46148
rect 6102 46092 6170 46148
rect 6226 46092 6294 46148
rect 6350 46092 6418 46148
rect 6474 46092 6542 46148
rect 6598 46092 6666 46148
rect 6722 46092 6790 46148
rect 6846 46092 6914 46148
rect 6970 46092 7038 46148
rect 7094 46092 7104 46148
rect 5168 46024 7104 46092
rect 5168 45968 5178 46024
rect 5234 45968 5302 46024
rect 5358 45968 5426 46024
rect 5482 45968 5550 46024
rect 5606 45968 5674 46024
rect 5730 45968 5798 46024
rect 5854 45968 5922 46024
rect 5978 45968 6046 46024
rect 6102 45968 6170 46024
rect 6226 45968 6294 46024
rect 6350 45968 6418 46024
rect 6474 45968 6542 46024
rect 6598 45968 6666 46024
rect 6722 45968 6790 46024
rect 6846 45968 6914 46024
rect 6970 45968 7038 46024
rect 7094 45968 7104 46024
rect 5168 45900 7104 45968
rect 5168 45844 5178 45900
rect 5234 45844 5302 45900
rect 5358 45844 5426 45900
rect 5482 45844 5550 45900
rect 5606 45844 5674 45900
rect 5730 45844 5798 45900
rect 5854 45844 5922 45900
rect 5978 45844 6046 45900
rect 6102 45844 6170 45900
rect 6226 45844 6294 45900
rect 6350 45844 6418 45900
rect 6474 45844 6542 45900
rect 6598 45844 6666 45900
rect 6722 45844 6790 45900
rect 6846 45844 6914 45900
rect 6970 45844 7038 45900
rect 7094 45844 7104 45900
rect 5168 45776 7104 45844
rect 5168 45720 5178 45776
rect 5234 45720 5302 45776
rect 5358 45720 5426 45776
rect 5482 45720 5550 45776
rect 5606 45720 5674 45776
rect 5730 45720 5798 45776
rect 5854 45720 5922 45776
rect 5978 45720 6046 45776
rect 6102 45720 6170 45776
rect 6226 45720 6294 45776
rect 6350 45720 6418 45776
rect 6474 45720 6542 45776
rect 6598 45720 6666 45776
rect 6722 45720 6790 45776
rect 6846 45720 6914 45776
rect 6970 45720 7038 45776
rect 7094 45720 7104 45776
rect 5168 45652 7104 45720
rect 5168 45596 5178 45652
rect 5234 45596 5302 45652
rect 5358 45596 5426 45652
rect 5482 45596 5550 45652
rect 5606 45596 5674 45652
rect 5730 45596 5798 45652
rect 5854 45596 5922 45652
rect 5978 45596 6046 45652
rect 6102 45596 6170 45652
rect 6226 45596 6294 45652
rect 6350 45596 6418 45652
rect 6474 45596 6542 45652
rect 6598 45596 6666 45652
rect 6722 45596 6790 45652
rect 6846 45596 6914 45652
rect 6970 45596 7038 45652
rect 7094 45596 7104 45652
rect 5168 45528 7104 45596
rect 5168 45472 5178 45528
rect 5234 45472 5302 45528
rect 5358 45472 5426 45528
rect 5482 45472 5550 45528
rect 5606 45472 5674 45528
rect 5730 45472 5798 45528
rect 5854 45472 5922 45528
rect 5978 45472 6046 45528
rect 6102 45472 6170 45528
rect 6226 45472 6294 45528
rect 6350 45472 6418 45528
rect 6474 45472 6542 45528
rect 6598 45472 6666 45528
rect 6722 45472 6790 45528
rect 6846 45472 6914 45528
rect 6970 45472 7038 45528
rect 7094 45472 7104 45528
rect 5168 45404 7104 45472
rect 5168 45348 5178 45404
rect 5234 45348 5302 45404
rect 5358 45348 5426 45404
rect 5482 45348 5550 45404
rect 5606 45348 5674 45404
rect 5730 45348 5798 45404
rect 5854 45348 5922 45404
rect 5978 45348 6046 45404
rect 6102 45348 6170 45404
rect 6226 45348 6294 45404
rect 6350 45348 6418 45404
rect 6474 45348 6542 45404
rect 6598 45348 6666 45404
rect 6722 45348 6790 45404
rect 6846 45348 6914 45404
rect 6970 45348 7038 45404
rect 7094 45348 7104 45404
rect 5168 45280 7104 45348
rect 5168 45224 5178 45280
rect 5234 45224 5302 45280
rect 5358 45224 5426 45280
rect 5482 45224 5550 45280
rect 5606 45224 5674 45280
rect 5730 45224 5798 45280
rect 5854 45224 5922 45280
rect 5978 45224 6046 45280
rect 6102 45224 6170 45280
rect 6226 45224 6294 45280
rect 6350 45224 6418 45280
rect 6474 45224 6542 45280
rect 6598 45224 6666 45280
rect 6722 45224 6790 45280
rect 6846 45224 6914 45280
rect 6970 45224 7038 45280
rect 7094 45224 7104 45280
rect 5168 45156 7104 45224
rect 5168 45100 5178 45156
rect 5234 45100 5302 45156
rect 5358 45100 5426 45156
rect 5482 45100 5550 45156
rect 5606 45100 5674 45156
rect 5730 45100 5798 45156
rect 5854 45100 5922 45156
rect 5978 45100 6046 45156
rect 6102 45100 6170 45156
rect 6226 45100 6294 45156
rect 6350 45100 6418 45156
rect 6474 45100 6542 45156
rect 6598 45100 6666 45156
rect 6722 45100 6790 45156
rect 6846 45100 6914 45156
rect 6970 45100 7038 45156
rect 7094 45100 7104 45156
rect 5168 45032 7104 45100
rect 5168 44976 5178 45032
rect 5234 44976 5302 45032
rect 5358 44976 5426 45032
rect 5482 44976 5550 45032
rect 5606 44976 5674 45032
rect 5730 44976 5798 45032
rect 5854 44976 5922 45032
rect 5978 44976 6046 45032
rect 6102 44976 6170 45032
rect 6226 44976 6294 45032
rect 6350 44976 6418 45032
rect 6474 44976 6542 45032
rect 6598 44976 6666 45032
rect 6722 44976 6790 45032
rect 6846 44976 6914 45032
rect 6970 44976 7038 45032
rect 7094 44976 7104 45032
rect 5168 44908 7104 44976
rect 5168 44852 5178 44908
rect 5234 44852 5302 44908
rect 5358 44852 5426 44908
rect 5482 44852 5550 44908
rect 5606 44852 5674 44908
rect 5730 44852 5798 44908
rect 5854 44852 5922 44908
rect 5978 44852 6046 44908
rect 6102 44852 6170 44908
rect 6226 44852 6294 44908
rect 6350 44852 6418 44908
rect 6474 44852 6542 44908
rect 6598 44852 6666 44908
rect 6722 44852 6790 44908
rect 6846 44852 6914 44908
rect 6970 44852 7038 44908
rect 7094 44852 7104 44908
rect 5168 44842 7104 44852
rect 7874 46148 9810 46158
rect 7874 46092 7884 46148
rect 7940 46092 8008 46148
rect 8064 46092 8132 46148
rect 8188 46092 8256 46148
rect 8312 46092 8380 46148
rect 8436 46092 8504 46148
rect 8560 46092 8628 46148
rect 8684 46092 8752 46148
rect 8808 46092 8876 46148
rect 8932 46092 9000 46148
rect 9056 46092 9124 46148
rect 9180 46092 9248 46148
rect 9304 46092 9372 46148
rect 9428 46092 9496 46148
rect 9552 46092 9620 46148
rect 9676 46092 9744 46148
rect 9800 46092 9810 46148
rect 7874 46024 9810 46092
rect 7874 45968 7884 46024
rect 7940 45968 8008 46024
rect 8064 45968 8132 46024
rect 8188 45968 8256 46024
rect 8312 45968 8380 46024
rect 8436 45968 8504 46024
rect 8560 45968 8628 46024
rect 8684 45968 8752 46024
rect 8808 45968 8876 46024
rect 8932 45968 9000 46024
rect 9056 45968 9124 46024
rect 9180 45968 9248 46024
rect 9304 45968 9372 46024
rect 9428 45968 9496 46024
rect 9552 45968 9620 46024
rect 9676 45968 9744 46024
rect 9800 45968 9810 46024
rect 7874 45900 9810 45968
rect 7874 45844 7884 45900
rect 7940 45844 8008 45900
rect 8064 45844 8132 45900
rect 8188 45844 8256 45900
rect 8312 45844 8380 45900
rect 8436 45844 8504 45900
rect 8560 45844 8628 45900
rect 8684 45844 8752 45900
rect 8808 45844 8876 45900
rect 8932 45844 9000 45900
rect 9056 45844 9124 45900
rect 9180 45844 9248 45900
rect 9304 45844 9372 45900
rect 9428 45844 9496 45900
rect 9552 45844 9620 45900
rect 9676 45844 9744 45900
rect 9800 45844 9810 45900
rect 7874 45776 9810 45844
rect 7874 45720 7884 45776
rect 7940 45720 8008 45776
rect 8064 45720 8132 45776
rect 8188 45720 8256 45776
rect 8312 45720 8380 45776
rect 8436 45720 8504 45776
rect 8560 45720 8628 45776
rect 8684 45720 8752 45776
rect 8808 45720 8876 45776
rect 8932 45720 9000 45776
rect 9056 45720 9124 45776
rect 9180 45720 9248 45776
rect 9304 45720 9372 45776
rect 9428 45720 9496 45776
rect 9552 45720 9620 45776
rect 9676 45720 9744 45776
rect 9800 45720 9810 45776
rect 7874 45652 9810 45720
rect 7874 45596 7884 45652
rect 7940 45596 8008 45652
rect 8064 45596 8132 45652
rect 8188 45596 8256 45652
rect 8312 45596 8380 45652
rect 8436 45596 8504 45652
rect 8560 45596 8628 45652
rect 8684 45596 8752 45652
rect 8808 45596 8876 45652
rect 8932 45596 9000 45652
rect 9056 45596 9124 45652
rect 9180 45596 9248 45652
rect 9304 45596 9372 45652
rect 9428 45596 9496 45652
rect 9552 45596 9620 45652
rect 9676 45596 9744 45652
rect 9800 45596 9810 45652
rect 7874 45528 9810 45596
rect 7874 45472 7884 45528
rect 7940 45472 8008 45528
rect 8064 45472 8132 45528
rect 8188 45472 8256 45528
rect 8312 45472 8380 45528
rect 8436 45472 8504 45528
rect 8560 45472 8628 45528
rect 8684 45472 8752 45528
rect 8808 45472 8876 45528
rect 8932 45472 9000 45528
rect 9056 45472 9124 45528
rect 9180 45472 9248 45528
rect 9304 45472 9372 45528
rect 9428 45472 9496 45528
rect 9552 45472 9620 45528
rect 9676 45472 9744 45528
rect 9800 45472 9810 45528
rect 7874 45404 9810 45472
rect 7874 45348 7884 45404
rect 7940 45348 8008 45404
rect 8064 45348 8132 45404
rect 8188 45348 8256 45404
rect 8312 45348 8380 45404
rect 8436 45348 8504 45404
rect 8560 45348 8628 45404
rect 8684 45348 8752 45404
rect 8808 45348 8876 45404
rect 8932 45348 9000 45404
rect 9056 45348 9124 45404
rect 9180 45348 9248 45404
rect 9304 45348 9372 45404
rect 9428 45348 9496 45404
rect 9552 45348 9620 45404
rect 9676 45348 9744 45404
rect 9800 45348 9810 45404
rect 7874 45280 9810 45348
rect 7874 45224 7884 45280
rect 7940 45224 8008 45280
rect 8064 45224 8132 45280
rect 8188 45224 8256 45280
rect 8312 45224 8380 45280
rect 8436 45224 8504 45280
rect 8560 45224 8628 45280
rect 8684 45224 8752 45280
rect 8808 45224 8876 45280
rect 8932 45224 9000 45280
rect 9056 45224 9124 45280
rect 9180 45224 9248 45280
rect 9304 45224 9372 45280
rect 9428 45224 9496 45280
rect 9552 45224 9620 45280
rect 9676 45224 9744 45280
rect 9800 45224 9810 45280
rect 7874 45156 9810 45224
rect 7874 45100 7884 45156
rect 7940 45100 8008 45156
rect 8064 45100 8132 45156
rect 8188 45100 8256 45156
rect 8312 45100 8380 45156
rect 8436 45100 8504 45156
rect 8560 45100 8628 45156
rect 8684 45100 8752 45156
rect 8808 45100 8876 45156
rect 8932 45100 9000 45156
rect 9056 45100 9124 45156
rect 9180 45100 9248 45156
rect 9304 45100 9372 45156
rect 9428 45100 9496 45156
rect 9552 45100 9620 45156
rect 9676 45100 9744 45156
rect 9800 45100 9810 45156
rect 7874 45032 9810 45100
rect 7874 44976 7884 45032
rect 7940 44976 8008 45032
rect 8064 44976 8132 45032
rect 8188 44976 8256 45032
rect 8312 44976 8380 45032
rect 8436 44976 8504 45032
rect 8560 44976 8628 45032
rect 8684 44976 8752 45032
rect 8808 44976 8876 45032
rect 8932 44976 9000 45032
rect 9056 44976 9124 45032
rect 9180 44976 9248 45032
rect 9304 44976 9372 45032
rect 9428 44976 9496 45032
rect 9552 44976 9620 45032
rect 9676 44976 9744 45032
rect 9800 44976 9810 45032
rect 7874 44908 9810 44976
rect 7874 44852 7884 44908
rect 7940 44852 8008 44908
rect 8064 44852 8132 44908
rect 8188 44852 8256 44908
rect 8312 44852 8380 44908
rect 8436 44852 8504 44908
rect 8560 44852 8628 44908
rect 8684 44852 8752 44908
rect 8808 44852 8876 44908
rect 8932 44852 9000 44908
rect 9056 44852 9124 44908
rect 9180 44852 9248 44908
rect 9304 44852 9372 44908
rect 9428 44852 9496 44908
rect 9552 44852 9620 44908
rect 9676 44852 9744 44908
rect 9800 44852 9810 44908
rect 7874 44842 9810 44852
rect 10244 46148 12180 46158
rect 10244 46092 10254 46148
rect 10310 46092 10378 46148
rect 10434 46092 10502 46148
rect 10558 46092 10626 46148
rect 10682 46092 10750 46148
rect 10806 46092 10874 46148
rect 10930 46092 10998 46148
rect 11054 46092 11122 46148
rect 11178 46092 11246 46148
rect 11302 46092 11370 46148
rect 11426 46092 11494 46148
rect 11550 46092 11618 46148
rect 11674 46092 11742 46148
rect 11798 46092 11866 46148
rect 11922 46092 11990 46148
rect 12046 46092 12114 46148
rect 12170 46092 12180 46148
rect 10244 46024 12180 46092
rect 10244 45968 10254 46024
rect 10310 45968 10378 46024
rect 10434 45968 10502 46024
rect 10558 45968 10626 46024
rect 10682 45968 10750 46024
rect 10806 45968 10874 46024
rect 10930 45968 10998 46024
rect 11054 45968 11122 46024
rect 11178 45968 11246 46024
rect 11302 45968 11370 46024
rect 11426 45968 11494 46024
rect 11550 45968 11618 46024
rect 11674 45968 11742 46024
rect 11798 45968 11866 46024
rect 11922 45968 11990 46024
rect 12046 45968 12114 46024
rect 12170 45968 12180 46024
rect 10244 45900 12180 45968
rect 10244 45844 10254 45900
rect 10310 45844 10378 45900
rect 10434 45844 10502 45900
rect 10558 45844 10626 45900
rect 10682 45844 10750 45900
rect 10806 45844 10874 45900
rect 10930 45844 10998 45900
rect 11054 45844 11122 45900
rect 11178 45844 11246 45900
rect 11302 45844 11370 45900
rect 11426 45844 11494 45900
rect 11550 45844 11618 45900
rect 11674 45844 11742 45900
rect 11798 45844 11866 45900
rect 11922 45844 11990 45900
rect 12046 45844 12114 45900
rect 12170 45844 12180 45900
rect 10244 45776 12180 45844
rect 10244 45720 10254 45776
rect 10310 45720 10378 45776
rect 10434 45720 10502 45776
rect 10558 45720 10626 45776
rect 10682 45720 10750 45776
rect 10806 45720 10874 45776
rect 10930 45720 10998 45776
rect 11054 45720 11122 45776
rect 11178 45720 11246 45776
rect 11302 45720 11370 45776
rect 11426 45720 11494 45776
rect 11550 45720 11618 45776
rect 11674 45720 11742 45776
rect 11798 45720 11866 45776
rect 11922 45720 11990 45776
rect 12046 45720 12114 45776
rect 12170 45720 12180 45776
rect 10244 45652 12180 45720
rect 10244 45596 10254 45652
rect 10310 45596 10378 45652
rect 10434 45596 10502 45652
rect 10558 45596 10626 45652
rect 10682 45596 10750 45652
rect 10806 45596 10874 45652
rect 10930 45596 10998 45652
rect 11054 45596 11122 45652
rect 11178 45596 11246 45652
rect 11302 45596 11370 45652
rect 11426 45596 11494 45652
rect 11550 45596 11618 45652
rect 11674 45596 11742 45652
rect 11798 45596 11866 45652
rect 11922 45596 11990 45652
rect 12046 45596 12114 45652
rect 12170 45596 12180 45652
rect 10244 45528 12180 45596
rect 10244 45472 10254 45528
rect 10310 45472 10378 45528
rect 10434 45472 10502 45528
rect 10558 45472 10626 45528
rect 10682 45472 10750 45528
rect 10806 45472 10874 45528
rect 10930 45472 10998 45528
rect 11054 45472 11122 45528
rect 11178 45472 11246 45528
rect 11302 45472 11370 45528
rect 11426 45472 11494 45528
rect 11550 45472 11618 45528
rect 11674 45472 11742 45528
rect 11798 45472 11866 45528
rect 11922 45472 11990 45528
rect 12046 45472 12114 45528
rect 12170 45472 12180 45528
rect 10244 45404 12180 45472
rect 10244 45348 10254 45404
rect 10310 45348 10378 45404
rect 10434 45348 10502 45404
rect 10558 45348 10626 45404
rect 10682 45348 10750 45404
rect 10806 45348 10874 45404
rect 10930 45348 10998 45404
rect 11054 45348 11122 45404
rect 11178 45348 11246 45404
rect 11302 45348 11370 45404
rect 11426 45348 11494 45404
rect 11550 45348 11618 45404
rect 11674 45348 11742 45404
rect 11798 45348 11866 45404
rect 11922 45348 11990 45404
rect 12046 45348 12114 45404
rect 12170 45348 12180 45404
rect 10244 45280 12180 45348
rect 10244 45224 10254 45280
rect 10310 45224 10378 45280
rect 10434 45224 10502 45280
rect 10558 45224 10626 45280
rect 10682 45224 10750 45280
rect 10806 45224 10874 45280
rect 10930 45224 10998 45280
rect 11054 45224 11122 45280
rect 11178 45224 11246 45280
rect 11302 45224 11370 45280
rect 11426 45224 11494 45280
rect 11550 45224 11618 45280
rect 11674 45224 11742 45280
rect 11798 45224 11866 45280
rect 11922 45224 11990 45280
rect 12046 45224 12114 45280
rect 12170 45224 12180 45280
rect 10244 45156 12180 45224
rect 10244 45100 10254 45156
rect 10310 45100 10378 45156
rect 10434 45100 10502 45156
rect 10558 45100 10626 45156
rect 10682 45100 10750 45156
rect 10806 45100 10874 45156
rect 10930 45100 10998 45156
rect 11054 45100 11122 45156
rect 11178 45100 11246 45156
rect 11302 45100 11370 45156
rect 11426 45100 11494 45156
rect 11550 45100 11618 45156
rect 11674 45100 11742 45156
rect 11798 45100 11866 45156
rect 11922 45100 11990 45156
rect 12046 45100 12114 45156
rect 12170 45100 12180 45156
rect 10244 45032 12180 45100
rect 10244 44976 10254 45032
rect 10310 44976 10378 45032
rect 10434 44976 10502 45032
rect 10558 44976 10626 45032
rect 10682 44976 10750 45032
rect 10806 44976 10874 45032
rect 10930 44976 10998 45032
rect 11054 44976 11122 45032
rect 11178 44976 11246 45032
rect 11302 44976 11370 45032
rect 11426 44976 11494 45032
rect 11550 44976 11618 45032
rect 11674 44976 11742 45032
rect 11798 44976 11866 45032
rect 11922 44976 11990 45032
rect 12046 44976 12114 45032
rect 12170 44976 12180 45032
rect 10244 44908 12180 44976
rect 10244 44852 10254 44908
rect 10310 44852 10378 44908
rect 10434 44852 10502 44908
rect 10558 44852 10626 44908
rect 10682 44852 10750 44908
rect 10806 44852 10874 44908
rect 10930 44852 10998 44908
rect 11054 44852 11122 44908
rect 11178 44852 11246 44908
rect 11302 44852 11370 44908
rect 11426 44852 11494 44908
rect 11550 44852 11618 44908
rect 11674 44852 11742 44908
rect 11798 44852 11866 44908
rect 11922 44852 11990 44908
rect 12046 44852 12114 44908
rect 12170 44852 12180 44908
rect 10244 44842 12180 44852
rect 12861 46148 14673 46158
rect 12861 46092 12871 46148
rect 12927 46092 12995 46148
rect 13051 46092 13119 46148
rect 13175 46092 13243 46148
rect 13299 46092 13367 46148
rect 13423 46092 13491 46148
rect 13547 46092 13615 46148
rect 13671 46092 13739 46148
rect 13795 46092 13863 46148
rect 13919 46092 13987 46148
rect 14043 46092 14111 46148
rect 14167 46092 14235 46148
rect 14291 46092 14359 46148
rect 14415 46092 14483 46148
rect 14539 46092 14607 46148
rect 14663 46092 14673 46148
rect 12861 46024 14673 46092
rect 12861 45968 12871 46024
rect 12927 45968 12995 46024
rect 13051 45968 13119 46024
rect 13175 45968 13243 46024
rect 13299 45968 13367 46024
rect 13423 45968 13491 46024
rect 13547 45968 13615 46024
rect 13671 45968 13739 46024
rect 13795 45968 13863 46024
rect 13919 45968 13987 46024
rect 14043 45968 14111 46024
rect 14167 45968 14235 46024
rect 14291 45968 14359 46024
rect 14415 45968 14483 46024
rect 14539 45968 14607 46024
rect 14663 45968 14673 46024
rect 12861 45900 14673 45968
rect 12861 45844 12871 45900
rect 12927 45844 12995 45900
rect 13051 45844 13119 45900
rect 13175 45844 13243 45900
rect 13299 45844 13367 45900
rect 13423 45844 13491 45900
rect 13547 45844 13615 45900
rect 13671 45844 13739 45900
rect 13795 45844 13863 45900
rect 13919 45844 13987 45900
rect 14043 45844 14111 45900
rect 14167 45844 14235 45900
rect 14291 45844 14359 45900
rect 14415 45844 14483 45900
rect 14539 45844 14607 45900
rect 14663 45844 14673 45900
rect 12861 45776 14673 45844
rect 12861 45720 12871 45776
rect 12927 45720 12995 45776
rect 13051 45720 13119 45776
rect 13175 45720 13243 45776
rect 13299 45720 13367 45776
rect 13423 45720 13491 45776
rect 13547 45720 13615 45776
rect 13671 45720 13739 45776
rect 13795 45720 13863 45776
rect 13919 45720 13987 45776
rect 14043 45720 14111 45776
rect 14167 45720 14235 45776
rect 14291 45720 14359 45776
rect 14415 45720 14483 45776
rect 14539 45720 14607 45776
rect 14663 45720 14673 45776
rect 12861 45652 14673 45720
rect 12861 45596 12871 45652
rect 12927 45596 12995 45652
rect 13051 45596 13119 45652
rect 13175 45596 13243 45652
rect 13299 45596 13367 45652
rect 13423 45596 13491 45652
rect 13547 45596 13615 45652
rect 13671 45596 13739 45652
rect 13795 45596 13863 45652
rect 13919 45596 13987 45652
rect 14043 45596 14111 45652
rect 14167 45596 14235 45652
rect 14291 45596 14359 45652
rect 14415 45596 14483 45652
rect 14539 45596 14607 45652
rect 14663 45596 14673 45652
rect 12861 45528 14673 45596
rect 12861 45472 12871 45528
rect 12927 45472 12995 45528
rect 13051 45472 13119 45528
rect 13175 45472 13243 45528
rect 13299 45472 13367 45528
rect 13423 45472 13491 45528
rect 13547 45472 13615 45528
rect 13671 45472 13739 45528
rect 13795 45472 13863 45528
rect 13919 45472 13987 45528
rect 14043 45472 14111 45528
rect 14167 45472 14235 45528
rect 14291 45472 14359 45528
rect 14415 45472 14483 45528
rect 14539 45472 14607 45528
rect 14663 45472 14673 45528
rect 12861 45404 14673 45472
rect 12861 45348 12871 45404
rect 12927 45348 12995 45404
rect 13051 45348 13119 45404
rect 13175 45348 13243 45404
rect 13299 45348 13367 45404
rect 13423 45348 13491 45404
rect 13547 45348 13615 45404
rect 13671 45348 13739 45404
rect 13795 45348 13863 45404
rect 13919 45348 13987 45404
rect 14043 45348 14111 45404
rect 14167 45348 14235 45404
rect 14291 45348 14359 45404
rect 14415 45348 14483 45404
rect 14539 45348 14607 45404
rect 14663 45348 14673 45404
rect 12861 45280 14673 45348
rect 12861 45224 12871 45280
rect 12927 45224 12995 45280
rect 13051 45224 13119 45280
rect 13175 45224 13243 45280
rect 13299 45224 13367 45280
rect 13423 45224 13491 45280
rect 13547 45224 13615 45280
rect 13671 45224 13739 45280
rect 13795 45224 13863 45280
rect 13919 45224 13987 45280
rect 14043 45224 14111 45280
rect 14167 45224 14235 45280
rect 14291 45224 14359 45280
rect 14415 45224 14483 45280
rect 14539 45224 14607 45280
rect 14663 45224 14673 45280
rect 12861 45156 14673 45224
rect 12861 45100 12871 45156
rect 12927 45100 12995 45156
rect 13051 45100 13119 45156
rect 13175 45100 13243 45156
rect 13299 45100 13367 45156
rect 13423 45100 13491 45156
rect 13547 45100 13615 45156
rect 13671 45100 13739 45156
rect 13795 45100 13863 45156
rect 13919 45100 13987 45156
rect 14043 45100 14111 45156
rect 14167 45100 14235 45156
rect 14291 45100 14359 45156
rect 14415 45100 14483 45156
rect 14539 45100 14607 45156
rect 14663 45100 14673 45156
rect 12861 45032 14673 45100
rect 12861 44976 12871 45032
rect 12927 44976 12995 45032
rect 13051 44976 13119 45032
rect 13175 44976 13243 45032
rect 13299 44976 13367 45032
rect 13423 44976 13491 45032
rect 13547 44976 13615 45032
rect 13671 44976 13739 45032
rect 13795 44976 13863 45032
rect 13919 44976 13987 45032
rect 14043 44976 14111 45032
rect 14167 44976 14235 45032
rect 14291 44976 14359 45032
rect 14415 44976 14483 45032
rect 14539 44976 14607 45032
rect 14663 44976 14673 45032
rect 12861 44908 14673 44976
rect 12861 44852 12871 44908
rect 12927 44852 12995 44908
rect 13051 44852 13119 44908
rect 13175 44852 13243 44908
rect 13299 44852 13367 44908
rect 13423 44852 13491 44908
rect 13547 44852 13615 44908
rect 13671 44852 13739 44908
rect 13795 44852 13863 44908
rect 13919 44852 13987 44908
rect 14043 44852 14111 44908
rect 14167 44852 14235 44908
rect 14291 44852 14359 44908
rect 14415 44852 14483 44908
rect 14539 44852 14607 44908
rect 14663 44852 14673 44908
rect 12861 44842 14673 44852
rect 10 44814 86 44824
rect 14892 44824 14902 46176
rect 14958 44824 14968 46176
rect 14892 44814 14968 44824
rect 2481 44548 2681 44558
rect 2481 44492 2491 44548
rect 2547 44492 2615 44548
rect 2671 44492 2681 44548
rect 2481 44424 2681 44492
rect 2481 44368 2491 44424
rect 2547 44368 2615 44424
rect 2671 44368 2681 44424
rect 2481 44300 2681 44368
rect 2481 44244 2491 44300
rect 2547 44244 2615 44300
rect 2671 44244 2681 44300
rect 2481 44176 2681 44244
rect 2481 44120 2491 44176
rect 2547 44120 2615 44176
rect 2671 44120 2681 44176
rect 2481 44052 2681 44120
rect 2481 43996 2491 44052
rect 2547 43996 2615 44052
rect 2671 43996 2681 44052
rect 2481 43928 2681 43996
rect 2481 43872 2491 43928
rect 2547 43872 2615 43928
rect 2671 43872 2681 43928
rect 2481 43804 2681 43872
rect 2481 43748 2491 43804
rect 2547 43748 2615 43804
rect 2671 43748 2681 43804
rect 2481 43680 2681 43748
rect 2481 43624 2491 43680
rect 2547 43624 2615 43680
rect 2671 43624 2681 43680
rect 2481 43556 2681 43624
rect 2481 43500 2491 43556
rect 2547 43500 2615 43556
rect 2671 43500 2681 43556
rect 2481 43432 2681 43500
rect 2481 43376 2491 43432
rect 2547 43376 2615 43432
rect 2671 43376 2681 43432
rect 2481 43308 2681 43376
rect 2481 43252 2491 43308
rect 2547 43252 2615 43308
rect 2671 43252 2681 43308
rect 2481 43242 2681 43252
rect 4851 44548 5051 44558
rect 4851 44492 4861 44548
rect 4917 44492 4985 44548
rect 5041 44492 5051 44548
rect 4851 44424 5051 44492
rect 4851 44368 4861 44424
rect 4917 44368 4985 44424
rect 5041 44368 5051 44424
rect 4851 44300 5051 44368
rect 4851 44244 4861 44300
rect 4917 44244 4985 44300
rect 5041 44244 5051 44300
rect 4851 44176 5051 44244
rect 4851 44120 4861 44176
rect 4917 44120 4985 44176
rect 5041 44120 5051 44176
rect 4851 44052 5051 44120
rect 4851 43996 4861 44052
rect 4917 43996 4985 44052
rect 5041 43996 5051 44052
rect 4851 43928 5051 43996
rect 4851 43872 4861 43928
rect 4917 43872 4985 43928
rect 5041 43872 5051 43928
rect 4851 43804 5051 43872
rect 4851 43748 4861 43804
rect 4917 43748 4985 43804
rect 5041 43748 5051 43804
rect 4851 43680 5051 43748
rect 4851 43624 4861 43680
rect 4917 43624 4985 43680
rect 5041 43624 5051 43680
rect 4851 43556 5051 43624
rect 4851 43500 4861 43556
rect 4917 43500 4985 43556
rect 5041 43500 5051 43556
rect 4851 43432 5051 43500
rect 4851 43376 4861 43432
rect 4917 43376 4985 43432
rect 5041 43376 5051 43432
rect 4851 43308 5051 43376
rect 4851 43252 4861 43308
rect 4917 43252 4985 43308
rect 5041 43252 5051 43308
rect 4851 43242 5051 43252
rect 7265 44548 7713 44558
rect 7265 44492 7275 44548
rect 7331 44492 7399 44548
rect 7455 44492 7523 44548
rect 7579 44492 7647 44548
rect 7703 44492 7713 44548
rect 7265 44424 7713 44492
rect 7265 44368 7275 44424
rect 7331 44368 7399 44424
rect 7455 44368 7523 44424
rect 7579 44368 7647 44424
rect 7703 44368 7713 44424
rect 7265 44300 7713 44368
rect 7265 44244 7275 44300
rect 7331 44244 7399 44300
rect 7455 44244 7523 44300
rect 7579 44244 7647 44300
rect 7703 44244 7713 44300
rect 7265 44176 7713 44244
rect 7265 44120 7275 44176
rect 7331 44120 7399 44176
rect 7455 44120 7523 44176
rect 7579 44120 7647 44176
rect 7703 44120 7713 44176
rect 7265 44052 7713 44120
rect 7265 43996 7275 44052
rect 7331 43996 7399 44052
rect 7455 43996 7523 44052
rect 7579 43996 7647 44052
rect 7703 43996 7713 44052
rect 7265 43928 7713 43996
rect 7265 43872 7275 43928
rect 7331 43872 7399 43928
rect 7455 43872 7523 43928
rect 7579 43872 7647 43928
rect 7703 43872 7713 43928
rect 7265 43804 7713 43872
rect 7265 43748 7275 43804
rect 7331 43748 7399 43804
rect 7455 43748 7523 43804
rect 7579 43748 7647 43804
rect 7703 43748 7713 43804
rect 7265 43680 7713 43748
rect 7265 43624 7275 43680
rect 7331 43624 7399 43680
rect 7455 43624 7523 43680
rect 7579 43624 7647 43680
rect 7703 43624 7713 43680
rect 7265 43556 7713 43624
rect 7265 43500 7275 43556
rect 7331 43500 7399 43556
rect 7455 43500 7523 43556
rect 7579 43500 7647 43556
rect 7703 43500 7713 43556
rect 7265 43432 7713 43500
rect 7265 43376 7275 43432
rect 7331 43376 7399 43432
rect 7455 43376 7523 43432
rect 7579 43376 7647 43432
rect 7703 43376 7713 43432
rect 7265 43308 7713 43376
rect 7265 43252 7275 43308
rect 7331 43252 7399 43308
rect 7455 43252 7523 43308
rect 7579 43252 7647 43308
rect 7703 43252 7713 43308
rect 7265 43242 7713 43252
rect 9927 44548 10127 44558
rect 9927 44492 9937 44548
rect 9993 44492 10061 44548
rect 10117 44492 10127 44548
rect 9927 44424 10127 44492
rect 9927 44368 9937 44424
rect 9993 44368 10061 44424
rect 10117 44368 10127 44424
rect 9927 44300 10127 44368
rect 9927 44244 9937 44300
rect 9993 44244 10061 44300
rect 10117 44244 10127 44300
rect 9927 44176 10127 44244
rect 9927 44120 9937 44176
rect 9993 44120 10061 44176
rect 10117 44120 10127 44176
rect 9927 44052 10127 44120
rect 9927 43996 9937 44052
rect 9993 43996 10061 44052
rect 10117 43996 10127 44052
rect 9927 43928 10127 43996
rect 9927 43872 9937 43928
rect 9993 43872 10061 43928
rect 10117 43872 10127 43928
rect 9927 43804 10127 43872
rect 9927 43748 9937 43804
rect 9993 43748 10061 43804
rect 10117 43748 10127 43804
rect 9927 43680 10127 43748
rect 9927 43624 9937 43680
rect 9993 43624 10061 43680
rect 10117 43624 10127 43680
rect 9927 43556 10127 43624
rect 9927 43500 9937 43556
rect 9993 43500 10061 43556
rect 10117 43500 10127 43556
rect 9927 43432 10127 43500
rect 9927 43376 9937 43432
rect 9993 43376 10061 43432
rect 10117 43376 10127 43432
rect 9927 43308 10127 43376
rect 9927 43252 9937 43308
rect 9993 43252 10061 43308
rect 10117 43252 10127 43308
rect 9927 43242 10127 43252
rect 12297 44548 12497 44558
rect 12297 44492 12307 44548
rect 12363 44492 12431 44548
rect 12487 44492 12497 44548
rect 12297 44424 12497 44492
rect 12297 44368 12307 44424
rect 12363 44368 12431 44424
rect 12487 44368 12497 44424
rect 12297 44300 12497 44368
rect 12297 44244 12307 44300
rect 12363 44244 12431 44300
rect 12487 44244 12497 44300
rect 12297 44176 12497 44244
rect 12297 44120 12307 44176
rect 12363 44120 12431 44176
rect 12487 44120 12497 44176
rect 12297 44052 12497 44120
rect 12297 43996 12307 44052
rect 12363 43996 12431 44052
rect 12487 43996 12497 44052
rect 12297 43928 12497 43996
rect 12297 43872 12307 43928
rect 12363 43872 12431 43928
rect 12487 43872 12497 43928
rect 12297 43804 12497 43872
rect 12297 43748 12307 43804
rect 12363 43748 12431 43804
rect 12487 43748 12497 43804
rect 12297 43680 12497 43748
rect 12297 43624 12307 43680
rect 12363 43624 12431 43680
rect 12487 43624 12497 43680
rect 12297 43556 12497 43624
rect 12297 43500 12307 43556
rect 12363 43500 12431 43556
rect 12487 43500 12497 43556
rect 12297 43432 12497 43500
rect 12297 43376 12307 43432
rect 12363 43376 12431 43432
rect 12487 43376 12497 43432
rect 12297 43308 12497 43376
rect 12297 43252 12307 43308
rect 12363 43252 12431 43308
rect 12487 43252 12497 43308
rect 12297 43242 12497 43252
rect 2481 42948 2681 42958
rect 2481 42892 2491 42948
rect 2547 42892 2615 42948
rect 2671 42892 2681 42948
rect 2481 42824 2681 42892
rect 2481 42768 2491 42824
rect 2547 42768 2615 42824
rect 2671 42768 2681 42824
rect 2481 42700 2681 42768
rect 2481 42644 2491 42700
rect 2547 42644 2615 42700
rect 2671 42644 2681 42700
rect 2481 42576 2681 42644
rect 2481 42520 2491 42576
rect 2547 42520 2615 42576
rect 2671 42520 2681 42576
rect 2481 42452 2681 42520
rect 2481 42396 2491 42452
rect 2547 42396 2615 42452
rect 2671 42396 2681 42452
rect 2481 42328 2681 42396
rect 2481 42272 2491 42328
rect 2547 42272 2615 42328
rect 2671 42272 2681 42328
rect 2481 42204 2681 42272
rect 2481 42148 2491 42204
rect 2547 42148 2615 42204
rect 2671 42148 2681 42204
rect 2481 42080 2681 42148
rect 2481 42024 2491 42080
rect 2547 42024 2615 42080
rect 2671 42024 2681 42080
rect 2481 41956 2681 42024
rect 2481 41900 2491 41956
rect 2547 41900 2615 41956
rect 2671 41900 2681 41956
rect 2481 41832 2681 41900
rect 2481 41776 2491 41832
rect 2547 41776 2615 41832
rect 2671 41776 2681 41832
rect 2481 41708 2681 41776
rect 2481 41652 2491 41708
rect 2547 41652 2615 41708
rect 2671 41652 2681 41708
rect 2481 41642 2681 41652
rect 4851 42948 5051 42958
rect 4851 42892 4861 42948
rect 4917 42892 4985 42948
rect 5041 42892 5051 42948
rect 4851 42824 5051 42892
rect 4851 42768 4861 42824
rect 4917 42768 4985 42824
rect 5041 42768 5051 42824
rect 4851 42700 5051 42768
rect 4851 42644 4861 42700
rect 4917 42644 4985 42700
rect 5041 42644 5051 42700
rect 4851 42576 5051 42644
rect 4851 42520 4861 42576
rect 4917 42520 4985 42576
rect 5041 42520 5051 42576
rect 4851 42452 5051 42520
rect 4851 42396 4861 42452
rect 4917 42396 4985 42452
rect 5041 42396 5051 42452
rect 4851 42328 5051 42396
rect 4851 42272 4861 42328
rect 4917 42272 4985 42328
rect 5041 42272 5051 42328
rect 4851 42204 5051 42272
rect 4851 42148 4861 42204
rect 4917 42148 4985 42204
rect 5041 42148 5051 42204
rect 4851 42080 5051 42148
rect 4851 42024 4861 42080
rect 4917 42024 4985 42080
rect 5041 42024 5051 42080
rect 4851 41956 5051 42024
rect 4851 41900 4861 41956
rect 4917 41900 4985 41956
rect 5041 41900 5051 41956
rect 4851 41832 5051 41900
rect 4851 41776 4861 41832
rect 4917 41776 4985 41832
rect 5041 41776 5051 41832
rect 4851 41708 5051 41776
rect 4851 41652 4861 41708
rect 4917 41652 4985 41708
rect 5041 41652 5051 41708
rect 4851 41642 5051 41652
rect 7265 42948 7713 42958
rect 7265 42892 7275 42948
rect 7331 42892 7399 42948
rect 7455 42892 7523 42948
rect 7579 42892 7647 42948
rect 7703 42892 7713 42948
rect 7265 42824 7713 42892
rect 7265 42768 7275 42824
rect 7331 42768 7399 42824
rect 7455 42768 7523 42824
rect 7579 42768 7647 42824
rect 7703 42768 7713 42824
rect 7265 42700 7713 42768
rect 7265 42644 7275 42700
rect 7331 42644 7399 42700
rect 7455 42644 7523 42700
rect 7579 42644 7647 42700
rect 7703 42644 7713 42700
rect 7265 42576 7713 42644
rect 7265 42520 7275 42576
rect 7331 42520 7399 42576
rect 7455 42520 7523 42576
rect 7579 42520 7647 42576
rect 7703 42520 7713 42576
rect 7265 42452 7713 42520
rect 7265 42396 7275 42452
rect 7331 42396 7399 42452
rect 7455 42396 7523 42452
rect 7579 42396 7647 42452
rect 7703 42396 7713 42452
rect 7265 42328 7713 42396
rect 7265 42272 7275 42328
rect 7331 42272 7399 42328
rect 7455 42272 7523 42328
rect 7579 42272 7647 42328
rect 7703 42272 7713 42328
rect 7265 42204 7713 42272
rect 7265 42148 7275 42204
rect 7331 42148 7399 42204
rect 7455 42148 7523 42204
rect 7579 42148 7647 42204
rect 7703 42148 7713 42204
rect 7265 42080 7713 42148
rect 7265 42024 7275 42080
rect 7331 42024 7399 42080
rect 7455 42024 7523 42080
rect 7579 42024 7647 42080
rect 7703 42024 7713 42080
rect 7265 41956 7713 42024
rect 7265 41900 7275 41956
rect 7331 41900 7399 41956
rect 7455 41900 7523 41956
rect 7579 41900 7647 41956
rect 7703 41900 7713 41956
rect 7265 41832 7713 41900
rect 7265 41776 7275 41832
rect 7331 41776 7399 41832
rect 7455 41776 7523 41832
rect 7579 41776 7647 41832
rect 7703 41776 7713 41832
rect 7265 41708 7713 41776
rect 7265 41652 7275 41708
rect 7331 41652 7399 41708
rect 7455 41652 7523 41708
rect 7579 41652 7647 41708
rect 7703 41652 7713 41708
rect 7265 41642 7713 41652
rect 9927 42948 10127 42958
rect 9927 42892 9937 42948
rect 9993 42892 10061 42948
rect 10117 42892 10127 42948
rect 9927 42824 10127 42892
rect 9927 42768 9937 42824
rect 9993 42768 10061 42824
rect 10117 42768 10127 42824
rect 9927 42700 10127 42768
rect 9927 42644 9937 42700
rect 9993 42644 10061 42700
rect 10117 42644 10127 42700
rect 9927 42576 10127 42644
rect 9927 42520 9937 42576
rect 9993 42520 10061 42576
rect 10117 42520 10127 42576
rect 9927 42452 10127 42520
rect 9927 42396 9937 42452
rect 9993 42396 10061 42452
rect 10117 42396 10127 42452
rect 9927 42328 10127 42396
rect 9927 42272 9937 42328
rect 9993 42272 10061 42328
rect 10117 42272 10127 42328
rect 9927 42204 10127 42272
rect 9927 42148 9937 42204
rect 9993 42148 10061 42204
rect 10117 42148 10127 42204
rect 9927 42080 10127 42148
rect 9927 42024 9937 42080
rect 9993 42024 10061 42080
rect 10117 42024 10127 42080
rect 9927 41956 10127 42024
rect 9927 41900 9937 41956
rect 9993 41900 10061 41956
rect 10117 41900 10127 41956
rect 9927 41832 10127 41900
rect 9927 41776 9937 41832
rect 9993 41776 10061 41832
rect 10117 41776 10127 41832
rect 9927 41708 10127 41776
rect 9927 41652 9937 41708
rect 9993 41652 10061 41708
rect 10117 41652 10127 41708
rect 9927 41642 10127 41652
rect 12297 42948 12497 42958
rect 12297 42892 12307 42948
rect 12363 42892 12431 42948
rect 12487 42892 12497 42948
rect 12297 42824 12497 42892
rect 12297 42768 12307 42824
rect 12363 42768 12431 42824
rect 12487 42768 12497 42824
rect 12297 42700 12497 42768
rect 12297 42644 12307 42700
rect 12363 42644 12431 42700
rect 12487 42644 12497 42700
rect 12297 42576 12497 42644
rect 12297 42520 12307 42576
rect 12363 42520 12431 42576
rect 12487 42520 12497 42576
rect 12297 42452 12497 42520
rect 12297 42396 12307 42452
rect 12363 42396 12431 42452
rect 12487 42396 12497 42452
rect 12297 42328 12497 42396
rect 12297 42272 12307 42328
rect 12363 42272 12431 42328
rect 12487 42272 12497 42328
rect 12297 42204 12497 42272
rect 12297 42148 12307 42204
rect 12363 42148 12431 42204
rect 12487 42148 12497 42204
rect 12297 42080 12497 42148
rect 12297 42024 12307 42080
rect 12363 42024 12431 42080
rect 12487 42024 12497 42080
rect 12297 41956 12497 42024
rect 12297 41900 12307 41956
rect 12363 41900 12431 41956
rect 12487 41900 12497 41956
rect 12297 41832 12497 41900
rect 12297 41776 12307 41832
rect 12363 41776 12431 41832
rect 12487 41776 12497 41832
rect 12297 41708 12497 41776
rect 12297 41652 12307 41708
rect 12363 41652 12431 41708
rect 12487 41652 12497 41708
rect 12297 41642 12497 41652
rect 2481 41348 2681 41358
rect 2481 41292 2491 41348
rect 2547 41292 2615 41348
rect 2671 41292 2681 41348
rect 2481 41224 2681 41292
rect 2481 41168 2491 41224
rect 2547 41168 2615 41224
rect 2671 41168 2681 41224
rect 2481 41100 2681 41168
rect 2481 41044 2491 41100
rect 2547 41044 2615 41100
rect 2671 41044 2681 41100
rect 2481 40976 2681 41044
rect 2481 40920 2491 40976
rect 2547 40920 2615 40976
rect 2671 40920 2681 40976
rect 2481 40852 2681 40920
rect 2481 40796 2491 40852
rect 2547 40796 2615 40852
rect 2671 40796 2681 40852
rect 2481 40728 2681 40796
rect 2481 40672 2491 40728
rect 2547 40672 2615 40728
rect 2671 40672 2681 40728
rect 2481 40604 2681 40672
rect 2481 40548 2491 40604
rect 2547 40548 2615 40604
rect 2671 40548 2681 40604
rect 2481 40480 2681 40548
rect 2481 40424 2491 40480
rect 2547 40424 2615 40480
rect 2671 40424 2681 40480
rect 2481 40356 2681 40424
rect 2481 40300 2491 40356
rect 2547 40300 2615 40356
rect 2671 40300 2681 40356
rect 2481 40232 2681 40300
rect 2481 40176 2491 40232
rect 2547 40176 2615 40232
rect 2671 40176 2681 40232
rect 2481 40108 2681 40176
rect 2481 40052 2491 40108
rect 2547 40052 2615 40108
rect 2671 40052 2681 40108
rect 2481 40042 2681 40052
rect 4851 41348 5051 41358
rect 4851 41292 4861 41348
rect 4917 41292 4985 41348
rect 5041 41292 5051 41348
rect 4851 41224 5051 41292
rect 4851 41168 4861 41224
rect 4917 41168 4985 41224
rect 5041 41168 5051 41224
rect 4851 41100 5051 41168
rect 4851 41044 4861 41100
rect 4917 41044 4985 41100
rect 5041 41044 5051 41100
rect 4851 40976 5051 41044
rect 4851 40920 4861 40976
rect 4917 40920 4985 40976
rect 5041 40920 5051 40976
rect 4851 40852 5051 40920
rect 4851 40796 4861 40852
rect 4917 40796 4985 40852
rect 5041 40796 5051 40852
rect 4851 40728 5051 40796
rect 4851 40672 4861 40728
rect 4917 40672 4985 40728
rect 5041 40672 5051 40728
rect 4851 40604 5051 40672
rect 4851 40548 4861 40604
rect 4917 40548 4985 40604
rect 5041 40548 5051 40604
rect 4851 40480 5051 40548
rect 4851 40424 4861 40480
rect 4917 40424 4985 40480
rect 5041 40424 5051 40480
rect 4851 40356 5051 40424
rect 4851 40300 4861 40356
rect 4917 40300 4985 40356
rect 5041 40300 5051 40356
rect 4851 40232 5051 40300
rect 4851 40176 4861 40232
rect 4917 40176 4985 40232
rect 5041 40176 5051 40232
rect 4851 40108 5051 40176
rect 4851 40052 4861 40108
rect 4917 40052 4985 40108
rect 5041 40052 5051 40108
rect 4851 40042 5051 40052
rect 7265 41348 7713 41358
rect 7265 41292 7275 41348
rect 7331 41292 7399 41348
rect 7455 41292 7523 41348
rect 7579 41292 7647 41348
rect 7703 41292 7713 41348
rect 7265 41224 7713 41292
rect 7265 41168 7275 41224
rect 7331 41168 7399 41224
rect 7455 41168 7523 41224
rect 7579 41168 7647 41224
rect 7703 41168 7713 41224
rect 7265 41100 7713 41168
rect 7265 41044 7275 41100
rect 7331 41044 7399 41100
rect 7455 41044 7523 41100
rect 7579 41044 7647 41100
rect 7703 41044 7713 41100
rect 7265 40976 7713 41044
rect 7265 40920 7275 40976
rect 7331 40920 7399 40976
rect 7455 40920 7523 40976
rect 7579 40920 7647 40976
rect 7703 40920 7713 40976
rect 7265 40852 7713 40920
rect 7265 40796 7275 40852
rect 7331 40796 7399 40852
rect 7455 40796 7523 40852
rect 7579 40796 7647 40852
rect 7703 40796 7713 40852
rect 7265 40728 7713 40796
rect 7265 40672 7275 40728
rect 7331 40672 7399 40728
rect 7455 40672 7523 40728
rect 7579 40672 7647 40728
rect 7703 40672 7713 40728
rect 7265 40604 7713 40672
rect 7265 40548 7275 40604
rect 7331 40548 7399 40604
rect 7455 40548 7523 40604
rect 7579 40548 7647 40604
rect 7703 40548 7713 40604
rect 7265 40480 7713 40548
rect 7265 40424 7275 40480
rect 7331 40424 7399 40480
rect 7455 40424 7523 40480
rect 7579 40424 7647 40480
rect 7703 40424 7713 40480
rect 7265 40356 7713 40424
rect 7265 40300 7275 40356
rect 7331 40300 7399 40356
rect 7455 40300 7523 40356
rect 7579 40300 7647 40356
rect 7703 40300 7713 40356
rect 7265 40232 7713 40300
rect 7265 40176 7275 40232
rect 7331 40176 7399 40232
rect 7455 40176 7523 40232
rect 7579 40176 7647 40232
rect 7703 40176 7713 40232
rect 7265 40108 7713 40176
rect 7265 40052 7275 40108
rect 7331 40052 7399 40108
rect 7455 40052 7523 40108
rect 7579 40052 7647 40108
rect 7703 40052 7713 40108
rect 7265 40042 7713 40052
rect 9927 41348 10127 41358
rect 9927 41292 9937 41348
rect 9993 41292 10061 41348
rect 10117 41292 10127 41348
rect 9927 41224 10127 41292
rect 9927 41168 9937 41224
rect 9993 41168 10061 41224
rect 10117 41168 10127 41224
rect 9927 41100 10127 41168
rect 9927 41044 9937 41100
rect 9993 41044 10061 41100
rect 10117 41044 10127 41100
rect 9927 40976 10127 41044
rect 9927 40920 9937 40976
rect 9993 40920 10061 40976
rect 10117 40920 10127 40976
rect 9927 40852 10127 40920
rect 9927 40796 9937 40852
rect 9993 40796 10061 40852
rect 10117 40796 10127 40852
rect 9927 40728 10127 40796
rect 9927 40672 9937 40728
rect 9993 40672 10061 40728
rect 10117 40672 10127 40728
rect 9927 40604 10127 40672
rect 9927 40548 9937 40604
rect 9993 40548 10061 40604
rect 10117 40548 10127 40604
rect 9927 40480 10127 40548
rect 9927 40424 9937 40480
rect 9993 40424 10061 40480
rect 10117 40424 10127 40480
rect 9927 40356 10127 40424
rect 9927 40300 9937 40356
rect 9993 40300 10061 40356
rect 10117 40300 10127 40356
rect 9927 40232 10127 40300
rect 9927 40176 9937 40232
rect 9993 40176 10061 40232
rect 10117 40176 10127 40232
rect 9927 40108 10127 40176
rect 9927 40052 9937 40108
rect 9993 40052 10061 40108
rect 10117 40052 10127 40108
rect 9927 40042 10127 40052
rect 12297 41348 12497 41358
rect 12297 41292 12307 41348
rect 12363 41292 12431 41348
rect 12487 41292 12497 41348
rect 12297 41224 12497 41292
rect 12297 41168 12307 41224
rect 12363 41168 12431 41224
rect 12487 41168 12497 41224
rect 12297 41100 12497 41168
rect 12297 41044 12307 41100
rect 12363 41044 12431 41100
rect 12487 41044 12497 41100
rect 12297 40976 12497 41044
rect 12297 40920 12307 40976
rect 12363 40920 12431 40976
rect 12487 40920 12497 40976
rect 12297 40852 12497 40920
rect 12297 40796 12307 40852
rect 12363 40796 12431 40852
rect 12487 40796 12497 40852
rect 12297 40728 12497 40796
rect 12297 40672 12307 40728
rect 12363 40672 12431 40728
rect 12487 40672 12497 40728
rect 12297 40604 12497 40672
rect 12297 40548 12307 40604
rect 12363 40548 12431 40604
rect 12487 40548 12497 40604
rect 12297 40480 12497 40548
rect 12297 40424 12307 40480
rect 12363 40424 12431 40480
rect 12487 40424 12497 40480
rect 12297 40356 12497 40424
rect 12297 40300 12307 40356
rect 12363 40300 12431 40356
rect 12487 40300 12497 40356
rect 12297 40232 12497 40300
rect 12297 40176 12307 40232
rect 12363 40176 12431 40232
rect 12487 40176 12497 40232
rect 12297 40108 12497 40176
rect 12297 40052 12307 40108
rect 12363 40052 12431 40108
rect 12487 40052 12497 40108
rect 12297 40042 12497 40052
rect 2292 39727 2368 39737
rect 2292 39671 2302 39727
rect 2358 39671 2368 39727
rect 2292 39595 2368 39671
rect 2292 39539 2302 39595
rect 2358 39539 2368 39595
rect 2292 39463 2368 39539
rect 2292 39407 2302 39463
rect 2358 39407 2368 39463
rect 2292 39331 2368 39407
rect 2292 39275 2302 39331
rect 2358 39275 2368 39331
rect 2292 39199 2368 39275
rect 2292 39143 2302 39199
rect 2358 39143 2368 39199
rect 2292 39067 2368 39143
rect 2292 39011 2302 39067
rect 2358 39011 2368 39067
rect 2292 38935 2368 39011
rect 2292 38879 2302 38935
rect 2358 38879 2368 38935
rect 2292 38803 2368 38879
rect 2292 38747 2302 38803
rect 2358 38747 2368 38803
rect 2292 38671 2368 38747
rect 2292 38615 2302 38671
rect 2358 38615 2368 38671
rect 2292 38539 2368 38615
rect 2292 38483 2302 38539
rect 2358 38483 2368 38539
rect 2292 38473 2368 38483
rect 10 38176 86 38186
rect 10 36824 20 38176
rect 76 36824 86 38176
rect 14892 38176 14968 38186
rect 305 38148 2117 38158
rect 305 38092 315 38148
rect 371 38092 439 38148
rect 495 38092 563 38148
rect 619 38092 687 38148
rect 743 38092 811 38148
rect 867 38092 935 38148
rect 991 38092 1059 38148
rect 1115 38092 1183 38148
rect 1239 38092 1307 38148
rect 1363 38092 1431 38148
rect 1487 38092 1555 38148
rect 1611 38092 1679 38148
rect 1735 38092 1803 38148
rect 1859 38092 1927 38148
rect 1983 38092 2051 38148
rect 2107 38092 2117 38148
rect 305 38024 2117 38092
rect 305 37968 315 38024
rect 371 37968 439 38024
rect 495 37968 563 38024
rect 619 37968 687 38024
rect 743 37968 811 38024
rect 867 37968 935 38024
rect 991 37968 1059 38024
rect 1115 37968 1183 38024
rect 1239 37968 1307 38024
rect 1363 37968 1431 38024
rect 1487 37968 1555 38024
rect 1611 37968 1679 38024
rect 1735 37968 1803 38024
rect 1859 37968 1927 38024
rect 1983 37968 2051 38024
rect 2107 37968 2117 38024
rect 305 37900 2117 37968
rect 305 37844 315 37900
rect 371 37844 439 37900
rect 495 37844 563 37900
rect 619 37844 687 37900
rect 743 37844 811 37900
rect 867 37844 935 37900
rect 991 37844 1059 37900
rect 1115 37844 1183 37900
rect 1239 37844 1307 37900
rect 1363 37844 1431 37900
rect 1487 37844 1555 37900
rect 1611 37844 1679 37900
rect 1735 37844 1803 37900
rect 1859 37844 1927 37900
rect 1983 37844 2051 37900
rect 2107 37844 2117 37900
rect 305 37776 2117 37844
rect 305 37720 315 37776
rect 371 37720 439 37776
rect 495 37720 563 37776
rect 619 37720 687 37776
rect 743 37720 811 37776
rect 867 37720 935 37776
rect 991 37720 1059 37776
rect 1115 37720 1183 37776
rect 1239 37720 1307 37776
rect 1363 37720 1431 37776
rect 1487 37720 1555 37776
rect 1611 37720 1679 37776
rect 1735 37720 1803 37776
rect 1859 37720 1927 37776
rect 1983 37720 2051 37776
rect 2107 37720 2117 37776
rect 305 37652 2117 37720
rect 305 37596 315 37652
rect 371 37596 439 37652
rect 495 37596 563 37652
rect 619 37596 687 37652
rect 743 37596 811 37652
rect 867 37596 935 37652
rect 991 37596 1059 37652
rect 1115 37596 1183 37652
rect 1239 37596 1307 37652
rect 1363 37596 1431 37652
rect 1487 37596 1555 37652
rect 1611 37596 1679 37652
rect 1735 37596 1803 37652
rect 1859 37596 1927 37652
rect 1983 37596 2051 37652
rect 2107 37596 2117 37652
rect 305 37528 2117 37596
rect 305 37472 315 37528
rect 371 37472 439 37528
rect 495 37472 563 37528
rect 619 37472 687 37528
rect 743 37472 811 37528
rect 867 37472 935 37528
rect 991 37472 1059 37528
rect 1115 37472 1183 37528
rect 1239 37472 1307 37528
rect 1363 37472 1431 37528
rect 1487 37472 1555 37528
rect 1611 37472 1679 37528
rect 1735 37472 1803 37528
rect 1859 37472 1927 37528
rect 1983 37472 2051 37528
rect 2107 37472 2117 37528
rect 305 37404 2117 37472
rect 305 37348 315 37404
rect 371 37348 439 37404
rect 495 37348 563 37404
rect 619 37348 687 37404
rect 743 37348 811 37404
rect 867 37348 935 37404
rect 991 37348 1059 37404
rect 1115 37348 1183 37404
rect 1239 37348 1307 37404
rect 1363 37348 1431 37404
rect 1487 37348 1555 37404
rect 1611 37348 1679 37404
rect 1735 37348 1803 37404
rect 1859 37348 1927 37404
rect 1983 37348 2051 37404
rect 2107 37348 2117 37404
rect 305 37280 2117 37348
rect 305 37224 315 37280
rect 371 37224 439 37280
rect 495 37224 563 37280
rect 619 37224 687 37280
rect 743 37224 811 37280
rect 867 37224 935 37280
rect 991 37224 1059 37280
rect 1115 37224 1183 37280
rect 1239 37224 1307 37280
rect 1363 37224 1431 37280
rect 1487 37224 1555 37280
rect 1611 37224 1679 37280
rect 1735 37224 1803 37280
rect 1859 37224 1927 37280
rect 1983 37224 2051 37280
rect 2107 37224 2117 37280
rect 305 37156 2117 37224
rect 305 37100 315 37156
rect 371 37100 439 37156
rect 495 37100 563 37156
rect 619 37100 687 37156
rect 743 37100 811 37156
rect 867 37100 935 37156
rect 991 37100 1059 37156
rect 1115 37100 1183 37156
rect 1239 37100 1307 37156
rect 1363 37100 1431 37156
rect 1487 37100 1555 37156
rect 1611 37100 1679 37156
rect 1735 37100 1803 37156
rect 1859 37100 1927 37156
rect 1983 37100 2051 37156
rect 2107 37100 2117 37156
rect 305 37032 2117 37100
rect 305 36976 315 37032
rect 371 36976 439 37032
rect 495 36976 563 37032
rect 619 36976 687 37032
rect 743 36976 811 37032
rect 867 36976 935 37032
rect 991 36976 1059 37032
rect 1115 36976 1183 37032
rect 1239 36976 1307 37032
rect 1363 36976 1431 37032
rect 1487 36976 1555 37032
rect 1611 36976 1679 37032
rect 1735 36976 1803 37032
rect 1859 36976 1927 37032
rect 1983 36976 2051 37032
rect 2107 36976 2117 37032
rect 305 36908 2117 36976
rect 305 36852 315 36908
rect 371 36852 439 36908
rect 495 36852 563 36908
rect 619 36852 687 36908
rect 743 36852 811 36908
rect 867 36852 935 36908
rect 991 36852 1059 36908
rect 1115 36852 1183 36908
rect 1239 36852 1307 36908
rect 1363 36852 1431 36908
rect 1487 36852 1555 36908
rect 1611 36852 1679 36908
rect 1735 36852 1803 36908
rect 1859 36852 1927 36908
rect 1983 36852 2051 36908
rect 2107 36852 2117 36908
rect 305 36842 2117 36852
rect 2798 38148 4734 38158
rect 2798 38092 2808 38148
rect 2864 38092 2932 38148
rect 2988 38092 3056 38148
rect 3112 38092 3180 38148
rect 3236 38092 3304 38148
rect 3360 38092 3428 38148
rect 3484 38092 3552 38148
rect 3608 38092 3676 38148
rect 3732 38092 3800 38148
rect 3856 38092 3924 38148
rect 3980 38092 4048 38148
rect 4104 38092 4172 38148
rect 4228 38092 4296 38148
rect 4352 38092 4420 38148
rect 4476 38092 4544 38148
rect 4600 38092 4668 38148
rect 4724 38092 4734 38148
rect 2798 38024 4734 38092
rect 2798 37968 2808 38024
rect 2864 37968 2932 38024
rect 2988 37968 3056 38024
rect 3112 37968 3180 38024
rect 3236 37968 3304 38024
rect 3360 37968 3428 38024
rect 3484 37968 3552 38024
rect 3608 37968 3676 38024
rect 3732 37968 3800 38024
rect 3856 37968 3924 38024
rect 3980 37968 4048 38024
rect 4104 37968 4172 38024
rect 4228 37968 4296 38024
rect 4352 37968 4420 38024
rect 4476 37968 4544 38024
rect 4600 37968 4668 38024
rect 4724 37968 4734 38024
rect 2798 37900 4734 37968
rect 2798 37844 2808 37900
rect 2864 37844 2932 37900
rect 2988 37844 3056 37900
rect 3112 37844 3180 37900
rect 3236 37844 3304 37900
rect 3360 37844 3428 37900
rect 3484 37844 3552 37900
rect 3608 37844 3676 37900
rect 3732 37844 3800 37900
rect 3856 37844 3924 37900
rect 3980 37844 4048 37900
rect 4104 37844 4172 37900
rect 4228 37844 4296 37900
rect 4352 37844 4420 37900
rect 4476 37844 4544 37900
rect 4600 37844 4668 37900
rect 4724 37844 4734 37900
rect 2798 37776 4734 37844
rect 2798 37720 2808 37776
rect 2864 37720 2932 37776
rect 2988 37720 3056 37776
rect 3112 37720 3180 37776
rect 3236 37720 3304 37776
rect 3360 37720 3428 37776
rect 3484 37720 3552 37776
rect 3608 37720 3676 37776
rect 3732 37720 3800 37776
rect 3856 37720 3924 37776
rect 3980 37720 4048 37776
rect 4104 37720 4172 37776
rect 4228 37720 4296 37776
rect 4352 37720 4420 37776
rect 4476 37720 4544 37776
rect 4600 37720 4668 37776
rect 4724 37720 4734 37776
rect 2798 37652 4734 37720
rect 2798 37596 2808 37652
rect 2864 37596 2932 37652
rect 2988 37596 3056 37652
rect 3112 37596 3180 37652
rect 3236 37596 3304 37652
rect 3360 37596 3428 37652
rect 3484 37596 3552 37652
rect 3608 37596 3676 37652
rect 3732 37596 3800 37652
rect 3856 37596 3924 37652
rect 3980 37596 4048 37652
rect 4104 37596 4172 37652
rect 4228 37596 4296 37652
rect 4352 37596 4420 37652
rect 4476 37596 4544 37652
rect 4600 37596 4668 37652
rect 4724 37596 4734 37652
rect 2798 37528 4734 37596
rect 2798 37472 2808 37528
rect 2864 37472 2932 37528
rect 2988 37472 3056 37528
rect 3112 37472 3180 37528
rect 3236 37472 3304 37528
rect 3360 37472 3428 37528
rect 3484 37472 3552 37528
rect 3608 37472 3676 37528
rect 3732 37472 3800 37528
rect 3856 37472 3924 37528
rect 3980 37472 4048 37528
rect 4104 37472 4172 37528
rect 4228 37472 4296 37528
rect 4352 37472 4420 37528
rect 4476 37472 4544 37528
rect 4600 37472 4668 37528
rect 4724 37472 4734 37528
rect 2798 37404 4734 37472
rect 2798 37348 2808 37404
rect 2864 37348 2932 37404
rect 2988 37348 3056 37404
rect 3112 37348 3180 37404
rect 3236 37348 3304 37404
rect 3360 37348 3428 37404
rect 3484 37348 3552 37404
rect 3608 37348 3676 37404
rect 3732 37348 3800 37404
rect 3856 37348 3924 37404
rect 3980 37348 4048 37404
rect 4104 37348 4172 37404
rect 4228 37348 4296 37404
rect 4352 37348 4420 37404
rect 4476 37348 4544 37404
rect 4600 37348 4668 37404
rect 4724 37348 4734 37404
rect 2798 37280 4734 37348
rect 2798 37224 2808 37280
rect 2864 37224 2932 37280
rect 2988 37224 3056 37280
rect 3112 37224 3180 37280
rect 3236 37224 3304 37280
rect 3360 37224 3428 37280
rect 3484 37224 3552 37280
rect 3608 37224 3676 37280
rect 3732 37224 3800 37280
rect 3856 37224 3924 37280
rect 3980 37224 4048 37280
rect 4104 37224 4172 37280
rect 4228 37224 4296 37280
rect 4352 37224 4420 37280
rect 4476 37224 4544 37280
rect 4600 37224 4668 37280
rect 4724 37224 4734 37280
rect 2798 37156 4734 37224
rect 2798 37100 2808 37156
rect 2864 37100 2932 37156
rect 2988 37100 3056 37156
rect 3112 37100 3180 37156
rect 3236 37100 3304 37156
rect 3360 37100 3428 37156
rect 3484 37100 3552 37156
rect 3608 37100 3676 37156
rect 3732 37100 3800 37156
rect 3856 37100 3924 37156
rect 3980 37100 4048 37156
rect 4104 37100 4172 37156
rect 4228 37100 4296 37156
rect 4352 37100 4420 37156
rect 4476 37100 4544 37156
rect 4600 37100 4668 37156
rect 4724 37100 4734 37156
rect 2798 37032 4734 37100
rect 2798 36976 2808 37032
rect 2864 36976 2932 37032
rect 2988 36976 3056 37032
rect 3112 36976 3180 37032
rect 3236 36976 3304 37032
rect 3360 36976 3428 37032
rect 3484 36976 3552 37032
rect 3608 36976 3676 37032
rect 3732 36976 3800 37032
rect 3856 36976 3924 37032
rect 3980 36976 4048 37032
rect 4104 36976 4172 37032
rect 4228 36976 4296 37032
rect 4352 36976 4420 37032
rect 4476 36976 4544 37032
rect 4600 36976 4668 37032
rect 4724 36976 4734 37032
rect 2798 36908 4734 36976
rect 2798 36852 2808 36908
rect 2864 36852 2932 36908
rect 2988 36852 3056 36908
rect 3112 36852 3180 36908
rect 3236 36852 3304 36908
rect 3360 36852 3428 36908
rect 3484 36852 3552 36908
rect 3608 36852 3676 36908
rect 3732 36852 3800 36908
rect 3856 36852 3924 36908
rect 3980 36852 4048 36908
rect 4104 36852 4172 36908
rect 4228 36852 4296 36908
rect 4352 36852 4420 36908
rect 4476 36852 4544 36908
rect 4600 36852 4668 36908
rect 4724 36852 4734 36908
rect 2798 36842 4734 36852
rect 5168 38148 7104 38158
rect 5168 38092 5178 38148
rect 5234 38092 5302 38148
rect 5358 38092 5426 38148
rect 5482 38092 5550 38148
rect 5606 38092 5674 38148
rect 5730 38092 5798 38148
rect 5854 38092 5922 38148
rect 5978 38092 6046 38148
rect 6102 38092 6170 38148
rect 6226 38092 6294 38148
rect 6350 38092 6418 38148
rect 6474 38092 6542 38148
rect 6598 38092 6666 38148
rect 6722 38092 6790 38148
rect 6846 38092 6914 38148
rect 6970 38092 7038 38148
rect 7094 38092 7104 38148
rect 5168 38024 7104 38092
rect 5168 37968 5178 38024
rect 5234 37968 5302 38024
rect 5358 37968 5426 38024
rect 5482 37968 5550 38024
rect 5606 37968 5674 38024
rect 5730 37968 5798 38024
rect 5854 37968 5922 38024
rect 5978 37968 6046 38024
rect 6102 37968 6170 38024
rect 6226 37968 6294 38024
rect 6350 37968 6418 38024
rect 6474 37968 6542 38024
rect 6598 37968 6666 38024
rect 6722 37968 6790 38024
rect 6846 37968 6914 38024
rect 6970 37968 7038 38024
rect 7094 37968 7104 38024
rect 5168 37900 7104 37968
rect 5168 37844 5178 37900
rect 5234 37844 5302 37900
rect 5358 37844 5426 37900
rect 5482 37844 5550 37900
rect 5606 37844 5674 37900
rect 5730 37844 5798 37900
rect 5854 37844 5922 37900
rect 5978 37844 6046 37900
rect 6102 37844 6170 37900
rect 6226 37844 6294 37900
rect 6350 37844 6418 37900
rect 6474 37844 6542 37900
rect 6598 37844 6666 37900
rect 6722 37844 6790 37900
rect 6846 37844 6914 37900
rect 6970 37844 7038 37900
rect 7094 37844 7104 37900
rect 5168 37776 7104 37844
rect 5168 37720 5178 37776
rect 5234 37720 5302 37776
rect 5358 37720 5426 37776
rect 5482 37720 5550 37776
rect 5606 37720 5674 37776
rect 5730 37720 5798 37776
rect 5854 37720 5922 37776
rect 5978 37720 6046 37776
rect 6102 37720 6170 37776
rect 6226 37720 6294 37776
rect 6350 37720 6418 37776
rect 6474 37720 6542 37776
rect 6598 37720 6666 37776
rect 6722 37720 6790 37776
rect 6846 37720 6914 37776
rect 6970 37720 7038 37776
rect 7094 37720 7104 37776
rect 5168 37652 7104 37720
rect 5168 37596 5178 37652
rect 5234 37596 5302 37652
rect 5358 37596 5426 37652
rect 5482 37596 5550 37652
rect 5606 37596 5674 37652
rect 5730 37596 5798 37652
rect 5854 37596 5922 37652
rect 5978 37596 6046 37652
rect 6102 37596 6170 37652
rect 6226 37596 6294 37652
rect 6350 37596 6418 37652
rect 6474 37596 6542 37652
rect 6598 37596 6666 37652
rect 6722 37596 6790 37652
rect 6846 37596 6914 37652
rect 6970 37596 7038 37652
rect 7094 37596 7104 37652
rect 5168 37528 7104 37596
rect 5168 37472 5178 37528
rect 5234 37472 5302 37528
rect 5358 37472 5426 37528
rect 5482 37472 5550 37528
rect 5606 37472 5674 37528
rect 5730 37472 5798 37528
rect 5854 37472 5922 37528
rect 5978 37472 6046 37528
rect 6102 37472 6170 37528
rect 6226 37472 6294 37528
rect 6350 37472 6418 37528
rect 6474 37472 6542 37528
rect 6598 37472 6666 37528
rect 6722 37472 6790 37528
rect 6846 37472 6914 37528
rect 6970 37472 7038 37528
rect 7094 37472 7104 37528
rect 5168 37404 7104 37472
rect 5168 37348 5178 37404
rect 5234 37348 5302 37404
rect 5358 37348 5426 37404
rect 5482 37348 5550 37404
rect 5606 37348 5674 37404
rect 5730 37348 5798 37404
rect 5854 37348 5922 37404
rect 5978 37348 6046 37404
rect 6102 37348 6170 37404
rect 6226 37348 6294 37404
rect 6350 37348 6418 37404
rect 6474 37348 6542 37404
rect 6598 37348 6666 37404
rect 6722 37348 6790 37404
rect 6846 37348 6914 37404
rect 6970 37348 7038 37404
rect 7094 37348 7104 37404
rect 5168 37280 7104 37348
rect 5168 37224 5178 37280
rect 5234 37224 5302 37280
rect 5358 37224 5426 37280
rect 5482 37224 5550 37280
rect 5606 37224 5674 37280
rect 5730 37224 5798 37280
rect 5854 37224 5922 37280
rect 5978 37224 6046 37280
rect 6102 37224 6170 37280
rect 6226 37224 6294 37280
rect 6350 37224 6418 37280
rect 6474 37224 6542 37280
rect 6598 37224 6666 37280
rect 6722 37224 6790 37280
rect 6846 37224 6914 37280
rect 6970 37224 7038 37280
rect 7094 37224 7104 37280
rect 5168 37156 7104 37224
rect 5168 37100 5178 37156
rect 5234 37100 5302 37156
rect 5358 37100 5426 37156
rect 5482 37100 5550 37156
rect 5606 37100 5674 37156
rect 5730 37100 5798 37156
rect 5854 37100 5922 37156
rect 5978 37100 6046 37156
rect 6102 37100 6170 37156
rect 6226 37100 6294 37156
rect 6350 37100 6418 37156
rect 6474 37100 6542 37156
rect 6598 37100 6666 37156
rect 6722 37100 6790 37156
rect 6846 37100 6914 37156
rect 6970 37100 7038 37156
rect 7094 37100 7104 37156
rect 5168 37032 7104 37100
rect 5168 36976 5178 37032
rect 5234 36976 5302 37032
rect 5358 36976 5426 37032
rect 5482 36976 5550 37032
rect 5606 36976 5674 37032
rect 5730 36976 5798 37032
rect 5854 36976 5922 37032
rect 5978 36976 6046 37032
rect 6102 36976 6170 37032
rect 6226 36976 6294 37032
rect 6350 36976 6418 37032
rect 6474 36976 6542 37032
rect 6598 36976 6666 37032
rect 6722 36976 6790 37032
rect 6846 36976 6914 37032
rect 6970 36976 7038 37032
rect 7094 36976 7104 37032
rect 5168 36908 7104 36976
rect 5168 36852 5178 36908
rect 5234 36852 5302 36908
rect 5358 36852 5426 36908
rect 5482 36852 5550 36908
rect 5606 36852 5674 36908
rect 5730 36852 5798 36908
rect 5854 36852 5922 36908
rect 5978 36852 6046 36908
rect 6102 36852 6170 36908
rect 6226 36852 6294 36908
rect 6350 36852 6418 36908
rect 6474 36852 6542 36908
rect 6598 36852 6666 36908
rect 6722 36852 6790 36908
rect 6846 36852 6914 36908
rect 6970 36852 7038 36908
rect 7094 36852 7104 36908
rect 5168 36842 7104 36852
rect 7874 38148 9810 38158
rect 7874 38092 7884 38148
rect 7940 38092 8008 38148
rect 8064 38092 8132 38148
rect 8188 38092 8256 38148
rect 8312 38092 8380 38148
rect 8436 38092 8504 38148
rect 8560 38092 8628 38148
rect 8684 38092 8752 38148
rect 8808 38092 8876 38148
rect 8932 38092 9000 38148
rect 9056 38092 9124 38148
rect 9180 38092 9248 38148
rect 9304 38092 9372 38148
rect 9428 38092 9496 38148
rect 9552 38092 9620 38148
rect 9676 38092 9744 38148
rect 9800 38092 9810 38148
rect 7874 38024 9810 38092
rect 7874 37968 7884 38024
rect 7940 37968 8008 38024
rect 8064 37968 8132 38024
rect 8188 37968 8256 38024
rect 8312 37968 8380 38024
rect 8436 37968 8504 38024
rect 8560 37968 8628 38024
rect 8684 37968 8752 38024
rect 8808 37968 8876 38024
rect 8932 37968 9000 38024
rect 9056 37968 9124 38024
rect 9180 37968 9248 38024
rect 9304 37968 9372 38024
rect 9428 37968 9496 38024
rect 9552 37968 9620 38024
rect 9676 37968 9744 38024
rect 9800 37968 9810 38024
rect 7874 37900 9810 37968
rect 7874 37844 7884 37900
rect 7940 37844 8008 37900
rect 8064 37844 8132 37900
rect 8188 37844 8256 37900
rect 8312 37844 8380 37900
rect 8436 37844 8504 37900
rect 8560 37844 8628 37900
rect 8684 37844 8752 37900
rect 8808 37844 8876 37900
rect 8932 37844 9000 37900
rect 9056 37844 9124 37900
rect 9180 37844 9248 37900
rect 9304 37844 9372 37900
rect 9428 37844 9496 37900
rect 9552 37844 9620 37900
rect 9676 37844 9744 37900
rect 9800 37844 9810 37900
rect 7874 37776 9810 37844
rect 7874 37720 7884 37776
rect 7940 37720 8008 37776
rect 8064 37720 8132 37776
rect 8188 37720 8256 37776
rect 8312 37720 8380 37776
rect 8436 37720 8504 37776
rect 8560 37720 8628 37776
rect 8684 37720 8752 37776
rect 8808 37720 8876 37776
rect 8932 37720 9000 37776
rect 9056 37720 9124 37776
rect 9180 37720 9248 37776
rect 9304 37720 9372 37776
rect 9428 37720 9496 37776
rect 9552 37720 9620 37776
rect 9676 37720 9744 37776
rect 9800 37720 9810 37776
rect 7874 37652 9810 37720
rect 7874 37596 7884 37652
rect 7940 37596 8008 37652
rect 8064 37596 8132 37652
rect 8188 37596 8256 37652
rect 8312 37596 8380 37652
rect 8436 37596 8504 37652
rect 8560 37596 8628 37652
rect 8684 37596 8752 37652
rect 8808 37596 8876 37652
rect 8932 37596 9000 37652
rect 9056 37596 9124 37652
rect 9180 37596 9248 37652
rect 9304 37596 9372 37652
rect 9428 37596 9496 37652
rect 9552 37596 9620 37652
rect 9676 37596 9744 37652
rect 9800 37596 9810 37652
rect 7874 37528 9810 37596
rect 7874 37472 7884 37528
rect 7940 37472 8008 37528
rect 8064 37472 8132 37528
rect 8188 37472 8256 37528
rect 8312 37472 8380 37528
rect 8436 37472 8504 37528
rect 8560 37472 8628 37528
rect 8684 37472 8752 37528
rect 8808 37472 8876 37528
rect 8932 37472 9000 37528
rect 9056 37472 9124 37528
rect 9180 37472 9248 37528
rect 9304 37472 9372 37528
rect 9428 37472 9496 37528
rect 9552 37472 9620 37528
rect 9676 37472 9744 37528
rect 9800 37472 9810 37528
rect 7874 37404 9810 37472
rect 7874 37348 7884 37404
rect 7940 37348 8008 37404
rect 8064 37348 8132 37404
rect 8188 37348 8256 37404
rect 8312 37348 8380 37404
rect 8436 37348 8504 37404
rect 8560 37348 8628 37404
rect 8684 37348 8752 37404
rect 8808 37348 8876 37404
rect 8932 37348 9000 37404
rect 9056 37348 9124 37404
rect 9180 37348 9248 37404
rect 9304 37348 9372 37404
rect 9428 37348 9496 37404
rect 9552 37348 9620 37404
rect 9676 37348 9744 37404
rect 9800 37348 9810 37404
rect 7874 37280 9810 37348
rect 7874 37224 7884 37280
rect 7940 37224 8008 37280
rect 8064 37224 8132 37280
rect 8188 37224 8256 37280
rect 8312 37224 8380 37280
rect 8436 37224 8504 37280
rect 8560 37224 8628 37280
rect 8684 37224 8752 37280
rect 8808 37224 8876 37280
rect 8932 37224 9000 37280
rect 9056 37224 9124 37280
rect 9180 37224 9248 37280
rect 9304 37224 9372 37280
rect 9428 37224 9496 37280
rect 9552 37224 9620 37280
rect 9676 37224 9744 37280
rect 9800 37224 9810 37280
rect 7874 37156 9810 37224
rect 7874 37100 7884 37156
rect 7940 37100 8008 37156
rect 8064 37100 8132 37156
rect 8188 37100 8256 37156
rect 8312 37100 8380 37156
rect 8436 37100 8504 37156
rect 8560 37100 8628 37156
rect 8684 37100 8752 37156
rect 8808 37100 8876 37156
rect 8932 37100 9000 37156
rect 9056 37100 9124 37156
rect 9180 37100 9248 37156
rect 9304 37100 9372 37156
rect 9428 37100 9496 37156
rect 9552 37100 9620 37156
rect 9676 37100 9744 37156
rect 9800 37100 9810 37156
rect 7874 37032 9810 37100
rect 7874 36976 7884 37032
rect 7940 36976 8008 37032
rect 8064 36976 8132 37032
rect 8188 36976 8256 37032
rect 8312 36976 8380 37032
rect 8436 36976 8504 37032
rect 8560 36976 8628 37032
rect 8684 36976 8752 37032
rect 8808 36976 8876 37032
rect 8932 36976 9000 37032
rect 9056 36976 9124 37032
rect 9180 36976 9248 37032
rect 9304 36976 9372 37032
rect 9428 36976 9496 37032
rect 9552 36976 9620 37032
rect 9676 36976 9744 37032
rect 9800 36976 9810 37032
rect 7874 36908 9810 36976
rect 7874 36852 7884 36908
rect 7940 36852 8008 36908
rect 8064 36852 8132 36908
rect 8188 36852 8256 36908
rect 8312 36852 8380 36908
rect 8436 36852 8504 36908
rect 8560 36852 8628 36908
rect 8684 36852 8752 36908
rect 8808 36852 8876 36908
rect 8932 36852 9000 36908
rect 9056 36852 9124 36908
rect 9180 36852 9248 36908
rect 9304 36852 9372 36908
rect 9428 36852 9496 36908
rect 9552 36852 9620 36908
rect 9676 36852 9744 36908
rect 9800 36852 9810 36908
rect 7874 36842 9810 36852
rect 10244 38148 12180 38158
rect 10244 38092 10254 38148
rect 10310 38092 10378 38148
rect 10434 38092 10502 38148
rect 10558 38092 10626 38148
rect 10682 38092 10750 38148
rect 10806 38092 10874 38148
rect 10930 38092 10998 38148
rect 11054 38092 11122 38148
rect 11178 38092 11246 38148
rect 11302 38092 11370 38148
rect 11426 38092 11494 38148
rect 11550 38092 11618 38148
rect 11674 38092 11742 38148
rect 11798 38092 11866 38148
rect 11922 38092 11990 38148
rect 12046 38092 12114 38148
rect 12170 38092 12180 38148
rect 10244 38024 12180 38092
rect 10244 37968 10254 38024
rect 10310 37968 10378 38024
rect 10434 37968 10502 38024
rect 10558 37968 10626 38024
rect 10682 37968 10750 38024
rect 10806 37968 10874 38024
rect 10930 37968 10998 38024
rect 11054 37968 11122 38024
rect 11178 37968 11246 38024
rect 11302 37968 11370 38024
rect 11426 37968 11494 38024
rect 11550 37968 11618 38024
rect 11674 37968 11742 38024
rect 11798 37968 11866 38024
rect 11922 37968 11990 38024
rect 12046 37968 12114 38024
rect 12170 37968 12180 38024
rect 10244 37900 12180 37968
rect 10244 37844 10254 37900
rect 10310 37844 10378 37900
rect 10434 37844 10502 37900
rect 10558 37844 10626 37900
rect 10682 37844 10750 37900
rect 10806 37844 10874 37900
rect 10930 37844 10998 37900
rect 11054 37844 11122 37900
rect 11178 37844 11246 37900
rect 11302 37844 11370 37900
rect 11426 37844 11494 37900
rect 11550 37844 11618 37900
rect 11674 37844 11742 37900
rect 11798 37844 11866 37900
rect 11922 37844 11990 37900
rect 12046 37844 12114 37900
rect 12170 37844 12180 37900
rect 10244 37776 12180 37844
rect 10244 37720 10254 37776
rect 10310 37720 10378 37776
rect 10434 37720 10502 37776
rect 10558 37720 10626 37776
rect 10682 37720 10750 37776
rect 10806 37720 10874 37776
rect 10930 37720 10998 37776
rect 11054 37720 11122 37776
rect 11178 37720 11246 37776
rect 11302 37720 11370 37776
rect 11426 37720 11494 37776
rect 11550 37720 11618 37776
rect 11674 37720 11742 37776
rect 11798 37720 11866 37776
rect 11922 37720 11990 37776
rect 12046 37720 12114 37776
rect 12170 37720 12180 37776
rect 10244 37652 12180 37720
rect 10244 37596 10254 37652
rect 10310 37596 10378 37652
rect 10434 37596 10502 37652
rect 10558 37596 10626 37652
rect 10682 37596 10750 37652
rect 10806 37596 10874 37652
rect 10930 37596 10998 37652
rect 11054 37596 11122 37652
rect 11178 37596 11246 37652
rect 11302 37596 11370 37652
rect 11426 37596 11494 37652
rect 11550 37596 11618 37652
rect 11674 37596 11742 37652
rect 11798 37596 11866 37652
rect 11922 37596 11990 37652
rect 12046 37596 12114 37652
rect 12170 37596 12180 37652
rect 10244 37528 12180 37596
rect 10244 37472 10254 37528
rect 10310 37472 10378 37528
rect 10434 37472 10502 37528
rect 10558 37472 10626 37528
rect 10682 37472 10750 37528
rect 10806 37472 10874 37528
rect 10930 37472 10998 37528
rect 11054 37472 11122 37528
rect 11178 37472 11246 37528
rect 11302 37472 11370 37528
rect 11426 37472 11494 37528
rect 11550 37472 11618 37528
rect 11674 37472 11742 37528
rect 11798 37472 11866 37528
rect 11922 37472 11990 37528
rect 12046 37472 12114 37528
rect 12170 37472 12180 37528
rect 10244 37404 12180 37472
rect 10244 37348 10254 37404
rect 10310 37348 10378 37404
rect 10434 37348 10502 37404
rect 10558 37348 10626 37404
rect 10682 37348 10750 37404
rect 10806 37348 10874 37404
rect 10930 37348 10998 37404
rect 11054 37348 11122 37404
rect 11178 37348 11246 37404
rect 11302 37348 11370 37404
rect 11426 37348 11494 37404
rect 11550 37348 11618 37404
rect 11674 37348 11742 37404
rect 11798 37348 11866 37404
rect 11922 37348 11990 37404
rect 12046 37348 12114 37404
rect 12170 37348 12180 37404
rect 10244 37280 12180 37348
rect 10244 37224 10254 37280
rect 10310 37224 10378 37280
rect 10434 37224 10502 37280
rect 10558 37224 10626 37280
rect 10682 37224 10750 37280
rect 10806 37224 10874 37280
rect 10930 37224 10998 37280
rect 11054 37224 11122 37280
rect 11178 37224 11246 37280
rect 11302 37224 11370 37280
rect 11426 37224 11494 37280
rect 11550 37224 11618 37280
rect 11674 37224 11742 37280
rect 11798 37224 11866 37280
rect 11922 37224 11990 37280
rect 12046 37224 12114 37280
rect 12170 37224 12180 37280
rect 10244 37156 12180 37224
rect 10244 37100 10254 37156
rect 10310 37100 10378 37156
rect 10434 37100 10502 37156
rect 10558 37100 10626 37156
rect 10682 37100 10750 37156
rect 10806 37100 10874 37156
rect 10930 37100 10998 37156
rect 11054 37100 11122 37156
rect 11178 37100 11246 37156
rect 11302 37100 11370 37156
rect 11426 37100 11494 37156
rect 11550 37100 11618 37156
rect 11674 37100 11742 37156
rect 11798 37100 11866 37156
rect 11922 37100 11990 37156
rect 12046 37100 12114 37156
rect 12170 37100 12180 37156
rect 10244 37032 12180 37100
rect 10244 36976 10254 37032
rect 10310 36976 10378 37032
rect 10434 36976 10502 37032
rect 10558 36976 10626 37032
rect 10682 36976 10750 37032
rect 10806 36976 10874 37032
rect 10930 36976 10998 37032
rect 11054 36976 11122 37032
rect 11178 36976 11246 37032
rect 11302 36976 11370 37032
rect 11426 36976 11494 37032
rect 11550 36976 11618 37032
rect 11674 36976 11742 37032
rect 11798 36976 11866 37032
rect 11922 36976 11990 37032
rect 12046 36976 12114 37032
rect 12170 36976 12180 37032
rect 10244 36908 12180 36976
rect 10244 36852 10254 36908
rect 10310 36852 10378 36908
rect 10434 36852 10502 36908
rect 10558 36852 10626 36908
rect 10682 36852 10750 36908
rect 10806 36852 10874 36908
rect 10930 36852 10998 36908
rect 11054 36852 11122 36908
rect 11178 36852 11246 36908
rect 11302 36852 11370 36908
rect 11426 36852 11494 36908
rect 11550 36852 11618 36908
rect 11674 36852 11742 36908
rect 11798 36852 11866 36908
rect 11922 36852 11990 36908
rect 12046 36852 12114 36908
rect 12170 36852 12180 36908
rect 10244 36842 12180 36852
rect 12861 38148 14673 38158
rect 12861 38092 12871 38148
rect 12927 38092 12995 38148
rect 13051 38092 13119 38148
rect 13175 38092 13243 38148
rect 13299 38092 13367 38148
rect 13423 38092 13491 38148
rect 13547 38092 13615 38148
rect 13671 38092 13739 38148
rect 13795 38092 13863 38148
rect 13919 38092 13987 38148
rect 14043 38092 14111 38148
rect 14167 38092 14235 38148
rect 14291 38092 14359 38148
rect 14415 38092 14483 38148
rect 14539 38092 14607 38148
rect 14663 38092 14673 38148
rect 12861 38024 14673 38092
rect 12861 37968 12871 38024
rect 12927 37968 12995 38024
rect 13051 37968 13119 38024
rect 13175 37968 13243 38024
rect 13299 37968 13367 38024
rect 13423 37968 13491 38024
rect 13547 37968 13615 38024
rect 13671 37968 13739 38024
rect 13795 37968 13863 38024
rect 13919 37968 13987 38024
rect 14043 37968 14111 38024
rect 14167 37968 14235 38024
rect 14291 37968 14359 38024
rect 14415 37968 14483 38024
rect 14539 37968 14607 38024
rect 14663 37968 14673 38024
rect 12861 37900 14673 37968
rect 12861 37844 12871 37900
rect 12927 37844 12995 37900
rect 13051 37844 13119 37900
rect 13175 37844 13243 37900
rect 13299 37844 13367 37900
rect 13423 37844 13491 37900
rect 13547 37844 13615 37900
rect 13671 37844 13739 37900
rect 13795 37844 13863 37900
rect 13919 37844 13987 37900
rect 14043 37844 14111 37900
rect 14167 37844 14235 37900
rect 14291 37844 14359 37900
rect 14415 37844 14483 37900
rect 14539 37844 14607 37900
rect 14663 37844 14673 37900
rect 12861 37776 14673 37844
rect 12861 37720 12871 37776
rect 12927 37720 12995 37776
rect 13051 37720 13119 37776
rect 13175 37720 13243 37776
rect 13299 37720 13367 37776
rect 13423 37720 13491 37776
rect 13547 37720 13615 37776
rect 13671 37720 13739 37776
rect 13795 37720 13863 37776
rect 13919 37720 13987 37776
rect 14043 37720 14111 37776
rect 14167 37720 14235 37776
rect 14291 37720 14359 37776
rect 14415 37720 14483 37776
rect 14539 37720 14607 37776
rect 14663 37720 14673 37776
rect 12861 37652 14673 37720
rect 12861 37596 12871 37652
rect 12927 37596 12995 37652
rect 13051 37596 13119 37652
rect 13175 37596 13243 37652
rect 13299 37596 13367 37652
rect 13423 37596 13491 37652
rect 13547 37596 13615 37652
rect 13671 37596 13739 37652
rect 13795 37596 13863 37652
rect 13919 37596 13987 37652
rect 14043 37596 14111 37652
rect 14167 37596 14235 37652
rect 14291 37596 14359 37652
rect 14415 37596 14483 37652
rect 14539 37596 14607 37652
rect 14663 37596 14673 37652
rect 12861 37528 14673 37596
rect 12861 37472 12871 37528
rect 12927 37472 12995 37528
rect 13051 37472 13119 37528
rect 13175 37472 13243 37528
rect 13299 37472 13367 37528
rect 13423 37472 13491 37528
rect 13547 37472 13615 37528
rect 13671 37472 13739 37528
rect 13795 37472 13863 37528
rect 13919 37472 13987 37528
rect 14043 37472 14111 37528
rect 14167 37472 14235 37528
rect 14291 37472 14359 37528
rect 14415 37472 14483 37528
rect 14539 37472 14607 37528
rect 14663 37472 14673 37528
rect 12861 37404 14673 37472
rect 12861 37348 12871 37404
rect 12927 37348 12995 37404
rect 13051 37348 13119 37404
rect 13175 37348 13243 37404
rect 13299 37348 13367 37404
rect 13423 37348 13491 37404
rect 13547 37348 13615 37404
rect 13671 37348 13739 37404
rect 13795 37348 13863 37404
rect 13919 37348 13987 37404
rect 14043 37348 14111 37404
rect 14167 37348 14235 37404
rect 14291 37348 14359 37404
rect 14415 37348 14483 37404
rect 14539 37348 14607 37404
rect 14663 37348 14673 37404
rect 12861 37280 14673 37348
rect 12861 37224 12871 37280
rect 12927 37224 12995 37280
rect 13051 37224 13119 37280
rect 13175 37224 13243 37280
rect 13299 37224 13367 37280
rect 13423 37224 13491 37280
rect 13547 37224 13615 37280
rect 13671 37224 13739 37280
rect 13795 37224 13863 37280
rect 13919 37224 13987 37280
rect 14043 37224 14111 37280
rect 14167 37224 14235 37280
rect 14291 37224 14359 37280
rect 14415 37224 14483 37280
rect 14539 37224 14607 37280
rect 14663 37224 14673 37280
rect 12861 37156 14673 37224
rect 12861 37100 12871 37156
rect 12927 37100 12995 37156
rect 13051 37100 13119 37156
rect 13175 37100 13243 37156
rect 13299 37100 13367 37156
rect 13423 37100 13491 37156
rect 13547 37100 13615 37156
rect 13671 37100 13739 37156
rect 13795 37100 13863 37156
rect 13919 37100 13987 37156
rect 14043 37100 14111 37156
rect 14167 37100 14235 37156
rect 14291 37100 14359 37156
rect 14415 37100 14483 37156
rect 14539 37100 14607 37156
rect 14663 37100 14673 37156
rect 12861 37032 14673 37100
rect 12861 36976 12871 37032
rect 12927 36976 12995 37032
rect 13051 36976 13119 37032
rect 13175 36976 13243 37032
rect 13299 36976 13367 37032
rect 13423 36976 13491 37032
rect 13547 36976 13615 37032
rect 13671 36976 13739 37032
rect 13795 36976 13863 37032
rect 13919 36976 13987 37032
rect 14043 36976 14111 37032
rect 14167 36976 14235 37032
rect 14291 36976 14359 37032
rect 14415 36976 14483 37032
rect 14539 36976 14607 37032
rect 14663 36976 14673 37032
rect 12861 36908 14673 36976
rect 12861 36852 12871 36908
rect 12927 36852 12995 36908
rect 13051 36852 13119 36908
rect 13175 36852 13243 36908
rect 13299 36852 13367 36908
rect 13423 36852 13491 36908
rect 13547 36852 13615 36908
rect 13671 36852 13739 36908
rect 13795 36852 13863 36908
rect 13919 36852 13987 36908
rect 14043 36852 14111 36908
rect 14167 36852 14235 36908
rect 14291 36852 14359 36908
rect 14415 36852 14483 36908
rect 14539 36852 14607 36908
rect 14663 36852 14673 36908
rect 12861 36842 14673 36852
rect 10 36814 86 36824
rect 14892 36824 14902 38176
rect 14958 36824 14968 38176
rect 14892 36814 14968 36824
rect 10 36586 86 36596
rect 10 33614 20 36586
rect 76 33614 86 36586
rect 14892 36586 14968 36596
rect 305 36554 2117 36564
rect 305 36498 315 36554
rect 371 36498 439 36554
rect 495 36498 563 36554
rect 619 36498 687 36554
rect 743 36498 811 36554
rect 867 36498 935 36554
rect 991 36498 1059 36554
rect 1115 36498 1183 36554
rect 1239 36498 1307 36554
rect 1363 36498 1431 36554
rect 1487 36498 1555 36554
rect 1611 36498 1679 36554
rect 1735 36498 1803 36554
rect 1859 36498 1927 36554
rect 1983 36498 2051 36554
rect 2107 36498 2117 36554
rect 305 36430 2117 36498
rect 305 36374 315 36430
rect 371 36374 439 36430
rect 495 36374 563 36430
rect 619 36374 687 36430
rect 743 36374 811 36430
rect 867 36374 935 36430
rect 991 36374 1059 36430
rect 1115 36374 1183 36430
rect 1239 36374 1307 36430
rect 1363 36374 1431 36430
rect 1487 36374 1555 36430
rect 1611 36374 1679 36430
rect 1735 36374 1803 36430
rect 1859 36374 1927 36430
rect 1983 36374 2051 36430
rect 2107 36374 2117 36430
rect 305 36306 2117 36374
rect 305 36250 315 36306
rect 371 36250 439 36306
rect 495 36250 563 36306
rect 619 36250 687 36306
rect 743 36250 811 36306
rect 867 36250 935 36306
rect 991 36250 1059 36306
rect 1115 36250 1183 36306
rect 1239 36250 1307 36306
rect 1363 36250 1431 36306
rect 1487 36250 1555 36306
rect 1611 36250 1679 36306
rect 1735 36250 1803 36306
rect 1859 36250 1927 36306
rect 1983 36250 2051 36306
rect 2107 36250 2117 36306
rect 305 36182 2117 36250
rect 305 36126 315 36182
rect 371 36126 439 36182
rect 495 36126 563 36182
rect 619 36126 687 36182
rect 743 36126 811 36182
rect 867 36126 935 36182
rect 991 36126 1059 36182
rect 1115 36126 1183 36182
rect 1239 36126 1307 36182
rect 1363 36126 1431 36182
rect 1487 36126 1555 36182
rect 1611 36126 1679 36182
rect 1735 36126 1803 36182
rect 1859 36126 1927 36182
rect 1983 36126 2051 36182
rect 2107 36126 2117 36182
rect 305 36058 2117 36126
rect 305 36002 315 36058
rect 371 36002 439 36058
rect 495 36002 563 36058
rect 619 36002 687 36058
rect 743 36002 811 36058
rect 867 36002 935 36058
rect 991 36002 1059 36058
rect 1115 36002 1183 36058
rect 1239 36002 1307 36058
rect 1363 36002 1431 36058
rect 1487 36002 1555 36058
rect 1611 36002 1679 36058
rect 1735 36002 1803 36058
rect 1859 36002 1927 36058
rect 1983 36002 2051 36058
rect 2107 36002 2117 36058
rect 305 35934 2117 36002
rect 305 35878 315 35934
rect 371 35878 439 35934
rect 495 35878 563 35934
rect 619 35878 687 35934
rect 743 35878 811 35934
rect 867 35878 935 35934
rect 991 35878 1059 35934
rect 1115 35878 1183 35934
rect 1239 35878 1307 35934
rect 1363 35878 1431 35934
rect 1487 35878 1555 35934
rect 1611 35878 1679 35934
rect 1735 35878 1803 35934
rect 1859 35878 1927 35934
rect 1983 35878 2051 35934
rect 2107 35878 2117 35934
rect 305 35810 2117 35878
rect 305 35754 315 35810
rect 371 35754 439 35810
rect 495 35754 563 35810
rect 619 35754 687 35810
rect 743 35754 811 35810
rect 867 35754 935 35810
rect 991 35754 1059 35810
rect 1115 35754 1183 35810
rect 1239 35754 1307 35810
rect 1363 35754 1431 35810
rect 1487 35754 1555 35810
rect 1611 35754 1679 35810
rect 1735 35754 1803 35810
rect 1859 35754 1927 35810
rect 1983 35754 2051 35810
rect 2107 35754 2117 35810
rect 305 35686 2117 35754
rect 305 35630 315 35686
rect 371 35630 439 35686
rect 495 35630 563 35686
rect 619 35630 687 35686
rect 743 35630 811 35686
rect 867 35630 935 35686
rect 991 35630 1059 35686
rect 1115 35630 1183 35686
rect 1239 35630 1307 35686
rect 1363 35630 1431 35686
rect 1487 35630 1555 35686
rect 1611 35630 1679 35686
rect 1735 35630 1803 35686
rect 1859 35630 1927 35686
rect 1983 35630 2051 35686
rect 2107 35630 2117 35686
rect 305 35562 2117 35630
rect 305 35506 315 35562
rect 371 35506 439 35562
rect 495 35506 563 35562
rect 619 35506 687 35562
rect 743 35506 811 35562
rect 867 35506 935 35562
rect 991 35506 1059 35562
rect 1115 35506 1183 35562
rect 1239 35506 1307 35562
rect 1363 35506 1431 35562
rect 1487 35506 1555 35562
rect 1611 35506 1679 35562
rect 1735 35506 1803 35562
rect 1859 35506 1927 35562
rect 1983 35506 2051 35562
rect 2107 35506 2117 35562
rect 305 35438 2117 35506
rect 305 35382 315 35438
rect 371 35382 439 35438
rect 495 35382 563 35438
rect 619 35382 687 35438
rect 743 35382 811 35438
rect 867 35382 935 35438
rect 991 35382 1059 35438
rect 1115 35382 1183 35438
rect 1239 35382 1307 35438
rect 1363 35382 1431 35438
rect 1487 35382 1555 35438
rect 1611 35382 1679 35438
rect 1735 35382 1803 35438
rect 1859 35382 1927 35438
rect 1983 35382 2051 35438
rect 2107 35382 2117 35438
rect 305 35314 2117 35382
rect 305 35258 315 35314
rect 371 35258 439 35314
rect 495 35258 563 35314
rect 619 35258 687 35314
rect 743 35258 811 35314
rect 867 35258 935 35314
rect 991 35258 1059 35314
rect 1115 35258 1183 35314
rect 1239 35258 1307 35314
rect 1363 35258 1431 35314
rect 1487 35258 1555 35314
rect 1611 35258 1679 35314
rect 1735 35258 1803 35314
rect 1859 35258 1927 35314
rect 1983 35258 2051 35314
rect 2107 35258 2117 35314
rect 305 35190 2117 35258
rect 305 35134 315 35190
rect 371 35134 439 35190
rect 495 35134 563 35190
rect 619 35134 687 35190
rect 743 35134 811 35190
rect 867 35134 935 35190
rect 991 35134 1059 35190
rect 1115 35134 1183 35190
rect 1239 35134 1307 35190
rect 1363 35134 1431 35190
rect 1487 35134 1555 35190
rect 1611 35134 1679 35190
rect 1735 35134 1803 35190
rect 1859 35134 1927 35190
rect 1983 35134 2051 35190
rect 2107 35134 2117 35190
rect 305 35066 2117 35134
rect 305 35010 315 35066
rect 371 35010 439 35066
rect 495 35010 563 35066
rect 619 35010 687 35066
rect 743 35010 811 35066
rect 867 35010 935 35066
rect 991 35010 1059 35066
rect 1115 35010 1183 35066
rect 1239 35010 1307 35066
rect 1363 35010 1431 35066
rect 1487 35010 1555 35066
rect 1611 35010 1679 35066
rect 1735 35010 1803 35066
rect 1859 35010 1927 35066
rect 1983 35010 2051 35066
rect 2107 35010 2117 35066
rect 305 34942 2117 35010
rect 305 34886 315 34942
rect 371 34886 439 34942
rect 495 34886 563 34942
rect 619 34886 687 34942
rect 743 34886 811 34942
rect 867 34886 935 34942
rect 991 34886 1059 34942
rect 1115 34886 1183 34942
rect 1239 34886 1307 34942
rect 1363 34886 1431 34942
rect 1487 34886 1555 34942
rect 1611 34886 1679 34942
rect 1735 34886 1803 34942
rect 1859 34886 1927 34942
rect 1983 34886 2051 34942
rect 2107 34886 2117 34942
rect 305 34818 2117 34886
rect 305 34762 315 34818
rect 371 34762 439 34818
rect 495 34762 563 34818
rect 619 34762 687 34818
rect 743 34762 811 34818
rect 867 34762 935 34818
rect 991 34762 1059 34818
rect 1115 34762 1183 34818
rect 1239 34762 1307 34818
rect 1363 34762 1431 34818
rect 1487 34762 1555 34818
rect 1611 34762 1679 34818
rect 1735 34762 1803 34818
rect 1859 34762 1927 34818
rect 1983 34762 2051 34818
rect 2107 34762 2117 34818
rect 305 34694 2117 34762
rect 305 34638 315 34694
rect 371 34638 439 34694
rect 495 34638 563 34694
rect 619 34638 687 34694
rect 743 34638 811 34694
rect 867 34638 935 34694
rect 991 34638 1059 34694
rect 1115 34638 1183 34694
rect 1239 34638 1307 34694
rect 1363 34638 1431 34694
rect 1487 34638 1555 34694
rect 1611 34638 1679 34694
rect 1735 34638 1803 34694
rect 1859 34638 1927 34694
rect 1983 34638 2051 34694
rect 2107 34638 2117 34694
rect 305 34570 2117 34638
rect 305 34514 315 34570
rect 371 34514 439 34570
rect 495 34514 563 34570
rect 619 34514 687 34570
rect 743 34514 811 34570
rect 867 34514 935 34570
rect 991 34514 1059 34570
rect 1115 34514 1183 34570
rect 1239 34514 1307 34570
rect 1363 34514 1431 34570
rect 1487 34514 1555 34570
rect 1611 34514 1679 34570
rect 1735 34514 1803 34570
rect 1859 34514 1927 34570
rect 1983 34514 2051 34570
rect 2107 34514 2117 34570
rect 305 34446 2117 34514
rect 305 34390 315 34446
rect 371 34390 439 34446
rect 495 34390 563 34446
rect 619 34390 687 34446
rect 743 34390 811 34446
rect 867 34390 935 34446
rect 991 34390 1059 34446
rect 1115 34390 1183 34446
rect 1239 34390 1307 34446
rect 1363 34390 1431 34446
rect 1487 34390 1555 34446
rect 1611 34390 1679 34446
rect 1735 34390 1803 34446
rect 1859 34390 1927 34446
rect 1983 34390 2051 34446
rect 2107 34390 2117 34446
rect 305 34322 2117 34390
rect 305 34266 315 34322
rect 371 34266 439 34322
rect 495 34266 563 34322
rect 619 34266 687 34322
rect 743 34266 811 34322
rect 867 34266 935 34322
rect 991 34266 1059 34322
rect 1115 34266 1183 34322
rect 1239 34266 1307 34322
rect 1363 34266 1431 34322
rect 1487 34266 1555 34322
rect 1611 34266 1679 34322
rect 1735 34266 1803 34322
rect 1859 34266 1927 34322
rect 1983 34266 2051 34322
rect 2107 34266 2117 34322
rect 305 34198 2117 34266
rect 305 34142 315 34198
rect 371 34142 439 34198
rect 495 34142 563 34198
rect 619 34142 687 34198
rect 743 34142 811 34198
rect 867 34142 935 34198
rect 991 34142 1059 34198
rect 1115 34142 1183 34198
rect 1239 34142 1307 34198
rect 1363 34142 1431 34198
rect 1487 34142 1555 34198
rect 1611 34142 1679 34198
rect 1735 34142 1803 34198
rect 1859 34142 1927 34198
rect 1983 34142 2051 34198
rect 2107 34142 2117 34198
rect 305 34074 2117 34142
rect 305 34018 315 34074
rect 371 34018 439 34074
rect 495 34018 563 34074
rect 619 34018 687 34074
rect 743 34018 811 34074
rect 867 34018 935 34074
rect 991 34018 1059 34074
rect 1115 34018 1183 34074
rect 1239 34018 1307 34074
rect 1363 34018 1431 34074
rect 1487 34018 1555 34074
rect 1611 34018 1679 34074
rect 1735 34018 1803 34074
rect 1859 34018 1927 34074
rect 1983 34018 2051 34074
rect 2107 34018 2117 34074
rect 305 33950 2117 34018
rect 305 33894 315 33950
rect 371 33894 439 33950
rect 495 33894 563 33950
rect 619 33894 687 33950
rect 743 33894 811 33950
rect 867 33894 935 33950
rect 991 33894 1059 33950
rect 1115 33894 1183 33950
rect 1239 33894 1307 33950
rect 1363 33894 1431 33950
rect 1487 33894 1555 33950
rect 1611 33894 1679 33950
rect 1735 33894 1803 33950
rect 1859 33894 1927 33950
rect 1983 33894 2051 33950
rect 2107 33894 2117 33950
rect 305 33826 2117 33894
rect 305 33770 315 33826
rect 371 33770 439 33826
rect 495 33770 563 33826
rect 619 33770 687 33826
rect 743 33770 811 33826
rect 867 33770 935 33826
rect 991 33770 1059 33826
rect 1115 33770 1183 33826
rect 1239 33770 1307 33826
rect 1363 33770 1431 33826
rect 1487 33770 1555 33826
rect 1611 33770 1679 33826
rect 1735 33770 1803 33826
rect 1859 33770 1927 33826
rect 1983 33770 2051 33826
rect 2107 33770 2117 33826
rect 305 33702 2117 33770
rect 305 33646 315 33702
rect 371 33646 439 33702
rect 495 33646 563 33702
rect 619 33646 687 33702
rect 743 33646 811 33702
rect 867 33646 935 33702
rect 991 33646 1059 33702
rect 1115 33646 1183 33702
rect 1239 33646 1307 33702
rect 1363 33646 1431 33702
rect 1487 33646 1555 33702
rect 1611 33646 1679 33702
rect 1735 33646 1803 33702
rect 1859 33646 1927 33702
rect 1983 33646 2051 33702
rect 2107 33646 2117 33702
rect 305 33636 2117 33646
rect 2798 36554 4734 36564
rect 2798 36498 2808 36554
rect 2864 36498 2932 36554
rect 2988 36498 3056 36554
rect 3112 36498 3180 36554
rect 3236 36498 3304 36554
rect 3360 36498 3428 36554
rect 3484 36498 3552 36554
rect 3608 36498 3676 36554
rect 3732 36498 3800 36554
rect 3856 36498 3924 36554
rect 3980 36498 4048 36554
rect 4104 36498 4172 36554
rect 4228 36498 4296 36554
rect 4352 36498 4420 36554
rect 4476 36498 4544 36554
rect 4600 36498 4668 36554
rect 4724 36498 4734 36554
rect 2798 36430 4734 36498
rect 2798 36374 2808 36430
rect 2864 36374 2932 36430
rect 2988 36374 3056 36430
rect 3112 36374 3180 36430
rect 3236 36374 3304 36430
rect 3360 36374 3428 36430
rect 3484 36374 3552 36430
rect 3608 36374 3676 36430
rect 3732 36374 3800 36430
rect 3856 36374 3924 36430
rect 3980 36374 4048 36430
rect 4104 36374 4172 36430
rect 4228 36374 4296 36430
rect 4352 36374 4420 36430
rect 4476 36374 4544 36430
rect 4600 36374 4668 36430
rect 4724 36374 4734 36430
rect 2798 36306 4734 36374
rect 2798 36250 2808 36306
rect 2864 36250 2932 36306
rect 2988 36250 3056 36306
rect 3112 36250 3180 36306
rect 3236 36250 3304 36306
rect 3360 36250 3428 36306
rect 3484 36250 3552 36306
rect 3608 36250 3676 36306
rect 3732 36250 3800 36306
rect 3856 36250 3924 36306
rect 3980 36250 4048 36306
rect 4104 36250 4172 36306
rect 4228 36250 4296 36306
rect 4352 36250 4420 36306
rect 4476 36250 4544 36306
rect 4600 36250 4668 36306
rect 4724 36250 4734 36306
rect 2798 36182 4734 36250
rect 2798 36126 2808 36182
rect 2864 36126 2932 36182
rect 2988 36126 3056 36182
rect 3112 36126 3180 36182
rect 3236 36126 3304 36182
rect 3360 36126 3428 36182
rect 3484 36126 3552 36182
rect 3608 36126 3676 36182
rect 3732 36126 3800 36182
rect 3856 36126 3924 36182
rect 3980 36126 4048 36182
rect 4104 36126 4172 36182
rect 4228 36126 4296 36182
rect 4352 36126 4420 36182
rect 4476 36126 4544 36182
rect 4600 36126 4668 36182
rect 4724 36126 4734 36182
rect 2798 36058 4734 36126
rect 2798 36002 2808 36058
rect 2864 36002 2932 36058
rect 2988 36002 3056 36058
rect 3112 36002 3180 36058
rect 3236 36002 3304 36058
rect 3360 36002 3428 36058
rect 3484 36002 3552 36058
rect 3608 36002 3676 36058
rect 3732 36002 3800 36058
rect 3856 36002 3924 36058
rect 3980 36002 4048 36058
rect 4104 36002 4172 36058
rect 4228 36002 4296 36058
rect 4352 36002 4420 36058
rect 4476 36002 4544 36058
rect 4600 36002 4668 36058
rect 4724 36002 4734 36058
rect 2798 35934 4734 36002
rect 2798 35878 2808 35934
rect 2864 35878 2932 35934
rect 2988 35878 3056 35934
rect 3112 35878 3180 35934
rect 3236 35878 3304 35934
rect 3360 35878 3428 35934
rect 3484 35878 3552 35934
rect 3608 35878 3676 35934
rect 3732 35878 3800 35934
rect 3856 35878 3924 35934
rect 3980 35878 4048 35934
rect 4104 35878 4172 35934
rect 4228 35878 4296 35934
rect 4352 35878 4420 35934
rect 4476 35878 4544 35934
rect 4600 35878 4668 35934
rect 4724 35878 4734 35934
rect 2798 35810 4734 35878
rect 2798 35754 2808 35810
rect 2864 35754 2932 35810
rect 2988 35754 3056 35810
rect 3112 35754 3180 35810
rect 3236 35754 3304 35810
rect 3360 35754 3428 35810
rect 3484 35754 3552 35810
rect 3608 35754 3676 35810
rect 3732 35754 3800 35810
rect 3856 35754 3924 35810
rect 3980 35754 4048 35810
rect 4104 35754 4172 35810
rect 4228 35754 4296 35810
rect 4352 35754 4420 35810
rect 4476 35754 4544 35810
rect 4600 35754 4668 35810
rect 4724 35754 4734 35810
rect 2798 35686 4734 35754
rect 2798 35630 2808 35686
rect 2864 35630 2932 35686
rect 2988 35630 3056 35686
rect 3112 35630 3180 35686
rect 3236 35630 3304 35686
rect 3360 35630 3428 35686
rect 3484 35630 3552 35686
rect 3608 35630 3676 35686
rect 3732 35630 3800 35686
rect 3856 35630 3924 35686
rect 3980 35630 4048 35686
rect 4104 35630 4172 35686
rect 4228 35630 4296 35686
rect 4352 35630 4420 35686
rect 4476 35630 4544 35686
rect 4600 35630 4668 35686
rect 4724 35630 4734 35686
rect 2798 35562 4734 35630
rect 2798 35506 2808 35562
rect 2864 35506 2932 35562
rect 2988 35506 3056 35562
rect 3112 35506 3180 35562
rect 3236 35506 3304 35562
rect 3360 35506 3428 35562
rect 3484 35506 3552 35562
rect 3608 35506 3676 35562
rect 3732 35506 3800 35562
rect 3856 35506 3924 35562
rect 3980 35506 4048 35562
rect 4104 35506 4172 35562
rect 4228 35506 4296 35562
rect 4352 35506 4420 35562
rect 4476 35506 4544 35562
rect 4600 35506 4668 35562
rect 4724 35506 4734 35562
rect 2798 35438 4734 35506
rect 2798 35382 2808 35438
rect 2864 35382 2932 35438
rect 2988 35382 3056 35438
rect 3112 35382 3180 35438
rect 3236 35382 3304 35438
rect 3360 35382 3428 35438
rect 3484 35382 3552 35438
rect 3608 35382 3676 35438
rect 3732 35382 3800 35438
rect 3856 35382 3924 35438
rect 3980 35382 4048 35438
rect 4104 35382 4172 35438
rect 4228 35382 4296 35438
rect 4352 35382 4420 35438
rect 4476 35382 4544 35438
rect 4600 35382 4668 35438
rect 4724 35382 4734 35438
rect 2798 35314 4734 35382
rect 2798 35258 2808 35314
rect 2864 35258 2932 35314
rect 2988 35258 3056 35314
rect 3112 35258 3180 35314
rect 3236 35258 3304 35314
rect 3360 35258 3428 35314
rect 3484 35258 3552 35314
rect 3608 35258 3676 35314
rect 3732 35258 3800 35314
rect 3856 35258 3924 35314
rect 3980 35258 4048 35314
rect 4104 35258 4172 35314
rect 4228 35258 4296 35314
rect 4352 35258 4420 35314
rect 4476 35258 4544 35314
rect 4600 35258 4668 35314
rect 4724 35258 4734 35314
rect 2798 35190 4734 35258
rect 2798 35134 2808 35190
rect 2864 35134 2932 35190
rect 2988 35134 3056 35190
rect 3112 35134 3180 35190
rect 3236 35134 3304 35190
rect 3360 35134 3428 35190
rect 3484 35134 3552 35190
rect 3608 35134 3676 35190
rect 3732 35134 3800 35190
rect 3856 35134 3924 35190
rect 3980 35134 4048 35190
rect 4104 35134 4172 35190
rect 4228 35134 4296 35190
rect 4352 35134 4420 35190
rect 4476 35134 4544 35190
rect 4600 35134 4668 35190
rect 4724 35134 4734 35190
rect 2798 35066 4734 35134
rect 2798 35010 2808 35066
rect 2864 35010 2932 35066
rect 2988 35010 3056 35066
rect 3112 35010 3180 35066
rect 3236 35010 3304 35066
rect 3360 35010 3428 35066
rect 3484 35010 3552 35066
rect 3608 35010 3676 35066
rect 3732 35010 3800 35066
rect 3856 35010 3924 35066
rect 3980 35010 4048 35066
rect 4104 35010 4172 35066
rect 4228 35010 4296 35066
rect 4352 35010 4420 35066
rect 4476 35010 4544 35066
rect 4600 35010 4668 35066
rect 4724 35010 4734 35066
rect 2798 34942 4734 35010
rect 2798 34886 2808 34942
rect 2864 34886 2932 34942
rect 2988 34886 3056 34942
rect 3112 34886 3180 34942
rect 3236 34886 3304 34942
rect 3360 34886 3428 34942
rect 3484 34886 3552 34942
rect 3608 34886 3676 34942
rect 3732 34886 3800 34942
rect 3856 34886 3924 34942
rect 3980 34886 4048 34942
rect 4104 34886 4172 34942
rect 4228 34886 4296 34942
rect 4352 34886 4420 34942
rect 4476 34886 4544 34942
rect 4600 34886 4668 34942
rect 4724 34886 4734 34942
rect 2798 34818 4734 34886
rect 2798 34762 2808 34818
rect 2864 34762 2932 34818
rect 2988 34762 3056 34818
rect 3112 34762 3180 34818
rect 3236 34762 3304 34818
rect 3360 34762 3428 34818
rect 3484 34762 3552 34818
rect 3608 34762 3676 34818
rect 3732 34762 3800 34818
rect 3856 34762 3924 34818
rect 3980 34762 4048 34818
rect 4104 34762 4172 34818
rect 4228 34762 4296 34818
rect 4352 34762 4420 34818
rect 4476 34762 4544 34818
rect 4600 34762 4668 34818
rect 4724 34762 4734 34818
rect 2798 34694 4734 34762
rect 2798 34638 2808 34694
rect 2864 34638 2932 34694
rect 2988 34638 3056 34694
rect 3112 34638 3180 34694
rect 3236 34638 3304 34694
rect 3360 34638 3428 34694
rect 3484 34638 3552 34694
rect 3608 34638 3676 34694
rect 3732 34638 3800 34694
rect 3856 34638 3924 34694
rect 3980 34638 4048 34694
rect 4104 34638 4172 34694
rect 4228 34638 4296 34694
rect 4352 34638 4420 34694
rect 4476 34638 4544 34694
rect 4600 34638 4668 34694
rect 4724 34638 4734 34694
rect 2798 34570 4734 34638
rect 2798 34514 2808 34570
rect 2864 34514 2932 34570
rect 2988 34514 3056 34570
rect 3112 34514 3180 34570
rect 3236 34514 3304 34570
rect 3360 34514 3428 34570
rect 3484 34514 3552 34570
rect 3608 34514 3676 34570
rect 3732 34514 3800 34570
rect 3856 34514 3924 34570
rect 3980 34514 4048 34570
rect 4104 34514 4172 34570
rect 4228 34514 4296 34570
rect 4352 34514 4420 34570
rect 4476 34514 4544 34570
rect 4600 34514 4668 34570
rect 4724 34514 4734 34570
rect 2798 34446 4734 34514
rect 2798 34390 2808 34446
rect 2864 34390 2932 34446
rect 2988 34390 3056 34446
rect 3112 34390 3180 34446
rect 3236 34390 3304 34446
rect 3360 34390 3428 34446
rect 3484 34390 3552 34446
rect 3608 34390 3676 34446
rect 3732 34390 3800 34446
rect 3856 34390 3924 34446
rect 3980 34390 4048 34446
rect 4104 34390 4172 34446
rect 4228 34390 4296 34446
rect 4352 34390 4420 34446
rect 4476 34390 4544 34446
rect 4600 34390 4668 34446
rect 4724 34390 4734 34446
rect 2798 34322 4734 34390
rect 2798 34266 2808 34322
rect 2864 34266 2932 34322
rect 2988 34266 3056 34322
rect 3112 34266 3180 34322
rect 3236 34266 3304 34322
rect 3360 34266 3428 34322
rect 3484 34266 3552 34322
rect 3608 34266 3676 34322
rect 3732 34266 3800 34322
rect 3856 34266 3924 34322
rect 3980 34266 4048 34322
rect 4104 34266 4172 34322
rect 4228 34266 4296 34322
rect 4352 34266 4420 34322
rect 4476 34266 4544 34322
rect 4600 34266 4668 34322
rect 4724 34266 4734 34322
rect 2798 34198 4734 34266
rect 2798 34142 2808 34198
rect 2864 34142 2932 34198
rect 2988 34142 3056 34198
rect 3112 34142 3180 34198
rect 3236 34142 3304 34198
rect 3360 34142 3428 34198
rect 3484 34142 3552 34198
rect 3608 34142 3676 34198
rect 3732 34142 3800 34198
rect 3856 34142 3924 34198
rect 3980 34142 4048 34198
rect 4104 34142 4172 34198
rect 4228 34142 4296 34198
rect 4352 34142 4420 34198
rect 4476 34142 4544 34198
rect 4600 34142 4668 34198
rect 4724 34142 4734 34198
rect 2798 34074 4734 34142
rect 2798 34018 2808 34074
rect 2864 34018 2932 34074
rect 2988 34018 3056 34074
rect 3112 34018 3180 34074
rect 3236 34018 3304 34074
rect 3360 34018 3428 34074
rect 3484 34018 3552 34074
rect 3608 34018 3676 34074
rect 3732 34018 3800 34074
rect 3856 34018 3924 34074
rect 3980 34018 4048 34074
rect 4104 34018 4172 34074
rect 4228 34018 4296 34074
rect 4352 34018 4420 34074
rect 4476 34018 4544 34074
rect 4600 34018 4668 34074
rect 4724 34018 4734 34074
rect 2798 33950 4734 34018
rect 2798 33894 2808 33950
rect 2864 33894 2932 33950
rect 2988 33894 3056 33950
rect 3112 33894 3180 33950
rect 3236 33894 3304 33950
rect 3360 33894 3428 33950
rect 3484 33894 3552 33950
rect 3608 33894 3676 33950
rect 3732 33894 3800 33950
rect 3856 33894 3924 33950
rect 3980 33894 4048 33950
rect 4104 33894 4172 33950
rect 4228 33894 4296 33950
rect 4352 33894 4420 33950
rect 4476 33894 4544 33950
rect 4600 33894 4668 33950
rect 4724 33894 4734 33950
rect 2798 33826 4734 33894
rect 2798 33770 2808 33826
rect 2864 33770 2932 33826
rect 2988 33770 3056 33826
rect 3112 33770 3180 33826
rect 3236 33770 3304 33826
rect 3360 33770 3428 33826
rect 3484 33770 3552 33826
rect 3608 33770 3676 33826
rect 3732 33770 3800 33826
rect 3856 33770 3924 33826
rect 3980 33770 4048 33826
rect 4104 33770 4172 33826
rect 4228 33770 4296 33826
rect 4352 33770 4420 33826
rect 4476 33770 4544 33826
rect 4600 33770 4668 33826
rect 4724 33770 4734 33826
rect 2798 33702 4734 33770
rect 2798 33646 2808 33702
rect 2864 33646 2932 33702
rect 2988 33646 3056 33702
rect 3112 33646 3180 33702
rect 3236 33646 3304 33702
rect 3360 33646 3428 33702
rect 3484 33646 3552 33702
rect 3608 33646 3676 33702
rect 3732 33646 3800 33702
rect 3856 33646 3924 33702
rect 3980 33646 4048 33702
rect 4104 33646 4172 33702
rect 4228 33646 4296 33702
rect 4352 33646 4420 33702
rect 4476 33646 4544 33702
rect 4600 33646 4668 33702
rect 4724 33646 4734 33702
rect 2798 33636 4734 33646
rect 5168 36554 7104 36564
rect 5168 36498 5178 36554
rect 5234 36498 5302 36554
rect 5358 36498 5426 36554
rect 5482 36498 5550 36554
rect 5606 36498 5674 36554
rect 5730 36498 5798 36554
rect 5854 36498 5922 36554
rect 5978 36498 6046 36554
rect 6102 36498 6170 36554
rect 6226 36498 6294 36554
rect 6350 36498 6418 36554
rect 6474 36498 6542 36554
rect 6598 36498 6666 36554
rect 6722 36498 6790 36554
rect 6846 36498 6914 36554
rect 6970 36498 7038 36554
rect 7094 36498 7104 36554
rect 5168 36430 7104 36498
rect 5168 36374 5178 36430
rect 5234 36374 5302 36430
rect 5358 36374 5426 36430
rect 5482 36374 5550 36430
rect 5606 36374 5674 36430
rect 5730 36374 5798 36430
rect 5854 36374 5922 36430
rect 5978 36374 6046 36430
rect 6102 36374 6170 36430
rect 6226 36374 6294 36430
rect 6350 36374 6418 36430
rect 6474 36374 6542 36430
rect 6598 36374 6666 36430
rect 6722 36374 6790 36430
rect 6846 36374 6914 36430
rect 6970 36374 7038 36430
rect 7094 36374 7104 36430
rect 5168 36306 7104 36374
rect 5168 36250 5178 36306
rect 5234 36250 5302 36306
rect 5358 36250 5426 36306
rect 5482 36250 5550 36306
rect 5606 36250 5674 36306
rect 5730 36250 5798 36306
rect 5854 36250 5922 36306
rect 5978 36250 6046 36306
rect 6102 36250 6170 36306
rect 6226 36250 6294 36306
rect 6350 36250 6418 36306
rect 6474 36250 6542 36306
rect 6598 36250 6666 36306
rect 6722 36250 6790 36306
rect 6846 36250 6914 36306
rect 6970 36250 7038 36306
rect 7094 36250 7104 36306
rect 5168 36182 7104 36250
rect 5168 36126 5178 36182
rect 5234 36126 5302 36182
rect 5358 36126 5426 36182
rect 5482 36126 5550 36182
rect 5606 36126 5674 36182
rect 5730 36126 5798 36182
rect 5854 36126 5922 36182
rect 5978 36126 6046 36182
rect 6102 36126 6170 36182
rect 6226 36126 6294 36182
rect 6350 36126 6418 36182
rect 6474 36126 6542 36182
rect 6598 36126 6666 36182
rect 6722 36126 6790 36182
rect 6846 36126 6914 36182
rect 6970 36126 7038 36182
rect 7094 36126 7104 36182
rect 5168 36058 7104 36126
rect 5168 36002 5178 36058
rect 5234 36002 5302 36058
rect 5358 36002 5426 36058
rect 5482 36002 5550 36058
rect 5606 36002 5674 36058
rect 5730 36002 5798 36058
rect 5854 36002 5922 36058
rect 5978 36002 6046 36058
rect 6102 36002 6170 36058
rect 6226 36002 6294 36058
rect 6350 36002 6418 36058
rect 6474 36002 6542 36058
rect 6598 36002 6666 36058
rect 6722 36002 6790 36058
rect 6846 36002 6914 36058
rect 6970 36002 7038 36058
rect 7094 36002 7104 36058
rect 5168 35934 7104 36002
rect 5168 35878 5178 35934
rect 5234 35878 5302 35934
rect 5358 35878 5426 35934
rect 5482 35878 5550 35934
rect 5606 35878 5674 35934
rect 5730 35878 5798 35934
rect 5854 35878 5922 35934
rect 5978 35878 6046 35934
rect 6102 35878 6170 35934
rect 6226 35878 6294 35934
rect 6350 35878 6418 35934
rect 6474 35878 6542 35934
rect 6598 35878 6666 35934
rect 6722 35878 6790 35934
rect 6846 35878 6914 35934
rect 6970 35878 7038 35934
rect 7094 35878 7104 35934
rect 5168 35810 7104 35878
rect 5168 35754 5178 35810
rect 5234 35754 5302 35810
rect 5358 35754 5426 35810
rect 5482 35754 5550 35810
rect 5606 35754 5674 35810
rect 5730 35754 5798 35810
rect 5854 35754 5922 35810
rect 5978 35754 6046 35810
rect 6102 35754 6170 35810
rect 6226 35754 6294 35810
rect 6350 35754 6418 35810
rect 6474 35754 6542 35810
rect 6598 35754 6666 35810
rect 6722 35754 6790 35810
rect 6846 35754 6914 35810
rect 6970 35754 7038 35810
rect 7094 35754 7104 35810
rect 5168 35686 7104 35754
rect 5168 35630 5178 35686
rect 5234 35630 5302 35686
rect 5358 35630 5426 35686
rect 5482 35630 5550 35686
rect 5606 35630 5674 35686
rect 5730 35630 5798 35686
rect 5854 35630 5922 35686
rect 5978 35630 6046 35686
rect 6102 35630 6170 35686
rect 6226 35630 6294 35686
rect 6350 35630 6418 35686
rect 6474 35630 6542 35686
rect 6598 35630 6666 35686
rect 6722 35630 6790 35686
rect 6846 35630 6914 35686
rect 6970 35630 7038 35686
rect 7094 35630 7104 35686
rect 5168 35562 7104 35630
rect 5168 35506 5178 35562
rect 5234 35506 5302 35562
rect 5358 35506 5426 35562
rect 5482 35506 5550 35562
rect 5606 35506 5674 35562
rect 5730 35506 5798 35562
rect 5854 35506 5922 35562
rect 5978 35506 6046 35562
rect 6102 35506 6170 35562
rect 6226 35506 6294 35562
rect 6350 35506 6418 35562
rect 6474 35506 6542 35562
rect 6598 35506 6666 35562
rect 6722 35506 6790 35562
rect 6846 35506 6914 35562
rect 6970 35506 7038 35562
rect 7094 35506 7104 35562
rect 5168 35438 7104 35506
rect 5168 35382 5178 35438
rect 5234 35382 5302 35438
rect 5358 35382 5426 35438
rect 5482 35382 5550 35438
rect 5606 35382 5674 35438
rect 5730 35382 5798 35438
rect 5854 35382 5922 35438
rect 5978 35382 6046 35438
rect 6102 35382 6170 35438
rect 6226 35382 6294 35438
rect 6350 35382 6418 35438
rect 6474 35382 6542 35438
rect 6598 35382 6666 35438
rect 6722 35382 6790 35438
rect 6846 35382 6914 35438
rect 6970 35382 7038 35438
rect 7094 35382 7104 35438
rect 5168 35314 7104 35382
rect 5168 35258 5178 35314
rect 5234 35258 5302 35314
rect 5358 35258 5426 35314
rect 5482 35258 5550 35314
rect 5606 35258 5674 35314
rect 5730 35258 5798 35314
rect 5854 35258 5922 35314
rect 5978 35258 6046 35314
rect 6102 35258 6170 35314
rect 6226 35258 6294 35314
rect 6350 35258 6418 35314
rect 6474 35258 6542 35314
rect 6598 35258 6666 35314
rect 6722 35258 6790 35314
rect 6846 35258 6914 35314
rect 6970 35258 7038 35314
rect 7094 35258 7104 35314
rect 5168 35190 7104 35258
rect 5168 35134 5178 35190
rect 5234 35134 5302 35190
rect 5358 35134 5426 35190
rect 5482 35134 5550 35190
rect 5606 35134 5674 35190
rect 5730 35134 5798 35190
rect 5854 35134 5922 35190
rect 5978 35134 6046 35190
rect 6102 35134 6170 35190
rect 6226 35134 6294 35190
rect 6350 35134 6418 35190
rect 6474 35134 6542 35190
rect 6598 35134 6666 35190
rect 6722 35134 6790 35190
rect 6846 35134 6914 35190
rect 6970 35134 7038 35190
rect 7094 35134 7104 35190
rect 5168 35066 7104 35134
rect 5168 35010 5178 35066
rect 5234 35010 5302 35066
rect 5358 35010 5426 35066
rect 5482 35010 5550 35066
rect 5606 35010 5674 35066
rect 5730 35010 5798 35066
rect 5854 35010 5922 35066
rect 5978 35010 6046 35066
rect 6102 35010 6170 35066
rect 6226 35010 6294 35066
rect 6350 35010 6418 35066
rect 6474 35010 6542 35066
rect 6598 35010 6666 35066
rect 6722 35010 6790 35066
rect 6846 35010 6914 35066
rect 6970 35010 7038 35066
rect 7094 35010 7104 35066
rect 5168 34942 7104 35010
rect 5168 34886 5178 34942
rect 5234 34886 5302 34942
rect 5358 34886 5426 34942
rect 5482 34886 5550 34942
rect 5606 34886 5674 34942
rect 5730 34886 5798 34942
rect 5854 34886 5922 34942
rect 5978 34886 6046 34942
rect 6102 34886 6170 34942
rect 6226 34886 6294 34942
rect 6350 34886 6418 34942
rect 6474 34886 6542 34942
rect 6598 34886 6666 34942
rect 6722 34886 6790 34942
rect 6846 34886 6914 34942
rect 6970 34886 7038 34942
rect 7094 34886 7104 34942
rect 5168 34818 7104 34886
rect 5168 34762 5178 34818
rect 5234 34762 5302 34818
rect 5358 34762 5426 34818
rect 5482 34762 5550 34818
rect 5606 34762 5674 34818
rect 5730 34762 5798 34818
rect 5854 34762 5922 34818
rect 5978 34762 6046 34818
rect 6102 34762 6170 34818
rect 6226 34762 6294 34818
rect 6350 34762 6418 34818
rect 6474 34762 6542 34818
rect 6598 34762 6666 34818
rect 6722 34762 6790 34818
rect 6846 34762 6914 34818
rect 6970 34762 7038 34818
rect 7094 34762 7104 34818
rect 5168 34694 7104 34762
rect 5168 34638 5178 34694
rect 5234 34638 5302 34694
rect 5358 34638 5426 34694
rect 5482 34638 5550 34694
rect 5606 34638 5674 34694
rect 5730 34638 5798 34694
rect 5854 34638 5922 34694
rect 5978 34638 6046 34694
rect 6102 34638 6170 34694
rect 6226 34638 6294 34694
rect 6350 34638 6418 34694
rect 6474 34638 6542 34694
rect 6598 34638 6666 34694
rect 6722 34638 6790 34694
rect 6846 34638 6914 34694
rect 6970 34638 7038 34694
rect 7094 34638 7104 34694
rect 5168 34570 7104 34638
rect 5168 34514 5178 34570
rect 5234 34514 5302 34570
rect 5358 34514 5426 34570
rect 5482 34514 5550 34570
rect 5606 34514 5674 34570
rect 5730 34514 5798 34570
rect 5854 34514 5922 34570
rect 5978 34514 6046 34570
rect 6102 34514 6170 34570
rect 6226 34514 6294 34570
rect 6350 34514 6418 34570
rect 6474 34514 6542 34570
rect 6598 34514 6666 34570
rect 6722 34514 6790 34570
rect 6846 34514 6914 34570
rect 6970 34514 7038 34570
rect 7094 34514 7104 34570
rect 5168 34446 7104 34514
rect 5168 34390 5178 34446
rect 5234 34390 5302 34446
rect 5358 34390 5426 34446
rect 5482 34390 5550 34446
rect 5606 34390 5674 34446
rect 5730 34390 5798 34446
rect 5854 34390 5922 34446
rect 5978 34390 6046 34446
rect 6102 34390 6170 34446
rect 6226 34390 6294 34446
rect 6350 34390 6418 34446
rect 6474 34390 6542 34446
rect 6598 34390 6666 34446
rect 6722 34390 6790 34446
rect 6846 34390 6914 34446
rect 6970 34390 7038 34446
rect 7094 34390 7104 34446
rect 5168 34322 7104 34390
rect 5168 34266 5178 34322
rect 5234 34266 5302 34322
rect 5358 34266 5426 34322
rect 5482 34266 5550 34322
rect 5606 34266 5674 34322
rect 5730 34266 5798 34322
rect 5854 34266 5922 34322
rect 5978 34266 6046 34322
rect 6102 34266 6170 34322
rect 6226 34266 6294 34322
rect 6350 34266 6418 34322
rect 6474 34266 6542 34322
rect 6598 34266 6666 34322
rect 6722 34266 6790 34322
rect 6846 34266 6914 34322
rect 6970 34266 7038 34322
rect 7094 34266 7104 34322
rect 5168 34198 7104 34266
rect 5168 34142 5178 34198
rect 5234 34142 5302 34198
rect 5358 34142 5426 34198
rect 5482 34142 5550 34198
rect 5606 34142 5674 34198
rect 5730 34142 5798 34198
rect 5854 34142 5922 34198
rect 5978 34142 6046 34198
rect 6102 34142 6170 34198
rect 6226 34142 6294 34198
rect 6350 34142 6418 34198
rect 6474 34142 6542 34198
rect 6598 34142 6666 34198
rect 6722 34142 6790 34198
rect 6846 34142 6914 34198
rect 6970 34142 7038 34198
rect 7094 34142 7104 34198
rect 5168 34074 7104 34142
rect 5168 34018 5178 34074
rect 5234 34018 5302 34074
rect 5358 34018 5426 34074
rect 5482 34018 5550 34074
rect 5606 34018 5674 34074
rect 5730 34018 5798 34074
rect 5854 34018 5922 34074
rect 5978 34018 6046 34074
rect 6102 34018 6170 34074
rect 6226 34018 6294 34074
rect 6350 34018 6418 34074
rect 6474 34018 6542 34074
rect 6598 34018 6666 34074
rect 6722 34018 6790 34074
rect 6846 34018 6914 34074
rect 6970 34018 7038 34074
rect 7094 34018 7104 34074
rect 5168 33950 7104 34018
rect 5168 33894 5178 33950
rect 5234 33894 5302 33950
rect 5358 33894 5426 33950
rect 5482 33894 5550 33950
rect 5606 33894 5674 33950
rect 5730 33894 5798 33950
rect 5854 33894 5922 33950
rect 5978 33894 6046 33950
rect 6102 33894 6170 33950
rect 6226 33894 6294 33950
rect 6350 33894 6418 33950
rect 6474 33894 6542 33950
rect 6598 33894 6666 33950
rect 6722 33894 6790 33950
rect 6846 33894 6914 33950
rect 6970 33894 7038 33950
rect 7094 33894 7104 33950
rect 5168 33826 7104 33894
rect 5168 33770 5178 33826
rect 5234 33770 5302 33826
rect 5358 33770 5426 33826
rect 5482 33770 5550 33826
rect 5606 33770 5674 33826
rect 5730 33770 5798 33826
rect 5854 33770 5922 33826
rect 5978 33770 6046 33826
rect 6102 33770 6170 33826
rect 6226 33770 6294 33826
rect 6350 33770 6418 33826
rect 6474 33770 6542 33826
rect 6598 33770 6666 33826
rect 6722 33770 6790 33826
rect 6846 33770 6914 33826
rect 6970 33770 7038 33826
rect 7094 33770 7104 33826
rect 5168 33702 7104 33770
rect 5168 33646 5178 33702
rect 5234 33646 5302 33702
rect 5358 33646 5426 33702
rect 5482 33646 5550 33702
rect 5606 33646 5674 33702
rect 5730 33646 5798 33702
rect 5854 33646 5922 33702
rect 5978 33646 6046 33702
rect 6102 33646 6170 33702
rect 6226 33646 6294 33702
rect 6350 33646 6418 33702
rect 6474 33646 6542 33702
rect 6598 33646 6666 33702
rect 6722 33646 6790 33702
rect 6846 33646 6914 33702
rect 6970 33646 7038 33702
rect 7094 33646 7104 33702
rect 5168 33636 7104 33646
rect 7874 36554 9810 36564
rect 7874 36498 7884 36554
rect 7940 36498 8008 36554
rect 8064 36498 8132 36554
rect 8188 36498 8256 36554
rect 8312 36498 8380 36554
rect 8436 36498 8504 36554
rect 8560 36498 8628 36554
rect 8684 36498 8752 36554
rect 8808 36498 8876 36554
rect 8932 36498 9000 36554
rect 9056 36498 9124 36554
rect 9180 36498 9248 36554
rect 9304 36498 9372 36554
rect 9428 36498 9496 36554
rect 9552 36498 9620 36554
rect 9676 36498 9744 36554
rect 9800 36498 9810 36554
rect 7874 36430 9810 36498
rect 7874 36374 7884 36430
rect 7940 36374 8008 36430
rect 8064 36374 8132 36430
rect 8188 36374 8256 36430
rect 8312 36374 8380 36430
rect 8436 36374 8504 36430
rect 8560 36374 8628 36430
rect 8684 36374 8752 36430
rect 8808 36374 8876 36430
rect 8932 36374 9000 36430
rect 9056 36374 9124 36430
rect 9180 36374 9248 36430
rect 9304 36374 9372 36430
rect 9428 36374 9496 36430
rect 9552 36374 9620 36430
rect 9676 36374 9744 36430
rect 9800 36374 9810 36430
rect 7874 36306 9810 36374
rect 7874 36250 7884 36306
rect 7940 36250 8008 36306
rect 8064 36250 8132 36306
rect 8188 36250 8256 36306
rect 8312 36250 8380 36306
rect 8436 36250 8504 36306
rect 8560 36250 8628 36306
rect 8684 36250 8752 36306
rect 8808 36250 8876 36306
rect 8932 36250 9000 36306
rect 9056 36250 9124 36306
rect 9180 36250 9248 36306
rect 9304 36250 9372 36306
rect 9428 36250 9496 36306
rect 9552 36250 9620 36306
rect 9676 36250 9744 36306
rect 9800 36250 9810 36306
rect 7874 36182 9810 36250
rect 7874 36126 7884 36182
rect 7940 36126 8008 36182
rect 8064 36126 8132 36182
rect 8188 36126 8256 36182
rect 8312 36126 8380 36182
rect 8436 36126 8504 36182
rect 8560 36126 8628 36182
rect 8684 36126 8752 36182
rect 8808 36126 8876 36182
rect 8932 36126 9000 36182
rect 9056 36126 9124 36182
rect 9180 36126 9248 36182
rect 9304 36126 9372 36182
rect 9428 36126 9496 36182
rect 9552 36126 9620 36182
rect 9676 36126 9744 36182
rect 9800 36126 9810 36182
rect 7874 36058 9810 36126
rect 7874 36002 7884 36058
rect 7940 36002 8008 36058
rect 8064 36002 8132 36058
rect 8188 36002 8256 36058
rect 8312 36002 8380 36058
rect 8436 36002 8504 36058
rect 8560 36002 8628 36058
rect 8684 36002 8752 36058
rect 8808 36002 8876 36058
rect 8932 36002 9000 36058
rect 9056 36002 9124 36058
rect 9180 36002 9248 36058
rect 9304 36002 9372 36058
rect 9428 36002 9496 36058
rect 9552 36002 9620 36058
rect 9676 36002 9744 36058
rect 9800 36002 9810 36058
rect 7874 35934 9810 36002
rect 7874 35878 7884 35934
rect 7940 35878 8008 35934
rect 8064 35878 8132 35934
rect 8188 35878 8256 35934
rect 8312 35878 8380 35934
rect 8436 35878 8504 35934
rect 8560 35878 8628 35934
rect 8684 35878 8752 35934
rect 8808 35878 8876 35934
rect 8932 35878 9000 35934
rect 9056 35878 9124 35934
rect 9180 35878 9248 35934
rect 9304 35878 9372 35934
rect 9428 35878 9496 35934
rect 9552 35878 9620 35934
rect 9676 35878 9744 35934
rect 9800 35878 9810 35934
rect 7874 35810 9810 35878
rect 7874 35754 7884 35810
rect 7940 35754 8008 35810
rect 8064 35754 8132 35810
rect 8188 35754 8256 35810
rect 8312 35754 8380 35810
rect 8436 35754 8504 35810
rect 8560 35754 8628 35810
rect 8684 35754 8752 35810
rect 8808 35754 8876 35810
rect 8932 35754 9000 35810
rect 9056 35754 9124 35810
rect 9180 35754 9248 35810
rect 9304 35754 9372 35810
rect 9428 35754 9496 35810
rect 9552 35754 9620 35810
rect 9676 35754 9744 35810
rect 9800 35754 9810 35810
rect 7874 35686 9810 35754
rect 7874 35630 7884 35686
rect 7940 35630 8008 35686
rect 8064 35630 8132 35686
rect 8188 35630 8256 35686
rect 8312 35630 8380 35686
rect 8436 35630 8504 35686
rect 8560 35630 8628 35686
rect 8684 35630 8752 35686
rect 8808 35630 8876 35686
rect 8932 35630 9000 35686
rect 9056 35630 9124 35686
rect 9180 35630 9248 35686
rect 9304 35630 9372 35686
rect 9428 35630 9496 35686
rect 9552 35630 9620 35686
rect 9676 35630 9744 35686
rect 9800 35630 9810 35686
rect 7874 35562 9810 35630
rect 7874 35506 7884 35562
rect 7940 35506 8008 35562
rect 8064 35506 8132 35562
rect 8188 35506 8256 35562
rect 8312 35506 8380 35562
rect 8436 35506 8504 35562
rect 8560 35506 8628 35562
rect 8684 35506 8752 35562
rect 8808 35506 8876 35562
rect 8932 35506 9000 35562
rect 9056 35506 9124 35562
rect 9180 35506 9248 35562
rect 9304 35506 9372 35562
rect 9428 35506 9496 35562
rect 9552 35506 9620 35562
rect 9676 35506 9744 35562
rect 9800 35506 9810 35562
rect 7874 35438 9810 35506
rect 7874 35382 7884 35438
rect 7940 35382 8008 35438
rect 8064 35382 8132 35438
rect 8188 35382 8256 35438
rect 8312 35382 8380 35438
rect 8436 35382 8504 35438
rect 8560 35382 8628 35438
rect 8684 35382 8752 35438
rect 8808 35382 8876 35438
rect 8932 35382 9000 35438
rect 9056 35382 9124 35438
rect 9180 35382 9248 35438
rect 9304 35382 9372 35438
rect 9428 35382 9496 35438
rect 9552 35382 9620 35438
rect 9676 35382 9744 35438
rect 9800 35382 9810 35438
rect 7874 35314 9810 35382
rect 7874 35258 7884 35314
rect 7940 35258 8008 35314
rect 8064 35258 8132 35314
rect 8188 35258 8256 35314
rect 8312 35258 8380 35314
rect 8436 35258 8504 35314
rect 8560 35258 8628 35314
rect 8684 35258 8752 35314
rect 8808 35258 8876 35314
rect 8932 35258 9000 35314
rect 9056 35258 9124 35314
rect 9180 35258 9248 35314
rect 9304 35258 9372 35314
rect 9428 35258 9496 35314
rect 9552 35258 9620 35314
rect 9676 35258 9744 35314
rect 9800 35258 9810 35314
rect 7874 35190 9810 35258
rect 7874 35134 7884 35190
rect 7940 35134 8008 35190
rect 8064 35134 8132 35190
rect 8188 35134 8256 35190
rect 8312 35134 8380 35190
rect 8436 35134 8504 35190
rect 8560 35134 8628 35190
rect 8684 35134 8752 35190
rect 8808 35134 8876 35190
rect 8932 35134 9000 35190
rect 9056 35134 9124 35190
rect 9180 35134 9248 35190
rect 9304 35134 9372 35190
rect 9428 35134 9496 35190
rect 9552 35134 9620 35190
rect 9676 35134 9744 35190
rect 9800 35134 9810 35190
rect 7874 35066 9810 35134
rect 7874 35010 7884 35066
rect 7940 35010 8008 35066
rect 8064 35010 8132 35066
rect 8188 35010 8256 35066
rect 8312 35010 8380 35066
rect 8436 35010 8504 35066
rect 8560 35010 8628 35066
rect 8684 35010 8752 35066
rect 8808 35010 8876 35066
rect 8932 35010 9000 35066
rect 9056 35010 9124 35066
rect 9180 35010 9248 35066
rect 9304 35010 9372 35066
rect 9428 35010 9496 35066
rect 9552 35010 9620 35066
rect 9676 35010 9744 35066
rect 9800 35010 9810 35066
rect 7874 34942 9810 35010
rect 7874 34886 7884 34942
rect 7940 34886 8008 34942
rect 8064 34886 8132 34942
rect 8188 34886 8256 34942
rect 8312 34886 8380 34942
rect 8436 34886 8504 34942
rect 8560 34886 8628 34942
rect 8684 34886 8752 34942
rect 8808 34886 8876 34942
rect 8932 34886 9000 34942
rect 9056 34886 9124 34942
rect 9180 34886 9248 34942
rect 9304 34886 9372 34942
rect 9428 34886 9496 34942
rect 9552 34886 9620 34942
rect 9676 34886 9744 34942
rect 9800 34886 9810 34942
rect 7874 34818 9810 34886
rect 7874 34762 7884 34818
rect 7940 34762 8008 34818
rect 8064 34762 8132 34818
rect 8188 34762 8256 34818
rect 8312 34762 8380 34818
rect 8436 34762 8504 34818
rect 8560 34762 8628 34818
rect 8684 34762 8752 34818
rect 8808 34762 8876 34818
rect 8932 34762 9000 34818
rect 9056 34762 9124 34818
rect 9180 34762 9248 34818
rect 9304 34762 9372 34818
rect 9428 34762 9496 34818
rect 9552 34762 9620 34818
rect 9676 34762 9744 34818
rect 9800 34762 9810 34818
rect 7874 34694 9810 34762
rect 7874 34638 7884 34694
rect 7940 34638 8008 34694
rect 8064 34638 8132 34694
rect 8188 34638 8256 34694
rect 8312 34638 8380 34694
rect 8436 34638 8504 34694
rect 8560 34638 8628 34694
rect 8684 34638 8752 34694
rect 8808 34638 8876 34694
rect 8932 34638 9000 34694
rect 9056 34638 9124 34694
rect 9180 34638 9248 34694
rect 9304 34638 9372 34694
rect 9428 34638 9496 34694
rect 9552 34638 9620 34694
rect 9676 34638 9744 34694
rect 9800 34638 9810 34694
rect 7874 34570 9810 34638
rect 7874 34514 7884 34570
rect 7940 34514 8008 34570
rect 8064 34514 8132 34570
rect 8188 34514 8256 34570
rect 8312 34514 8380 34570
rect 8436 34514 8504 34570
rect 8560 34514 8628 34570
rect 8684 34514 8752 34570
rect 8808 34514 8876 34570
rect 8932 34514 9000 34570
rect 9056 34514 9124 34570
rect 9180 34514 9248 34570
rect 9304 34514 9372 34570
rect 9428 34514 9496 34570
rect 9552 34514 9620 34570
rect 9676 34514 9744 34570
rect 9800 34514 9810 34570
rect 7874 34446 9810 34514
rect 7874 34390 7884 34446
rect 7940 34390 8008 34446
rect 8064 34390 8132 34446
rect 8188 34390 8256 34446
rect 8312 34390 8380 34446
rect 8436 34390 8504 34446
rect 8560 34390 8628 34446
rect 8684 34390 8752 34446
rect 8808 34390 8876 34446
rect 8932 34390 9000 34446
rect 9056 34390 9124 34446
rect 9180 34390 9248 34446
rect 9304 34390 9372 34446
rect 9428 34390 9496 34446
rect 9552 34390 9620 34446
rect 9676 34390 9744 34446
rect 9800 34390 9810 34446
rect 7874 34322 9810 34390
rect 7874 34266 7884 34322
rect 7940 34266 8008 34322
rect 8064 34266 8132 34322
rect 8188 34266 8256 34322
rect 8312 34266 8380 34322
rect 8436 34266 8504 34322
rect 8560 34266 8628 34322
rect 8684 34266 8752 34322
rect 8808 34266 8876 34322
rect 8932 34266 9000 34322
rect 9056 34266 9124 34322
rect 9180 34266 9248 34322
rect 9304 34266 9372 34322
rect 9428 34266 9496 34322
rect 9552 34266 9620 34322
rect 9676 34266 9744 34322
rect 9800 34266 9810 34322
rect 7874 34198 9810 34266
rect 7874 34142 7884 34198
rect 7940 34142 8008 34198
rect 8064 34142 8132 34198
rect 8188 34142 8256 34198
rect 8312 34142 8380 34198
rect 8436 34142 8504 34198
rect 8560 34142 8628 34198
rect 8684 34142 8752 34198
rect 8808 34142 8876 34198
rect 8932 34142 9000 34198
rect 9056 34142 9124 34198
rect 9180 34142 9248 34198
rect 9304 34142 9372 34198
rect 9428 34142 9496 34198
rect 9552 34142 9620 34198
rect 9676 34142 9744 34198
rect 9800 34142 9810 34198
rect 7874 34074 9810 34142
rect 7874 34018 7884 34074
rect 7940 34018 8008 34074
rect 8064 34018 8132 34074
rect 8188 34018 8256 34074
rect 8312 34018 8380 34074
rect 8436 34018 8504 34074
rect 8560 34018 8628 34074
rect 8684 34018 8752 34074
rect 8808 34018 8876 34074
rect 8932 34018 9000 34074
rect 9056 34018 9124 34074
rect 9180 34018 9248 34074
rect 9304 34018 9372 34074
rect 9428 34018 9496 34074
rect 9552 34018 9620 34074
rect 9676 34018 9744 34074
rect 9800 34018 9810 34074
rect 7874 33950 9810 34018
rect 7874 33894 7884 33950
rect 7940 33894 8008 33950
rect 8064 33894 8132 33950
rect 8188 33894 8256 33950
rect 8312 33894 8380 33950
rect 8436 33894 8504 33950
rect 8560 33894 8628 33950
rect 8684 33894 8752 33950
rect 8808 33894 8876 33950
rect 8932 33894 9000 33950
rect 9056 33894 9124 33950
rect 9180 33894 9248 33950
rect 9304 33894 9372 33950
rect 9428 33894 9496 33950
rect 9552 33894 9620 33950
rect 9676 33894 9744 33950
rect 9800 33894 9810 33950
rect 7874 33826 9810 33894
rect 7874 33770 7884 33826
rect 7940 33770 8008 33826
rect 8064 33770 8132 33826
rect 8188 33770 8256 33826
rect 8312 33770 8380 33826
rect 8436 33770 8504 33826
rect 8560 33770 8628 33826
rect 8684 33770 8752 33826
rect 8808 33770 8876 33826
rect 8932 33770 9000 33826
rect 9056 33770 9124 33826
rect 9180 33770 9248 33826
rect 9304 33770 9372 33826
rect 9428 33770 9496 33826
rect 9552 33770 9620 33826
rect 9676 33770 9744 33826
rect 9800 33770 9810 33826
rect 7874 33702 9810 33770
rect 7874 33646 7884 33702
rect 7940 33646 8008 33702
rect 8064 33646 8132 33702
rect 8188 33646 8256 33702
rect 8312 33646 8380 33702
rect 8436 33646 8504 33702
rect 8560 33646 8628 33702
rect 8684 33646 8752 33702
rect 8808 33646 8876 33702
rect 8932 33646 9000 33702
rect 9056 33646 9124 33702
rect 9180 33646 9248 33702
rect 9304 33646 9372 33702
rect 9428 33646 9496 33702
rect 9552 33646 9620 33702
rect 9676 33646 9744 33702
rect 9800 33646 9810 33702
rect 7874 33636 9810 33646
rect 10244 36554 12180 36564
rect 10244 36498 10254 36554
rect 10310 36498 10378 36554
rect 10434 36498 10502 36554
rect 10558 36498 10626 36554
rect 10682 36498 10750 36554
rect 10806 36498 10874 36554
rect 10930 36498 10998 36554
rect 11054 36498 11122 36554
rect 11178 36498 11246 36554
rect 11302 36498 11370 36554
rect 11426 36498 11494 36554
rect 11550 36498 11618 36554
rect 11674 36498 11742 36554
rect 11798 36498 11866 36554
rect 11922 36498 11990 36554
rect 12046 36498 12114 36554
rect 12170 36498 12180 36554
rect 10244 36430 12180 36498
rect 10244 36374 10254 36430
rect 10310 36374 10378 36430
rect 10434 36374 10502 36430
rect 10558 36374 10626 36430
rect 10682 36374 10750 36430
rect 10806 36374 10874 36430
rect 10930 36374 10998 36430
rect 11054 36374 11122 36430
rect 11178 36374 11246 36430
rect 11302 36374 11370 36430
rect 11426 36374 11494 36430
rect 11550 36374 11618 36430
rect 11674 36374 11742 36430
rect 11798 36374 11866 36430
rect 11922 36374 11990 36430
rect 12046 36374 12114 36430
rect 12170 36374 12180 36430
rect 10244 36306 12180 36374
rect 10244 36250 10254 36306
rect 10310 36250 10378 36306
rect 10434 36250 10502 36306
rect 10558 36250 10626 36306
rect 10682 36250 10750 36306
rect 10806 36250 10874 36306
rect 10930 36250 10998 36306
rect 11054 36250 11122 36306
rect 11178 36250 11246 36306
rect 11302 36250 11370 36306
rect 11426 36250 11494 36306
rect 11550 36250 11618 36306
rect 11674 36250 11742 36306
rect 11798 36250 11866 36306
rect 11922 36250 11990 36306
rect 12046 36250 12114 36306
rect 12170 36250 12180 36306
rect 10244 36182 12180 36250
rect 10244 36126 10254 36182
rect 10310 36126 10378 36182
rect 10434 36126 10502 36182
rect 10558 36126 10626 36182
rect 10682 36126 10750 36182
rect 10806 36126 10874 36182
rect 10930 36126 10998 36182
rect 11054 36126 11122 36182
rect 11178 36126 11246 36182
rect 11302 36126 11370 36182
rect 11426 36126 11494 36182
rect 11550 36126 11618 36182
rect 11674 36126 11742 36182
rect 11798 36126 11866 36182
rect 11922 36126 11990 36182
rect 12046 36126 12114 36182
rect 12170 36126 12180 36182
rect 10244 36058 12180 36126
rect 10244 36002 10254 36058
rect 10310 36002 10378 36058
rect 10434 36002 10502 36058
rect 10558 36002 10626 36058
rect 10682 36002 10750 36058
rect 10806 36002 10874 36058
rect 10930 36002 10998 36058
rect 11054 36002 11122 36058
rect 11178 36002 11246 36058
rect 11302 36002 11370 36058
rect 11426 36002 11494 36058
rect 11550 36002 11618 36058
rect 11674 36002 11742 36058
rect 11798 36002 11866 36058
rect 11922 36002 11990 36058
rect 12046 36002 12114 36058
rect 12170 36002 12180 36058
rect 10244 35934 12180 36002
rect 10244 35878 10254 35934
rect 10310 35878 10378 35934
rect 10434 35878 10502 35934
rect 10558 35878 10626 35934
rect 10682 35878 10750 35934
rect 10806 35878 10874 35934
rect 10930 35878 10998 35934
rect 11054 35878 11122 35934
rect 11178 35878 11246 35934
rect 11302 35878 11370 35934
rect 11426 35878 11494 35934
rect 11550 35878 11618 35934
rect 11674 35878 11742 35934
rect 11798 35878 11866 35934
rect 11922 35878 11990 35934
rect 12046 35878 12114 35934
rect 12170 35878 12180 35934
rect 10244 35810 12180 35878
rect 10244 35754 10254 35810
rect 10310 35754 10378 35810
rect 10434 35754 10502 35810
rect 10558 35754 10626 35810
rect 10682 35754 10750 35810
rect 10806 35754 10874 35810
rect 10930 35754 10998 35810
rect 11054 35754 11122 35810
rect 11178 35754 11246 35810
rect 11302 35754 11370 35810
rect 11426 35754 11494 35810
rect 11550 35754 11618 35810
rect 11674 35754 11742 35810
rect 11798 35754 11866 35810
rect 11922 35754 11990 35810
rect 12046 35754 12114 35810
rect 12170 35754 12180 35810
rect 10244 35686 12180 35754
rect 10244 35630 10254 35686
rect 10310 35630 10378 35686
rect 10434 35630 10502 35686
rect 10558 35630 10626 35686
rect 10682 35630 10750 35686
rect 10806 35630 10874 35686
rect 10930 35630 10998 35686
rect 11054 35630 11122 35686
rect 11178 35630 11246 35686
rect 11302 35630 11370 35686
rect 11426 35630 11494 35686
rect 11550 35630 11618 35686
rect 11674 35630 11742 35686
rect 11798 35630 11866 35686
rect 11922 35630 11990 35686
rect 12046 35630 12114 35686
rect 12170 35630 12180 35686
rect 10244 35562 12180 35630
rect 10244 35506 10254 35562
rect 10310 35506 10378 35562
rect 10434 35506 10502 35562
rect 10558 35506 10626 35562
rect 10682 35506 10750 35562
rect 10806 35506 10874 35562
rect 10930 35506 10998 35562
rect 11054 35506 11122 35562
rect 11178 35506 11246 35562
rect 11302 35506 11370 35562
rect 11426 35506 11494 35562
rect 11550 35506 11618 35562
rect 11674 35506 11742 35562
rect 11798 35506 11866 35562
rect 11922 35506 11990 35562
rect 12046 35506 12114 35562
rect 12170 35506 12180 35562
rect 10244 35438 12180 35506
rect 10244 35382 10254 35438
rect 10310 35382 10378 35438
rect 10434 35382 10502 35438
rect 10558 35382 10626 35438
rect 10682 35382 10750 35438
rect 10806 35382 10874 35438
rect 10930 35382 10998 35438
rect 11054 35382 11122 35438
rect 11178 35382 11246 35438
rect 11302 35382 11370 35438
rect 11426 35382 11494 35438
rect 11550 35382 11618 35438
rect 11674 35382 11742 35438
rect 11798 35382 11866 35438
rect 11922 35382 11990 35438
rect 12046 35382 12114 35438
rect 12170 35382 12180 35438
rect 10244 35314 12180 35382
rect 10244 35258 10254 35314
rect 10310 35258 10378 35314
rect 10434 35258 10502 35314
rect 10558 35258 10626 35314
rect 10682 35258 10750 35314
rect 10806 35258 10874 35314
rect 10930 35258 10998 35314
rect 11054 35258 11122 35314
rect 11178 35258 11246 35314
rect 11302 35258 11370 35314
rect 11426 35258 11494 35314
rect 11550 35258 11618 35314
rect 11674 35258 11742 35314
rect 11798 35258 11866 35314
rect 11922 35258 11990 35314
rect 12046 35258 12114 35314
rect 12170 35258 12180 35314
rect 10244 35190 12180 35258
rect 10244 35134 10254 35190
rect 10310 35134 10378 35190
rect 10434 35134 10502 35190
rect 10558 35134 10626 35190
rect 10682 35134 10750 35190
rect 10806 35134 10874 35190
rect 10930 35134 10998 35190
rect 11054 35134 11122 35190
rect 11178 35134 11246 35190
rect 11302 35134 11370 35190
rect 11426 35134 11494 35190
rect 11550 35134 11618 35190
rect 11674 35134 11742 35190
rect 11798 35134 11866 35190
rect 11922 35134 11990 35190
rect 12046 35134 12114 35190
rect 12170 35134 12180 35190
rect 10244 35066 12180 35134
rect 10244 35010 10254 35066
rect 10310 35010 10378 35066
rect 10434 35010 10502 35066
rect 10558 35010 10626 35066
rect 10682 35010 10750 35066
rect 10806 35010 10874 35066
rect 10930 35010 10998 35066
rect 11054 35010 11122 35066
rect 11178 35010 11246 35066
rect 11302 35010 11370 35066
rect 11426 35010 11494 35066
rect 11550 35010 11618 35066
rect 11674 35010 11742 35066
rect 11798 35010 11866 35066
rect 11922 35010 11990 35066
rect 12046 35010 12114 35066
rect 12170 35010 12180 35066
rect 10244 34942 12180 35010
rect 10244 34886 10254 34942
rect 10310 34886 10378 34942
rect 10434 34886 10502 34942
rect 10558 34886 10626 34942
rect 10682 34886 10750 34942
rect 10806 34886 10874 34942
rect 10930 34886 10998 34942
rect 11054 34886 11122 34942
rect 11178 34886 11246 34942
rect 11302 34886 11370 34942
rect 11426 34886 11494 34942
rect 11550 34886 11618 34942
rect 11674 34886 11742 34942
rect 11798 34886 11866 34942
rect 11922 34886 11990 34942
rect 12046 34886 12114 34942
rect 12170 34886 12180 34942
rect 10244 34818 12180 34886
rect 10244 34762 10254 34818
rect 10310 34762 10378 34818
rect 10434 34762 10502 34818
rect 10558 34762 10626 34818
rect 10682 34762 10750 34818
rect 10806 34762 10874 34818
rect 10930 34762 10998 34818
rect 11054 34762 11122 34818
rect 11178 34762 11246 34818
rect 11302 34762 11370 34818
rect 11426 34762 11494 34818
rect 11550 34762 11618 34818
rect 11674 34762 11742 34818
rect 11798 34762 11866 34818
rect 11922 34762 11990 34818
rect 12046 34762 12114 34818
rect 12170 34762 12180 34818
rect 10244 34694 12180 34762
rect 10244 34638 10254 34694
rect 10310 34638 10378 34694
rect 10434 34638 10502 34694
rect 10558 34638 10626 34694
rect 10682 34638 10750 34694
rect 10806 34638 10874 34694
rect 10930 34638 10998 34694
rect 11054 34638 11122 34694
rect 11178 34638 11246 34694
rect 11302 34638 11370 34694
rect 11426 34638 11494 34694
rect 11550 34638 11618 34694
rect 11674 34638 11742 34694
rect 11798 34638 11866 34694
rect 11922 34638 11990 34694
rect 12046 34638 12114 34694
rect 12170 34638 12180 34694
rect 10244 34570 12180 34638
rect 10244 34514 10254 34570
rect 10310 34514 10378 34570
rect 10434 34514 10502 34570
rect 10558 34514 10626 34570
rect 10682 34514 10750 34570
rect 10806 34514 10874 34570
rect 10930 34514 10998 34570
rect 11054 34514 11122 34570
rect 11178 34514 11246 34570
rect 11302 34514 11370 34570
rect 11426 34514 11494 34570
rect 11550 34514 11618 34570
rect 11674 34514 11742 34570
rect 11798 34514 11866 34570
rect 11922 34514 11990 34570
rect 12046 34514 12114 34570
rect 12170 34514 12180 34570
rect 10244 34446 12180 34514
rect 10244 34390 10254 34446
rect 10310 34390 10378 34446
rect 10434 34390 10502 34446
rect 10558 34390 10626 34446
rect 10682 34390 10750 34446
rect 10806 34390 10874 34446
rect 10930 34390 10998 34446
rect 11054 34390 11122 34446
rect 11178 34390 11246 34446
rect 11302 34390 11370 34446
rect 11426 34390 11494 34446
rect 11550 34390 11618 34446
rect 11674 34390 11742 34446
rect 11798 34390 11866 34446
rect 11922 34390 11990 34446
rect 12046 34390 12114 34446
rect 12170 34390 12180 34446
rect 10244 34322 12180 34390
rect 10244 34266 10254 34322
rect 10310 34266 10378 34322
rect 10434 34266 10502 34322
rect 10558 34266 10626 34322
rect 10682 34266 10750 34322
rect 10806 34266 10874 34322
rect 10930 34266 10998 34322
rect 11054 34266 11122 34322
rect 11178 34266 11246 34322
rect 11302 34266 11370 34322
rect 11426 34266 11494 34322
rect 11550 34266 11618 34322
rect 11674 34266 11742 34322
rect 11798 34266 11866 34322
rect 11922 34266 11990 34322
rect 12046 34266 12114 34322
rect 12170 34266 12180 34322
rect 10244 34198 12180 34266
rect 10244 34142 10254 34198
rect 10310 34142 10378 34198
rect 10434 34142 10502 34198
rect 10558 34142 10626 34198
rect 10682 34142 10750 34198
rect 10806 34142 10874 34198
rect 10930 34142 10998 34198
rect 11054 34142 11122 34198
rect 11178 34142 11246 34198
rect 11302 34142 11370 34198
rect 11426 34142 11494 34198
rect 11550 34142 11618 34198
rect 11674 34142 11742 34198
rect 11798 34142 11866 34198
rect 11922 34142 11990 34198
rect 12046 34142 12114 34198
rect 12170 34142 12180 34198
rect 10244 34074 12180 34142
rect 10244 34018 10254 34074
rect 10310 34018 10378 34074
rect 10434 34018 10502 34074
rect 10558 34018 10626 34074
rect 10682 34018 10750 34074
rect 10806 34018 10874 34074
rect 10930 34018 10998 34074
rect 11054 34018 11122 34074
rect 11178 34018 11246 34074
rect 11302 34018 11370 34074
rect 11426 34018 11494 34074
rect 11550 34018 11618 34074
rect 11674 34018 11742 34074
rect 11798 34018 11866 34074
rect 11922 34018 11990 34074
rect 12046 34018 12114 34074
rect 12170 34018 12180 34074
rect 10244 33950 12180 34018
rect 10244 33894 10254 33950
rect 10310 33894 10378 33950
rect 10434 33894 10502 33950
rect 10558 33894 10626 33950
rect 10682 33894 10750 33950
rect 10806 33894 10874 33950
rect 10930 33894 10998 33950
rect 11054 33894 11122 33950
rect 11178 33894 11246 33950
rect 11302 33894 11370 33950
rect 11426 33894 11494 33950
rect 11550 33894 11618 33950
rect 11674 33894 11742 33950
rect 11798 33894 11866 33950
rect 11922 33894 11990 33950
rect 12046 33894 12114 33950
rect 12170 33894 12180 33950
rect 10244 33826 12180 33894
rect 10244 33770 10254 33826
rect 10310 33770 10378 33826
rect 10434 33770 10502 33826
rect 10558 33770 10626 33826
rect 10682 33770 10750 33826
rect 10806 33770 10874 33826
rect 10930 33770 10998 33826
rect 11054 33770 11122 33826
rect 11178 33770 11246 33826
rect 11302 33770 11370 33826
rect 11426 33770 11494 33826
rect 11550 33770 11618 33826
rect 11674 33770 11742 33826
rect 11798 33770 11866 33826
rect 11922 33770 11990 33826
rect 12046 33770 12114 33826
rect 12170 33770 12180 33826
rect 10244 33702 12180 33770
rect 10244 33646 10254 33702
rect 10310 33646 10378 33702
rect 10434 33646 10502 33702
rect 10558 33646 10626 33702
rect 10682 33646 10750 33702
rect 10806 33646 10874 33702
rect 10930 33646 10998 33702
rect 11054 33646 11122 33702
rect 11178 33646 11246 33702
rect 11302 33646 11370 33702
rect 11426 33646 11494 33702
rect 11550 33646 11618 33702
rect 11674 33646 11742 33702
rect 11798 33646 11866 33702
rect 11922 33646 11990 33702
rect 12046 33646 12114 33702
rect 12170 33646 12180 33702
rect 10244 33636 12180 33646
rect 12861 36554 14673 36564
rect 12861 36498 12871 36554
rect 12927 36498 12995 36554
rect 13051 36498 13119 36554
rect 13175 36498 13243 36554
rect 13299 36498 13367 36554
rect 13423 36498 13491 36554
rect 13547 36498 13615 36554
rect 13671 36498 13739 36554
rect 13795 36498 13863 36554
rect 13919 36498 13987 36554
rect 14043 36498 14111 36554
rect 14167 36498 14235 36554
rect 14291 36498 14359 36554
rect 14415 36498 14483 36554
rect 14539 36498 14607 36554
rect 14663 36498 14673 36554
rect 12861 36430 14673 36498
rect 12861 36374 12871 36430
rect 12927 36374 12995 36430
rect 13051 36374 13119 36430
rect 13175 36374 13243 36430
rect 13299 36374 13367 36430
rect 13423 36374 13491 36430
rect 13547 36374 13615 36430
rect 13671 36374 13739 36430
rect 13795 36374 13863 36430
rect 13919 36374 13987 36430
rect 14043 36374 14111 36430
rect 14167 36374 14235 36430
rect 14291 36374 14359 36430
rect 14415 36374 14483 36430
rect 14539 36374 14607 36430
rect 14663 36374 14673 36430
rect 12861 36306 14673 36374
rect 12861 36250 12871 36306
rect 12927 36250 12995 36306
rect 13051 36250 13119 36306
rect 13175 36250 13243 36306
rect 13299 36250 13367 36306
rect 13423 36250 13491 36306
rect 13547 36250 13615 36306
rect 13671 36250 13739 36306
rect 13795 36250 13863 36306
rect 13919 36250 13987 36306
rect 14043 36250 14111 36306
rect 14167 36250 14235 36306
rect 14291 36250 14359 36306
rect 14415 36250 14483 36306
rect 14539 36250 14607 36306
rect 14663 36250 14673 36306
rect 12861 36182 14673 36250
rect 12861 36126 12871 36182
rect 12927 36126 12995 36182
rect 13051 36126 13119 36182
rect 13175 36126 13243 36182
rect 13299 36126 13367 36182
rect 13423 36126 13491 36182
rect 13547 36126 13615 36182
rect 13671 36126 13739 36182
rect 13795 36126 13863 36182
rect 13919 36126 13987 36182
rect 14043 36126 14111 36182
rect 14167 36126 14235 36182
rect 14291 36126 14359 36182
rect 14415 36126 14483 36182
rect 14539 36126 14607 36182
rect 14663 36126 14673 36182
rect 12861 36058 14673 36126
rect 12861 36002 12871 36058
rect 12927 36002 12995 36058
rect 13051 36002 13119 36058
rect 13175 36002 13243 36058
rect 13299 36002 13367 36058
rect 13423 36002 13491 36058
rect 13547 36002 13615 36058
rect 13671 36002 13739 36058
rect 13795 36002 13863 36058
rect 13919 36002 13987 36058
rect 14043 36002 14111 36058
rect 14167 36002 14235 36058
rect 14291 36002 14359 36058
rect 14415 36002 14483 36058
rect 14539 36002 14607 36058
rect 14663 36002 14673 36058
rect 12861 35934 14673 36002
rect 12861 35878 12871 35934
rect 12927 35878 12995 35934
rect 13051 35878 13119 35934
rect 13175 35878 13243 35934
rect 13299 35878 13367 35934
rect 13423 35878 13491 35934
rect 13547 35878 13615 35934
rect 13671 35878 13739 35934
rect 13795 35878 13863 35934
rect 13919 35878 13987 35934
rect 14043 35878 14111 35934
rect 14167 35878 14235 35934
rect 14291 35878 14359 35934
rect 14415 35878 14483 35934
rect 14539 35878 14607 35934
rect 14663 35878 14673 35934
rect 12861 35810 14673 35878
rect 12861 35754 12871 35810
rect 12927 35754 12995 35810
rect 13051 35754 13119 35810
rect 13175 35754 13243 35810
rect 13299 35754 13367 35810
rect 13423 35754 13491 35810
rect 13547 35754 13615 35810
rect 13671 35754 13739 35810
rect 13795 35754 13863 35810
rect 13919 35754 13987 35810
rect 14043 35754 14111 35810
rect 14167 35754 14235 35810
rect 14291 35754 14359 35810
rect 14415 35754 14483 35810
rect 14539 35754 14607 35810
rect 14663 35754 14673 35810
rect 12861 35686 14673 35754
rect 12861 35630 12871 35686
rect 12927 35630 12995 35686
rect 13051 35630 13119 35686
rect 13175 35630 13243 35686
rect 13299 35630 13367 35686
rect 13423 35630 13491 35686
rect 13547 35630 13615 35686
rect 13671 35630 13739 35686
rect 13795 35630 13863 35686
rect 13919 35630 13987 35686
rect 14043 35630 14111 35686
rect 14167 35630 14235 35686
rect 14291 35630 14359 35686
rect 14415 35630 14483 35686
rect 14539 35630 14607 35686
rect 14663 35630 14673 35686
rect 12861 35562 14673 35630
rect 12861 35506 12871 35562
rect 12927 35506 12995 35562
rect 13051 35506 13119 35562
rect 13175 35506 13243 35562
rect 13299 35506 13367 35562
rect 13423 35506 13491 35562
rect 13547 35506 13615 35562
rect 13671 35506 13739 35562
rect 13795 35506 13863 35562
rect 13919 35506 13987 35562
rect 14043 35506 14111 35562
rect 14167 35506 14235 35562
rect 14291 35506 14359 35562
rect 14415 35506 14483 35562
rect 14539 35506 14607 35562
rect 14663 35506 14673 35562
rect 12861 35438 14673 35506
rect 12861 35382 12871 35438
rect 12927 35382 12995 35438
rect 13051 35382 13119 35438
rect 13175 35382 13243 35438
rect 13299 35382 13367 35438
rect 13423 35382 13491 35438
rect 13547 35382 13615 35438
rect 13671 35382 13739 35438
rect 13795 35382 13863 35438
rect 13919 35382 13987 35438
rect 14043 35382 14111 35438
rect 14167 35382 14235 35438
rect 14291 35382 14359 35438
rect 14415 35382 14483 35438
rect 14539 35382 14607 35438
rect 14663 35382 14673 35438
rect 12861 35314 14673 35382
rect 12861 35258 12871 35314
rect 12927 35258 12995 35314
rect 13051 35258 13119 35314
rect 13175 35258 13243 35314
rect 13299 35258 13367 35314
rect 13423 35258 13491 35314
rect 13547 35258 13615 35314
rect 13671 35258 13739 35314
rect 13795 35258 13863 35314
rect 13919 35258 13987 35314
rect 14043 35258 14111 35314
rect 14167 35258 14235 35314
rect 14291 35258 14359 35314
rect 14415 35258 14483 35314
rect 14539 35258 14607 35314
rect 14663 35258 14673 35314
rect 12861 35190 14673 35258
rect 12861 35134 12871 35190
rect 12927 35134 12995 35190
rect 13051 35134 13119 35190
rect 13175 35134 13243 35190
rect 13299 35134 13367 35190
rect 13423 35134 13491 35190
rect 13547 35134 13615 35190
rect 13671 35134 13739 35190
rect 13795 35134 13863 35190
rect 13919 35134 13987 35190
rect 14043 35134 14111 35190
rect 14167 35134 14235 35190
rect 14291 35134 14359 35190
rect 14415 35134 14483 35190
rect 14539 35134 14607 35190
rect 14663 35134 14673 35190
rect 12861 35066 14673 35134
rect 12861 35010 12871 35066
rect 12927 35010 12995 35066
rect 13051 35010 13119 35066
rect 13175 35010 13243 35066
rect 13299 35010 13367 35066
rect 13423 35010 13491 35066
rect 13547 35010 13615 35066
rect 13671 35010 13739 35066
rect 13795 35010 13863 35066
rect 13919 35010 13987 35066
rect 14043 35010 14111 35066
rect 14167 35010 14235 35066
rect 14291 35010 14359 35066
rect 14415 35010 14483 35066
rect 14539 35010 14607 35066
rect 14663 35010 14673 35066
rect 12861 34942 14673 35010
rect 12861 34886 12871 34942
rect 12927 34886 12995 34942
rect 13051 34886 13119 34942
rect 13175 34886 13243 34942
rect 13299 34886 13367 34942
rect 13423 34886 13491 34942
rect 13547 34886 13615 34942
rect 13671 34886 13739 34942
rect 13795 34886 13863 34942
rect 13919 34886 13987 34942
rect 14043 34886 14111 34942
rect 14167 34886 14235 34942
rect 14291 34886 14359 34942
rect 14415 34886 14483 34942
rect 14539 34886 14607 34942
rect 14663 34886 14673 34942
rect 12861 34818 14673 34886
rect 12861 34762 12871 34818
rect 12927 34762 12995 34818
rect 13051 34762 13119 34818
rect 13175 34762 13243 34818
rect 13299 34762 13367 34818
rect 13423 34762 13491 34818
rect 13547 34762 13615 34818
rect 13671 34762 13739 34818
rect 13795 34762 13863 34818
rect 13919 34762 13987 34818
rect 14043 34762 14111 34818
rect 14167 34762 14235 34818
rect 14291 34762 14359 34818
rect 14415 34762 14483 34818
rect 14539 34762 14607 34818
rect 14663 34762 14673 34818
rect 12861 34694 14673 34762
rect 12861 34638 12871 34694
rect 12927 34638 12995 34694
rect 13051 34638 13119 34694
rect 13175 34638 13243 34694
rect 13299 34638 13367 34694
rect 13423 34638 13491 34694
rect 13547 34638 13615 34694
rect 13671 34638 13739 34694
rect 13795 34638 13863 34694
rect 13919 34638 13987 34694
rect 14043 34638 14111 34694
rect 14167 34638 14235 34694
rect 14291 34638 14359 34694
rect 14415 34638 14483 34694
rect 14539 34638 14607 34694
rect 14663 34638 14673 34694
rect 12861 34570 14673 34638
rect 12861 34514 12871 34570
rect 12927 34514 12995 34570
rect 13051 34514 13119 34570
rect 13175 34514 13243 34570
rect 13299 34514 13367 34570
rect 13423 34514 13491 34570
rect 13547 34514 13615 34570
rect 13671 34514 13739 34570
rect 13795 34514 13863 34570
rect 13919 34514 13987 34570
rect 14043 34514 14111 34570
rect 14167 34514 14235 34570
rect 14291 34514 14359 34570
rect 14415 34514 14483 34570
rect 14539 34514 14607 34570
rect 14663 34514 14673 34570
rect 12861 34446 14673 34514
rect 12861 34390 12871 34446
rect 12927 34390 12995 34446
rect 13051 34390 13119 34446
rect 13175 34390 13243 34446
rect 13299 34390 13367 34446
rect 13423 34390 13491 34446
rect 13547 34390 13615 34446
rect 13671 34390 13739 34446
rect 13795 34390 13863 34446
rect 13919 34390 13987 34446
rect 14043 34390 14111 34446
rect 14167 34390 14235 34446
rect 14291 34390 14359 34446
rect 14415 34390 14483 34446
rect 14539 34390 14607 34446
rect 14663 34390 14673 34446
rect 12861 34322 14673 34390
rect 12861 34266 12871 34322
rect 12927 34266 12995 34322
rect 13051 34266 13119 34322
rect 13175 34266 13243 34322
rect 13299 34266 13367 34322
rect 13423 34266 13491 34322
rect 13547 34266 13615 34322
rect 13671 34266 13739 34322
rect 13795 34266 13863 34322
rect 13919 34266 13987 34322
rect 14043 34266 14111 34322
rect 14167 34266 14235 34322
rect 14291 34266 14359 34322
rect 14415 34266 14483 34322
rect 14539 34266 14607 34322
rect 14663 34266 14673 34322
rect 12861 34198 14673 34266
rect 12861 34142 12871 34198
rect 12927 34142 12995 34198
rect 13051 34142 13119 34198
rect 13175 34142 13243 34198
rect 13299 34142 13367 34198
rect 13423 34142 13491 34198
rect 13547 34142 13615 34198
rect 13671 34142 13739 34198
rect 13795 34142 13863 34198
rect 13919 34142 13987 34198
rect 14043 34142 14111 34198
rect 14167 34142 14235 34198
rect 14291 34142 14359 34198
rect 14415 34142 14483 34198
rect 14539 34142 14607 34198
rect 14663 34142 14673 34198
rect 12861 34074 14673 34142
rect 12861 34018 12871 34074
rect 12927 34018 12995 34074
rect 13051 34018 13119 34074
rect 13175 34018 13243 34074
rect 13299 34018 13367 34074
rect 13423 34018 13491 34074
rect 13547 34018 13615 34074
rect 13671 34018 13739 34074
rect 13795 34018 13863 34074
rect 13919 34018 13987 34074
rect 14043 34018 14111 34074
rect 14167 34018 14235 34074
rect 14291 34018 14359 34074
rect 14415 34018 14483 34074
rect 14539 34018 14607 34074
rect 14663 34018 14673 34074
rect 12861 33950 14673 34018
rect 12861 33894 12871 33950
rect 12927 33894 12995 33950
rect 13051 33894 13119 33950
rect 13175 33894 13243 33950
rect 13299 33894 13367 33950
rect 13423 33894 13491 33950
rect 13547 33894 13615 33950
rect 13671 33894 13739 33950
rect 13795 33894 13863 33950
rect 13919 33894 13987 33950
rect 14043 33894 14111 33950
rect 14167 33894 14235 33950
rect 14291 33894 14359 33950
rect 14415 33894 14483 33950
rect 14539 33894 14607 33950
rect 14663 33894 14673 33950
rect 12861 33826 14673 33894
rect 12861 33770 12871 33826
rect 12927 33770 12995 33826
rect 13051 33770 13119 33826
rect 13175 33770 13243 33826
rect 13299 33770 13367 33826
rect 13423 33770 13491 33826
rect 13547 33770 13615 33826
rect 13671 33770 13739 33826
rect 13795 33770 13863 33826
rect 13919 33770 13987 33826
rect 14043 33770 14111 33826
rect 14167 33770 14235 33826
rect 14291 33770 14359 33826
rect 14415 33770 14483 33826
rect 14539 33770 14607 33826
rect 14663 33770 14673 33826
rect 12861 33702 14673 33770
rect 12861 33646 12871 33702
rect 12927 33646 12995 33702
rect 13051 33646 13119 33702
rect 13175 33646 13243 33702
rect 13299 33646 13367 33702
rect 13423 33646 13491 33702
rect 13547 33646 13615 33702
rect 13671 33646 13739 33702
rect 13795 33646 13863 33702
rect 13919 33646 13987 33702
rect 14043 33646 14111 33702
rect 14167 33646 14235 33702
rect 14291 33646 14359 33702
rect 14415 33646 14483 33702
rect 14539 33646 14607 33702
rect 14663 33646 14673 33702
rect 12861 33636 14673 33646
rect 10 33604 86 33614
rect 14892 33614 14902 36586
rect 14958 33614 14968 36586
rect 14892 33604 14968 33614
rect 2481 33354 2681 33364
rect 2481 33298 2491 33354
rect 2547 33298 2615 33354
rect 2671 33298 2681 33354
rect 2481 33230 2681 33298
rect 2481 33174 2491 33230
rect 2547 33174 2615 33230
rect 2671 33174 2681 33230
rect 2481 33106 2681 33174
rect 2481 33050 2491 33106
rect 2547 33050 2615 33106
rect 2671 33050 2681 33106
rect 2481 32982 2681 33050
rect 2481 32926 2491 32982
rect 2547 32926 2615 32982
rect 2671 32926 2681 32982
rect 2481 32858 2681 32926
rect 2481 32802 2491 32858
rect 2547 32802 2615 32858
rect 2671 32802 2681 32858
rect 2481 32734 2681 32802
rect 2481 32678 2491 32734
rect 2547 32678 2615 32734
rect 2671 32678 2681 32734
rect 2481 32610 2681 32678
rect 2481 32554 2491 32610
rect 2547 32554 2615 32610
rect 2671 32554 2681 32610
rect 2481 32486 2681 32554
rect 2481 32430 2491 32486
rect 2547 32430 2615 32486
rect 2671 32430 2681 32486
rect 2481 32362 2681 32430
rect 2481 32306 2491 32362
rect 2547 32306 2615 32362
rect 2671 32306 2681 32362
rect 2481 32238 2681 32306
rect 2481 32182 2491 32238
rect 2547 32182 2615 32238
rect 2671 32182 2681 32238
rect 2481 32114 2681 32182
rect 2481 32058 2491 32114
rect 2547 32058 2615 32114
rect 2671 32058 2681 32114
rect 2481 31990 2681 32058
rect 2481 31934 2491 31990
rect 2547 31934 2615 31990
rect 2671 31934 2681 31990
rect 2481 31866 2681 31934
rect 2481 31810 2491 31866
rect 2547 31810 2615 31866
rect 2671 31810 2681 31866
rect 2481 31742 2681 31810
rect 2481 31686 2491 31742
rect 2547 31686 2615 31742
rect 2671 31686 2681 31742
rect 2481 31618 2681 31686
rect 2481 31562 2491 31618
rect 2547 31562 2615 31618
rect 2671 31562 2681 31618
rect 2481 31494 2681 31562
rect 2481 31438 2491 31494
rect 2547 31438 2615 31494
rect 2671 31438 2681 31494
rect 2481 31370 2681 31438
rect 2481 31314 2491 31370
rect 2547 31314 2615 31370
rect 2671 31314 2681 31370
rect 2481 31246 2681 31314
rect 2481 31190 2491 31246
rect 2547 31190 2615 31246
rect 2671 31190 2681 31246
rect 2481 31122 2681 31190
rect 2481 31066 2491 31122
rect 2547 31066 2615 31122
rect 2671 31066 2681 31122
rect 2481 30998 2681 31066
rect 2481 30942 2491 30998
rect 2547 30942 2615 30998
rect 2671 30942 2681 30998
rect 2481 30874 2681 30942
rect 2481 30818 2491 30874
rect 2547 30818 2615 30874
rect 2671 30818 2681 30874
rect 2481 30750 2681 30818
rect 2481 30694 2491 30750
rect 2547 30694 2615 30750
rect 2671 30694 2681 30750
rect 2481 30626 2681 30694
rect 2481 30570 2491 30626
rect 2547 30570 2615 30626
rect 2671 30570 2681 30626
rect 2481 30502 2681 30570
rect 2481 30446 2491 30502
rect 2547 30446 2615 30502
rect 2671 30446 2681 30502
rect 2481 30436 2681 30446
rect 4851 33354 5051 33364
rect 4851 33298 4861 33354
rect 4917 33298 4985 33354
rect 5041 33298 5051 33354
rect 4851 33230 5051 33298
rect 4851 33174 4861 33230
rect 4917 33174 4985 33230
rect 5041 33174 5051 33230
rect 4851 33106 5051 33174
rect 4851 33050 4861 33106
rect 4917 33050 4985 33106
rect 5041 33050 5051 33106
rect 4851 32982 5051 33050
rect 4851 32926 4861 32982
rect 4917 32926 4985 32982
rect 5041 32926 5051 32982
rect 4851 32858 5051 32926
rect 4851 32802 4861 32858
rect 4917 32802 4985 32858
rect 5041 32802 5051 32858
rect 4851 32734 5051 32802
rect 4851 32678 4861 32734
rect 4917 32678 4985 32734
rect 5041 32678 5051 32734
rect 4851 32610 5051 32678
rect 4851 32554 4861 32610
rect 4917 32554 4985 32610
rect 5041 32554 5051 32610
rect 4851 32486 5051 32554
rect 4851 32430 4861 32486
rect 4917 32430 4985 32486
rect 5041 32430 5051 32486
rect 4851 32362 5051 32430
rect 4851 32306 4861 32362
rect 4917 32306 4985 32362
rect 5041 32306 5051 32362
rect 4851 32238 5051 32306
rect 4851 32182 4861 32238
rect 4917 32182 4985 32238
rect 5041 32182 5051 32238
rect 4851 32114 5051 32182
rect 4851 32058 4861 32114
rect 4917 32058 4985 32114
rect 5041 32058 5051 32114
rect 4851 31990 5051 32058
rect 4851 31934 4861 31990
rect 4917 31934 4985 31990
rect 5041 31934 5051 31990
rect 4851 31866 5051 31934
rect 4851 31810 4861 31866
rect 4917 31810 4985 31866
rect 5041 31810 5051 31866
rect 4851 31742 5051 31810
rect 4851 31686 4861 31742
rect 4917 31686 4985 31742
rect 5041 31686 5051 31742
rect 4851 31618 5051 31686
rect 4851 31562 4861 31618
rect 4917 31562 4985 31618
rect 5041 31562 5051 31618
rect 4851 31494 5051 31562
rect 4851 31438 4861 31494
rect 4917 31438 4985 31494
rect 5041 31438 5051 31494
rect 4851 31370 5051 31438
rect 4851 31314 4861 31370
rect 4917 31314 4985 31370
rect 5041 31314 5051 31370
rect 4851 31246 5051 31314
rect 4851 31190 4861 31246
rect 4917 31190 4985 31246
rect 5041 31190 5051 31246
rect 4851 31122 5051 31190
rect 4851 31066 4861 31122
rect 4917 31066 4985 31122
rect 5041 31066 5051 31122
rect 4851 30998 5051 31066
rect 4851 30942 4861 30998
rect 4917 30942 4985 30998
rect 5041 30942 5051 30998
rect 4851 30874 5051 30942
rect 4851 30818 4861 30874
rect 4917 30818 4985 30874
rect 5041 30818 5051 30874
rect 4851 30750 5051 30818
rect 4851 30694 4861 30750
rect 4917 30694 4985 30750
rect 5041 30694 5051 30750
rect 4851 30626 5051 30694
rect 4851 30570 4861 30626
rect 4917 30570 4985 30626
rect 5041 30570 5051 30626
rect 4851 30502 5051 30570
rect 4851 30446 4861 30502
rect 4917 30446 4985 30502
rect 5041 30446 5051 30502
rect 4851 30436 5051 30446
rect 7265 33354 7713 33364
rect 7265 33298 7275 33354
rect 7331 33298 7399 33354
rect 7455 33298 7523 33354
rect 7579 33298 7647 33354
rect 7703 33298 7713 33354
rect 7265 33230 7713 33298
rect 7265 33174 7275 33230
rect 7331 33174 7399 33230
rect 7455 33174 7523 33230
rect 7579 33174 7647 33230
rect 7703 33174 7713 33230
rect 7265 33106 7713 33174
rect 7265 33050 7275 33106
rect 7331 33050 7399 33106
rect 7455 33050 7523 33106
rect 7579 33050 7647 33106
rect 7703 33050 7713 33106
rect 7265 32982 7713 33050
rect 7265 32926 7275 32982
rect 7331 32926 7399 32982
rect 7455 32926 7523 32982
rect 7579 32926 7647 32982
rect 7703 32926 7713 32982
rect 7265 32858 7713 32926
rect 7265 32802 7275 32858
rect 7331 32802 7399 32858
rect 7455 32802 7523 32858
rect 7579 32802 7647 32858
rect 7703 32802 7713 32858
rect 7265 32734 7713 32802
rect 7265 32678 7275 32734
rect 7331 32678 7399 32734
rect 7455 32678 7523 32734
rect 7579 32678 7647 32734
rect 7703 32678 7713 32734
rect 7265 32610 7713 32678
rect 7265 32554 7275 32610
rect 7331 32554 7399 32610
rect 7455 32554 7523 32610
rect 7579 32554 7647 32610
rect 7703 32554 7713 32610
rect 7265 32486 7713 32554
rect 7265 32430 7275 32486
rect 7331 32430 7399 32486
rect 7455 32430 7523 32486
rect 7579 32430 7647 32486
rect 7703 32430 7713 32486
rect 7265 32362 7713 32430
rect 7265 32306 7275 32362
rect 7331 32306 7399 32362
rect 7455 32306 7523 32362
rect 7579 32306 7647 32362
rect 7703 32306 7713 32362
rect 7265 32238 7713 32306
rect 7265 32182 7275 32238
rect 7331 32182 7399 32238
rect 7455 32182 7523 32238
rect 7579 32182 7647 32238
rect 7703 32182 7713 32238
rect 7265 32114 7713 32182
rect 7265 32058 7275 32114
rect 7331 32058 7399 32114
rect 7455 32058 7523 32114
rect 7579 32058 7647 32114
rect 7703 32058 7713 32114
rect 7265 31990 7713 32058
rect 7265 31934 7275 31990
rect 7331 31934 7399 31990
rect 7455 31934 7523 31990
rect 7579 31934 7647 31990
rect 7703 31934 7713 31990
rect 7265 31866 7713 31934
rect 7265 31810 7275 31866
rect 7331 31810 7399 31866
rect 7455 31810 7523 31866
rect 7579 31810 7647 31866
rect 7703 31810 7713 31866
rect 7265 31742 7713 31810
rect 7265 31686 7275 31742
rect 7331 31686 7399 31742
rect 7455 31686 7523 31742
rect 7579 31686 7647 31742
rect 7703 31686 7713 31742
rect 7265 31618 7713 31686
rect 7265 31562 7275 31618
rect 7331 31562 7399 31618
rect 7455 31562 7523 31618
rect 7579 31562 7647 31618
rect 7703 31562 7713 31618
rect 7265 31494 7713 31562
rect 7265 31438 7275 31494
rect 7331 31438 7399 31494
rect 7455 31438 7523 31494
rect 7579 31438 7647 31494
rect 7703 31438 7713 31494
rect 7265 31370 7713 31438
rect 7265 31314 7275 31370
rect 7331 31314 7399 31370
rect 7455 31314 7523 31370
rect 7579 31314 7647 31370
rect 7703 31314 7713 31370
rect 7265 31246 7713 31314
rect 7265 31190 7275 31246
rect 7331 31190 7399 31246
rect 7455 31190 7523 31246
rect 7579 31190 7647 31246
rect 7703 31190 7713 31246
rect 7265 31122 7713 31190
rect 7265 31066 7275 31122
rect 7331 31066 7399 31122
rect 7455 31066 7523 31122
rect 7579 31066 7647 31122
rect 7703 31066 7713 31122
rect 7265 30998 7713 31066
rect 7265 30942 7275 30998
rect 7331 30942 7399 30998
rect 7455 30942 7523 30998
rect 7579 30942 7647 30998
rect 7703 30942 7713 30998
rect 7265 30874 7713 30942
rect 7265 30818 7275 30874
rect 7331 30818 7399 30874
rect 7455 30818 7523 30874
rect 7579 30818 7647 30874
rect 7703 30818 7713 30874
rect 7265 30750 7713 30818
rect 7265 30694 7275 30750
rect 7331 30694 7399 30750
rect 7455 30694 7523 30750
rect 7579 30694 7647 30750
rect 7703 30694 7713 30750
rect 7265 30626 7713 30694
rect 7265 30570 7275 30626
rect 7331 30570 7399 30626
rect 7455 30570 7523 30626
rect 7579 30570 7647 30626
rect 7703 30570 7713 30626
rect 7265 30502 7713 30570
rect 7265 30446 7275 30502
rect 7331 30446 7399 30502
rect 7455 30446 7523 30502
rect 7579 30446 7647 30502
rect 7703 30446 7713 30502
rect 7265 30436 7713 30446
rect 9927 33354 10127 33364
rect 9927 33298 9937 33354
rect 9993 33298 10061 33354
rect 10117 33298 10127 33354
rect 9927 33230 10127 33298
rect 9927 33174 9937 33230
rect 9993 33174 10061 33230
rect 10117 33174 10127 33230
rect 9927 33106 10127 33174
rect 9927 33050 9937 33106
rect 9993 33050 10061 33106
rect 10117 33050 10127 33106
rect 9927 32982 10127 33050
rect 9927 32926 9937 32982
rect 9993 32926 10061 32982
rect 10117 32926 10127 32982
rect 9927 32858 10127 32926
rect 9927 32802 9937 32858
rect 9993 32802 10061 32858
rect 10117 32802 10127 32858
rect 9927 32734 10127 32802
rect 9927 32678 9937 32734
rect 9993 32678 10061 32734
rect 10117 32678 10127 32734
rect 9927 32610 10127 32678
rect 9927 32554 9937 32610
rect 9993 32554 10061 32610
rect 10117 32554 10127 32610
rect 9927 32486 10127 32554
rect 9927 32430 9937 32486
rect 9993 32430 10061 32486
rect 10117 32430 10127 32486
rect 9927 32362 10127 32430
rect 9927 32306 9937 32362
rect 9993 32306 10061 32362
rect 10117 32306 10127 32362
rect 9927 32238 10127 32306
rect 9927 32182 9937 32238
rect 9993 32182 10061 32238
rect 10117 32182 10127 32238
rect 9927 32114 10127 32182
rect 9927 32058 9937 32114
rect 9993 32058 10061 32114
rect 10117 32058 10127 32114
rect 9927 31990 10127 32058
rect 9927 31934 9937 31990
rect 9993 31934 10061 31990
rect 10117 31934 10127 31990
rect 9927 31866 10127 31934
rect 9927 31810 9937 31866
rect 9993 31810 10061 31866
rect 10117 31810 10127 31866
rect 9927 31742 10127 31810
rect 9927 31686 9937 31742
rect 9993 31686 10061 31742
rect 10117 31686 10127 31742
rect 9927 31618 10127 31686
rect 9927 31562 9937 31618
rect 9993 31562 10061 31618
rect 10117 31562 10127 31618
rect 9927 31494 10127 31562
rect 9927 31438 9937 31494
rect 9993 31438 10061 31494
rect 10117 31438 10127 31494
rect 9927 31370 10127 31438
rect 9927 31314 9937 31370
rect 9993 31314 10061 31370
rect 10117 31314 10127 31370
rect 9927 31246 10127 31314
rect 9927 31190 9937 31246
rect 9993 31190 10061 31246
rect 10117 31190 10127 31246
rect 9927 31122 10127 31190
rect 9927 31066 9937 31122
rect 9993 31066 10061 31122
rect 10117 31066 10127 31122
rect 9927 30998 10127 31066
rect 9927 30942 9937 30998
rect 9993 30942 10061 30998
rect 10117 30942 10127 30998
rect 9927 30874 10127 30942
rect 9927 30818 9937 30874
rect 9993 30818 10061 30874
rect 10117 30818 10127 30874
rect 9927 30750 10127 30818
rect 9927 30694 9937 30750
rect 9993 30694 10061 30750
rect 10117 30694 10127 30750
rect 9927 30626 10127 30694
rect 9927 30570 9937 30626
rect 9993 30570 10061 30626
rect 10117 30570 10127 30626
rect 9927 30502 10127 30570
rect 9927 30446 9937 30502
rect 9993 30446 10061 30502
rect 10117 30446 10127 30502
rect 9927 30436 10127 30446
rect 12297 33354 12497 33364
rect 12297 33298 12307 33354
rect 12363 33298 12431 33354
rect 12487 33298 12497 33354
rect 12297 33230 12497 33298
rect 12297 33174 12307 33230
rect 12363 33174 12431 33230
rect 12487 33174 12497 33230
rect 12297 33106 12497 33174
rect 12297 33050 12307 33106
rect 12363 33050 12431 33106
rect 12487 33050 12497 33106
rect 12297 32982 12497 33050
rect 12297 32926 12307 32982
rect 12363 32926 12431 32982
rect 12487 32926 12497 32982
rect 12297 32858 12497 32926
rect 12297 32802 12307 32858
rect 12363 32802 12431 32858
rect 12487 32802 12497 32858
rect 12297 32734 12497 32802
rect 12297 32678 12307 32734
rect 12363 32678 12431 32734
rect 12487 32678 12497 32734
rect 12297 32610 12497 32678
rect 12297 32554 12307 32610
rect 12363 32554 12431 32610
rect 12487 32554 12497 32610
rect 12297 32486 12497 32554
rect 12297 32430 12307 32486
rect 12363 32430 12431 32486
rect 12487 32430 12497 32486
rect 12297 32362 12497 32430
rect 12297 32306 12307 32362
rect 12363 32306 12431 32362
rect 12487 32306 12497 32362
rect 12297 32238 12497 32306
rect 12297 32182 12307 32238
rect 12363 32182 12431 32238
rect 12487 32182 12497 32238
rect 12297 32114 12497 32182
rect 12297 32058 12307 32114
rect 12363 32058 12431 32114
rect 12487 32058 12497 32114
rect 12297 31990 12497 32058
rect 12297 31934 12307 31990
rect 12363 31934 12431 31990
rect 12487 31934 12497 31990
rect 12297 31866 12497 31934
rect 12297 31810 12307 31866
rect 12363 31810 12431 31866
rect 12487 31810 12497 31866
rect 12297 31742 12497 31810
rect 12297 31686 12307 31742
rect 12363 31686 12431 31742
rect 12487 31686 12497 31742
rect 12297 31618 12497 31686
rect 12297 31562 12307 31618
rect 12363 31562 12431 31618
rect 12487 31562 12497 31618
rect 12297 31494 12497 31562
rect 12297 31438 12307 31494
rect 12363 31438 12431 31494
rect 12487 31438 12497 31494
rect 12297 31370 12497 31438
rect 12297 31314 12307 31370
rect 12363 31314 12431 31370
rect 12487 31314 12497 31370
rect 12297 31246 12497 31314
rect 12297 31190 12307 31246
rect 12363 31190 12431 31246
rect 12487 31190 12497 31246
rect 12297 31122 12497 31190
rect 12297 31066 12307 31122
rect 12363 31066 12431 31122
rect 12487 31066 12497 31122
rect 12297 30998 12497 31066
rect 12297 30942 12307 30998
rect 12363 30942 12431 30998
rect 12487 30942 12497 30998
rect 12297 30874 12497 30942
rect 12297 30818 12307 30874
rect 12363 30818 12431 30874
rect 12487 30818 12497 30874
rect 12297 30750 12497 30818
rect 12297 30694 12307 30750
rect 12363 30694 12431 30750
rect 12487 30694 12497 30750
rect 12297 30626 12497 30694
rect 12297 30570 12307 30626
rect 12363 30570 12431 30626
rect 12487 30570 12497 30626
rect 12297 30502 12497 30570
rect 12297 30446 12307 30502
rect 12363 30446 12431 30502
rect 12487 30446 12497 30502
rect 12297 30436 12497 30446
rect 2481 30148 2681 30158
rect 2481 30092 2491 30148
rect 2547 30092 2615 30148
rect 2671 30092 2681 30148
rect 2481 30024 2681 30092
rect 2481 29968 2491 30024
rect 2547 29968 2615 30024
rect 2671 29968 2681 30024
rect 2481 29900 2681 29968
rect 2481 29844 2491 29900
rect 2547 29844 2615 29900
rect 2671 29844 2681 29900
rect 2481 29776 2681 29844
rect 2481 29720 2491 29776
rect 2547 29720 2615 29776
rect 2671 29720 2681 29776
rect 2481 29652 2681 29720
rect 2481 29596 2491 29652
rect 2547 29596 2615 29652
rect 2671 29596 2681 29652
rect 2481 29528 2681 29596
rect 2481 29472 2491 29528
rect 2547 29472 2615 29528
rect 2671 29472 2681 29528
rect 2481 29404 2681 29472
rect 2481 29348 2491 29404
rect 2547 29348 2615 29404
rect 2671 29348 2681 29404
rect 2481 29280 2681 29348
rect 2481 29224 2491 29280
rect 2547 29224 2615 29280
rect 2671 29224 2681 29280
rect 2481 29156 2681 29224
rect 2481 29100 2491 29156
rect 2547 29100 2615 29156
rect 2671 29100 2681 29156
rect 2481 29032 2681 29100
rect 2481 28976 2491 29032
rect 2547 28976 2615 29032
rect 2671 28976 2681 29032
rect 2481 28908 2681 28976
rect 2481 28852 2491 28908
rect 2547 28852 2615 28908
rect 2671 28852 2681 28908
rect 2481 28842 2681 28852
rect 4851 30148 5051 30158
rect 4851 30092 4861 30148
rect 4917 30092 4985 30148
rect 5041 30092 5051 30148
rect 4851 30024 5051 30092
rect 4851 29968 4861 30024
rect 4917 29968 4985 30024
rect 5041 29968 5051 30024
rect 4851 29900 5051 29968
rect 4851 29844 4861 29900
rect 4917 29844 4985 29900
rect 5041 29844 5051 29900
rect 4851 29776 5051 29844
rect 4851 29720 4861 29776
rect 4917 29720 4985 29776
rect 5041 29720 5051 29776
rect 4851 29652 5051 29720
rect 4851 29596 4861 29652
rect 4917 29596 4985 29652
rect 5041 29596 5051 29652
rect 4851 29528 5051 29596
rect 4851 29472 4861 29528
rect 4917 29472 4985 29528
rect 5041 29472 5051 29528
rect 4851 29404 5051 29472
rect 4851 29348 4861 29404
rect 4917 29348 4985 29404
rect 5041 29348 5051 29404
rect 4851 29280 5051 29348
rect 4851 29224 4861 29280
rect 4917 29224 4985 29280
rect 5041 29224 5051 29280
rect 4851 29156 5051 29224
rect 4851 29100 4861 29156
rect 4917 29100 4985 29156
rect 5041 29100 5051 29156
rect 4851 29032 5051 29100
rect 4851 28976 4861 29032
rect 4917 28976 4985 29032
rect 5041 28976 5051 29032
rect 4851 28908 5051 28976
rect 4851 28852 4861 28908
rect 4917 28852 4985 28908
rect 5041 28852 5051 28908
rect 4851 28842 5051 28852
rect 7265 30148 7713 30158
rect 7265 30092 7275 30148
rect 7331 30092 7399 30148
rect 7455 30092 7523 30148
rect 7579 30092 7647 30148
rect 7703 30092 7713 30148
rect 7265 30024 7713 30092
rect 7265 29968 7275 30024
rect 7331 29968 7399 30024
rect 7455 29968 7523 30024
rect 7579 29968 7647 30024
rect 7703 29968 7713 30024
rect 7265 29900 7713 29968
rect 7265 29844 7275 29900
rect 7331 29844 7399 29900
rect 7455 29844 7523 29900
rect 7579 29844 7647 29900
rect 7703 29844 7713 29900
rect 7265 29776 7713 29844
rect 7265 29720 7275 29776
rect 7331 29720 7399 29776
rect 7455 29720 7523 29776
rect 7579 29720 7647 29776
rect 7703 29720 7713 29776
rect 7265 29652 7713 29720
rect 7265 29596 7275 29652
rect 7331 29596 7399 29652
rect 7455 29596 7523 29652
rect 7579 29596 7647 29652
rect 7703 29596 7713 29652
rect 7265 29528 7713 29596
rect 7265 29472 7275 29528
rect 7331 29472 7399 29528
rect 7455 29472 7523 29528
rect 7579 29472 7647 29528
rect 7703 29472 7713 29528
rect 7265 29404 7713 29472
rect 7265 29348 7275 29404
rect 7331 29348 7399 29404
rect 7455 29348 7523 29404
rect 7579 29348 7647 29404
rect 7703 29348 7713 29404
rect 7265 29280 7713 29348
rect 7265 29224 7275 29280
rect 7331 29224 7399 29280
rect 7455 29224 7523 29280
rect 7579 29224 7647 29280
rect 7703 29224 7713 29280
rect 7265 29156 7713 29224
rect 7265 29100 7275 29156
rect 7331 29100 7399 29156
rect 7455 29100 7523 29156
rect 7579 29100 7647 29156
rect 7703 29100 7713 29156
rect 7265 29032 7713 29100
rect 7265 28976 7275 29032
rect 7331 28976 7399 29032
rect 7455 28976 7523 29032
rect 7579 28976 7647 29032
rect 7703 28976 7713 29032
rect 7265 28908 7713 28976
rect 7265 28852 7275 28908
rect 7331 28852 7399 28908
rect 7455 28852 7523 28908
rect 7579 28852 7647 28908
rect 7703 28852 7713 28908
rect 7265 28842 7713 28852
rect 9927 30148 10127 30158
rect 9927 30092 9937 30148
rect 9993 30092 10061 30148
rect 10117 30092 10127 30148
rect 9927 30024 10127 30092
rect 9927 29968 9937 30024
rect 9993 29968 10061 30024
rect 10117 29968 10127 30024
rect 9927 29900 10127 29968
rect 9927 29844 9937 29900
rect 9993 29844 10061 29900
rect 10117 29844 10127 29900
rect 9927 29776 10127 29844
rect 9927 29720 9937 29776
rect 9993 29720 10061 29776
rect 10117 29720 10127 29776
rect 9927 29652 10127 29720
rect 9927 29596 9937 29652
rect 9993 29596 10061 29652
rect 10117 29596 10127 29652
rect 9927 29528 10127 29596
rect 9927 29472 9937 29528
rect 9993 29472 10061 29528
rect 10117 29472 10127 29528
rect 9927 29404 10127 29472
rect 9927 29348 9937 29404
rect 9993 29348 10061 29404
rect 10117 29348 10127 29404
rect 9927 29280 10127 29348
rect 9927 29224 9937 29280
rect 9993 29224 10061 29280
rect 10117 29224 10127 29280
rect 9927 29156 10127 29224
rect 9927 29100 9937 29156
rect 9993 29100 10061 29156
rect 10117 29100 10127 29156
rect 9927 29032 10127 29100
rect 9927 28976 9937 29032
rect 9993 28976 10061 29032
rect 10117 28976 10127 29032
rect 9927 28908 10127 28976
rect 9927 28852 9937 28908
rect 9993 28852 10061 28908
rect 10117 28852 10127 28908
rect 9927 28842 10127 28852
rect 12297 30148 12497 30158
rect 12297 30092 12307 30148
rect 12363 30092 12431 30148
rect 12487 30092 12497 30148
rect 12297 30024 12497 30092
rect 12297 29968 12307 30024
rect 12363 29968 12431 30024
rect 12487 29968 12497 30024
rect 12297 29900 12497 29968
rect 12297 29844 12307 29900
rect 12363 29844 12431 29900
rect 12487 29844 12497 29900
rect 12297 29776 12497 29844
rect 12297 29720 12307 29776
rect 12363 29720 12431 29776
rect 12487 29720 12497 29776
rect 12297 29652 12497 29720
rect 12297 29596 12307 29652
rect 12363 29596 12431 29652
rect 12487 29596 12497 29652
rect 12297 29528 12497 29596
rect 12297 29472 12307 29528
rect 12363 29472 12431 29528
rect 12487 29472 12497 29528
rect 12297 29404 12497 29472
rect 12297 29348 12307 29404
rect 12363 29348 12431 29404
rect 12487 29348 12497 29404
rect 12297 29280 12497 29348
rect 12297 29224 12307 29280
rect 12363 29224 12431 29280
rect 12487 29224 12497 29280
rect 12297 29156 12497 29224
rect 12297 29100 12307 29156
rect 12363 29100 12431 29156
rect 12487 29100 12497 29156
rect 12297 29032 12497 29100
rect 12297 28976 12307 29032
rect 12363 28976 12431 29032
rect 12487 28976 12497 29032
rect 12297 28908 12497 28976
rect 12297 28852 12307 28908
rect 12363 28852 12431 28908
rect 12487 28852 12497 28908
rect 12297 28842 12497 28852
rect 10 28576 86 28586
rect 10 27224 20 28576
rect 76 27224 86 28576
rect 14892 28576 14968 28586
rect 305 28548 2117 28558
rect 305 28492 315 28548
rect 371 28492 439 28548
rect 495 28492 563 28548
rect 619 28492 687 28548
rect 743 28492 811 28548
rect 867 28492 935 28548
rect 991 28492 1059 28548
rect 1115 28492 1183 28548
rect 1239 28492 1307 28548
rect 1363 28492 1431 28548
rect 1487 28492 1555 28548
rect 1611 28492 1679 28548
rect 1735 28492 1803 28548
rect 1859 28492 1927 28548
rect 1983 28492 2051 28548
rect 2107 28492 2117 28548
rect 305 28424 2117 28492
rect 305 28368 315 28424
rect 371 28368 439 28424
rect 495 28368 563 28424
rect 619 28368 687 28424
rect 743 28368 811 28424
rect 867 28368 935 28424
rect 991 28368 1059 28424
rect 1115 28368 1183 28424
rect 1239 28368 1307 28424
rect 1363 28368 1431 28424
rect 1487 28368 1555 28424
rect 1611 28368 1679 28424
rect 1735 28368 1803 28424
rect 1859 28368 1927 28424
rect 1983 28368 2051 28424
rect 2107 28368 2117 28424
rect 305 28300 2117 28368
rect 305 28244 315 28300
rect 371 28244 439 28300
rect 495 28244 563 28300
rect 619 28244 687 28300
rect 743 28244 811 28300
rect 867 28244 935 28300
rect 991 28244 1059 28300
rect 1115 28244 1183 28300
rect 1239 28244 1307 28300
rect 1363 28244 1431 28300
rect 1487 28244 1555 28300
rect 1611 28244 1679 28300
rect 1735 28244 1803 28300
rect 1859 28244 1927 28300
rect 1983 28244 2051 28300
rect 2107 28244 2117 28300
rect 305 28176 2117 28244
rect 305 28120 315 28176
rect 371 28120 439 28176
rect 495 28120 563 28176
rect 619 28120 687 28176
rect 743 28120 811 28176
rect 867 28120 935 28176
rect 991 28120 1059 28176
rect 1115 28120 1183 28176
rect 1239 28120 1307 28176
rect 1363 28120 1431 28176
rect 1487 28120 1555 28176
rect 1611 28120 1679 28176
rect 1735 28120 1803 28176
rect 1859 28120 1927 28176
rect 1983 28120 2051 28176
rect 2107 28120 2117 28176
rect 305 28052 2117 28120
rect 305 27996 315 28052
rect 371 27996 439 28052
rect 495 27996 563 28052
rect 619 27996 687 28052
rect 743 27996 811 28052
rect 867 27996 935 28052
rect 991 27996 1059 28052
rect 1115 27996 1183 28052
rect 1239 27996 1307 28052
rect 1363 27996 1431 28052
rect 1487 27996 1555 28052
rect 1611 27996 1679 28052
rect 1735 27996 1803 28052
rect 1859 27996 1927 28052
rect 1983 27996 2051 28052
rect 2107 27996 2117 28052
rect 305 27928 2117 27996
rect 305 27872 315 27928
rect 371 27872 439 27928
rect 495 27872 563 27928
rect 619 27872 687 27928
rect 743 27872 811 27928
rect 867 27872 935 27928
rect 991 27872 1059 27928
rect 1115 27872 1183 27928
rect 1239 27872 1307 27928
rect 1363 27872 1431 27928
rect 1487 27872 1555 27928
rect 1611 27872 1679 27928
rect 1735 27872 1803 27928
rect 1859 27872 1927 27928
rect 1983 27872 2051 27928
rect 2107 27872 2117 27928
rect 305 27804 2117 27872
rect 305 27748 315 27804
rect 371 27748 439 27804
rect 495 27748 563 27804
rect 619 27748 687 27804
rect 743 27748 811 27804
rect 867 27748 935 27804
rect 991 27748 1059 27804
rect 1115 27748 1183 27804
rect 1239 27748 1307 27804
rect 1363 27748 1431 27804
rect 1487 27748 1555 27804
rect 1611 27748 1679 27804
rect 1735 27748 1803 27804
rect 1859 27748 1927 27804
rect 1983 27748 2051 27804
rect 2107 27748 2117 27804
rect 305 27680 2117 27748
rect 305 27624 315 27680
rect 371 27624 439 27680
rect 495 27624 563 27680
rect 619 27624 687 27680
rect 743 27624 811 27680
rect 867 27624 935 27680
rect 991 27624 1059 27680
rect 1115 27624 1183 27680
rect 1239 27624 1307 27680
rect 1363 27624 1431 27680
rect 1487 27624 1555 27680
rect 1611 27624 1679 27680
rect 1735 27624 1803 27680
rect 1859 27624 1927 27680
rect 1983 27624 2051 27680
rect 2107 27624 2117 27680
rect 305 27556 2117 27624
rect 305 27500 315 27556
rect 371 27500 439 27556
rect 495 27500 563 27556
rect 619 27500 687 27556
rect 743 27500 811 27556
rect 867 27500 935 27556
rect 991 27500 1059 27556
rect 1115 27500 1183 27556
rect 1239 27500 1307 27556
rect 1363 27500 1431 27556
rect 1487 27500 1555 27556
rect 1611 27500 1679 27556
rect 1735 27500 1803 27556
rect 1859 27500 1927 27556
rect 1983 27500 2051 27556
rect 2107 27500 2117 27556
rect 305 27432 2117 27500
rect 305 27376 315 27432
rect 371 27376 439 27432
rect 495 27376 563 27432
rect 619 27376 687 27432
rect 743 27376 811 27432
rect 867 27376 935 27432
rect 991 27376 1059 27432
rect 1115 27376 1183 27432
rect 1239 27376 1307 27432
rect 1363 27376 1431 27432
rect 1487 27376 1555 27432
rect 1611 27376 1679 27432
rect 1735 27376 1803 27432
rect 1859 27376 1927 27432
rect 1983 27376 2051 27432
rect 2107 27376 2117 27432
rect 305 27308 2117 27376
rect 305 27252 315 27308
rect 371 27252 439 27308
rect 495 27252 563 27308
rect 619 27252 687 27308
rect 743 27252 811 27308
rect 867 27252 935 27308
rect 991 27252 1059 27308
rect 1115 27252 1183 27308
rect 1239 27252 1307 27308
rect 1363 27252 1431 27308
rect 1487 27252 1555 27308
rect 1611 27252 1679 27308
rect 1735 27252 1803 27308
rect 1859 27252 1927 27308
rect 1983 27252 2051 27308
rect 2107 27252 2117 27308
rect 305 27242 2117 27252
rect 2798 28548 4734 28558
rect 2798 28492 2808 28548
rect 2864 28492 2932 28548
rect 2988 28492 3056 28548
rect 3112 28492 3180 28548
rect 3236 28492 3304 28548
rect 3360 28492 3428 28548
rect 3484 28492 3552 28548
rect 3608 28492 3676 28548
rect 3732 28492 3800 28548
rect 3856 28492 3924 28548
rect 3980 28492 4048 28548
rect 4104 28492 4172 28548
rect 4228 28492 4296 28548
rect 4352 28492 4420 28548
rect 4476 28492 4544 28548
rect 4600 28492 4668 28548
rect 4724 28492 4734 28548
rect 2798 28424 4734 28492
rect 2798 28368 2808 28424
rect 2864 28368 2932 28424
rect 2988 28368 3056 28424
rect 3112 28368 3180 28424
rect 3236 28368 3304 28424
rect 3360 28368 3428 28424
rect 3484 28368 3552 28424
rect 3608 28368 3676 28424
rect 3732 28368 3800 28424
rect 3856 28368 3924 28424
rect 3980 28368 4048 28424
rect 4104 28368 4172 28424
rect 4228 28368 4296 28424
rect 4352 28368 4420 28424
rect 4476 28368 4544 28424
rect 4600 28368 4668 28424
rect 4724 28368 4734 28424
rect 2798 28300 4734 28368
rect 2798 28244 2808 28300
rect 2864 28244 2932 28300
rect 2988 28244 3056 28300
rect 3112 28244 3180 28300
rect 3236 28244 3304 28300
rect 3360 28244 3428 28300
rect 3484 28244 3552 28300
rect 3608 28244 3676 28300
rect 3732 28244 3800 28300
rect 3856 28244 3924 28300
rect 3980 28244 4048 28300
rect 4104 28244 4172 28300
rect 4228 28244 4296 28300
rect 4352 28244 4420 28300
rect 4476 28244 4544 28300
rect 4600 28244 4668 28300
rect 4724 28244 4734 28300
rect 2798 28176 4734 28244
rect 2798 28120 2808 28176
rect 2864 28120 2932 28176
rect 2988 28120 3056 28176
rect 3112 28120 3180 28176
rect 3236 28120 3304 28176
rect 3360 28120 3428 28176
rect 3484 28120 3552 28176
rect 3608 28120 3676 28176
rect 3732 28120 3800 28176
rect 3856 28120 3924 28176
rect 3980 28120 4048 28176
rect 4104 28120 4172 28176
rect 4228 28120 4296 28176
rect 4352 28120 4420 28176
rect 4476 28120 4544 28176
rect 4600 28120 4668 28176
rect 4724 28120 4734 28176
rect 2798 28052 4734 28120
rect 2798 27996 2808 28052
rect 2864 27996 2932 28052
rect 2988 27996 3056 28052
rect 3112 27996 3180 28052
rect 3236 27996 3304 28052
rect 3360 27996 3428 28052
rect 3484 27996 3552 28052
rect 3608 27996 3676 28052
rect 3732 27996 3800 28052
rect 3856 27996 3924 28052
rect 3980 27996 4048 28052
rect 4104 27996 4172 28052
rect 4228 27996 4296 28052
rect 4352 27996 4420 28052
rect 4476 27996 4544 28052
rect 4600 27996 4668 28052
rect 4724 27996 4734 28052
rect 2798 27928 4734 27996
rect 2798 27872 2808 27928
rect 2864 27872 2932 27928
rect 2988 27872 3056 27928
rect 3112 27872 3180 27928
rect 3236 27872 3304 27928
rect 3360 27872 3428 27928
rect 3484 27872 3552 27928
rect 3608 27872 3676 27928
rect 3732 27872 3800 27928
rect 3856 27872 3924 27928
rect 3980 27872 4048 27928
rect 4104 27872 4172 27928
rect 4228 27872 4296 27928
rect 4352 27872 4420 27928
rect 4476 27872 4544 27928
rect 4600 27872 4668 27928
rect 4724 27872 4734 27928
rect 2798 27804 4734 27872
rect 2798 27748 2808 27804
rect 2864 27748 2932 27804
rect 2988 27748 3056 27804
rect 3112 27748 3180 27804
rect 3236 27748 3304 27804
rect 3360 27748 3428 27804
rect 3484 27748 3552 27804
rect 3608 27748 3676 27804
rect 3732 27748 3800 27804
rect 3856 27748 3924 27804
rect 3980 27748 4048 27804
rect 4104 27748 4172 27804
rect 4228 27748 4296 27804
rect 4352 27748 4420 27804
rect 4476 27748 4544 27804
rect 4600 27748 4668 27804
rect 4724 27748 4734 27804
rect 2798 27680 4734 27748
rect 2798 27624 2808 27680
rect 2864 27624 2932 27680
rect 2988 27624 3056 27680
rect 3112 27624 3180 27680
rect 3236 27624 3304 27680
rect 3360 27624 3428 27680
rect 3484 27624 3552 27680
rect 3608 27624 3676 27680
rect 3732 27624 3800 27680
rect 3856 27624 3924 27680
rect 3980 27624 4048 27680
rect 4104 27624 4172 27680
rect 4228 27624 4296 27680
rect 4352 27624 4420 27680
rect 4476 27624 4544 27680
rect 4600 27624 4668 27680
rect 4724 27624 4734 27680
rect 2798 27556 4734 27624
rect 2798 27500 2808 27556
rect 2864 27500 2932 27556
rect 2988 27500 3056 27556
rect 3112 27500 3180 27556
rect 3236 27500 3304 27556
rect 3360 27500 3428 27556
rect 3484 27500 3552 27556
rect 3608 27500 3676 27556
rect 3732 27500 3800 27556
rect 3856 27500 3924 27556
rect 3980 27500 4048 27556
rect 4104 27500 4172 27556
rect 4228 27500 4296 27556
rect 4352 27500 4420 27556
rect 4476 27500 4544 27556
rect 4600 27500 4668 27556
rect 4724 27500 4734 27556
rect 2798 27432 4734 27500
rect 2798 27376 2808 27432
rect 2864 27376 2932 27432
rect 2988 27376 3056 27432
rect 3112 27376 3180 27432
rect 3236 27376 3304 27432
rect 3360 27376 3428 27432
rect 3484 27376 3552 27432
rect 3608 27376 3676 27432
rect 3732 27376 3800 27432
rect 3856 27376 3924 27432
rect 3980 27376 4048 27432
rect 4104 27376 4172 27432
rect 4228 27376 4296 27432
rect 4352 27376 4420 27432
rect 4476 27376 4544 27432
rect 4600 27376 4668 27432
rect 4724 27376 4734 27432
rect 2798 27308 4734 27376
rect 2798 27252 2808 27308
rect 2864 27252 2932 27308
rect 2988 27252 3056 27308
rect 3112 27252 3180 27308
rect 3236 27252 3304 27308
rect 3360 27252 3428 27308
rect 3484 27252 3552 27308
rect 3608 27252 3676 27308
rect 3732 27252 3800 27308
rect 3856 27252 3924 27308
rect 3980 27252 4048 27308
rect 4104 27252 4172 27308
rect 4228 27252 4296 27308
rect 4352 27252 4420 27308
rect 4476 27252 4544 27308
rect 4600 27252 4668 27308
rect 4724 27252 4734 27308
rect 2798 27242 4734 27252
rect 5168 28548 7104 28558
rect 5168 28492 5178 28548
rect 5234 28492 5302 28548
rect 5358 28492 5426 28548
rect 5482 28492 5550 28548
rect 5606 28492 5674 28548
rect 5730 28492 5798 28548
rect 5854 28492 5922 28548
rect 5978 28492 6046 28548
rect 6102 28492 6170 28548
rect 6226 28492 6294 28548
rect 6350 28492 6418 28548
rect 6474 28492 6542 28548
rect 6598 28492 6666 28548
rect 6722 28492 6790 28548
rect 6846 28492 6914 28548
rect 6970 28492 7038 28548
rect 7094 28492 7104 28548
rect 5168 28424 7104 28492
rect 5168 28368 5178 28424
rect 5234 28368 5302 28424
rect 5358 28368 5426 28424
rect 5482 28368 5550 28424
rect 5606 28368 5674 28424
rect 5730 28368 5798 28424
rect 5854 28368 5922 28424
rect 5978 28368 6046 28424
rect 6102 28368 6170 28424
rect 6226 28368 6294 28424
rect 6350 28368 6418 28424
rect 6474 28368 6542 28424
rect 6598 28368 6666 28424
rect 6722 28368 6790 28424
rect 6846 28368 6914 28424
rect 6970 28368 7038 28424
rect 7094 28368 7104 28424
rect 5168 28300 7104 28368
rect 5168 28244 5178 28300
rect 5234 28244 5302 28300
rect 5358 28244 5426 28300
rect 5482 28244 5550 28300
rect 5606 28244 5674 28300
rect 5730 28244 5798 28300
rect 5854 28244 5922 28300
rect 5978 28244 6046 28300
rect 6102 28244 6170 28300
rect 6226 28244 6294 28300
rect 6350 28244 6418 28300
rect 6474 28244 6542 28300
rect 6598 28244 6666 28300
rect 6722 28244 6790 28300
rect 6846 28244 6914 28300
rect 6970 28244 7038 28300
rect 7094 28244 7104 28300
rect 5168 28176 7104 28244
rect 5168 28120 5178 28176
rect 5234 28120 5302 28176
rect 5358 28120 5426 28176
rect 5482 28120 5550 28176
rect 5606 28120 5674 28176
rect 5730 28120 5798 28176
rect 5854 28120 5922 28176
rect 5978 28120 6046 28176
rect 6102 28120 6170 28176
rect 6226 28120 6294 28176
rect 6350 28120 6418 28176
rect 6474 28120 6542 28176
rect 6598 28120 6666 28176
rect 6722 28120 6790 28176
rect 6846 28120 6914 28176
rect 6970 28120 7038 28176
rect 7094 28120 7104 28176
rect 5168 28052 7104 28120
rect 5168 27996 5178 28052
rect 5234 27996 5302 28052
rect 5358 27996 5426 28052
rect 5482 27996 5550 28052
rect 5606 27996 5674 28052
rect 5730 27996 5798 28052
rect 5854 27996 5922 28052
rect 5978 27996 6046 28052
rect 6102 27996 6170 28052
rect 6226 27996 6294 28052
rect 6350 27996 6418 28052
rect 6474 27996 6542 28052
rect 6598 27996 6666 28052
rect 6722 27996 6790 28052
rect 6846 27996 6914 28052
rect 6970 27996 7038 28052
rect 7094 27996 7104 28052
rect 5168 27928 7104 27996
rect 5168 27872 5178 27928
rect 5234 27872 5302 27928
rect 5358 27872 5426 27928
rect 5482 27872 5550 27928
rect 5606 27872 5674 27928
rect 5730 27872 5798 27928
rect 5854 27872 5922 27928
rect 5978 27872 6046 27928
rect 6102 27872 6170 27928
rect 6226 27872 6294 27928
rect 6350 27872 6418 27928
rect 6474 27872 6542 27928
rect 6598 27872 6666 27928
rect 6722 27872 6790 27928
rect 6846 27872 6914 27928
rect 6970 27872 7038 27928
rect 7094 27872 7104 27928
rect 5168 27804 7104 27872
rect 5168 27748 5178 27804
rect 5234 27748 5302 27804
rect 5358 27748 5426 27804
rect 5482 27748 5550 27804
rect 5606 27748 5674 27804
rect 5730 27748 5798 27804
rect 5854 27748 5922 27804
rect 5978 27748 6046 27804
rect 6102 27748 6170 27804
rect 6226 27748 6294 27804
rect 6350 27748 6418 27804
rect 6474 27748 6542 27804
rect 6598 27748 6666 27804
rect 6722 27748 6790 27804
rect 6846 27748 6914 27804
rect 6970 27748 7038 27804
rect 7094 27748 7104 27804
rect 5168 27680 7104 27748
rect 5168 27624 5178 27680
rect 5234 27624 5302 27680
rect 5358 27624 5426 27680
rect 5482 27624 5550 27680
rect 5606 27624 5674 27680
rect 5730 27624 5798 27680
rect 5854 27624 5922 27680
rect 5978 27624 6046 27680
rect 6102 27624 6170 27680
rect 6226 27624 6294 27680
rect 6350 27624 6418 27680
rect 6474 27624 6542 27680
rect 6598 27624 6666 27680
rect 6722 27624 6790 27680
rect 6846 27624 6914 27680
rect 6970 27624 7038 27680
rect 7094 27624 7104 27680
rect 5168 27556 7104 27624
rect 5168 27500 5178 27556
rect 5234 27500 5302 27556
rect 5358 27500 5426 27556
rect 5482 27500 5550 27556
rect 5606 27500 5674 27556
rect 5730 27500 5798 27556
rect 5854 27500 5922 27556
rect 5978 27500 6046 27556
rect 6102 27500 6170 27556
rect 6226 27500 6294 27556
rect 6350 27500 6418 27556
rect 6474 27500 6542 27556
rect 6598 27500 6666 27556
rect 6722 27500 6790 27556
rect 6846 27500 6914 27556
rect 6970 27500 7038 27556
rect 7094 27500 7104 27556
rect 5168 27432 7104 27500
rect 5168 27376 5178 27432
rect 5234 27376 5302 27432
rect 5358 27376 5426 27432
rect 5482 27376 5550 27432
rect 5606 27376 5674 27432
rect 5730 27376 5798 27432
rect 5854 27376 5922 27432
rect 5978 27376 6046 27432
rect 6102 27376 6170 27432
rect 6226 27376 6294 27432
rect 6350 27376 6418 27432
rect 6474 27376 6542 27432
rect 6598 27376 6666 27432
rect 6722 27376 6790 27432
rect 6846 27376 6914 27432
rect 6970 27376 7038 27432
rect 7094 27376 7104 27432
rect 5168 27308 7104 27376
rect 5168 27252 5178 27308
rect 5234 27252 5302 27308
rect 5358 27252 5426 27308
rect 5482 27252 5550 27308
rect 5606 27252 5674 27308
rect 5730 27252 5798 27308
rect 5854 27252 5922 27308
rect 5978 27252 6046 27308
rect 6102 27252 6170 27308
rect 6226 27252 6294 27308
rect 6350 27252 6418 27308
rect 6474 27252 6542 27308
rect 6598 27252 6666 27308
rect 6722 27252 6790 27308
rect 6846 27252 6914 27308
rect 6970 27252 7038 27308
rect 7094 27252 7104 27308
rect 5168 27242 7104 27252
rect 7874 28548 9810 28558
rect 7874 28492 7884 28548
rect 7940 28492 8008 28548
rect 8064 28492 8132 28548
rect 8188 28492 8256 28548
rect 8312 28492 8380 28548
rect 8436 28492 8504 28548
rect 8560 28492 8628 28548
rect 8684 28492 8752 28548
rect 8808 28492 8876 28548
rect 8932 28492 9000 28548
rect 9056 28492 9124 28548
rect 9180 28492 9248 28548
rect 9304 28492 9372 28548
rect 9428 28492 9496 28548
rect 9552 28492 9620 28548
rect 9676 28492 9744 28548
rect 9800 28492 9810 28548
rect 7874 28424 9810 28492
rect 7874 28368 7884 28424
rect 7940 28368 8008 28424
rect 8064 28368 8132 28424
rect 8188 28368 8256 28424
rect 8312 28368 8380 28424
rect 8436 28368 8504 28424
rect 8560 28368 8628 28424
rect 8684 28368 8752 28424
rect 8808 28368 8876 28424
rect 8932 28368 9000 28424
rect 9056 28368 9124 28424
rect 9180 28368 9248 28424
rect 9304 28368 9372 28424
rect 9428 28368 9496 28424
rect 9552 28368 9620 28424
rect 9676 28368 9744 28424
rect 9800 28368 9810 28424
rect 7874 28300 9810 28368
rect 7874 28244 7884 28300
rect 7940 28244 8008 28300
rect 8064 28244 8132 28300
rect 8188 28244 8256 28300
rect 8312 28244 8380 28300
rect 8436 28244 8504 28300
rect 8560 28244 8628 28300
rect 8684 28244 8752 28300
rect 8808 28244 8876 28300
rect 8932 28244 9000 28300
rect 9056 28244 9124 28300
rect 9180 28244 9248 28300
rect 9304 28244 9372 28300
rect 9428 28244 9496 28300
rect 9552 28244 9620 28300
rect 9676 28244 9744 28300
rect 9800 28244 9810 28300
rect 7874 28176 9810 28244
rect 7874 28120 7884 28176
rect 7940 28120 8008 28176
rect 8064 28120 8132 28176
rect 8188 28120 8256 28176
rect 8312 28120 8380 28176
rect 8436 28120 8504 28176
rect 8560 28120 8628 28176
rect 8684 28120 8752 28176
rect 8808 28120 8876 28176
rect 8932 28120 9000 28176
rect 9056 28120 9124 28176
rect 9180 28120 9248 28176
rect 9304 28120 9372 28176
rect 9428 28120 9496 28176
rect 9552 28120 9620 28176
rect 9676 28120 9744 28176
rect 9800 28120 9810 28176
rect 7874 28052 9810 28120
rect 7874 27996 7884 28052
rect 7940 27996 8008 28052
rect 8064 27996 8132 28052
rect 8188 27996 8256 28052
rect 8312 27996 8380 28052
rect 8436 27996 8504 28052
rect 8560 27996 8628 28052
rect 8684 27996 8752 28052
rect 8808 27996 8876 28052
rect 8932 27996 9000 28052
rect 9056 27996 9124 28052
rect 9180 27996 9248 28052
rect 9304 27996 9372 28052
rect 9428 27996 9496 28052
rect 9552 27996 9620 28052
rect 9676 27996 9744 28052
rect 9800 27996 9810 28052
rect 7874 27928 9810 27996
rect 7874 27872 7884 27928
rect 7940 27872 8008 27928
rect 8064 27872 8132 27928
rect 8188 27872 8256 27928
rect 8312 27872 8380 27928
rect 8436 27872 8504 27928
rect 8560 27872 8628 27928
rect 8684 27872 8752 27928
rect 8808 27872 8876 27928
rect 8932 27872 9000 27928
rect 9056 27872 9124 27928
rect 9180 27872 9248 27928
rect 9304 27872 9372 27928
rect 9428 27872 9496 27928
rect 9552 27872 9620 27928
rect 9676 27872 9744 27928
rect 9800 27872 9810 27928
rect 7874 27804 9810 27872
rect 7874 27748 7884 27804
rect 7940 27748 8008 27804
rect 8064 27748 8132 27804
rect 8188 27748 8256 27804
rect 8312 27748 8380 27804
rect 8436 27748 8504 27804
rect 8560 27748 8628 27804
rect 8684 27748 8752 27804
rect 8808 27748 8876 27804
rect 8932 27748 9000 27804
rect 9056 27748 9124 27804
rect 9180 27748 9248 27804
rect 9304 27748 9372 27804
rect 9428 27748 9496 27804
rect 9552 27748 9620 27804
rect 9676 27748 9744 27804
rect 9800 27748 9810 27804
rect 7874 27680 9810 27748
rect 7874 27624 7884 27680
rect 7940 27624 8008 27680
rect 8064 27624 8132 27680
rect 8188 27624 8256 27680
rect 8312 27624 8380 27680
rect 8436 27624 8504 27680
rect 8560 27624 8628 27680
rect 8684 27624 8752 27680
rect 8808 27624 8876 27680
rect 8932 27624 9000 27680
rect 9056 27624 9124 27680
rect 9180 27624 9248 27680
rect 9304 27624 9372 27680
rect 9428 27624 9496 27680
rect 9552 27624 9620 27680
rect 9676 27624 9744 27680
rect 9800 27624 9810 27680
rect 7874 27556 9810 27624
rect 7874 27500 7884 27556
rect 7940 27500 8008 27556
rect 8064 27500 8132 27556
rect 8188 27500 8256 27556
rect 8312 27500 8380 27556
rect 8436 27500 8504 27556
rect 8560 27500 8628 27556
rect 8684 27500 8752 27556
rect 8808 27500 8876 27556
rect 8932 27500 9000 27556
rect 9056 27500 9124 27556
rect 9180 27500 9248 27556
rect 9304 27500 9372 27556
rect 9428 27500 9496 27556
rect 9552 27500 9620 27556
rect 9676 27500 9744 27556
rect 9800 27500 9810 27556
rect 7874 27432 9810 27500
rect 7874 27376 7884 27432
rect 7940 27376 8008 27432
rect 8064 27376 8132 27432
rect 8188 27376 8256 27432
rect 8312 27376 8380 27432
rect 8436 27376 8504 27432
rect 8560 27376 8628 27432
rect 8684 27376 8752 27432
rect 8808 27376 8876 27432
rect 8932 27376 9000 27432
rect 9056 27376 9124 27432
rect 9180 27376 9248 27432
rect 9304 27376 9372 27432
rect 9428 27376 9496 27432
rect 9552 27376 9620 27432
rect 9676 27376 9744 27432
rect 9800 27376 9810 27432
rect 7874 27308 9810 27376
rect 7874 27252 7884 27308
rect 7940 27252 8008 27308
rect 8064 27252 8132 27308
rect 8188 27252 8256 27308
rect 8312 27252 8380 27308
rect 8436 27252 8504 27308
rect 8560 27252 8628 27308
rect 8684 27252 8752 27308
rect 8808 27252 8876 27308
rect 8932 27252 9000 27308
rect 9056 27252 9124 27308
rect 9180 27252 9248 27308
rect 9304 27252 9372 27308
rect 9428 27252 9496 27308
rect 9552 27252 9620 27308
rect 9676 27252 9744 27308
rect 9800 27252 9810 27308
rect 7874 27242 9810 27252
rect 10244 28548 12180 28558
rect 10244 28492 10254 28548
rect 10310 28492 10378 28548
rect 10434 28492 10502 28548
rect 10558 28492 10626 28548
rect 10682 28492 10750 28548
rect 10806 28492 10874 28548
rect 10930 28492 10998 28548
rect 11054 28492 11122 28548
rect 11178 28492 11246 28548
rect 11302 28492 11370 28548
rect 11426 28492 11494 28548
rect 11550 28492 11618 28548
rect 11674 28492 11742 28548
rect 11798 28492 11866 28548
rect 11922 28492 11990 28548
rect 12046 28492 12114 28548
rect 12170 28492 12180 28548
rect 10244 28424 12180 28492
rect 10244 28368 10254 28424
rect 10310 28368 10378 28424
rect 10434 28368 10502 28424
rect 10558 28368 10626 28424
rect 10682 28368 10750 28424
rect 10806 28368 10874 28424
rect 10930 28368 10998 28424
rect 11054 28368 11122 28424
rect 11178 28368 11246 28424
rect 11302 28368 11370 28424
rect 11426 28368 11494 28424
rect 11550 28368 11618 28424
rect 11674 28368 11742 28424
rect 11798 28368 11866 28424
rect 11922 28368 11990 28424
rect 12046 28368 12114 28424
rect 12170 28368 12180 28424
rect 10244 28300 12180 28368
rect 10244 28244 10254 28300
rect 10310 28244 10378 28300
rect 10434 28244 10502 28300
rect 10558 28244 10626 28300
rect 10682 28244 10750 28300
rect 10806 28244 10874 28300
rect 10930 28244 10998 28300
rect 11054 28244 11122 28300
rect 11178 28244 11246 28300
rect 11302 28244 11370 28300
rect 11426 28244 11494 28300
rect 11550 28244 11618 28300
rect 11674 28244 11742 28300
rect 11798 28244 11866 28300
rect 11922 28244 11990 28300
rect 12046 28244 12114 28300
rect 12170 28244 12180 28300
rect 10244 28176 12180 28244
rect 10244 28120 10254 28176
rect 10310 28120 10378 28176
rect 10434 28120 10502 28176
rect 10558 28120 10626 28176
rect 10682 28120 10750 28176
rect 10806 28120 10874 28176
rect 10930 28120 10998 28176
rect 11054 28120 11122 28176
rect 11178 28120 11246 28176
rect 11302 28120 11370 28176
rect 11426 28120 11494 28176
rect 11550 28120 11618 28176
rect 11674 28120 11742 28176
rect 11798 28120 11866 28176
rect 11922 28120 11990 28176
rect 12046 28120 12114 28176
rect 12170 28120 12180 28176
rect 10244 28052 12180 28120
rect 10244 27996 10254 28052
rect 10310 27996 10378 28052
rect 10434 27996 10502 28052
rect 10558 27996 10626 28052
rect 10682 27996 10750 28052
rect 10806 27996 10874 28052
rect 10930 27996 10998 28052
rect 11054 27996 11122 28052
rect 11178 27996 11246 28052
rect 11302 27996 11370 28052
rect 11426 27996 11494 28052
rect 11550 27996 11618 28052
rect 11674 27996 11742 28052
rect 11798 27996 11866 28052
rect 11922 27996 11990 28052
rect 12046 27996 12114 28052
rect 12170 27996 12180 28052
rect 10244 27928 12180 27996
rect 10244 27872 10254 27928
rect 10310 27872 10378 27928
rect 10434 27872 10502 27928
rect 10558 27872 10626 27928
rect 10682 27872 10750 27928
rect 10806 27872 10874 27928
rect 10930 27872 10998 27928
rect 11054 27872 11122 27928
rect 11178 27872 11246 27928
rect 11302 27872 11370 27928
rect 11426 27872 11494 27928
rect 11550 27872 11618 27928
rect 11674 27872 11742 27928
rect 11798 27872 11866 27928
rect 11922 27872 11990 27928
rect 12046 27872 12114 27928
rect 12170 27872 12180 27928
rect 10244 27804 12180 27872
rect 10244 27748 10254 27804
rect 10310 27748 10378 27804
rect 10434 27748 10502 27804
rect 10558 27748 10626 27804
rect 10682 27748 10750 27804
rect 10806 27748 10874 27804
rect 10930 27748 10998 27804
rect 11054 27748 11122 27804
rect 11178 27748 11246 27804
rect 11302 27748 11370 27804
rect 11426 27748 11494 27804
rect 11550 27748 11618 27804
rect 11674 27748 11742 27804
rect 11798 27748 11866 27804
rect 11922 27748 11990 27804
rect 12046 27748 12114 27804
rect 12170 27748 12180 27804
rect 10244 27680 12180 27748
rect 10244 27624 10254 27680
rect 10310 27624 10378 27680
rect 10434 27624 10502 27680
rect 10558 27624 10626 27680
rect 10682 27624 10750 27680
rect 10806 27624 10874 27680
rect 10930 27624 10998 27680
rect 11054 27624 11122 27680
rect 11178 27624 11246 27680
rect 11302 27624 11370 27680
rect 11426 27624 11494 27680
rect 11550 27624 11618 27680
rect 11674 27624 11742 27680
rect 11798 27624 11866 27680
rect 11922 27624 11990 27680
rect 12046 27624 12114 27680
rect 12170 27624 12180 27680
rect 10244 27556 12180 27624
rect 10244 27500 10254 27556
rect 10310 27500 10378 27556
rect 10434 27500 10502 27556
rect 10558 27500 10626 27556
rect 10682 27500 10750 27556
rect 10806 27500 10874 27556
rect 10930 27500 10998 27556
rect 11054 27500 11122 27556
rect 11178 27500 11246 27556
rect 11302 27500 11370 27556
rect 11426 27500 11494 27556
rect 11550 27500 11618 27556
rect 11674 27500 11742 27556
rect 11798 27500 11866 27556
rect 11922 27500 11990 27556
rect 12046 27500 12114 27556
rect 12170 27500 12180 27556
rect 10244 27432 12180 27500
rect 10244 27376 10254 27432
rect 10310 27376 10378 27432
rect 10434 27376 10502 27432
rect 10558 27376 10626 27432
rect 10682 27376 10750 27432
rect 10806 27376 10874 27432
rect 10930 27376 10998 27432
rect 11054 27376 11122 27432
rect 11178 27376 11246 27432
rect 11302 27376 11370 27432
rect 11426 27376 11494 27432
rect 11550 27376 11618 27432
rect 11674 27376 11742 27432
rect 11798 27376 11866 27432
rect 11922 27376 11990 27432
rect 12046 27376 12114 27432
rect 12170 27376 12180 27432
rect 10244 27308 12180 27376
rect 10244 27252 10254 27308
rect 10310 27252 10378 27308
rect 10434 27252 10502 27308
rect 10558 27252 10626 27308
rect 10682 27252 10750 27308
rect 10806 27252 10874 27308
rect 10930 27252 10998 27308
rect 11054 27252 11122 27308
rect 11178 27252 11246 27308
rect 11302 27252 11370 27308
rect 11426 27252 11494 27308
rect 11550 27252 11618 27308
rect 11674 27252 11742 27308
rect 11798 27252 11866 27308
rect 11922 27252 11990 27308
rect 12046 27252 12114 27308
rect 12170 27252 12180 27308
rect 10244 27242 12180 27252
rect 12861 28548 14673 28558
rect 12861 28492 12871 28548
rect 12927 28492 12995 28548
rect 13051 28492 13119 28548
rect 13175 28492 13243 28548
rect 13299 28492 13367 28548
rect 13423 28492 13491 28548
rect 13547 28492 13615 28548
rect 13671 28492 13739 28548
rect 13795 28492 13863 28548
rect 13919 28492 13987 28548
rect 14043 28492 14111 28548
rect 14167 28492 14235 28548
rect 14291 28492 14359 28548
rect 14415 28492 14483 28548
rect 14539 28492 14607 28548
rect 14663 28492 14673 28548
rect 12861 28424 14673 28492
rect 12861 28368 12871 28424
rect 12927 28368 12995 28424
rect 13051 28368 13119 28424
rect 13175 28368 13243 28424
rect 13299 28368 13367 28424
rect 13423 28368 13491 28424
rect 13547 28368 13615 28424
rect 13671 28368 13739 28424
rect 13795 28368 13863 28424
rect 13919 28368 13987 28424
rect 14043 28368 14111 28424
rect 14167 28368 14235 28424
rect 14291 28368 14359 28424
rect 14415 28368 14483 28424
rect 14539 28368 14607 28424
rect 14663 28368 14673 28424
rect 12861 28300 14673 28368
rect 12861 28244 12871 28300
rect 12927 28244 12995 28300
rect 13051 28244 13119 28300
rect 13175 28244 13243 28300
rect 13299 28244 13367 28300
rect 13423 28244 13491 28300
rect 13547 28244 13615 28300
rect 13671 28244 13739 28300
rect 13795 28244 13863 28300
rect 13919 28244 13987 28300
rect 14043 28244 14111 28300
rect 14167 28244 14235 28300
rect 14291 28244 14359 28300
rect 14415 28244 14483 28300
rect 14539 28244 14607 28300
rect 14663 28244 14673 28300
rect 12861 28176 14673 28244
rect 12861 28120 12871 28176
rect 12927 28120 12995 28176
rect 13051 28120 13119 28176
rect 13175 28120 13243 28176
rect 13299 28120 13367 28176
rect 13423 28120 13491 28176
rect 13547 28120 13615 28176
rect 13671 28120 13739 28176
rect 13795 28120 13863 28176
rect 13919 28120 13987 28176
rect 14043 28120 14111 28176
rect 14167 28120 14235 28176
rect 14291 28120 14359 28176
rect 14415 28120 14483 28176
rect 14539 28120 14607 28176
rect 14663 28120 14673 28176
rect 12861 28052 14673 28120
rect 12861 27996 12871 28052
rect 12927 27996 12995 28052
rect 13051 27996 13119 28052
rect 13175 27996 13243 28052
rect 13299 27996 13367 28052
rect 13423 27996 13491 28052
rect 13547 27996 13615 28052
rect 13671 27996 13739 28052
rect 13795 27996 13863 28052
rect 13919 27996 13987 28052
rect 14043 27996 14111 28052
rect 14167 27996 14235 28052
rect 14291 27996 14359 28052
rect 14415 27996 14483 28052
rect 14539 27996 14607 28052
rect 14663 27996 14673 28052
rect 12861 27928 14673 27996
rect 12861 27872 12871 27928
rect 12927 27872 12995 27928
rect 13051 27872 13119 27928
rect 13175 27872 13243 27928
rect 13299 27872 13367 27928
rect 13423 27872 13491 27928
rect 13547 27872 13615 27928
rect 13671 27872 13739 27928
rect 13795 27872 13863 27928
rect 13919 27872 13987 27928
rect 14043 27872 14111 27928
rect 14167 27872 14235 27928
rect 14291 27872 14359 27928
rect 14415 27872 14483 27928
rect 14539 27872 14607 27928
rect 14663 27872 14673 27928
rect 12861 27804 14673 27872
rect 12861 27748 12871 27804
rect 12927 27748 12995 27804
rect 13051 27748 13119 27804
rect 13175 27748 13243 27804
rect 13299 27748 13367 27804
rect 13423 27748 13491 27804
rect 13547 27748 13615 27804
rect 13671 27748 13739 27804
rect 13795 27748 13863 27804
rect 13919 27748 13987 27804
rect 14043 27748 14111 27804
rect 14167 27748 14235 27804
rect 14291 27748 14359 27804
rect 14415 27748 14483 27804
rect 14539 27748 14607 27804
rect 14663 27748 14673 27804
rect 12861 27680 14673 27748
rect 12861 27624 12871 27680
rect 12927 27624 12995 27680
rect 13051 27624 13119 27680
rect 13175 27624 13243 27680
rect 13299 27624 13367 27680
rect 13423 27624 13491 27680
rect 13547 27624 13615 27680
rect 13671 27624 13739 27680
rect 13795 27624 13863 27680
rect 13919 27624 13987 27680
rect 14043 27624 14111 27680
rect 14167 27624 14235 27680
rect 14291 27624 14359 27680
rect 14415 27624 14483 27680
rect 14539 27624 14607 27680
rect 14663 27624 14673 27680
rect 12861 27556 14673 27624
rect 12861 27500 12871 27556
rect 12927 27500 12995 27556
rect 13051 27500 13119 27556
rect 13175 27500 13243 27556
rect 13299 27500 13367 27556
rect 13423 27500 13491 27556
rect 13547 27500 13615 27556
rect 13671 27500 13739 27556
rect 13795 27500 13863 27556
rect 13919 27500 13987 27556
rect 14043 27500 14111 27556
rect 14167 27500 14235 27556
rect 14291 27500 14359 27556
rect 14415 27500 14483 27556
rect 14539 27500 14607 27556
rect 14663 27500 14673 27556
rect 12861 27432 14673 27500
rect 12861 27376 12871 27432
rect 12927 27376 12995 27432
rect 13051 27376 13119 27432
rect 13175 27376 13243 27432
rect 13299 27376 13367 27432
rect 13423 27376 13491 27432
rect 13547 27376 13615 27432
rect 13671 27376 13739 27432
rect 13795 27376 13863 27432
rect 13919 27376 13987 27432
rect 14043 27376 14111 27432
rect 14167 27376 14235 27432
rect 14291 27376 14359 27432
rect 14415 27376 14483 27432
rect 14539 27376 14607 27432
rect 14663 27376 14673 27432
rect 12861 27308 14673 27376
rect 12861 27252 12871 27308
rect 12927 27252 12995 27308
rect 13051 27252 13119 27308
rect 13175 27252 13243 27308
rect 13299 27252 13367 27308
rect 13423 27252 13491 27308
rect 13547 27252 13615 27308
rect 13671 27252 13739 27308
rect 13795 27252 13863 27308
rect 13919 27252 13987 27308
rect 14043 27252 14111 27308
rect 14167 27252 14235 27308
rect 14291 27252 14359 27308
rect 14415 27252 14483 27308
rect 14539 27252 14607 27308
rect 14663 27252 14673 27308
rect 12861 27242 14673 27252
rect 10 27214 86 27224
rect 14892 27224 14902 28576
rect 14958 27224 14968 28576
rect 14892 27214 14968 27224
rect 2481 26954 2681 26964
rect 2481 26898 2491 26954
rect 2547 26898 2615 26954
rect 2671 26898 2681 26954
rect 2481 26830 2681 26898
rect 2481 26774 2491 26830
rect 2547 26774 2615 26830
rect 2671 26774 2681 26830
rect 2481 26706 2681 26774
rect 2481 26650 2491 26706
rect 2547 26650 2615 26706
rect 2671 26650 2681 26706
rect 2481 26582 2681 26650
rect 2481 26526 2491 26582
rect 2547 26526 2615 26582
rect 2671 26526 2681 26582
rect 2481 26458 2681 26526
rect 2481 26402 2491 26458
rect 2547 26402 2615 26458
rect 2671 26402 2681 26458
rect 2481 26334 2681 26402
rect 2481 26278 2491 26334
rect 2547 26278 2615 26334
rect 2671 26278 2681 26334
rect 2481 26210 2681 26278
rect 2481 26154 2491 26210
rect 2547 26154 2615 26210
rect 2671 26154 2681 26210
rect 2481 26086 2681 26154
rect 2481 26030 2491 26086
rect 2547 26030 2615 26086
rect 2671 26030 2681 26086
rect 2481 25962 2681 26030
rect 2481 25906 2491 25962
rect 2547 25906 2615 25962
rect 2671 25906 2681 25962
rect 2481 25838 2681 25906
rect 2481 25782 2491 25838
rect 2547 25782 2615 25838
rect 2671 25782 2681 25838
rect 2481 25714 2681 25782
rect 2481 25658 2491 25714
rect 2547 25658 2615 25714
rect 2671 25658 2681 25714
rect 2481 25590 2681 25658
rect 2481 25534 2491 25590
rect 2547 25534 2615 25590
rect 2671 25534 2681 25590
rect 2481 25466 2681 25534
rect 2481 25410 2491 25466
rect 2547 25410 2615 25466
rect 2671 25410 2681 25466
rect 2481 25342 2681 25410
rect 2481 25286 2491 25342
rect 2547 25286 2615 25342
rect 2671 25286 2681 25342
rect 2481 25218 2681 25286
rect 2481 25162 2491 25218
rect 2547 25162 2615 25218
rect 2671 25162 2681 25218
rect 2481 25094 2681 25162
rect 2481 25038 2491 25094
rect 2547 25038 2615 25094
rect 2671 25038 2681 25094
rect 2481 24970 2681 25038
rect 2481 24914 2491 24970
rect 2547 24914 2615 24970
rect 2671 24914 2681 24970
rect 2481 24846 2681 24914
rect 2481 24790 2491 24846
rect 2547 24790 2615 24846
rect 2671 24790 2681 24846
rect 2481 24722 2681 24790
rect 2481 24666 2491 24722
rect 2547 24666 2615 24722
rect 2671 24666 2681 24722
rect 2481 24598 2681 24666
rect 2481 24542 2491 24598
rect 2547 24542 2615 24598
rect 2671 24542 2681 24598
rect 2481 24474 2681 24542
rect 2481 24418 2491 24474
rect 2547 24418 2615 24474
rect 2671 24418 2681 24474
rect 2481 24350 2681 24418
rect 2481 24294 2491 24350
rect 2547 24294 2615 24350
rect 2671 24294 2681 24350
rect 2481 24226 2681 24294
rect 2481 24170 2491 24226
rect 2547 24170 2615 24226
rect 2671 24170 2681 24226
rect 2481 24102 2681 24170
rect 2481 24046 2491 24102
rect 2547 24046 2615 24102
rect 2671 24046 2681 24102
rect 2481 24036 2681 24046
rect 4851 26954 5051 26964
rect 4851 26898 4861 26954
rect 4917 26898 4985 26954
rect 5041 26898 5051 26954
rect 4851 26830 5051 26898
rect 4851 26774 4861 26830
rect 4917 26774 4985 26830
rect 5041 26774 5051 26830
rect 4851 26706 5051 26774
rect 4851 26650 4861 26706
rect 4917 26650 4985 26706
rect 5041 26650 5051 26706
rect 4851 26582 5051 26650
rect 4851 26526 4861 26582
rect 4917 26526 4985 26582
rect 5041 26526 5051 26582
rect 4851 26458 5051 26526
rect 4851 26402 4861 26458
rect 4917 26402 4985 26458
rect 5041 26402 5051 26458
rect 4851 26334 5051 26402
rect 4851 26278 4861 26334
rect 4917 26278 4985 26334
rect 5041 26278 5051 26334
rect 4851 26210 5051 26278
rect 4851 26154 4861 26210
rect 4917 26154 4985 26210
rect 5041 26154 5051 26210
rect 4851 26086 5051 26154
rect 4851 26030 4861 26086
rect 4917 26030 4985 26086
rect 5041 26030 5051 26086
rect 4851 25962 5051 26030
rect 4851 25906 4861 25962
rect 4917 25906 4985 25962
rect 5041 25906 5051 25962
rect 4851 25838 5051 25906
rect 4851 25782 4861 25838
rect 4917 25782 4985 25838
rect 5041 25782 5051 25838
rect 4851 25714 5051 25782
rect 4851 25658 4861 25714
rect 4917 25658 4985 25714
rect 5041 25658 5051 25714
rect 4851 25590 5051 25658
rect 4851 25534 4861 25590
rect 4917 25534 4985 25590
rect 5041 25534 5051 25590
rect 4851 25466 5051 25534
rect 4851 25410 4861 25466
rect 4917 25410 4985 25466
rect 5041 25410 5051 25466
rect 4851 25342 5051 25410
rect 4851 25286 4861 25342
rect 4917 25286 4985 25342
rect 5041 25286 5051 25342
rect 4851 25218 5051 25286
rect 4851 25162 4861 25218
rect 4917 25162 4985 25218
rect 5041 25162 5051 25218
rect 4851 25094 5051 25162
rect 4851 25038 4861 25094
rect 4917 25038 4985 25094
rect 5041 25038 5051 25094
rect 4851 24970 5051 25038
rect 4851 24914 4861 24970
rect 4917 24914 4985 24970
rect 5041 24914 5051 24970
rect 4851 24846 5051 24914
rect 4851 24790 4861 24846
rect 4917 24790 4985 24846
rect 5041 24790 5051 24846
rect 4851 24722 5051 24790
rect 4851 24666 4861 24722
rect 4917 24666 4985 24722
rect 5041 24666 5051 24722
rect 4851 24598 5051 24666
rect 4851 24542 4861 24598
rect 4917 24542 4985 24598
rect 5041 24542 5051 24598
rect 4851 24474 5051 24542
rect 4851 24418 4861 24474
rect 4917 24418 4985 24474
rect 5041 24418 5051 24474
rect 4851 24350 5051 24418
rect 4851 24294 4861 24350
rect 4917 24294 4985 24350
rect 5041 24294 5051 24350
rect 4851 24226 5051 24294
rect 4851 24170 4861 24226
rect 4917 24170 4985 24226
rect 5041 24170 5051 24226
rect 4851 24102 5051 24170
rect 4851 24046 4861 24102
rect 4917 24046 4985 24102
rect 5041 24046 5051 24102
rect 4851 24036 5051 24046
rect 7265 26954 7713 26964
rect 7265 26898 7275 26954
rect 7331 26898 7399 26954
rect 7455 26898 7523 26954
rect 7579 26898 7647 26954
rect 7703 26898 7713 26954
rect 7265 26830 7713 26898
rect 7265 26774 7275 26830
rect 7331 26774 7399 26830
rect 7455 26774 7523 26830
rect 7579 26774 7647 26830
rect 7703 26774 7713 26830
rect 7265 26706 7713 26774
rect 7265 26650 7275 26706
rect 7331 26650 7399 26706
rect 7455 26650 7523 26706
rect 7579 26650 7647 26706
rect 7703 26650 7713 26706
rect 7265 26582 7713 26650
rect 7265 26526 7275 26582
rect 7331 26526 7399 26582
rect 7455 26526 7523 26582
rect 7579 26526 7647 26582
rect 7703 26526 7713 26582
rect 7265 26458 7713 26526
rect 7265 26402 7275 26458
rect 7331 26402 7399 26458
rect 7455 26402 7523 26458
rect 7579 26402 7647 26458
rect 7703 26402 7713 26458
rect 7265 26334 7713 26402
rect 7265 26278 7275 26334
rect 7331 26278 7399 26334
rect 7455 26278 7523 26334
rect 7579 26278 7647 26334
rect 7703 26278 7713 26334
rect 7265 26210 7713 26278
rect 7265 26154 7275 26210
rect 7331 26154 7399 26210
rect 7455 26154 7523 26210
rect 7579 26154 7647 26210
rect 7703 26154 7713 26210
rect 7265 26086 7713 26154
rect 7265 26030 7275 26086
rect 7331 26030 7399 26086
rect 7455 26030 7523 26086
rect 7579 26030 7647 26086
rect 7703 26030 7713 26086
rect 7265 25962 7713 26030
rect 7265 25906 7275 25962
rect 7331 25906 7399 25962
rect 7455 25906 7523 25962
rect 7579 25906 7647 25962
rect 7703 25906 7713 25962
rect 7265 25838 7713 25906
rect 7265 25782 7275 25838
rect 7331 25782 7399 25838
rect 7455 25782 7523 25838
rect 7579 25782 7647 25838
rect 7703 25782 7713 25838
rect 7265 25714 7713 25782
rect 7265 25658 7275 25714
rect 7331 25658 7399 25714
rect 7455 25658 7523 25714
rect 7579 25658 7647 25714
rect 7703 25658 7713 25714
rect 7265 25590 7713 25658
rect 7265 25534 7275 25590
rect 7331 25534 7399 25590
rect 7455 25534 7523 25590
rect 7579 25534 7647 25590
rect 7703 25534 7713 25590
rect 7265 25466 7713 25534
rect 7265 25410 7275 25466
rect 7331 25410 7399 25466
rect 7455 25410 7523 25466
rect 7579 25410 7647 25466
rect 7703 25410 7713 25466
rect 7265 25342 7713 25410
rect 7265 25286 7275 25342
rect 7331 25286 7399 25342
rect 7455 25286 7523 25342
rect 7579 25286 7647 25342
rect 7703 25286 7713 25342
rect 7265 25218 7713 25286
rect 7265 25162 7275 25218
rect 7331 25162 7399 25218
rect 7455 25162 7523 25218
rect 7579 25162 7647 25218
rect 7703 25162 7713 25218
rect 7265 25094 7713 25162
rect 7265 25038 7275 25094
rect 7331 25038 7399 25094
rect 7455 25038 7523 25094
rect 7579 25038 7647 25094
rect 7703 25038 7713 25094
rect 7265 24970 7713 25038
rect 7265 24914 7275 24970
rect 7331 24914 7399 24970
rect 7455 24914 7523 24970
rect 7579 24914 7647 24970
rect 7703 24914 7713 24970
rect 7265 24846 7713 24914
rect 7265 24790 7275 24846
rect 7331 24790 7399 24846
rect 7455 24790 7523 24846
rect 7579 24790 7647 24846
rect 7703 24790 7713 24846
rect 7265 24722 7713 24790
rect 7265 24666 7275 24722
rect 7331 24666 7399 24722
rect 7455 24666 7523 24722
rect 7579 24666 7647 24722
rect 7703 24666 7713 24722
rect 7265 24598 7713 24666
rect 7265 24542 7275 24598
rect 7331 24542 7399 24598
rect 7455 24542 7523 24598
rect 7579 24542 7647 24598
rect 7703 24542 7713 24598
rect 7265 24474 7713 24542
rect 7265 24418 7275 24474
rect 7331 24418 7399 24474
rect 7455 24418 7523 24474
rect 7579 24418 7647 24474
rect 7703 24418 7713 24474
rect 7265 24350 7713 24418
rect 7265 24294 7275 24350
rect 7331 24294 7399 24350
rect 7455 24294 7523 24350
rect 7579 24294 7647 24350
rect 7703 24294 7713 24350
rect 7265 24226 7713 24294
rect 7265 24170 7275 24226
rect 7331 24170 7399 24226
rect 7455 24170 7523 24226
rect 7579 24170 7647 24226
rect 7703 24170 7713 24226
rect 7265 24102 7713 24170
rect 7265 24046 7275 24102
rect 7331 24046 7399 24102
rect 7455 24046 7523 24102
rect 7579 24046 7647 24102
rect 7703 24046 7713 24102
rect 7265 24036 7713 24046
rect 9927 26954 10127 26964
rect 9927 26898 9937 26954
rect 9993 26898 10061 26954
rect 10117 26898 10127 26954
rect 9927 26830 10127 26898
rect 9927 26774 9937 26830
rect 9993 26774 10061 26830
rect 10117 26774 10127 26830
rect 9927 26706 10127 26774
rect 9927 26650 9937 26706
rect 9993 26650 10061 26706
rect 10117 26650 10127 26706
rect 9927 26582 10127 26650
rect 9927 26526 9937 26582
rect 9993 26526 10061 26582
rect 10117 26526 10127 26582
rect 9927 26458 10127 26526
rect 9927 26402 9937 26458
rect 9993 26402 10061 26458
rect 10117 26402 10127 26458
rect 9927 26334 10127 26402
rect 9927 26278 9937 26334
rect 9993 26278 10061 26334
rect 10117 26278 10127 26334
rect 9927 26210 10127 26278
rect 9927 26154 9937 26210
rect 9993 26154 10061 26210
rect 10117 26154 10127 26210
rect 9927 26086 10127 26154
rect 9927 26030 9937 26086
rect 9993 26030 10061 26086
rect 10117 26030 10127 26086
rect 9927 25962 10127 26030
rect 9927 25906 9937 25962
rect 9993 25906 10061 25962
rect 10117 25906 10127 25962
rect 9927 25838 10127 25906
rect 9927 25782 9937 25838
rect 9993 25782 10061 25838
rect 10117 25782 10127 25838
rect 9927 25714 10127 25782
rect 9927 25658 9937 25714
rect 9993 25658 10061 25714
rect 10117 25658 10127 25714
rect 9927 25590 10127 25658
rect 9927 25534 9937 25590
rect 9993 25534 10061 25590
rect 10117 25534 10127 25590
rect 9927 25466 10127 25534
rect 9927 25410 9937 25466
rect 9993 25410 10061 25466
rect 10117 25410 10127 25466
rect 9927 25342 10127 25410
rect 9927 25286 9937 25342
rect 9993 25286 10061 25342
rect 10117 25286 10127 25342
rect 9927 25218 10127 25286
rect 9927 25162 9937 25218
rect 9993 25162 10061 25218
rect 10117 25162 10127 25218
rect 9927 25094 10127 25162
rect 9927 25038 9937 25094
rect 9993 25038 10061 25094
rect 10117 25038 10127 25094
rect 9927 24970 10127 25038
rect 9927 24914 9937 24970
rect 9993 24914 10061 24970
rect 10117 24914 10127 24970
rect 9927 24846 10127 24914
rect 9927 24790 9937 24846
rect 9993 24790 10061 24846
rect 10117 24790 10127 24846
rect 9927 24722 10127 24790
rect 9927 24666 9937 24722
rect 9993 24666 10061 24722
rect 10117 24666 10127 24722
rect 9927 24598 10127 24666
rect 9927 24542 9937 24598
rect 9993 24542 10061 24598
rect 10117 24542 10127 24598
rect 9927 24474 10127 24542
rect 9927 24418 9937 24474
rect 9993 24418 10061 24474
rect 10117 24418 10127 24474
rect 9927 24350 10127 24418
rect 9927 24294 9937 24350
rect 9993 24294 10061 24350
rect 10117 24294 10127 24350
rect 9927 24226 10127 24294
rect 9927 24170 9937 24226
rect 9993 24170 10061 24226
rect 10117 24170 10127 24226
rect 9927 24102 10127 24170
rect 9927 24046 9937 24102
rect 9993 24046 10061 24102
rect 10117 24046 10127 24102
rect 9927 24036 10127 24046
rect 12297 26954 12497 26964
rect 12297 26898 12307 26954
rect 12363 26898 12431 26954
rect 12487 26898 12497 26954
rect 12297 26830 12497 26898
rect 12297 26774 12307 26830
rect 12363 26774 12431 26830
rect 12487 26774 12497 26830
rect 12297 26706 12497 26774
rect 12297 26650 12307 26706
rect 12363 26650 12431 26706
rect 12487 26650 12497 26706
rect 12297 26582 12497 26650
rect 12297 26526 12307 26582
rect 12363 26526 12431 26582
rect 12487 26526 12497 26582
rect 12297 26458 12497 26526
rect 12297 26402 12307 26458
rect 12363 26402 12431 26458
rect 12487 26402 12497 26458
rect 12297 26334 12497 26402
rect 12297 26278 12307 26334
rect 12363 26278 12431 26334
rect 12487 26278 12497 26334
rect 12297 26210 12497 26278
rect 12297 26154 12307 26210
rect 12363 26154 12431 26210
rect 12487 26154 12497 26210
rect 12297 26086 12497 26154
rect 12297 26030 12307 26086
rect 12363 26030 12431 26086
rect 12487 26030 12497 26086
rect 12297 25962 12497 26030
rect 12297 25906 12307 25962
rect 12363 25906 12431 25962
rect 12487 25906 12497 25962
rect 12297 25838 12497 25906
rect 12297 25782 12307 25838
rect 12363 25782 12431 25838
rect 12487 25782 12497 25838
rect 12297 25714 12497 25782
rect 12297 25658 12307 25714
rect 12363 25658 12431 25714
rect 12487 25658 12497 25714
rect 12297 25590 12497 25658
rect 12297 25534 12307 25590
rect 12363 25534 12431 25590
rect 12487 25534 12497 25590
rect 12297 25466 12497 25534
rect 12297 25410 12307 25466
rect 12363 25410 12431 25466
rect 12487 25410 12497 25466
rect 12297 25342 12497 25410
rect 12297 25286 12307 25342
rect 12363 25286 12431 25342
rect 12487 25286 12497 25342
rect 12297 25218 12497 25286
rect 12297 25162 12307 25218
rect 12363 25162 12431 25218
rect 12487 25162 12497 25218
rect 12297 25094 12497 25162
rect 12297 25038 12307 25094
rect 12363 25038 12431 25094
rect 12487 25038 12497 25094
rect 12297 24970 12497 25038
rect 12297 24914 12307 24970
rect 12363 24914 12431 24970
rect 12487 24914 12497 24970
rect 12297 24846 12497 24914
rect 12297 24790 12307 24846
rect 12363 24790 12431 24846
rect 12487 24790 12497 24846
rect 12297 24722 12497 24790
rect 12297 24666 12307 24722
rect 12363 24666 12431 24722
rect 12487 24666 12497 24722
rect 12297 24598 12497 24666
rect 12297 24542 12307 24598
rect 12363 24542 12431 24598
rect 12487 24542 12497 24598
rect 12297 24474 12497 24542
rect 12297 24418 12307 24474
rect 12363 24418 12431 24474
rect 12487 24418 12497 24474
rect 12297 24350 12497 24418
rect 12297 24294 12307 24350
rect 12363 24294 12431 24350
rect 12487 24294 12497 24350
rect 12297 24226 12497 24294
rect 12297 24170 12307 24226
rect 12363 24170 12431 24226
rect 12487 24170 12497 24226
rect 12297 24102 12497 24170
rect 12297 24046 12307 24102
rect 12363 24046 12431 24102
rect 12487 24046 12497 24102
rect 12297 24036 12497 24046
rect 2481 23754 2681 23764
rect 2481 23698 2491 23754
rect 2547 23698 2615 23754
rect 2671 23698 2681 23754
rect 2481 23630 2681 23698
rect 2481 23574 2491 23630
rect 2547 23574 2615 23630
rect 2671 23574 2681 23630
rect 2481 23506 2681 23574
rect 2481 23450 2491 23506
rect 2547 23450 2615 23506
rect 2671 23450 2681 23506
rect 2481 23382 2681 23450
rect 2481 23326 2491 23382
rect 2547 23326 2615 23382
rect 2671 23326 2681 23382
rect 2481 23258 2681 23326
rect 2481 23202 2491 23258
rect 2547 23202 2615 23258
rect 2671 23202 2681 23258
rect 2481 23134 2681 23202
rect 2481 23078 2491 23134
rect 2547 23078 2615 23134
rect 2671 23078 2681 23134
rect 2481 23010 2681 23078
rect 2481 22954 2491 23010
rect 2547 22954 2615 23010
rect 2671 22954 2681 23010
rect 2481 22886 2681 22954
rect 2481 22830 2491 22886
rect 2547 22830 2615 22886
rect 2671 22830 2681 22886
rect 2481 22762 2681 22830
rect 2481 22706 2491 22762
rect 2547 22706 2615 22762
rect 2671 22706 2681 22762
rect 2481 22638 2681 22706
rect 2481 22582 2491 22638
rect 2547 22582 2615 22638
rect 2671 22582 2681 22638
rect 2481 22514 2681 22582
rect 2481 22458 2491 22514
rect 2547 22458 2615 22514
rect 2671 22458 2681 22514
rect 2481 22390 2681 22458
rect 2481 22334 2491 22390
rect 2547 22334 2615 22390
rect 2671 22334 2681 22390
rect 2481 22266 2681 22334
rect 2481 22210 2491 22266
rect 2547 22210 2615 22266
rect 2671 22210 2681 22266
rect 2481 22142 2681 22210
rect 2481 22086 2491 22142
rect 2547 22086 2615 22142
rect 2671 22086 2681 22142
rect 2481 22018 2681 22086
rect 2481 21962 2491 22018
rect 2547 21962 2615 22018
rect 2671 21962 2681 22018
rect 2481 21894 2681 21962
rect 2481 21838 2491 21894
rect 2547 21838 2615 21894
rect 2671 21838 2681 21894
rect 2481 21770 2681 21838
rect 2481 21714 2491 21770
rect 2547 21714 2615 21770
rect 2671 21714 2681 21770
rect 2481 21646 2681 21714
rect 2481 21590 2491 21646
rect 2547 21590 2615 21646
rect 2671 21590 2681 21646
rect 2481 21522 2681 21590
rect 2481 21466 2491 21522
rect 2547 21466 2615 21522
rect 2671 21466 2681 21522
rect 2481 21398 2681 21466
rect 2481 21342 2491 21398
rect 2547 21342 2615 21398
rect 2671 21342 2681 21398
rect 2481 21274 2681 21342
rect 2481 21218 2491 21274
rect 2547 21218 2615 21274
rect 2671 21218 2681 21274
rect 2481 21150 2681 21218
rect 2481 21094 2491 21150
rect 2547 21094 2615 21150
rect 2671 21094 2681 21150
rect 2481 21026 2681 21094
rect 2481 20970 2491 21026
rect 2547 20970 2615 21026
rect 2671 20970 2681 21026
rect 2481 20902 2681 20970
rect 2481 20846 2491 20902
rect 2547 20846 2615 20902
rect 2671 20846 2681 20902
rect 2481 20836 2681 20846
rect 4851 23754 5051 23764
rect 4851 23698 4861 23754
rect 4917 23698 4985 23754
rect 5041 23698 5051 23754
rect 4851 23630 5051 23698
rect 4851 23574 4861 23630
rect 4917 23574 4985 23630
rect 5041 23574 5051 23630
rect 4851 23506 5051 23574
rect 4851 23450 4861 23506
rect 4917 23450 4985 23506
rect 5041 23450 5051 23506
rect 4851 23382 5051 23450
rect 4851 23326 4861 23382
rect 4917 23326 4985 23382
rect 5041 23326 5051 23382
rect 4851 23258 5051 23326
rect 4851 23202 4861 23258
rect 4917 23202 4985 23258
rect 5041 23202 5051 23258
rect 4851 23134 5051 23202
rect 4851 23078 4861 23134
rect 4917 23078 4985 23134
rect 5041 23078 5051 23134
rect 4851 23010 5051 23078
rect 4851 22954 4861 23010
rect 4917 22954 4985 23010
rect 5041 22954 5051 23010
rect 4851 22886 5051 22954
rect 4851 22830 4861 22886
rect 4917 22830 4985 22886
rect 5041 22830 5051 22886
rect 4851 22762 5051 22830
rect 4851 22706 4861 22762
rect 4917 22706 4985 22762
rect 5041 22706 5051 22762
rect 4851 22638 5051 22706
rect 4851 22582 4861 22638
rect 4917 22582 4985 22638
rect 5041 22582 5051 22638
rect 4851 22514 5051 22582
rect 4851 22458 4861 22514
rect 4917 22458 4985 22514
rect 5041 22458 5051 22514
rect 4851 22390 5051 22458
rect 4851 22334 4861 22390
rect 4917 22334 4985 22390
rect 5041 22334 5051 22390
rect 4851 22266 5051 22334
rect 4851 22210 4861 22266
rect 4917 22210 4985 22266
rect 5041 22210 5051 22266
rect 4851 22142 5051 22210
rect 4851 22086 4861 22142
rect 4917 22086 4985 22142
rect 5041 22086 5051 22142
rect 4851 22018 5051 22086
rect 4851 21962 4861 22018
rect 4917 21962 4985 22018
rect 5041 21962 5051 22018
rect 4851 21894 5051 21962
rect 4851 21838 4861 21894
rect 4917 21838 4985 21894
rect 5041 21838 5051 21894
rect 4851 21770 5051 21838
rect 4851 21714 4861 21770
rect 4917 21714 4985 21770
rect 5041 21714 5051 21770
rect 4851 21646 5051 21714
rect 4851 21590 4861 21646
rect 4917 21590 4985 21646
rect 5041 21590 5051 21646
rect 4851 21522 5051 21590
rect 4851 21466 4861 21522
rect 4917 21466 4985 21522
rect 5041 21466 5051 21522
rect 4851 21398 5051 21466
rect 4851 21342 4861 21398
rect 4917 21342 4985 21398
rect 5041 21342 5051 21398
rect 4851 21274 5051 21342
rect 4851 21218 4861 21274
rect 4917 21218 4985 21274
rect 5041 21218 5051 21274
rect 4851 21150 5051 21218
rect 4851 21094 4861 21150
rect 4917 21094 4985 21150
rect 5041 21094 5051 21150
rect 4851 21026 5051 21094
rect 4851 20970 4861 21026
rect 4917 20970 4985 21026
rect 5041 20970 5051 21026
rect 4851 20902 5051 20970
rect 4851 20846 4861 20902
rect 4917 20846 4985 20902
rect 5041 20846 5051 20902
rect 4851 20836 5051 20846
rect 7265 23754 7713 23764
rect 7265 23698 7275 23754
rect 7331 23698 7399 23754
rect 7455 23698 7523 23754
rect 7579 23698 7647 23754
rect 7703 23698 7713 23754
rect 7265 23630 7713 23698
rect 7265 23574 7275 23630
rect 7331 23574 7399 23630
rect 7455 23574 7523 23630
rect 7579 23574 7647 23630
rect 7703 23574 7713 23630
rect 7265 23506 7713 23574
rect 7265 23450 7275 23506
rect 7331 23450 7399 23506
rect 7455 23450 7523 23506
rect 7579 23450 7647 23506
rect 7703 23450 7713 23506
rect 7265 23382 7713 23450
rect 7265 23326 7275 23382
rect 7331 23326 7399 23382
rect 7455 23326 7523 23382
rect 7579 23326 7647 23382
rect 7703 23326 7713 23382
rect 7265 23258 7713 23326
rect 7265 23202 7275 23258
rect 7331 23202 7399 23258
rect 7455 23202 7523 23258
rect 7579 23202 7647 23258
rect 7703 23202 7713 23258
rect 7265 23134 7713 23202
rect 7265 23078 7275 23134
rect 7331 23078 7399 23134
rect 7455 23078 7523 23134
rect 7579 23078 7647 23134
rect 7703 23078 7713 23134
rect 7265 23010 7713 23078
rect 7265 22954 7275 23010
rect 7331 22954 7399 23010
rect 7455 22954 7523 23010
rect 7579 22954 7647 23010
rect 7703 22954 7713 23010
rect 7265 22886 7713 22954
rect 7265 22830 7275 22886
rect 7331 22830 7399 22886
rect 7455 22830 7523 22886
rect 7579 22830 7647 22886
rect 7703 22830 7713 22886
rect 7265 22762 7713 22830
rect 7265 22706 7275 22762
rect 7331 22706 7399 22762
rect 7455 22706 7523 22762
rect 7579 22706 7647 22762
rect 7703 22706 7713 22762
rect 7265 22638 7713 22706
rect 7265 22582 7275 22638
rect 7331 22582 7399 22638
rect 7455 22582 7523 22638
rect 7579 22582 7647 22638
rect 7703 22582 7713 22638
rect 7265 22514 7713 22582
rect 7265 22458 7275 22514
rect 7331 22458 7399 22514
rect 7455 22458 7523 22514
rect 7579 22458 7647 22514
rect 7703 22458 7713 22514
rect 7265 22390 7713 22458
rect 7265 22334 7275 22390
rect 7331 22334 7399 22390
rect 7455 22334 7523 22390
rect 7579 22334 7647 22390
rect 7703 22334 7713 22390
rect 7265 22266 7713 22334
rect 7265 22210 7275 22266
rect 7331 22210 7399 22266
rect 7455 22210 7523 22266
rect 7579 22210 7647 22266
rect 7703 22210 7713 22266
rect 7265 22142 7713 22210
rect 7265 22086 7275 22142
rect 7331 22086 7399 22142
rect 7455 22086 7523 22142
rect 7579 22086 7647 22142
rect 7703 22086 7713 22142
rect 7265 22018 7713 22086
rect 7265 21962 7275 22018
rect 7331 21962 7399 22018
rect 7455 21962 7523 22018
rect 7579 21962 7647 22018
rect 7703 21962 7713 22018
rect 7265 21894 7713 21962
rect 7265 21838 7275 21894
rect 7331 21838 7399 21894
rect 7455 21838 7523 21894
rect 7579 21838 7647 21894
rect 7703 21838 7713 21894
rect 7265 21770 7713 21838
rect 7265 21714 7275 21770
rect 7331 21714 7399 21770
rect 7455 21714 7523 21770
rect 7579 21714 7647 21770
rect 7703 21714 7713 21770
rect 7265 21646 7713 21714
rect 7265 21590 7275 21646
rect 7331 21590 7399 21646
rect 7455 21590 7523 21646
rect 7579 21590 7647 21646
rect 7703 21590 7713 21646
rect 7265 21522 7713 21590
rect 7265 21466 7275 21522
rect 7331 21466 7399 21522
rect 7455 21466 7523 21522
rect 7579 21466 7647 21522
rect 7703 21466 7713 21522
rect 7265 21398 7713 21466
rect 7265 21342 7275 21398
rect 7331 21342 7399 21398
rect 7455 21342 7523 21398
rect 7579 21342 7647 21398
rect 7703 21342 7713 21398
rect 7265 21274 7713 21342
rect 7265 21218 7275 21274
rect 7331 21218 7399 21274
rect 7455 21218 7523 21274
rect 7579 21218 7647 21274
rect 7703 21218 7713 21274
rect 7265 21150 7713 21218
rect 7265 21094 7275 21150
rect 7331 21094 7399 21150
rect 7455 21094 7523 21150
rect 7579 21094 7647 21150
rect 7703 21094 7713 21150
rect 7265 21026 7713 21094
rect 7265 20970 7275 21026
rect 7331 20970 7399 21026
rect 7455 20970 7523 21026
rect 7579 20970 7647 21026
rect 7703 20970 7713 21026
rect 7265 20902 7713 20970
rect 7265 20846 7275 20902
rect 7331 20846 7399 20902
rect 7455 20846 7523 20902
rect 7579 20846 7647 20902
rect 7703 20846 7713 20902
rect 7265 20836 7713 20846
rect 9927 23754 10127 23764
rect 9927 23698 9937 23754
rect 9993 23698 10061 23754
rect 10117 23698 10127 23754
rect 9927 23630 10127 23698
rect 9927 23574 9937 23630
rect 9993 23574 10061 23630
rect 10117 23574 10127 23630
rect 9927 23506 10127 23574
rect 9927 23450 9937 23506
rect 9993 23450 10061 23506
rect 10117 23450 10127 23506
rect 9927 23382 10127 23450
rect 9927 23326 9937 23382
rect 9993 23326 10061 23382
rect 10117 23326 10127 23382
rect 9927 23258 10127 23326
rect 9927 23202 9937 23258
rect 9993 23202 10061 23258
rect 10117 23202 10127 23258
rect 9927 23134 10127 23202
rect 9927 23078 9937 23134
rect 9993 23078 10061 23134
rect 10117 23078 10127 23134
rect 9927 23010 10127 23078
rect 9927 22954 9937 23010
rect 9993 22954 10061 23010
rect 10117 22954 10127 23010
rect 9927 22886 10127 22954
rect 9927 22830 9937 22886
rect 9993 22830 10061 22886
rect 10117 22830 10127 22886
rect 9927 22762 10127 22830
rect 9927 22706 9937 22762
rect 9993 22706 10061 22762
rect 10117 22706 10127 22762
rect 9927 22638 10127 22706
rect 9927 22582 9937 22638
rect 9993 22582 10061 22638
rect 10117 22582 10127 22638
rect 9927 22514 10127 22582
rect 9927 22458 9937 22514
rect 9993 22458 10061 22514
rect 10117 22458 10127 22514
rect 9927 22390 10127 22458
rect 9927 22334 9937 22390
rect 9993 22334 10061 22390
rect 10117 22334 10127 22390
rect 9927 22266 10127 22334
rect 9927 22210 9937 22266
rect 9993 22210 10061 22266
rect 10117 22210 10127 22266
rect 9927 22142 10127 22210
rect 9927 22086 9937 22142
rect 9993 22086 10061 22142
rect 10117 22086 10127 22142
rect 9927 22018 10127 22086
rect 9927 21962 9937 22018
rect 9993 21962 10061 22018
rect 10117 21962 10127 22018
rect 9927 21894 10127 21962
rect 9927 21838 9937 21894
rect 9993 21838 10061 21894
rect 10117 21838 10127 21894
rect 9927 21770 10127 21838
rect 9927 21714 9937 21770
rect 9993 21714 10061 21770
rect 10117 21714 10127 21770
rect 9927 21646 10127 21714
rect 9927 21590 9937 21646
rect 9993 21590 10061 21646
rect 10117 21590 10127 21646
rect 9927 21522 10127 21590
rect 9927 21466 9937 21522
rect 9993 21466 10061 21522
rect 10117 21466 10127 21522
rect 9927 21398 10127 21466
rect 9927 21342 9937 21398
rect 9993 21342 10061 21398
rect 10117 21342 10127 21398
rect 9927 21274 10127 21342
rect 9927 21218 9937 21274
rect 9993 21218 10061 21274
rect 10117 21218 10127 21274
rect 9927 21150 10127 21218
rect 9927 21094 9937 21150
rect 9993 21094 10061 21150
rect 10117 21094 10127 21150
rect 9927 21026 10127 21094
rect 9927 20970 9937 21026
rect 9993 20970 10061 21026
rect 10117 20970 10127 21026
rect 9927 20902 10127 20970
rect 9927 20846 9937 20902
rect 9993 20846 10061 20902
rect 10117 20846 10127 20902
rect 9927 20836 10127 20846
rect 12297 23754 12497 23764
rect 12297 23698 12307 23754
rect 12363 23698 12431 23754
rect 12487 23698 12497 23754
rect 12297 23630 12497 23698
rect 12297 23574 12307 23630
rect 12363 23574 12431 23630
rect 12487 23574 12497 23630
rect 12297 23506 12497 23574
rect 12297 23450 12307 23506
rect 12363 23450 12431 23506
rect 12487 23450 12497 23506
rect 12297 23382 12497 23450
rect 12297 23326 12307 23382
rect 12363 23326 12431 23382
rect 12487 23326 12497 23382
rect 12297 23258 12497 23326
rect 12297 23202 12307 23258
rect 12363 23202 12431 23258
rect 12487 23202 12497 23258
rect 12297 23134 12497 23202
rect 12297 23078 12307 23134
rect 12363 23078 12431 23134
rect 12487 23078 12497 23134
rect 12297 23010 12497 23078
rect 12297 22954 12307 23010
rect 12363 22954 12431 23010
rect 12487 22954 12497 23010
rect 12297 22886 12497 22954
rect 12297 22830 12307 22886
rect 12363 22830 12431 22886
rect 12487 22830 12497 22886
rect 12297 22762 12497 22830
rect 12297 22706 12307 22762
rect 12363 22706 12431 22762
rect 12487 22706 12497 22762
rect 12297 22638 12497 22706
rect 12297 22582 12307 22638
rect 12363 22582 12431 22638
rect 12487 22582 12497 22638
rect 12297 22514 12497 22582
rect 12297 22458 12307 22514
rect 12363 22458 12431 22514
rect 12487 22458 12497 22514
rect 12297 22390 12497 22458
rect 12297 22334 12307 22390
rect 12363 22334 12431 22390
rect 12487 22334 12497 22390
rect 12297 22266 12497 22334
rect 12297 22210 12307 22266
rect 12363 22210 12431 22266
rect 12487 22210 12497 22266
rect 12297 22142 12497 22210
rect 12297 22086 12307 22142
rect 12363 22086 12431 22142
rect 12487 22086 12497 22142
rect 12297 22018 12497 22086
rect 12297 21962 12307 22018
rect 12363 21962 12431 22018
rect 12487 21962 12497 22018
rect 12297 21894 12497 21962
rect 12297 21838 12307 21894
rect 12363 21838 12431 21894
rect 12487 21838 12497 21894
rect 12297 21770 12497 21838
rect 12297 21714 12307 21770
rect 12363 21714 12431 21770
rect 12487 21714 12497 21770
rect 12297 21646 12497 21714
rect 12297 21590 12307 21646
rect 12363 21590 12431 21646
rect 12487 21590 12497 21646
rect 12297 21522 12497 21590
rect 12297 21466 12307 21522
rect 12363 21466 12431 21522
rect 12487 21466 12497 21522
rect 12297 21398 12497 21466
rect 12297 21342 12307 21398
rect 12363 21342 12431 21398
rect 12487 21342 12497 21398
rect 12297 21274 12497 21342
rect 12297 21218 12307 21274
rect 12363 21218 12431 21274
rect 12487 21218 12497 21274
rect 12297 21150 12497 21218
rect 12297 21094 12307 21150
rect 12363 21094 12431 21150
rect 12487 21094 12497 21150
rect 12297 21026 12497 21094
rect 12297 20970 12307 21026
rect 12363 20970 12431 21026
rect 12487 20970 12497 21026
rect 12297 20902 12497 20970
rect 12297 20846 12307 20902
rect 12363 20846 12431 20902
rect 12487 20846 12497 20902
rect 12297 20836 12497 20846
rect 2481 20554 2681 20564
rect 2481 20498 2491 20554
rect 2547 20498 2615 20554
rect 2671 20498 2681 20554
rect 2481 20430 2681 20498
rect 2481 20374 2491 20430
rect 2547 20374 2615 20430
rect 2671 20374 2681 20430
rect 2481 20306 2681 20374
rect 2481 20250 2491 20306
rect 2547 20250 2615 20306
rect 2671 20250 2681 20306
rect 2481 20182 2681 20250
rect 2481 20126 2491 20182
rect 2547 20126 2615 20182
rect 2671 20126 2681 20182
rect 2481 20058 2681 20126
rect 2481 20002 2491 20058
rect 2547 20002 2615 20058
rect 2671 20002 2681 20058
rect 2481 19934 2681 20002
rect 2481 19878 2491 19934
rect 2547 19878 2615 19934
rect 2671 19878 2681 19934
rect 2481 19810 2681 19878
rect 2481 19754 2491 19810
rect 2547 19754 2615 19810
rect 2671 19754 2681 19810
rect 2481 19686 2681 19754
rect 2481 19630 2491 19686
rect 2547 19630 2615 19686
rect 2671 19630 2681 19686
rect 2481 19562 2681 19630
rect 2481 19506 2491 19562
rect 2547 19506 2615 19562
rect 2671 19506 2681 19562
rect 2481 19438 2681 19506
rect 2481 19382 2491 19438
rect 2547 19382 2615 19438
rect 2671 19382 2681 19438
rect 2481 19314 2681 19382
rect 2481 19258 2491 19314
rect 2547 19258 2615 19314
rect 2671 19258 2681 19314
rect 2481 19190 2681 19258
rect 2481 19134 2491 19190
rect 2547 19134 2615 19190
rect 2671 19134 2681 19190
rect 2481 19066 2681 19134
rect 2481 19010 2491 19066
rect 2547 19010 2615 19066
rect 2671 19010 2681 19066
rect 2481 18942 2681 19010
rect 2481 18886 2491 18942
rect 2547 18886 2615 18942
rect 2671 18886 2681 18942
rect 2481 18818 2681 18886
rect 2481 18762 2491 18818
rect 2547 18762 2615 18818
rect 2671 18762 2681 18818
rect 2481 18694 2681 18762
rect 2481 18638 2491 18694
rect 2547 18638 2615 18694
rect 2671 18638 2681 18694
rect 2481 18570 2681 18638
rect 2481 18514 2491 18570
rect 2547 18514 2615 18570
rect 2671 18514 2681 18570
rect 2481 18446 2681 18514
rect 2481 18390 2491 18446
rect 2547 18390 2615 18446
rect 2671 18390 2681 18446
rect 2481 18322 2681 18390
rect 2481 18266 2491 18322
rect 2547 18266 2615 18322
rect 2671 18266 2681 18322
rect 2481 18198 2681 18266
rect 2481 18142 2491 18198
rect 2547 18142 2615 18198
rect 2671 18142 2681 18198
rect 2481 18074 2681 18142
rect 2481 18018 2491 18074
rect 2547 18018 2615 18074
rect 2671 18018 2681 18074
rect 2481 17950 2681 18018
rect 2481 17894 2491 17950
rect 2547 17894 2615 17950
rect 2671 17894 2681 17950
rect 2481 17826 2681 17894
rect 2481 17770 2491 17826
rect 2547 17770 2615 17826
rect 2671 17770 2681 17826
rect 2481 17702 2681 17770
rect 2481 17646 2491 17702
rect 2547 17646 2615 17702
rect 2671 17646 2681 17702
rect 2481 17636 2681 17646
rect 4851 20554 5051 20564
rect 4851 20498 4861 20554
rect 4917 20498 4985 20554
rect 5041 20498 5051 20554
rect 4851 20430 5051 20498
rect 4851 20374 4861 20430
rect 4917 20374 4985 20430
rect 5041 20374 5051 20430
rect 4851 20306 5051 20374
rect 4851 20250 4861 20306
rect 4917 20250 4985 20306
rect 5041 20250 5051 20306
rect 4851 20182 5051 20250
rect 4851 20126 4861 20182
rect 4917 20126 4985 20182
rect 5041 20126 5051 20182
rect 4851 20058 5051 20126
rect 4851 20002 4861 20058
rect 4917 20002 4985 20058
rect 5041 20002 5051 20058
rect 4851 19934 5051 20002
rect 4851 19878 4861 19934
rect 4917 19878 4985 19934
rect 5041 19878 5051 19934
rect 4851 19810 5051 19878
rect 4851 19754 4861 19810
rect 4917 19754 4985 19810
rect 5041 19754 5051 19810
rect 4851 19686 5051 19754
rect 4851 19630 4861 19686
rect 4917 19630 4985 19686
rect 5041 19630 5051 19686
rect 4851 19562 5051 19630
rect 4851 19506 4861 19562
rect 4917 19506 4985 19562
rect 5041 19506 5051 19562
rect 4851 19438 5051 19506
rect 4851 19382 4861 19438
rect 4917 19382 4985 19438
rect 5041 19382 5051 19438
rect 4851 19314 5051 19382
rect 4851 19258 4861 19314
rect 4917 19258 4985 19314
rect 5041 19258 5051 19314
rect 4851 19190 5051 19258
rect 4851 19134 4861 19190
rect 4917 19134 4985 19190
rect 5041 19134 5051 19190
rect 4851 19066 5051 19134
rect 4851 19010 4861 19066
rect 4917 19010 4985 19066
rect 5041 19010 5051 19066
rect 4851 18942 5051 19010
rect 4851 18886 4861 18942
rect 4917 18886 4985 18942
rect 5041 18886 5051 18942
rect 4851 18818 5051 18886
rect 4851 18762 4861 18818
rect 4917 18762 4985 18818
rect 5041 18762 5051 18818
rect 4851 18694 5051 18762
rect 4851 18638 4861 18694
rect 4917 18638 4985 18694
rect 5041 18638 5051 18694
rect 4851 18570 5051 18638
rect 4851 18514 4861 18570
rect 4917 18514 4985 18570
rect 5041 18514 5051 18570
rect 4851 18446 5051 18514
rect 4851 18390 4861 18446
rect 4917 18390 4985 18446
rect 5041 18390 5051 18446
rect 4851 18322 5051 18390
rect 4851 18266 4861 18322
rect 4917 18266 4985 18322
rect 5041 18266 5051 18322
rect 4851 18198 5051 18266
rect 4851 18142 4861 18198
rect 4917 18142 4985 18198
rect 5041 18142 5051 18198
rect 4851 18074 5051 18142
rect 4851 18018 4861 18074
rect 4917 18018 4985 18074
rect 5041 18018 5051 18074
rect 4851 17950 5051 18018
rect 4851 17894 4861 17950
rect 4917 17894 4985 17950
rect 5041 17894 5051 17950
rect 4851 17826 5051 17894
rect 4851 17770 4861 17826
rect 4917 17770 4985 17826
rect 5041 17770 5051 17826
rect 4851 17702 5051 17770
rect 4851 17646 4861 17702
rect 4917 17646 4985 17702
rect 5041 17646 5051 17702
rect 4851 17636 5051 17646
rect 7265 20554 7713 20564
rect 7265 20498 7275 20554
rect 7331 20498 7399 20554
rect 7455 20498 7523 20554
rect 7579 20498 7647 20554
rect 7703 20498 7713 20554
rect 7265 20430 7713 20498
rect 7265 20374 7275 20430
rect 7331 20374 7399 20430
rect 7455 20374 7523 20430
rect 7579 20374 7647 20430
rect 7703 20374 7713 20430
rect 7265 20306 7713 20374
rect 7265 20250 7275 20306
rect 7331 20250 7399 20306
rect 7455 20250 7523 20306
rect 7579 20250 7647 20306
rect 7703 20250 7713 20306
rect 7265 20182 7713 20250
rect 7265 20126 7275 20182
rect 7331 20126 7399 20182
rect 7455 20126 7523 20182
rect 7579 20126 7647 20182
rect 7703 20126 7713 20182
rect 7265 20058 7713 20126
rect 7265 20002 7275 20058
rect 7331 20002 7399 20058
rect 7455 20002 7523 20058
rect 7579 20002 7647 20058
rect 7703 20002 7713 20058
rect 7265 19934 7713 20002
rect 7265 19878 7275 19934
rect 7331 19878 7399 19934
rect 7455 19878 7523 19934
rect 7579 19878 7647 19934
rect 7703 19878 7713 19934
rect 7265 19810 7713 19878
rect 7265 19754 7275 19810
rect 7331 19754 7399 19810
rect 7455 19754 7523 19810
rect 7579 19754 7647 19810
rect 7703 19754 7713 19810
rect 7265 19686 7713 19754
rect 7265 19630 7275 19686
rect 7331 19630 7399 19686
rect 7455 19630 7523 19686
rect 7579 19630 7647 19686
rect 7703 19630 7713 19686
rect 7265 19562 7713 19630
rect 7265 19506 7275 19562
rect 7331 19506 7399 19562
rect 7455 19506 7523 19562
rect 7579 19506 7647 19562
rect 7703 19506 7713 19562
rect 7265 19438 7713 19506
rect 7265 19382 7275 19438
rect 7331 19382 7399 19438
rect 7455 19382 7523 19438
rect 7579 19382 7647 19438
rect 7703 19382 7713 19438
rect 7265 19314 7713 19382
rect 7265 19258 7275 19314
rect 7331 19258 7399 19314
rect 7455 19258 7523 19314
rect 7579 19258 7647 19314
rect 7703 19258 7713 19314
rect 7265 19190 7713 19258
rect 7265 19134 7275 19190
rect 7331 19134 7399 19190
rect 7455 19134 7523 19190
rect 7579 19134 7647 19190
rect 7703 19134 7713 19190
rect 7265 19066 7713 19134
rect 7265 19010 7275 19066
rect 7331 19010 7399 19066
rect 7455 19010 7523 19066
rect 7579 19010 7647 19066
rect 7703 19010 7713 19066
rect 7265 18942 7713 19010
rect 7265 18886 7275 18942
rect 7331 18886 7399 18942
rect 7455 18886 7523 18942
rect 7579 18886 7647 18942
rect 7703 18886 7713 18942
rect 7265 18818 7713 18886
rect 7265 18762 7275 18818
rect 7331 18762 7399 18818
rect 7455 18762 7523 18818
rect 7579 18762 7647 18818
rect 7703 18762 7713 18818
rect 7265 18694 7713 18762
rect 7265 18638 7275 18694
rect 7331 18638 7399 18694
rect 7455 18638 7523 18694
rect 7579 18638 7647 18694
rect 7703 18638 7713 18694
rect 7265 18570 7713 18638
rect 7265 18514 7275 18570
rect 7331 18514 7399 18570
rect 7455 18514 7523 18570
rect 7579 18514 7647 18570
rect 7703 18514 7713 18570
rect 7265 18446 7713 18514
rect 7265 18390 7275 18446
rect 7331 18390 7399 18446
rect 7455 18390 7523 18446
rect 7579 18390 7647 18446
rect 7703 18390 7713 18446
rect 7265 18322 7713 18390
rect 7265 18266 7275 18322
rect 7331 18266 7399 18322
rect 7455 18266 7523 18322
rect 7579 18266 7647 18322
rect 7703 18266 7713 18322
rect 7265 18198 7713 18266
rect 7265 18142 7275 18198
rect 7331 18142 7399 18198
rect 7455 18142 7523 18198
rect 7579 18142 7647 18198
rect 7703 18142 7713 18198
rect 7265 18074 7713 18142
rect 7265 18018 7275 18074
rect 7331 18018 7399 18074
rect 7455 18018 7523 18074
rect 7579 18018 7647 18074
rect 7703 18018 7713 18074
rect 7265 17950 7713 18018
rect 7265 17894 7275 17950
rect 7331 17894 7399 17950
rect 7455 17894 7523 17950
rect 7579 17894 7647 17950
rect 7703 17894 7713 17950
rect 7265 17826 7713 17894
rect 7265 17770 7275 17826
rect 7331 17770 7399 17826
rect 7455 17770 7523 17826
rect 7579 17770 7647 17826
rect 7703 17770 7713 17826
rect 7265 17702 7713 17770
rect 7265 17646 7275 17702
rect 7331 17646 7399 17702
rect 7455 17646 7523 17702
rect 7579 17646 7647 17702
rect 7703 17646 7713 17702
rect 7265 17636 7713 17646
rect 9927 20554 10127 20564
rect 9927 20498 9937 20554
rect 9993 20498 10061 20554
rect 10117 20498 10127 20554
rect 9927 20430 10127 20498
rect 9927 20374 9937 20430
rect 9993 20374 10061 20430
rect 10117 20374 10127 20430
rect 9927 20306 10127 20374
rect 9927 20250 9937 20306
rect 9993 20250 10061 20306
rect 10117 20250 10127 20306
rect 9927 20182 10127 20250
rect 9927 20126 9937 20182
rect 9993 20126 10061 20182
rect 10117 20126 10127 20182
rect 9927 20058 10127 20126
rect 9927 20002 9937 20058
rect 9993 20002 10061 20058
rect 10117 20002 10127 20058
rect 9927 19934 10127 20002
rect 9927 19878 9937 19934
rect 9993 19878 10061 19934
rect 10117 19878 10127 19934
rect 9927 19810 10127 19878
rect 9927 19754 9937 19810
rect 9993 19754 10061 19810
rect 10117 19754 10127 19810
rect 9927 19686 10127 19754
rect 9927 19630 9937 19686
rect 9993 19630 10061 19686
rect 10117 19630 10127 19686
rect 9927 19562 10127 19630
rect 9927 19506 9937 19562
rect 9993 19506 10061 19562
rect 10117 19506 10127 19562
rect 9927 19438 10127 19506
rect 9927 19382 9937 19438
rect 9993 19382 10061 19438
rect 10117 19382 10127 19438
rect 9927 19314 10127 19382
rect 9927 19258 9937 19314
rect 9993 19258 10061 19314
rect 10117 19258 10127 19314
rect 9927 19190 10127 19258
rect 9927 19134 9937 19190
rect 9993 19134 10061 19190
rect 10117 19134 10127 19190
rect 9927 19066 10127 19134
rect 9927 19010 9937 19066
rect 9993 19010 10061 19066
rect 10117 19010 10127 19066
rect 9927 18942 10127 19010
rect 9927 18886 9937 18942
rect 9993 18886 10061 18942
rect 10117 18886 10127 18942
rect 9927 18818 10127 18886
rect 9927 18762 9937 18818
rect 9993 18762 10061 18818
rect 10117 18762 10127 18818
rect 9927 18694 10127 18762
rect 9927 18638 9937 18694
rect 9993 18638 10061 18694
rect 10117 18638 10127 18694
rect 9927 18570 10127 18638
rect 9927 18514 9937 18570
rect 9993 18514 10061 18570
rect 10117 18514 10127 18570
rect 9927 18446 10127 18514
rect 9927 18390 9937 18446
rect 9993 18390 10061 18446
rect 10117 18390 10127 18446
rect 9927 18322 10127 18390
rect 9927 18266 9937 18322
rect 9993 18266 10061 18322
rect 10117 18266 10127 18322
rect 9927 18198 10127 18266
rect 9927 18142 9937 18198
rect 9993 18142 10061 18198
rect 10117 18142 10127 18198
rect 9927 18074 10127 18142
rect 9927 18018 9937 18074
rect 9993 18018 10061 18074
rect 10117 18018 10127 18074
rect 9927 17950 10127 18018
rect 9927 17894 9937 17950
rect 9993 17894 10061 17950
rect 10117 17894 10127 17950
rect 9927 17826 10127 17894
rect 9927 17770 9937 17826
rect 9993 17770 10061 17826
rect 10117 17770 10127 17826
rect 9927 17702 10127 17770
rect 9927 17646 9937 17702
rect 9993 17646 10061 17702
rect 10117 17646 10127 17702
rect 9927 17636 10127 17646
rect 12297 20554 12497 20564
rect 12297 20498 12307 20554
rect 12363 20498 12431 20554
rect 12487 20498 12497 20554
rect 12297 20430 12497 20498
rect 12297 20374 12307 20430
rect 12363 20374 12431 20430
rect 12487 20374 12497 20430
rect 12297 20306 12497 20374
rect 12297 20250 12307 20306
rect 12363 20250 12431 20306
rect 12487 20250 12497 20306
rect 12297 20182 12497 20250
rect 12297 20126 12307 20182
rect 12363 20126 12431 20182
rect 12487 20126 12497 20182
rect 12297 20058 12497 20126
rect 12297 20002 12307 20058
rect 12363 20002 12431 20058
rect 12487 20002 12497 20058
rect 12297 19934 12497 20002
rect 12297 19878 12307 19934
rect 12363 19878 12431 19934
rect 12487 19878 12497 19934
rect 12297 19810 12497 19878
rect 12297 19754 12307 19810
rect 12363 19754 12431 19810
rect 12487 19754 12497 19810
rect 12297 19686 12497 19754
rect 12297 19630 12307 19686
rect 12363 19630 12431 19686
rect 12487 19630 12497 19686
rect 12297 19562 12497 19630
rect 12297 19506 12307 19562
rect 12363 19506 12431 19562
rect 12487 19506 12497 19562
rect 12297 19438 12497 19506
rect 12297 19382 12307 19438
rect 12363 19382 12431 19438
rect 12487 19382 12497 19438
rect 12297 19314 12497 19382
rect 12297 19258 12307 19314
rect 12363 19258 12431 19314
rect 12487 19258 12497 19314
rect 12297 19190 12497 19258
rect 12297 19134 12307 19190
rect 12363 19134 12431 19190
rect 12487 19134 12497 19190
rect 12297 19066 12497 19134
rect 12297 19010 12307 19066
rect 12363 19010 12431 19066
rect 12487 19010 12497 19066
rect 12297 18942 12497 19010
rect 12297 18886 12307 18942
rect 12363 18886 12431 18942
rect 12487 18886 12497 18942
rect 12297 18818 12497 18886
rect 12297 18762 12307 18818
rect 12363 18762 12431 18818
rect 12487 18762 12497 18818
rect 12297 18694 12497 18762
rect 12297 18638 12307 18694
rect 12363 18638 12431 18694
rect 12487 18638 12497 18694
rect 12297 18570 12497 18638
rect 12297 18514 12307 18570
rect 12363 18514 12431 18570
rect 12487 18514 12497 18570
rect 12297 18446 12497 18514
rect 12297 18390 12307 18446
rect 12363 18390 12431 18446
rect 12487 18390 12497 18446
rect 12297 18322 12497 18390
rect 12297 18266 12307 18322
rect 12363 18266 12431 18322
rect 12487 18266 12497 18322
rect 12297 18198 12497 18266
rect 12297 18142 12307 18198
rect 12363 18142 12431 18198
rect 12487 18142 12497 18198
rect 12297 18074 12497 18142
rect 12297 18018 12307 18074
rect 12363 18018 12431 18074
rect 12487 18018 12497 18074
rect 12297 17950 12497 18018
rect 12297 17894 12307 17950
rect 12363 17894 12431 17950
rect 12487 17894 12497 17950
rect 12297 17826 12497 17894
rect 12297 17770 12307 17826
rect 12363 17770 12431 17826
rect 12487 17770 12497 17826
rect 12297 17702 12497 17770
rect 12297 17646 12307 17702
rect 12363 17646 12431 17702
rect 12487 17646 12497 17702
rect 12297 17636 12497 17646
rect 2481 17354 2681 17364
rect 2481 17298 2491 17354
rect 2547 17298 2615 17354
rect 2671 17298 2681 17354
rect 2481 17230 2681 17298
rect 2481 17174 2491 17230
rect 2547 17174 2615 17230
rect 2671 17174 2681 17230
rect 2481 17106 2681 17174
rect 2481 17050 2491 17106
rect 2547 17050 2615 17106
rect 2671 17050 2681 17106
rect 2481 16982 2681 17050
rect 2481 16926 2491 16982
rect 2547 16926 2615 16982
rect 2671 16926 2681 16982
rect 2481 16858 2681 16926
rect 2481 16802 2491 16858
rect 2547 16802 2615 16858
rect 2671 16802 2681 16858
rect 2481 16734 2681 16802
rect 2481 16678 2491 16734
rect 2547 16678 2615 16734
rect 2671 16678 2681 16734
rect 2481 16610 2681 16678
rect 2481 16554 2491 16610
rect 2547 16554 2615 16610
rect 2671 16554 2681 16610
rect 2481 16486 2681 16554
rect 2481 16430 2491 16486
rect 2547 16430 2615 16486
rect 2671 16430 2681 16486
rect 2481 16362 2681 16430
rect 2481 16306 2491 16362
rect 2547 16306 2615 16362
rect 2671 16306 2681 16362
rect 2481 16238 2681 16306
rect 2481 16182 2491 16238
rect 2547 16182 2615 16238
rect 2671 16182 2681 16238
rect 2481 16114 2681 16182
rect 2481 16058 2491 16114
rect 2547 16058 2615 16114
rect 2671 16058 2681 16114
rect 2481 15990 2681 16058
rect 2481 15934 2491 15990
rect 2547 15934 2615 15990
rect 2671 15934 2681 15990
rect 2481 15866 2681 15934
rect 2481 15810 2491 15866
rect 2547 15810 2615 15866
rect 2671 15810 2681 15866
rect 2481 15742 2681 15810
rect 2481 15686 2491 15742
rect 2547 15686 2615 15742
rect 2671 15686 2681 15742
rect 2481 15618 2681 15686
rect 2481 15562 2491 15618
rect 2547 15562 2615 15618
rect 2671 15562 2681 15618
rect 2481 15494 2681 15562
rect 2481 15438 2491 15494
rect 2547 15438 2615 15494
rect 2671 15438 2681 15494
rect 2481 15370 2681 15438
rect 2481 15314 2491 15370
rect 2547 15314 2615 15370
rect 2671 15314 2681 15370
rect 2481 15246 2681 15314
rect 2481 15190 2491 15246
rect 2547 15190 2615 15246
rect 2671 15190 2681 15246
rect 2481 15122 2681 15190
rect 2481 15066 2491 15122
rect 2547 15066 2615 15122
rect 2671 15066 2681 15122
rect 2481 14998 2681 15066
rect 2481 14942 2491 14998
rect 2547 14942 2615 14998
rect 2671 14942 2681 14998
rect 2481 14874 2681 14942
rect 2481 14818 2491 14874
rect 2547 14818 2615 14874
rect 2671 14818 2681 14874
rect 2481 14750 2681 14818
rect 2481 14694 2491 14750
rect 2547 14694 2615 14750
rect 2671 14694 2681 14750
rect 2481 14626 2681 14694
rect 2481 14570 2491 14626
rect 2547 14570 2615 14626
rect 2671 14570 2681 14626
rect 2481 14502 2681 14570
rect 2481 14446 2491 14502
rect 2547 14446 2615 14502
rect 2671 14446 2681 14502
rect 2481 14436 2681 14446
rect 4851 17354 5051 17364
rect 4851 17298 4861 17354
rect 4917 17298 4985 17354
rect 5041 17298 5051 17354
rect 4851 17230 5051 17298
rect 4851 17174 4861 17230
rect 4917 17174 4985 17230
rect 5041 17174 5051 17230
rect 4851 17106 5051 17174
rect 4851 17050 4861 17106
rect 4917 17050 4985 17106
rect 5041 17050 5051 17106
rect 4851 16982 5051 17050
rect 4851 16926 4861 16982
rect 4917 16926 4985 16982
rect 5041 16926 5051 16982
rect 4851 16858 5051 16926
rect 4851 16802 4861 16858
rect 4917 16802 4985 16858
rect 5041 16802 5051 16858
rect 4851 16734 5051 16802
rect 4851 16678 4861 16734
rect 4917 16678 4985 16734
rect 5041 16678 5051 16734
rect 4851 16610 5051 16678
rect 4851 16554 4861 16610
rect 4917 16554 4985 16610
rect 5041 16554 5051 16610
rect 4851 16486 5051 16554
rect 4851 16430 4861 16486
rect 4917 16430 4985 16486
rect 5041 16430 5051 16486
rect 4851 16362 5051 16430
rect 4851 16306 4861 16362
rect 4917 16306 4985 16362
rect 5041 16306 5051 16362
rect 4851 16238 5051 16306
rect 4851 16182 4861 16238
rect 4917 16182 4985 16238
rect 5041 16182 5051 16238
rect 4851 16114 5051 16182
rect 4851 16058 4861 16114
rect 4917 16058 4985 16114
rect 5041 16058 5051 16114
rect 4851 15990 5051 16058
rect 4851 15934 4861 15990
rect 4917 15934 4985 15990
rect 5041 15934 5051 15990
rect 4851 15866 5051 15934
rect 4851 15810 4861 15866
rect 4917 15810 4985 15866
rect 5041 15810 5051 15866
rect 4851 15742 5051 15810
rect 4851 15686 4861 15742
rect 4917 15686 4985 15742
rect 5041 15686 5051 15742
rect 4851 15618 5051 15686
rect 4851 15562 4861 15618
rect 4917 15562 4985 15618
rect 5041 15562 5051 15618
rect 4851 15494 5051 15562
rect 4851 15438 4861 15494
rect 4917 15438 4985 15494
rect 5041 15438 5051 15494
rect 4851 15370 5051 15438
rect 4851 15314 4861 15370
rect 4917 15314 4985 15370
rect 5041 15314 5051 15370
rect 4851 15246 5051 15314
rect 4851 15190 4861 15246
rect 4917 15190 4985 15246
rect 5041 15190 5051 15246
rect 4851 15122 5051 15190
rect 4851 15066 4861 15122
rect 4917 15066 4985 15122
rect 5041 15066 5051 15122
rect 4851 14998 5051 15066
rect 4851 14942 4861 14998
rect 4917 14942 4985 14998
rect 5041 14942 5051 14998
rect 4851 14874 5051 14942
rect 4851 14818 4861 14874
rect 4917 14818 4985 14874
rect 5041 14818 5051 14874
rect 4851 14750 5051 14818
rect 4851 14694 4861 14750
rect 4917 14694 4985 14750
rect 5041 14694 5051 14750
rect 4851 14626 5051 14694
rect 4851 14570 4861 14626
rect 4917 14570 4985 14626
rect 5041 14570 5051 14626
rect 4851 14502 5051 14570
rect 4851 14446 4861 14502
rect 4917 14446 4985 14502
rect 5041 14446 5051 14502
rect 4851 14436 5051 14446
rect 7265 17354 7713 17364
rect 7265 17298 7275 17354
rect 7331 17298 7399 17354
rect 7455 17298 7523 17354
rect 7579 17298 7647 17354
rect 7703 17298 7713 17354
rect 7265 17230 7713 17298
rect 7265 17174 7275 17230
rect 7331 17174 7399 17230
rect 7455 17174 7523 17230
rect 7579 17174 7647 17230
rect 7703 17174 7713 17230
rect 7265 17106 7713 17174
rect 7265 17050 7275 17106
rect 7331 17050 7399 17106
rect 7455 17050 7523 17106
rect 7579 17050 7647 17106
rect 7703 17050 7713 17106
rect 7265 16982 7713 17050
rect 7265 16926 7275 16982
rect 7331 16926 7399 16982
rect 7455 16926 7523 16982
rect 7579 16926 7647 16982
rect 7703 16926 7713 16982
rect 7265 16858 7713 16926
rect 7265 16802 7275 16858
rect 7331 16802 7399 16858
rect 7455 16802 7523 16858
rect 7579 16802 7647 16858
rect 7703 16802 7713 16858
rect 7265 16734 7713 16802
rect 7265 16678 7275 16734
rect 7331 16678 7399 16734
rect 7455 16678 7523 16734
rect 7579 16678 7647 16734
rect 7703 16678 7713 16734
rect 7265 16610 7713 16678
rect 7265 16554 7275 16610
rect 7331 16554 7399 16610
rect 7455 16554 7523 16610
rect 7579 16554 7647 16610
rect 7703 16554 7713 16610
rect 7265 16486 7713 16554
rect 7265 16430 7275 16486
rect 7331 16430 7399 16486
rect 7455 16430 7523 16486
rect 7579 16430 7647 16486
rect 7703 16430 7713 16486
rect 7265 16362 7713 16430
rect 7265 16306 7275 16362
rect 7331 16306 7399 16362
rect 7455 16306 7523 16362
rect 7579 16306 7647 16362
rect 7703 16306 7713 16362
rect 7265 16238 7713 16306
rect 7265 16182 7275 16238
rect 7331 16182 7399 16238
rect 7455 16182 7523 16238
rect 7579 16182 7647 16238
rect 7703 16182 7713 16238
rect 7265 16114 7713 16182
rect 7265 16058 7275 16114
rect 7331 16058 7399 16114
rect 7455 16058 7523 16114
rect 7579 16058 7647 16114
rect 7703 16058 7713 16114
rect 7265 15990 7713 16058
rect 7265 15934 7275 15990
rect 7331 15934 7399 15990
rect 7455 15934 7523 15990
rect 7579 15934 7647 15990
rect 7703 15934 7713 15990
rect 7265 15866 7713 15934
rect 7265 15810 7275 15866
rect 7331 15810 7399 15866
rect 7455 15810 7523 15866
rect 7579 15810 7647 15866
rect 7703 15810 7713 15866
rect 7265 15742 7713 15810
rect 7265 15686 7275 15742
rect 7331 15686 7399 15742
rect 7455 15686 7523 15742
rect 7579 15686 7647 15742
rect 7703 15686 7713 15742
rect 7265 15618 7713 15686
rect 7265 15562 7275 15618
rect 7331 15562 7399 15618
rect 7455 15562 7523 15618
rect 7579 15562 7647 15618
rect 7703 15562 7713 15618
rect 7265 15494 7713 15562
rect 7265 15438 7275 15494
rect 7331 15438 7399 15494
rect 7455 15438 7523 15494
rect 7579 15438 7647 15494
rect 7703 15438 7713 15494
rect 7265 15370 7713 15438
rect 7265 15314 7275 15370
rect 7331 15314 7399 15370
rect 7455 15314 7523 15370
rect 7579 15314 7647 15370
rect 7703 15314 7713 15370
rect 7265 15246 7713 15314
rect 7265 15190 7275 15246
rect 7331 15190 7399 15246
rect 7455 15190 7523 15246
rect 7579 15190 7647 15246
rect 7703 15190 7713 15246
rect 7265 15122 7713 15190
rect 7265 15066 7275 15122
rect 7331 15066 7399 15122
rect 7455 15066 7523 15122
rect 7579 15066 7647 15122
rect 7703 15066 7713 15122
rect 7265 14998 7713 15066
rect 7265 14942 7275 14998
rect 7331 14942 7399 14998
rect 7455 14942 7523 14998
rect 7579 14942 7647 14998
rect 7703 14942 7713 14998
rect 7265 14874 7713 14942
rect 7265 14818 7275 14874
rect 7331 14818 7399 14874
rect 7455 14818 7523 14874
rect 7579 14818 7647 14874
rect 7703 14818 7713 14874
rect 7265 14750 7713 14818
rect 7265 14694 7275 14750
rect 7331 14694 7399 14750
rect 7455 14694 7523 14750
rect 7579 14694 7647 14750
rect 7703 14694 7713 14750
rect 7265 14626 7713 14694
rect 7265 14570 7275 14626
rect 7331 14570 7399 14626
rect 7455 14570 7523 14626
rect 7579 14570 7647 14626
rect 7703 14570 7713 14626
rect 7265 14502 7713 14570
rect 7265 14446 7275 14502
rect 7331 14446 7399 14502
rect 7455 14446 7523 14502
rect 7579 14446 7647 14502
rect 7703 14446 7713 14502
rect 7265 14436 7713 14446
rect 9927 17354 10127 17364
rect 9927 17298 9937 17354
rect 9993 17298 10061 17354
rect 10117 17298 10127 17354
rect 9927 17230 10127 17298
rect 9927 17174 9937 17230
rect 9993 17174 10061 17230
rect 10117 17174 10127 17230
rect 9927 17106 10127 17174
rect 9927 17050 9937 17106
rect 9993 17050 10061 17106
rect 10117 17050 10127 17106
rect 9927 16982 10127 17050
rect 9927 16926 9937 16982
rect 9993 16926 10061 16982
rect 10117 16926 10127 16982
rect 9927 16858 10127 16926
rect 9927 16802 9937 16858
rect 9993 16802 10061 16858
rect 10117 16802 10127 16858
rect 9927 16734 10127 16802
rect 9927 16678 9937 16734
rect 9993 16678 10061 16734
rect 10117 16678 10127 16734
rect 9927 16610 10127 16678
rect 9927 16554 9937 16610
rect 9993 16554 10061 16610
rect 10117 16554 10127 16610
rect 9927 16486 10127 16554
rect 9927 16430 9937 16486
rect 9993 16430 10061 16486
rect 10117 16430 10127 16486
rect 9927 16362 10127 16430
rect 9927 16306 9937 16362
rect 9993 16306 10061 16362
rect 10117 16306 10127 16362
rect 9927 16238 10127 16306
rect 9927 16182 9937 16238
rect 9993 16182 10061 16238
rect 10117 16182 10127 16238
rect 9927 16114 10127 16182
rect 9927 16058 9937 16114
rect 9993 16058 10061 16114
rect 10117 16058 10127 16114
rect 9927 15990 10127 16058
rect 9927 15934 9937 15990
rect 9993 15934 10061 15990
rect 10117 15934 10127 15990
rect 9927 15866 10127 15934
rect 9927 15810 9937 15866
rect 9993 15810 10061 15866
rect 10117 15810 10127 15866
rect 9927 15742 10127 15810
rect 9927 15686 9937 15742
rect 9993 15686 10061 15742
rect 10117 15686 10127 15742
rect 9927 15618 10127 15686
rect 9927 15562 9937 15618
rect 9993 15562 10061 15618
rect 10117 15562 10127 15618
rect 9927 15494 10127 15562
rect 9927 15438 9937 15494
rect 9993 15438 10061 15494
rect 10117 15438 10127 15494
rect 9927 15370 10127 15438
rect 9927 15314 9937 15370
rect 9993 15314 10061 15370
rect 10117 15314 10127 15370
rect 9927 15246 10127 15314
rect 9927 15190 9937 15246
rect 9993 15190 10061 15246
rect 10117 15190 10127 15246
rect 9927 15122 10127 15190
rect 9927 15066 9937 15122
rect 9993 15066 10061 15122
rect 10117 15066 10127 15122
rect 9927 14998 10127 15066
rect 9927 14942 9937 14998
rect 9993 14942 10061 14998
rect 10117 14942 10127 14998
rect 9927 14874 10127 14942
rect 9927 14818 9937 14874
rect 9993 14818 10061 14874
rect 10117 14818 10127 14874
rect 9927 14750 10127 14818
rect 9927 14694 9937 14750
rect 9993 14694 10061 14750
rect 10117 14694 10127 14750
rect 9927 14626 10127 14694
rect 9927 14570 9937 14626
rect 9993 14570 10061 14626
rect 10117 14570 10127 14626
rect 9927 14502 10127 14570
rect 9927 14446 9937 14502
rect 9993 14446 10061 14502
rect 10117 14446 10127 14502
rect 9927 14436 10127 14446
rect 12297 17354 12497 17364
rect 12297 17298 12307 17354
rect 12363 17298 12431 17354
rect 12487 17298 12497 17354
rect 12297 17230 12497 17298
rect 12297 17174 12307 17230
rect 12363 17174 12431 17230
rect 12487 17174 12497 17230
rect 12297 17106 12497 17174
rect 12297 17050 12307 17106
rect 12363 17050 12431 17106
rect 12487 17050 12497 17106
rect 12297 16982 12497 17050
rect 12297 16926 12307 16982
rect 12363 16926 12431 16982
rect 12487 16926 12497 16982
rect 12297 16858 12497 16926
rect 12297 16802 12307 16858
rect 12363 16802 12431 16858
rect 12487 16802 12497 16858
rect 12297 16734 12497 16802
rect 12297 16678 12307 16734
rect 12363 16678 12431 16734
rect 12487 16678 12497 16734
rect 12297 16610 12497 16678
rect 12297 16554 12307 16610
rect 12363 16554 12431 16610
rect 12487 16554 12497 16610
rect 12297 16486 12497 16554
rect 12297 16430 12307 16486
rect 12363 16430 12431 16486
rect 12487 16430 12497 16486
rect 12297 16362 12497 16430
rect 12297 16306 12307 16362
rect 12363 16306 12431 16362
rect 12487 16306 12497 16362
rect 12297 16238 12497 16306
rect 12297 16182 12307 16238
rect 12363 16182 12431 16238
rect 12487 16182 12497 16238
rect 12297 16114 12497 16182
rect 12297 16058 12307 16114
rect 12363 16058 12431 16114
rect 12487 16058 12497 16114
rect 12297 15990 12497 16058
rect 12297 15934 12307 15990
rect 12363 15934 12431 15990
rect 12487 15934 12497 15990
rect 12297 15866 12497 15934
rect 12297 15810 12307 15866
rect 12363 15810 12431 15866
rect 12487 15810 12497 15866
rect 12297 15742 12497 15810
rect 12297 15686 12307 15742
rect 12363 15686 12431 15742
rect 12487 15686 12497 15742
rect 12297 15618 12497 15686
rect 12297 15562 12307 15618
rect 12363 15562 12431 15618
rect 12487 15562 12497 15618
rect 12297 15494 12497 15562
rect 12297 15438 12307 15494
rect 12363 15438 12431 15494
rect 12487 15438 12497 15494
rect 12297 15370 12497 15438
rect 12297 15314 12307 15370
rect 12363 15314 12431 15370
rect 12487 15314 12497 15370
rect 12297 15246 12497 15314
rect 12297 15190 12307 15246
rect 12363 15190 12431 15246
rect 12487 15190 12497 15246
rect 12297 15122 12497 15190
rect 12297 15066 12307 15122
rect 12363 15066 12431 15122
rect 12487 15066 12497 15122
rect 12297 14998 12497 15066
rect 12297 14942 12307 14998
rect 12363 14942 12431 14998
rect 12487 14942 12497 14998
rect 12297 14874 12497 14942
rect 12297 14818 12307 14874
rect 12363 14818 12431 14874
rect 12487 14818 12497 14874
rect 12297 14750 12497 14818
rect 12297 14694 12307 14750
rect 12363 14694 12431 14750
rect 12487 14694 12497 14750
rect 12297 14626 12497 14694
rect 12297 14570 12307 14626
rect 12363 14570 12431 14626
rect 12487 14570 12497 14626
rect 12297 14502 12497 14570
rect 12297 14446 12307 14502
rect 12363 14446 12431 14502
rect 12487 14446 12497 14502
rect 12297 14436 12497 14446
rect 10 14176 86 14186
rect 10 12824 20 14176
rect 76 12824 86 14176
rect 14892 14176 14968 14186
rect 305 14148 2117 14158
rect 305 14092 315 14148
rect 371 14092 439 14148
rect 495 14092 563 14148
rect 619 14092 687 14148
rect 743 14092 811 14148
rect 867 14092 935 14148
rect 991 14092 1059 14148
rect 1115 14092 1183 14148
rect 1239 14092 1307 14148
rect 1363 14092 1431 14148
rect 1487 14092 1555 14148
rect 1611 14092 1679 14148
rect 1735 14092 1803 14148
rect 1859 14092 1927 14148
rect 1983 14092 2051 14148
rect 2107 14092 2117 14148
rect 305 14024 2117 14092
rect 305 13968 315 14024
rect 371 13968 439 14024
rect 495 13968 563 14024
rect 619 13968 687 14024
rect 743 13968 811 14024
rect 867 13968 935 14024
rect 991 13968 1059 14024
rect 1115 13968 1183 14024
rect 1239 13968 1307 14024
rect 1363 13968 1431 14024
rect 1487 13968 1555 14024
rect 1611 13968 1679 14024
rect 1735 13968 1803 14024
rect 1859 13968 1927 14024
rect 1983 13968 2051 14024
rect 2107 13968 2117 14024
rect 305 13900 2117 13968
rect 305 13844 315 13900
rect 371 13844 439 13900
rect 495 13844 563 13900
rect 619 13844 687 13900
rect 743 13844 811 13900
rect 867 13844 935 13900
rect 991 13844 1059 13900
rect 1115 13844 1183 13900
rect 1239 13844 1307 13900
rect 1363 13844 1431 13900
rect 1487 13844 1555 13900
rect 1611 13844 1679 13900
rect 1735 13844 1803 13900
rect 1859 13844 1927 13900
rect 1983 13844 2051 13900
rect 2107 13844 2117 13900
rect 305 13776 2117 13844
rect 305 13720 315 13776
rect 371 13720 439 13776
rect 495 13720 563 13776
rect 619 13720 687 13776
rect 743 13720 811 13776
rect 867 13720 935 13776
rect 991 13720 1059 13776
rect 1115 13720 1183 13776
rect 1239 13720 1307 13776
rect 1363 13720 1431 13776
rect 1487 13720 1555 13776
rect 1611 13720 1679 13776
rect 1735 13720 1803 13776
rect 1859 13720 1927 13776
rect 1983 13720 2051 13776
rect 2107 13720 2117 13776
rect 305 13652 2117 13720
rect 305 13596 315 13652
rect 371 13596 439 13652
rect 495 13596 563 13652
rect 619 13596 687 13652
rect 743 13596 811 13652
rect 867 13596 935 13652
rect 991 13596 1059 13652
rect 1115 13596 1183 13652
rect 1239 13596 1307 13652
rect 1363 13596 1431 13652
rect 1487 13596 1555 13652
rect 1611 13596 1679 13652
rect 1735 13596 1803 13652
rect 1859 13596 1927 13652
rect 1983 13596 2051 13652
rect 2107 13596 2117 13652
rect 305 13528 2117 13596
rect 305 13472 315 13528
rect 371 13472 439 13528
rect 495 13472 563 13528
rect 619 13472 687 13528
rect 743 13472 811 13528
rect 867 13472 935 13528
rect 991 13472 1059 13528
rect 1115 13472 1183 13528
rect 1239 13472 1307 13528
rect 1363 13472 1431 13528
rect 1487 13472 1555 13528
rect 1611 13472 1679 13528
rect 1735 13472 1803 13528
rect 1859 13472 1927 13528
rect 1983 13472 2051 13528
rect 2107 13472 2117 13528
rect 305 13404 2117 13472
rect 305 13348 315 13404
rect 371 13348 439 13404
rect 495 13348 563 13404
rect 619 13348 687 13404
rect 743 13348 811 13404
rect 867 13348 935 13404
rect 991 13348 1059 13404
rect 1115 13348 1183 13404
rect 1239 13348 1307 13404
rect 1363 13348 1431 13404
rect 1487 13348 1555 13404
rect 1611 13348 1679 13404
rect 1735 13348 1803 13404
rect 1859 13348 1927 13404
rect 1983 13348 2051 13404
rect 2107 13348 2117 13404
rect 305 13280 2117 13348
rect 305 13224 315 13280
rect 371 13224 439 13280
rect 495 13224 563 13280
rect 619 13224 687 13280
rect 743 13224 811 13280
rect 867 13224 935 13280
rect 991 13224 1059 13280
rect 1115 13224 1183 13280
rect 1239 13224 1307 13280
rect 1363 13224 1431 13280
rect 1487 13224 1555 13280
rect 1611 13224 1679 13280
rect 1735 13224 1803 13280
rect 1859 13224 1927 13280
rect 1983 13224 2051 13280
rect 2107 13224 2117 13280
rect 305 13156 2117 13224
rect 305 13100 315 13156
rect 371 13100 439 13156
rect 495 13100 563 13156
rect 619 13100 687 13156
rect 743 13100 811 13156
rect 867 13100 935 13156
rect 991 13100 1059 13156
rect 1115 13100 1183 13156
rect 1239 13100 1307 13156
rect 1363 13100 1431 13156
rect 1487 13100 1555 13156
rect 1611 13100 1679 13156
rect 1735 13100 1803 13156
rect 1859 13100 1927 13156
rect 1983 13100 2051 13156
rect 2107 13100 2117 13156
rect 305 13032 2117 13100
rect 305 12976 315 13032
rect 371 12976 439 13032
rect 495 12976 563 13032
rect 619 12976 687 13032
rect 743 12976 811 13032
rect 867 12976 935 13032
rect 991 12976 1059 13032
rect 1115 12976 1183 13032
rect 1239 12976 1307 13032
rect 1363 12976 1431 13032
rect 1487 12976 1555 13032
rect 1611 12976 1679 13032
rect 1735 12976 1803 13032
rect 1859 12976 1927 13032
rect 1983 12976 2051 13032
rect 2107 12976 2117 13032
rect 305 12908 2117 12976
rect 305 12852 315 12908
rect 371 12852 439 12908
rect 495 12852 563 12908
rect 619 12852 687 12908
rect 743 12852 811 12908
rect 867 12852 935 12908
rect 991 12852 1059 12908
rect 1115 12852 1183 12908
rect 1239 12852 1307 12908
rect 1363 12852 1431 12908
rect 1487 12852 1555 12908
rect 1611 12852 1679 12908
rect 1735 12852 1803 12908
rect 1859 12852 1927 12908
rect 1983 12852 2051 12908
rect 2107 12852 2117 12908
rect 305 12842 2117 12852
rect 2798 14148 4734 14158
rect 2798 14092 2808 14148
rect 2864 14092 2932 14148
rect 2988 14092 3056 14148
rect 3112 14092 3180 14148
rect 3236 14092 3304 14148
rect 3360 14092 3428 14148
rect 3484 14092 3552 14148
rect 3608 14092 3676 14148
rect 3732 14092 3800 14148
rect 3856 14092 3924 14148
rect 3980 14092 4048 14148
rect 4104 14092 4172 14148
rect 4228 14092 4296 14148
rect 4352 14092 4420 14148
rect 4476 14092 4544 14148
rect 4600 14092 4668 14148
rect 4724 14092 4734 14148
rect 2798 14024 4734 14092
rect 2798 13968 2808 14024
rect 2864 13968 2932 14024
rect 2988 13968 3056 14024
rect 3112 13968 3180 14024
rect 3236 13968 3304 14024
rect 3360 13968 3428 14024
rect 3484 13968 3552 14024
rect 3608 13968 3676 14024
rect 3732 13968 3800 14024
rect 3856 13968 3924 14024
rect 3980 13968 4048 14024
rect 4104 13968 4172 14024
rect 4228 13968 4296 14024
rect 4352 13968 4420 14024
rect 4476 13968 4544 14024
rect 4600 13968 4668 14024
rect 4724 13968 4734 14024
rect 2798 13900 4734 13968
rect 2798 13844 2808 13900
rect 2864 13844 2932 13900
rect 2988 13844 3056 13900
rect 3112 13844 3180 13900
rect 3236 13844 3304 13900
rect 3360 13844 3428 13900
rect 3484 13844 3552 13900
rect 3608 13844 3676 13900
rect 3732 13844 3800 13900
rect 3856 13844 3924 13900
rect 3980 13844 4048 13900
rect 4104 13844 4172 13900
rect 4228 13844 4296 13900
rect 4352 13844 4420 13900
rect 4476 13844 4544 13900
rect 4600 13844 4668 13900
rect 4724 13844 4734 13900
rect 2798 13776 4734 13844
rect 2798 13720 2808 13776
rect 2864 13720 2932 13776
rect 2988 13720 3056 13776
rect 3112 13720 3180 13776
rect 3236 13720 3304 13776
rect 3360 13720 3428 13776
rect 3484 13720 3552 13776
rect 3608 13720 3676 13776
rect 3732 13720 3800 13776
rect 3856 13720 3924 13776
rect 3980 13720 4048 13776
rect 4104 13720 4172 13776
rect 4228 13720 4296 13776
rect 4352 13720 4420 13776
rect 4476 13720 4544 13776
rect 4600 13720 4668 13776
rect 4724 13720 4734 13776
rect 2798 13652 4734 13720
rect 2798 13596 2808 13652
rect 2864 13596 2932 13652
rect 2988 13596 3056 13652
rect 3112 13596 3180 13652
rect 3236 13596 3304 13652
rect 3360 13596 3428 13652
rect 3484 13596 3552 13652
rect 3608 13596 3676 13652
rect 3732 13596 3800 13652
rect 3856 13596 3924 13652
rect 3980 13596 4048 13652
rect 4104 13596 4172 13652
rect 4228 13596 4296 13652
rect 4352 13596 4420 13652
rect 4476 13596 4544 13652
rect 4600 13596 4668 13652
rect 4724 13596 4734 13652
rect 2798 13528 4734 13596
rect 2798 13472 2808 13528
rect 2864 13472 2932 13528
rect 2988 13472 3056 13528
rect 3112 13472 3180 13528
rect 3236 13472 3304 13528
rect 3360 13472 3428 13528
rect 3484 13472 3552 13528
rect 3608 13472 3676 13528
rect 3732 13472 3800 13528
rect 3856 13472 3924 13528
rect 3980 13472 4048 13528
rect 4104 13472 4172 13528
rect 4228 13472 4296 13528
rect 4352 13472 4420 13528
rect 4476 13472 4544 13528
rect 4600 13472 4668 13528
rect 4724 13472 4734 13528
rect 2798 13404 4734 13472
rect 2798 13348 2808 13404
rect 2864 13348 2932 13404
rect 2988 13348 3056 13404
rect 3112 13348 3180 13404
rect 3236 13348 3304 13404
rect 3360 13348 3428 13404
rect 3484 13348 3552 13404
rect 3608 13348 3676 13404
rect 3732 13348 3800 13404
rect 3856 13348 3924 13404
rect 3980 13348 4048 13404
rect 4104 13348 4172 13404
rect 4228 13348 4296 13404
rect 4352 13348 4420 13404
rect 4476 13348 4544 13404
rect 4600 13348 4668 13404
rect 4724 13348 4734 13404
rect 2798 13280 4734 13348
rect 2798 13224 2808 13280
rect 2864 13224 2932 13280
rect 2988 13224 3056 13280
rect 3112 13224 3180 13280
rect 3236 13224 3304 13280
rect 3360 13224 3428 13280
rect 3484 13224 3552 13280
rect 3608 13224 3676 13280
rect 3732 13224 3800 13280
rect 3856 13224 3924 13280
rect 3980 13224 4048 13280
rect 4104 13224 4172 13280
rect 4228 13224 4296 13280
rect 4352 13224 4420 13280
rect 4476 13224 4544 13280
rect 4600 13224 4668 13280
rect 4724 13224 4734 13280
rect 2798 13156 4734 13224
rect 2798 13100 2808 13156
rect 2864 13100 2932 13156
rect 2988 13100 3056 13156
rect 3112 13100 3180 13156
rect 3236 13100 3304 13156
rect 3360 13100 3428 13156
rect 3484 13100 3552 13156
rect 3608 13100 3676 13156
rect 3732 13100 3800 13156
rect 3856 13100 3924 13156
rect 3980 13100 4048 13156
rect 4104 13100 4172 13156
rect 4228 13100 4296 13156
rect 4352 13100 4420 13156
rect 4476 13100 4544 13156
rect 4600 13100 4668 13156
rect 4724 13100 4734 13156
rect 2798 13032 4734 13100
rect 2798 12976 2808 13032
rect 2864 12976 2932 13032
rect 2988 12976 3056 13032
rect 3112 12976 3180 13032
rect 3236 12976 3304 13032
rect 3360 12976 3428 13032
rect 3484 12976 3552 13032
rect 3608 12976 3676 13032
rect 3732 12976 3800 13032
rect 3856 12976 3924 13032
rect 3980 12976 4048 13032
rect 4104 12976 4172 13032
rect 4228 12976 4296 13032
rect 4352 12976 4420 13032
rect 4476 12976 4544 13032
rect 4600 12976 4668 13032
rect 4724 12976 4734 13032
rect 2798 12908 4734 12976
rect 2798 12852 2808 12908
rect 2864 12852 2932 12908
rect 2988 12852 3056 12908
rect 3112 12852 3180 12908
rect 3236 12852 3304 12908
rect 3360 12852 3428 12908
rect 3484 12852 3552 12908
rect 3608 12852 3676 12908
rect 3732 12852 3800 12908
rect 3856 12852 3924 12908
rect 3980 12852 4048 12908
rect 4104 12852 4172 12908
rect 4228 12852 4296 12908
rect 4352 12852 4420 12908
rect 4476 12852 4544 12908
rect 4600 12852 4668 12908
rect 4724 12852 4734 12908
rect 2798 12842 4734 12852
rect 5168 14148 7104 14158
rect 5168 14092 5178 14148
rect 5234 14092 5302 14148
rect 5358 14092 5426 14148
rect 5482 14092 5550 14148
rect 5606 14092 5674 14148
rect 5730 14092 5798 14148
rect 5854 14092 5922 14148
rect 5978 14092 6046 14148
rect 6102 14092 6170 14148
rect 6226 14092 6294 14148
rect 6350 14092 6418 14148
rect 6474 14092 6542 14148
rect 6598 14092 6666 14148
rect 6722 14092 6790 14148
rect 6846 14092 6914 14148
rect 6970 14092 7038 14148
rect 7094 14092 7104 14148
rect 5168 14024 7104 14092
rect 5168 13968 5178 14024
rect 5234 13968 5302 14024
rect 5358 13968 5426 14024
rect 5482 13968 5550 14024
rect 5606 13968 5674 14024
rect 5730 13968 5798 14024
rect 5854 13968 5922 14024
rect 5978 13968 6046 14024
rect 6102 13968 6170 14024
rect 6226 13968 6294 14024
rect 6350 13968 6418 14024
rect 6474 13968 6542 14024
rect 6598 13968 6666 14024
rect 6722 13968 6790 14024
rect 6846 13968 6914 14024
rect 6970 13968 7038 14024
rect 7094 13968 7104 14024
rect 5168 13900 7104 13968
rect 5168 13844 5178 13900
rect 5234 13844 5302 13900
rect 5358 13844 5426 13900
rect 5482 13844 5550 13900
rect 5606 13844 5674 13900
rect 5730 13844 5798 13900
rect 5854 13844 5922 13900
rect 5978 13844 6046 13900
rect 6102 13844 6170 13900
rect 6226 13844 6294 13900
rect 6350 13844 6418 13900
rect 6474 13844 6542 13900
rect 6598 13844 6666 13900
rect 6722 13844 6790 13900
rect 6846 13844 6914 13900
rect 6970 13844 7038 13900
rect 7094 13844 7104 13900
rect 5168 13776 7104 13844
rect 5168 13720 5178 13776
rect 5234 13720 5302 13776
rect 5358 13720 5426 13776
rect 5482 13720 5550 13776
rect 5606 13720 5674 13776
rect 5730 13720 5798 13776
rect 5854 13720 5922 13776
rect 5978 13720 6046 13776
rect 6102 13720 6170 13776
rect 6226 13720 6294 13776
rect 6350 13720 6418 13776
rect 6474 13720 6542 13776
rect 6598 13720 6666 13776
rect 6722 13720 6790 13776
rect 6846 13720 6914 13776
rect 6970 13720 7038 13776
rect 7094 13720 7104 13776
rect 5168 13652 7104 13720
rect 5168 13596 5178 13652
rect 5234 13596 5302 13652
rect 5358 13596 5426 13652
rect 5482 13596 5550 13652
rect 5606 13596 5674 13652
rect 5730 13596 5798 13652
rect 5854 13596 5922 13652
rect 5978 13596 6046 13652
rect 6102 13596 6170 13652
rect 6226 13596 6294 13652
rect 6350 13596 6418 13652
rect 6474 13596 6542 13652
rect 6598 13596 6666 13652
rect 6722 13596 6790 13652
rect 6846 13596 6914 13652
rect 6970 13596 7038 13652
rect 7094 13596 7104 13652
rect 5168 13528 7104 13596
rect 5168 13472 5178 13528
rect 5234 13472 5302 13528
rect 5358 13472 5426 13528
rect 5482 13472 5550 13528
rect 5606 13472 5674 13528
rect 5730 13472 5798 13528
rect 5854 13472 5922 13528
rect 5978 13472 6046 13528
rect 6102 13472 6170 13528
rect 6226 13472 6294 13528
rect 6350 13472 6418 13528
rect 6474 13472 6542 13528
rect 6598 13472 6666 13528
rect 6722 13472 6790 13528
rect 6846 13472 6914 13528
rect 6970 13472 7038 13528
rect 7094 13472 7104 13528
rect 5168 13404 7104 13472
rect 5168 13348 5178 13404
rect 5234 13348 5302 13404
rect 5358 13348 5426 13404
rect 5482 13348 5550 13404
rect 5606 13348 5674 13404
rect 5730 13348 5798 13404
rect 5854 13348 5922 13404
rect 5978 13348 6046 13404
rect 6102 13348 6170 13404
rect 6226 13348 6294 13404
rect 6350 13348 6418 13404
rect 6474 13348 6542 13404
rect 6598 13348 6666 13404
rect 6722 13348 6790 13404
rect 6846 13348 6914 13404
rect 6970 13348 7038 13404
rect 7094 13348 7104 13404
rect 5168 13280 7104 13348
rect 5168 13224 5178 13280
rect 5234 13224 5302 13280
rect 5358 13224 5426 13280
rect 5482 13224 5550 13280
rect 5606 13224 5674 13280
rect 5730 13224 5798 13280
rect 5854 13224 5922 13280
rect 5978 13224 6046 13280
rect 6102 13224 6170 13280
rect 6226 13224 6294 13280
rect 6350 13224 6418 13280
rect 6474 13224 6542 13280
rect 6598 13224 6666 13280
rect 6722 13224 6790 13280
rect 6846 13224 6914 13280
rect 6970 13224 7038 13280
rect 7094 13224 7104 13280
rect 5168 13156 7104 13224
rect 5168 13100 5178 13156
rect 5234 13100 5302 13156
rect 5358 13100 5426 13156
rect 5482 13100 5550 13156
rect 5606 13100 5674 13156
rect 5730 13100 5798 13156
rect 5854 13100 5922 13156
rect 5978 13100 6046 13156
rect 6102 13100 6170 13156
rect 6226 13100 6294 13156
rect 6350 13100 6418 13156
rect 6474 13100 6542 13156
rect 6598 13100 6666 13156
rect 6722 13100 6790 13156
rect 6846 13100 6914 13156
rect 6970 13100 7038 13156
rect 7094 13100 7104 13156
rect 5168 13032 7104 13100
rect 5168 12976 5178 13032
rect 5234 12976 5302 13032
rect 5358 12976 5426 13032
rect 5482 12976 5550 13032
rect 5606 12976 5674 13032
rect 5730 12976 5798 13032
rect 5854 12976 5922 13032
rect 5978 12976 6046 13032
rect 6102 12976 6170 13032
rect 6226 12976 6294 13032
rect 6350 12976 6418 13032
rect 6474 12976 6542 13032
rect 6598 12976 6666 13032
rect 6722 12976 6790 13032
rect 6846 12976 6914 13032
rect 6970 12976 7038 13032
rect 7094 12976 7104 13032
rect 5168 12908 7104 12976
rect 5168 12852 5178 12908
rect 5234 12852 5302 12908
rect 5358 12852 5426 12908
rect 5482 12852 5550 12908
rect 5606 12852 5674 12908
rect 5730 12852 5798 12908
rect 5854 12852 5922 12908
rect 5978 12852 6046 12908
rect 6102 12852 6170 12908
rect 6226 12852 6294 12908
rect 6350 12852 6418 12908
rect 6474 12852 6542 12908
rect 6598 12852 6666 12908
rect 6722 12852 6790 12908
rect 6846 12852 6914 12908
rect 6970 12852 7038 12908
rect 7094 12852 7104 12908
rect 5168 12842 7104 12852
rect 7874 14148 9810 14158
rect 7874 14092 7884 14148
rect 7940 14092 8008 14148
rect 8064 14092 8132 14148
rect 8188 14092 8256 14148
rect 8312 14092 8380 14148
rect 8436 14092 8504 14148
rect 8560 14092 8628 14148
rect 8684 14092 8752 14148
rect 8808 14092 8876 14148
rect 8932 14092 9000 14148
rect 9056 14092 9124 14148
rect 9180 14092 9248 14148
rect 9304 14092 9372 14148
rect 9428 14092 9496 14148
rect 9552 14092 9620 14148
rect 9676 14092 9744 14148
rect 9800 14092 9810 14148
rect 7874 14024 9810 14092
rect 7874 13968 7884 14024
rect 7940 13968 8008 14024
rect 8064 13968 8132 14024
rect 8188 13968 8256 14024
rect 8312 13968 8380 14024
rect 8436 13968 8504 14024
rect 8560 13968 8628 14024
rect 8684 13968 8752 14024
rect 8808 13968 8876 14024
rect 8932 13968 9000 14024
rect 9056 13968 9124 14024
rect 9180 13968 9248 14024
rect 9304 13968 9372 14024
rect 9428 13968 9496 14024
rect 9552 13968 9620 14024
rect 9676 13968 9744 14024
rect 9800 13968 9810 14024
rect 7874 13900 9810 13968
rect 7874 13844 7884 13900
rect 7940 13844 8008 13900
rect 8064 13844 8132 13900
rect 8188 13844 8256 13900
rect 8312 13844 8380 13900
rect 8436 13844 8504 13900
rect 8560 13844 8628 13900
rect 8684 13844 8752 13900
rect 8808 13844 8876 13900
rect 8932 13844 9000 13900
rect 9056 13844 9124 13900
rect 9180 13844 9248 13900
rect 9304 13844 9372 13900
rect 9428 13844 9496 13900
rect 9552 13844 9620 13900
rect 9676 13844 9744 13900
rect 9800 13844 9810 13900
rect 7874 13776 9810 13844
rect 7874 13720 7884 13776
rect 7940 13720 8008 13776
rect 8064 13720 8132 13776
rect 8188 13720 8256 13776
rect 8312 13720 8380 13776
rect 8436 13720 8504 13776
rect 8560 13720 8628 13776
rect 8684 13720 8752 13776
rect 8808 13720 8876 13776
rect 8932 13720 9000 13776
rect 9056 13720 9124 13776
rect 9180 13720 9248 13776
rect 9304 13720 9372 13776
rect 9428 13720 9496 13776
rect 9552 13720 9620 13776
rect 9676 13720 9744 13776
rect 9800 13720 9810 13776
rect 7874 13652 9810 13720
rect 7874 13596 7884 13652
rect 7940 13596 8008 13652
rect 8064 13596 8132 13652
rect 8188 13596 8256 13652
rect 8312 13596 8380 13652
rect 8436 13596 8504 13652
rect 8560 13596 8628 13652
rect 8684 13596 8752 13652
rect 8808 13596 8876 13652
rect 8932 13596 9000 13652
rect 9056 13596 9124 13652
rect 9180 13596 9248 13652
rect 9304 13596 9372 13652
rect 9428 13596 9496 13652
rect 9552 13596 9620 13652
rect 9676 13596 9744 13652
rect 9800 13596 9810 13652
rect 7874 13528 9810 13596
rect 7874 13472 7884 13528
rect 7940 13472 8008 13528
rect 8064 13472 8132 13528
rect 8188 13472 8256 13528
rect 8312 13472 8380 13528
rect 8436 13472 8504 13528
rect 8560 13472 8628 13528
rect 8684 13472 8752 13528
rect 8808 13472 8876 13528
rect 8932 13472 9000 13528
rect 9056 13472 9124 13528
rect 9180 13472 9248 13528
rect 9304 13472 9372 13528
rect 9428 13472 9496 13528
rect 9552 13472 9620 13528
rect 9676 13472 9744 13528
rect 9800 13472 9810 13528
rect 7874 13404 9810 13472
rect 7874 13348 7884 13404
rect 7940 13348 8008 13404
rect 8064 13348 8132 13404
rect 8188 13348 8256 13404
rect 8312 13348 8380 13404
rect 8436 13348 8504 13404
rect 8560 13348 8628 13404
rect 8684 13348 8752 13404
rect 8808 13348 8876 13404
rect 8932 13348 9000 13404
rect 9056 13348 9124 13404
rect 9180 13348 9248 13404
rect 9304 13348 9372 13404
rect 9428 13348 9496 13404
rect 9552 13348 9620 13404
rect 9676 13348 9744 13404
rect 9800 13348 9810 13404
rect 7874 13280 9810 13348
rect 7874 13224 7884 13280
rect 7940 13224 8008 13280
rect 8064 13224 8132 13280
rect 8188 13224 8256 13280
rect 8312 13224 8380 13280
rect 8436 13224 8504 13280
rect 8560 13224 8628 13280
rect 8684 13224 8752 13280
rect 8808 13224 8876 13280
rect 8932 13224 9000 13280
rect 9056 13224 9124 13280
rect 9180 13224 9248 13280
rect 9304 13224 9372 13280
rect 9428 13224 9496 13280
rect 9552 13224 9620 13280
rect 9676 13224 9744 13280
rect 9800 13224 9810 13280
rect 7874 13156 9810 13224
rect 7874 13100 7884 13156
rect 7940 13100 8008 13156
rect 8064 13100 8132 13156
rect 8188 13100 8256 13156
rect 8312 13100 8380 13156
rect 8436 13100 8504 13156
rect 8560 13100 8628 13156
rect 8684 13100 8752 13156
rect 8808 13100 8876 13156
rect 8932 13100 9000 13156
rect 9056 13100 9124 13156
rect 9180 13100 9248 13156
rect 9304 13100 9372 13156
rect 9428 13100 9496 13156
rect 9552 13100 9620 13156
rect 9676 13100 9744 13156
rect 9800 13100 9810 13156
rect 7874 13032 9810 13100
rect 7874 12976 7884 13032
rect 7940 12976 8008 13032
rect 8064 12976 8132 13032
rect 8188 12976 8256 13032
rect 8312 12976 8380 13032
rect 8436 12976 8504 13032
rect 8560 12976 8628 13032
rect 8684 12976 8752 13032
rect 8808 12976 8876 13032
rect 8932 12976 9000 13032
rect 9056 12976 9124 13032
rect 9180 12976 9248 13032
rect 9304 12976 9372 13032
rect 9428 12976 9496 13032
rect 9552 12976 9620 13032
rect 9676 12976 9744 13032
rect 9800 12976 9810 13032
rect 7874 12908 9810 12976
rect 7874 12852 7884 12908
rect 7940 12852 8008 12908
rect 8064 12852 8132 12908
rect 8188 12852 8256 12908
rect 8312 12852 8380 12908
rect 8436 12852 8504 12908
rect 8560 12852 8628 12908
rect 8684 12852 8752 12908
rect 8808 12852 8876 12908
rect 8932 12852 9000 12908
rect 9056 12852 9124 12908
rect 9180 12852 9248 12908
rect 9304 12852 9372 12908
rect 9428 12852 9496 12908
rect 9552 12852 9620 12908
rect 9676 12852 9744 12908
rect 9800 12852 9810 12908
rect 7874 12842 9810 12852
rect 10244 14148 12180 14158
rect 10244 14092 10254 14148
rect 10310 14092 10378 14148
rect 10434 14092 10502 14148
rect 10558 14092 10626 14148
rect 10682 14092 10750 14148
rect 10806 14092 10874 14148
rect 10930 14092 10998 14148
rect 11054 14092 11122 14148
rect 11178 14092 11246 14148
rect 11302 14092 11370 14148
rect 11426 14092 11494 14148
rect 11550 14092 11618 14148
rect 11674 14092 11742 14148
rect 11798 14092 11866 14148
rect 11922 14092 11990 14148
rect 12046 14092 12114 14148
rect 12170 14092 12180 14148
rect 10244 14024 12180 14092
rect 10244 13968 10254 14024
rect 10310 13968 10378 14024
rect 10434 13968 10502 14024
rect 10558 13968 10626 14024
rect 10682 13968 10750 14024
rect 10806 13968 10874 14024
rect 10930 13968 10998 14024
rect 11054 13968 11122 14024
rect 11178 13968 11246 14024
rect 11302 13968 11370 14024
rect 11426 13968 11494 14024
rect 11550 13968 11618 14024
rect 11674 13968 11742 14024
rect 11798 13968 11866 14024
rect 11922 13968 11990 14024
rect 12046 13968 12114 14024
rect 12170 13968 12180 14024
rect 10244 13900 12180 13968
rect 10244 13844 10254 13900
rect 10310 13844 10378 13900
rect 10434 13844 10502 13900
rect 10558 13844 10626 13900
rect 10682 13844 10750 13900
rect 10806 13844 10874 13900
rect 10930 13844 10998 13900
rect 11054 13844 11122 13900
rect 11178 13844 11246 13900
rect 11302 13844 11370 13900
rect 11426 13844 11494 13900
rect 11550 13844 11618 13900
rect 11674 13844 11742 13900
rect 11798 13844 11866 13900
rect 11922 13844 11990 13900
rect 12046 13844 12114 13900
rect 12170 13844 12180 13900
rect 10244 13776 12180 13844
rect 10244 13720 10254 13776
rect 10310 13720 10378 13776
rect 10434 13720 10502 13776
rect 10558 13720 10626 13776
rect 10682 13720 10750 13776
rect 10806 13720 10874 13776
rect 10930 13720 10998 13776
rect 11054 13720 11122 13776
rect 11178 13720 11246 13776
rect 11302 13720 11370 13776
rect 11426 13720 11494 13776
rect 11550 13720 11618 13776
rect 11674 13720 11742 13776
rect 11798 13720 11866 13776
rect 11922 13720 11990 13776
rect 12046 13720 12114 13776
rect 12170 13720 12180 13776
rect 10244 13652 12180 13720
rect 10244 13596 10254 13652
rect 10310 13596 10378 13652
rect 10434 13596 10502 13652
rect 10558 13596 10626 13652
rect 10682 13596 10750 13652
rect 10806 13596 10874 13652
rect 10930 13596 10998 13652
rect 11054 13596 11122 13652
rect 11178 13596 11246 13652
rect 11302 13596 11370 13652
rect 11426 13596 11494 13652
rect 11550 13596 11618 13652
rect 11674 13596 11742 13652
rect 11798 13596 11866 13652
rect 11922 13596 11990 13652
rect 12046 13596 12114 13652
rect 12170 13596 12180 13652
rect 10244 13528 12180 13596
rect 10244 13472 10254 13528
rect 10310 13472 10378 13528
rect 10434 13472 10502 13528
rect 10558 13472 10626 13528
rect 10682 13472 10750 13528
rect 10806 13472 10874 13528
rect 10930 13472 10998 13528
rect 11054 13472 11122 13528
rect 11178 13472 11246 13528
rect 11302 13472 11370 13528
rect 11426 13472 11494 13528
rect 11550 13472 11618 13528
rect 11674 13472 11742 13528
rect 11798 13472 11866 13528
rect 11922 13472 11990 13528
rect 12046 13472 12114 13528
rect 12170 13472 12180 13528
rect 10244 13404 12180 13472
rect 10244 13348 10254 13404
rect 10310 13348 10378 13404
rect 10434 13348 10502 13404
rect 10558 13348 10626 13404
rect 10682 13348 10750 13404
rect 10806 13348 10874 13404
rect 10930 13348 10998 13404
rect 11054 13348 11122 13404
rect 11178 13348 11246 13404
rect 11302 13348 11370 13404
rect 11426 13348 11494 13404
rect 11550 13348 11618 13404
rect 11674 13348 11742 13404
rect 11798 13348 11866 13404
rect 11922 13348 11990 13404
rect 12046 13348 12114 13404
rect 12170 13348 12180 13404
rect 10244 13280 12180 13348
rect 10244 13224 10254 13280
rect 10310 13224 10378 13280
rect 10434 13224 10502 13280
rect 10558 13224 10626 13280
rect 10682 13224 10750 13280
rect 10806 13224 10874 13280
rect 10930 13224 10998 13280
rect 11054 13224 11122 13280
rect 11178 13224 11246 13280
rect 11302 13224 11370 13280
rect 11426 13224 11494 13280
rect 11550 13224 11618 13280
rect 11674 13224 11742 13280
rect 11798 13224 11866 13280
rect 11922 13224 11990 13280
rect 12046 13224 12114 13280
rect 12170 13224 12180 13280
rect 10244 13156 12180 13224
rect 10244 13100 10254 13156
rect 10310 13100 10378 13156
rect 10434 13100 10502 13156
rect 10558 13100 10626 13156
rect 10682 13100 10750 13156
rect 10806 13100 10874 13156
rect 10930 13100 10998 13156
rect 11054 13100 11122 13156
rect 11178 13100 11246 13156
rect 11302 13100 11370 13156
rect 11426 13100 11494 13156
rect 11550 13100 11618 13156
rect 11674 13100 11742 13156
rect 11798 13100 11866 13156
rect 11922 13100 11990 13156
rect 12046 13100 12114 13156
rect 12170 13100 12180 13156
rect 10244 13032 12180 13100
rect 10244 12976 10254 13032
rect 10310 12976 10378 13032
rect 10434 12976 10502 13032
rect 10558 12976 10626 13032
rect 10682 12976 10750 13032
rect 10806 12976 10874 13032
rect 10930 12976 10998 13032
rect 11054 12976 11122 13032
rect 11178 12976 11246 13032
rect 11302 12976 11370 13032
rect 11426 12976 11494 13032
rect 11550 12976 11618 13032
rect 11674 12976 11742 13032
rect 11798 12976 11866 13032
rect 11922 12976 11990 13032
rect 12046 12976 12114 13032
rect 12170 12976 12180 13032
rect 10244 12908 12180 12976
rect 10244 12852 10254 12908
rect 10310 12852 10378 12908
rect 10434 12852 10502 12908
rect 10558 12852 10626 12908
rect 10682 12852 10750 12908
rect 10806 12852 10874 12908
rect 10930 12852 10998 12908
rect 11054 12852 11122 12908
rect 11178 12852 11246 12908
rect 11302 12852 11370 12908
rect 11426 12852 11494 12908
rect 11550 12852 11618 12908
rect 11674 12852 11742 12908
rect 11798 12852 11866 12908
rect 11922 12852 11990 12908
rect 12046 12852 12114 12908
rect 12170 12852 12180 12908
rect 10244 12842 12180 12852
rect 12861 14148 14673 14158
rect 12861 14092 12871 14148
rect 12927 14092 12995 14148
rect 13051 14092 13119 14148
rect 13175 14092 13243 14148
rect 13299 14092 13367 14148
rect 13423 14092 13491 14148
rect 13547 14092 13615 14148
rect 13671 14092 13739 14148
rect 13795 14092 13863 14148
rect 13919 14092 13987 14148
rect 14043 14092 14111 14148
rect 14167 14092 14235 14148
rect 14291 14092 14359 14148
rect 14415 14092 14483 14148
rect 14539 14092 14607 14148
rect 14663 14092 14673 14148
rect 12861 14024 14673 14092
rect 12861 13968 12871 14024
rect 12927 13968 12995 14024
rect 13051 13968 13119 14024
rect 13175 13968 13243 14024
rect 13299 13968 13367 14024
rect 13423 13968 13491 14024
rect 13547 13968 13615 14024
rect 13671 13968 13739 14024
rect 13795 13968 13863 14024
rect 13919 13968 13987 14024
rect 14043 13968 14111 14024
rect 14167 13968 14235 14024
rect 14291 13968 14359 14024
rect 14415 13968 14483 14024
rect 14539 13968 14607 14024
rect 14663 13968 14673 14024
rect 12861 13900 14673 13968
rect 12861 13844 12871 13900
rect 12927 13844 12995 13900
rect 13051 13844 13119 13900
rect 13175 13844 13243 13900
rect 13299 13844 13367 13900
rect 13423 13844 13491 13900
rect 13547 13844 13615 13900
rect 13671 13844 13739 13900
rect 13795 13844 13863 13900
rect 13919 13844 13987 13900
rect 14043 13844 14111 13900
rect 14167 13844 14235 13900
rect 14291 13844 14359 13900
rect 14415 13844 14483 13900
rect 14539 13844 14607 13900
rect 14663 13844 14673 13900
rect 12861 13776 14673 13844
rect 12861 13720 12871 13776
rect 12927 13720 12995 13776
rect 13051 13720 13119 13776
rect 13175 13720 13243 13776
rect 13299 13720 13367 13776
rect 13423 13720 13491 13776
rect 13547 13720 13615 13776
rect 13671 13720 13739 13776
rect 13795 13720 13863 13776
rect 13919 13720 13987 13776
rect 14043 13720 14111 13776
rect 14167 13720 14235 13776
rect 14291 13720 14359 13776
rect 14415 13720 14483 13776
rect 14539 13720 14607 13776
rect 14663 13720 14673 13776
rect 12861 13652 14673 13720
rect 12861 13596 12871 13652
rect 12927 13596 12995 13652
rect 13051 13596 13119 13652
rect 13175 13596 13243 13652
rect 13299 13596 13367 13652
rect 13423 13596 13491 13652
rect 13547 13596 13615 13652
rect 13671 13596 13739 13652
rect 13795 13596 13863 13652
rect 13919 13596 13987 13652
rect 14043 13596 14111 13652
rect 14167 13596 14235 13652
rect 14291 13596 14359 13652
rect 14415 13596 14483 13652
rect 14539 13596 14607 13652
rect 14663 13596 14673 13652
rect 12861 13528 14673 13596
rect 12861 13472 12871 13528
rect 12927 13472 12995 13528
rect 13051 13472 13119 13528
rect 13175 13472 13243 13528
rect 13299 13472 13367 13528
rect 13423 13472 13491 13528
rect 13547 13472 13615 13528
rect 13671 13472 13739 13528
rect 13795 13472 13863 13528
rect 13919 13472 13987 13528
rect 14043 13472 14111 13528
rect 14167 13472 14235 13528
rect 14291 13472 14359 13528
rect 14415 13472 14483 13528
rect 14539 13472 14607 13528
rect 14663 13472 14673 13528
rect 12861 13404 14673 13472
rect 12861 13348 12871 13404
rect 12927 13348 12995 13404
rect 13051 13348 13119 13404
rect 13175 13348 13243 13404
rect 13299 13348 13367 13404
rect 13423 13348 13491 13404
rect 13547 13348 13615 13404
rect 13671 13348 13739 13404
rect 13795 13348 13863 13404
rect 13919 13348 13987 13404
rect 14043 13348 14111 13404
rect 14167 13348 14235 13404
rect 14291 13348 14359 13404
rect 14415 13348 14483 13404
rect 14539 13348 14607 13404
rect 14663 13348 14673 13404
rect 12861 13280 14673 13348
rect 12861 13224 12871 13280
rect 12927 13224 12995 13280
rect 13051 13224 13119 13280
rect 13175 13224 13243 13280
rect 13299 13224 13367 13280
rect 13423 13224 13491 13280
rect 13547 13224 13615 13280
rect 13671 13224 13739 13280
rect 13795 13224 13863 13280
rect 13919 13224 13987 13280
rect 14043 13224 14111 13280
rect 14167 13224 14235 13280
rect 14291 13224 14359 13280
rect 14415 13224 14483 13280
rect 14539 13224 14607 13280
rect 14663 13224 14673 13280
rect 12861 13156 14673 13224
rect 12861 13100 12871 13156
rect 12927 13100 12995 13156
rect 13051 13100 13119 13156
rect 13175 13100 13243 13156
rect 13299 13100 13367 13156
rect 13423 13100 13491 13156
rect 13547 13100 13615 13156
rect 13671 13100 13739 13156
rect 13795 13100 13863 13156
rect 13919 13100 13987 13156
rect 14043 13100 14111 13156
rect 14167 13100 14235 13156
rect 14291 13100 14359 13156
rect 14415 13100 14483 13156
rect 14539 13100 14607 13156
rect 14663 13100 14673 13156
rect 12861 13032 14673 13100
rect 12861 12976 12871 13032
rect 12927 12976 12995 13032
rect 13051 12976 13119 13032
rect 13175 12976 13243 13032
rect 13299 12976 13367 13032
rect 13423 12976 13491 13032
rect 13547 12976 13615 13032
rect 13671 12976 13739 13032
rect 13795 12976 13863 13032
rect 13919 12976 13987 13032
rect 14043 12976 14111 13032
rect 14167 12976 14235 13032
rect 14291 12976 14359 13032
rect 14415 12976 14483 13032
rect 14539 12976 14607 13032
rect 14663 12976 14673 13032
rect 12861 12908 14673 12976
rect 12861 12852 12871 12908
rect 12927 12852 12995 12908
rect 13051 12852 13119 12908
rect 13175 12852 13243 12908
rect 13299 12852 13367 12908
rect 13423 12852 13491 12908
rect 13547 12852 13615 12908
rect 13671 12852 13739 12908
rect 13795 12852 13863 12908
rect 13919 12852 13987 12908
rect 14043 12852 14111 12908
rect 14167 12852 14235 12908
rect 14291 12852 14359 12908
rect 14415 12852 14483 12908
rect 14539 12852 14607 12908
rect 14663 12852 14673 12908
rect 12861 12842 14673 12852
rect 10 12814 86 12824
rect 14892 12824 14902 14176
rect 14958 12824 14968 14176
rect 14892 12814 14968 12824
rect 2481 12548 2681 12558
rect 2481 12492 2491 12548
rect 2547 12492 2615 12548
rect 2671 12492 2681 12548
rect 2481 12424 2681 12492
rect 2481 12368 2491 12424
rect 2547 12368 2615 12424
rect 2671 12368 2681 12424
rect 2481 12300 2681 12368
rect 2481 12244 2491 12300
rect 2547 12244 2615 12300
rect 2671 12244 2681 12300
rect 2481 12176 2681 12244
rect 2481 12120 2491 12176
rect 2547 12120 2615 12176
rect 2671 12120 2681 12176
rect 2481 12052 2681 12120
rect 2481 11996 2491 12052
rect 2547 11996 2615 12052
rect 2671 11996 2681 12052
rect 2481 11928 2681 11996
rect 2481 11872 2491 11928
rect 2547 11872 2615 11928
rect 2671 11872 2681 11928
rect 2481 11804 2681 11872
rect 2481 11748 2491 11804
rect 2547 11748 2615 11804
rect 2671 11748 2681 11804
rect 2481 11680 2681 11748
rect 2481 11624 2491 11680
rect 2547 11624 2615 11680
rect 2671 11624 2681 11680
rect 2481 11556 2681 11624
rect 2481 11500 2491 11556
rect 2547 11500 2615 11556
rect 2671 11500 2681 11556
rect 2481 11432 2681 11500
rect 2481 11376 2491 11432
rect 2547 11376 2615 11432
rect 2671 11376 2681 11432
rect 2481 11308 2681 11376
rect 2481 11252 2491 11308
rect 2547 11252 2615 11308
rect 2671 11252 2681 11308
rect 2481 11242 2681 11252
rect 4851 12548 5051 12558
rect 4851 12492 4861 12548
rect 4917 12492 4985 12548
rect 5041 12492 5051 12548
rect 4851 12424 5051 12492
rect 4851 12368 4861 12424
rect 4917 12368 4985 12424
rect 5041 12368 5051 12424
rect 4851 12300 5051 12368
rect 4851 12244 4861 12300
rect 4917 12244 4985 12300
rect 5041 12244 5051 12300
rect 4851 12176 5051 12244
rect 4851 12120 4861 12176
rect 4917 12120 4985 12176
rect 5041 12120 5051 12176
rect 4851 12052 5051 12120
rect 4851 11996 4861 12052
rect 4917 11996 4985 12052
rect 5041 11996 5051 12052
rect 4851 11928 5051 11996
rect 4851 11872 4861 11928
rect 4917 11872 4985 11928
rect 5041 11872 5051 11928
rect 4851 11804 5051 11872
rect 4851 11748 4861 11804
rect 4917 11748 4985 11804
rect 5041 11748 5051 11804
rect 4851 11680 5051 11748
rect 4851 11624 4861 11680
rect 4917 11624 4985 11680
rect 5041 11624 5051 11680
rect 4851 11556 5051 11624
rect 4851 11500 4861 11556
rect 4917 11500 4985 11556
rect 5041 11500 5051 11556
rect 4851 11432 5051 11500
rect 4851 11376 4861 11432
rect 4917 11376 4985 11432
rect 5041 11376 5051 11432
rect 4851 11308 5051 11376
rect 4851 11252 4861 11308
rect 4917 11252 4985 11308
rect 5041 11252 5051 11308
rect 4851 11242 5051 11252
rect 7265 12548 7713 12558
rect 7265 12492 7275 12548
rect 7331 12492 7399 12548
rect 7455 12492 7523 12548
rect 7579 12492 7647 12548
rect 7703 12492 7713 12548
rect 7265 12424 7713 12492
rect 7265 12368 7275 12424
rect 7331 12368 7399 12424
rect 7455 12368 7523 12424
rect 7579 12368 7647 12424
rect 7703 12368 7713 12424
rect 7265 12300 7713 12368
rect 7265 12244 7275 12300
rect 7331 12244 7399 12300
rect 7455 12244 7523 12300
rect 7579 12244 7647 12300
rect 7703 12244 7713 12300
rect 7265 12176 7713 12244
rect 7265 12120 7275 12176
rect 7331 12120 7399 12176
rect 7455 12120 7523 12176
rect 7579 12120 7647 12176
rect 7703 12120 7713 12176
rect 7265 12052 7713 12120
rect 7265 11996 7275 12052
rect 7331 11996 7399 12052
rect 7455 11996 7523 12052
rect 7579 11996 7647 12052
rect 7703 11996 7713 12052
rect 7265 11928 7713 11996
rect 7265 11872 7275 11928
rect 7331 11872 7399 11928
rect 7455 11872 7523 11928
rect 7579 11872 7647 11928
rect 7703 11872 7713 11928
rect 7265 11804 7713 11872
rect 7265 11748 7275 11804
rect 7331 11748 7399 11804
rect 7455 11748 7523 11804
rect 7579 11748 7647 11804
rect 7703 11748 7713 11804
rect 7265 11680 7713 11748
rect 7265 11624 7275 11680
rect 7331 11624 7399 11680
rect 7455 11624 7523 11680
rect 7579 11624 7647 11680
rect 7703 11624 7713 11680
rect 7265 11556 7713 11624
rect 7265 11500 7275 11556
rect 7331 11500 7399 11556
rect 7455 11500 7523 11556
rect 7579 11500 7647 11556
rect 7703 11500 7713 11556
rect 7265 11432 7713 11500
rect 7265 11376 7275 11432
rect 7331 11376 7399 11432
rect 7455 11376 7523 11432
rect 7579 11376 7647 11432
rect 7703 11376 7713 11432
rect 7265 11308 7713 11376
rect 7265 11252 7275 11308
rect 7331 11252 7399 11308
rect 7455 11252 7523 11308
rect 7579 11252 7647 11308
rect 7703 11252 7713 11308
rect 7265 11242 7713 11252
rect 9927 12548 10127 12558
rect 9927 12492 9937 12548
rect 9993 12492 10061 12548
rect 10117 12492 10127 12548
rect 9927 12424 10127 12492
rect 9927 12368 9937 12424
rect 9993 12368 10061 12424
rect 10117 12368 10127 12424
rect 9927 12300 10127 12368
rect 9927 12244 9937 12300
rect 9993 12244 10061 12300
rect 10117 12244 10127 12300
rect 9927 12176 10127 12244
rect 9927 12120 9937 12176
rect 9993 12120 10061 12176
rect 10117 12120 10127 12176
rect 9927 12052 10127 12120
rect 9927 11996 9937 12052
rect 9993 11996 10061 12052
rect 10117 11996 10127 12052
rect 9927 11928 10127 11996
rect 9927 11872 9937 11928
rect 9993 11872 10061 11928
rect 10117 11872 10127 11928
rect 9927 11804 10127 11872
rect 9927 11748 9937 11804
rect 9993 11748 10061 11804
rect 10117 11748 10127 11804
rect 9927 11680 10127 11748
rect 9927 11624 9937 11680
rect 9993 11624 10061 11680
rect 10117 11624 10127 11680
rect 9927 11556 10127 11624
rect 9927 11500 9937 11556
rect 9993 11500 10061 11556
rect 10117 11500 10127 11556
rect 9927 11432 10127 11500
rect 9927 11376 9937 11432
rect 9993 11376 10061 11432
rect 10117 11376 10127 11432
rect 9927 11308 10127 11376
rect 9927 11252 9937 11308
rect 9993 11252 10061 11308
rect 10117 11252 10127 11308
rect 9927 11242 10127 11252
rect 12297 12548 12497 12558
rect 12297 12492 12307 12548
rect 12363 12492 12431 12548
rect 12487 12492 12497 12548
rect 12297 12424 12497 12492
rect 12297 12368 12307 12424
rect 12363 12368 12431 12424
rect 12487 12368 12497 12424
rect 12297 12300 12497 12368
rect 12297 12244 12307 12300
rect 12363 12244 12431 12300
rect 12487 12244 12497 12300
rect 12297 12176 12497 12244
rect 12297 12120 12307 12176
rect 12363 12120 12431 12176
rect 12487 12120 12497 12176
rect 12297 12052 12497 12120
rect 12297 11996 12307 12052
rect 12363 11996 12431 12052
rect 12487 11996 12497 12052
rect 12297 11928 12497 11996
rect 12297 11872 12307 11928
rect 12363 11872 12431 11928
rect 12487 11872 12497 11928
rect 12297 11804 12497 11872
rect 12297 11748 12307 11804
rect 12363 11748 12431 11804
rect 12487 11748 12497 11804
rect 12297 11680 12497 11748
rect 12297 11624 12307 11680
rect 12363 11624 12431 11680
rect 12487 11624 12497 11680
rect 12297 11556 12497 11624
rect 12297 11500 12307 11556
rect 12363 11500 12431 11556
rect 12487 11500 12497 11556
rect 12297 11432 12497 11500
rect 12297 11376 12307 11432
rect 12363 11376 12431 11432
rect 12487 11376 12497 11432
rect 12297 11308 12497 11376
rect 12297 11252 12307 11308
rect 12363 11252 12431 11308
rect 12487 11252 12497 11308
rect 12297 11242 12497 11252
rect 10 10986 86 10996
rect 10 8014 20 10986
rect 76 8014 86 10986
rect 14892 10986 14968 10996
rect 305 10954 2117 10964
rect 305 10898 315 10954
rect 371 10898 439 10954
rect 495 10898 563 10954
rect 619 10898 687 10954
rect 743 10898 811 10954
rect 867 10898 935 10954
rect 991 10898 1059 10954
rect 1115 10898 1183 10954
rect 1239 10898 1307 10954
rect 1363 10898 1431 10954
rect 1487 10898 1555 10954
rect 1611 10898 1679 10954
rect 1735 10898 1803 10954
rect 1859 10898 1927 10954
rect 1983 10898 2051 10954
rect 2107 10898 2117 10954
rect 305 10830 2117 10898
rect 305 10774 315 10830
rect 371 10774 439 10830
rect 495 10774 563 10830
rect 619 10774 687 10830
rect 743 10774 811 10830
rect 867 10774 935 10830
rect 991 10774 1059 10830
rect 1115 10774 1183 10830
rect 1239 10774 1307 10830
rect 1363 10774 1431 10830
rect 1487 10774 1555 10830
rect 1611 10774 1679 10830
rect 1735 10774 1803 10830
rect 1859 10774 1927 10830
rect 1983 10774 2051 10830
rect 2107 10774 2117 10830
rect 305 10706 2117 10774
rect 305 10650 315 10706
rect 371 10650 439 10706
rect 495 10650 563 10706
rect 619 10650 687 10706
rect 743 10650 811 10706
rect 867 10650 935 10706
rect 991 10650 1059 10706
rect 1115 10650 1183 10706
rect 1239 10650 1307 10706
rect 1363 10650 1431 10706
rect 1487 10650 1555 10706
rect 1611 10650 1679 10706
rect 1735 10650 1803 10706
rect 1859 10650 1927 10706
rect 1983 10650 2051 10706
rect 2107 10650 2117 10706
rect 305 10582 2117 10650
rect 305 10526 315 10582
rect 371 10526 439 10582
rect 495 10526 563 10582
rect 619 10526 687 10582
rect 743 10526 811 10582
rect 867 10526 935 10582
rect 991 10526 1059 10582
rect 1115 10526 1183 10582
rect 1239 10526 1307 10582
rect 1363 10526 1431 10582
rect 1487 10526 1555 10582
rect 1611 10526 1679 10582
rect 1735 10526 1803 10582
rect 1859 10526 1927 10582
rect 1983 10526 2051 10582
rect 2107 10526 2117 10582
rect 305 10458 2117 10526
rect 305 10402 315 10458
rect 371 10402 439 10458
rect 495 10402 563 10458
rect 619 10402 687 10458
rect 743 10402 811 10458
rect 867 10402 935 10458
rect 991 10402 1059 10458
rect 1115 10402 1183 10458
rect 1239 10402 1307 10458
rect 1363 10402 1431 10458
rect 1487 10402 1555 10458
rect 1611 10402 1679 10458
rect 1735 10402 1803 10458
rect 1859 10402 1927 10458
rect 1983 10402 2051 10458
rect 2107 10402 2117 10458
rect 305 10334 2117 10402
rect 305 10278 315 10334
rect 371 10278 439 10334
rect 495 10278 563 10334
rect 619 10278 687 10334
rect 743 10278 811 10334
rect 867 10278 935 10334
rect 991 10278 1059 10334
rect 1115 10278 1183 10334
rect 1239 10278 1307 10334
rect 1363 10278 1431 10334
rect 1487 10278 1555 10334
rect 1611 10278 1679 10334
rect 1735 10278 1803 10334
rect 1859 10278 1927 10334
rect 1983 10278 2051 10334
rect 2107 10278 2117 10334
rect 305 10210 2117 10278
rect 305 10154 315 10210
rect 371 10154 439 10210
rect 495 10154 563 10210
rect 619 10154 687 10210
rect 743 10154 811 10210
rect 867 10154 935 10210
rect 991 10154 1059 10210
rect 1115 10154 1183 10210
rect 1239 10154 1307 10210
rect 1363 10154 1431 10210
rect 1487 10154 1555 10210
rect 1611 10154 1679 10210
rect 1735 10154 1803 10210
rect 1859 10154 1927 10210
rect 1983 10154 2051 10210
rect 2107 10154 2117 10210
rect 305 10086 2117 10154
rect 305 10030 315 10086
rect 371 10030 439 10086
rect 495 10030 563 10086
rect 619 10030 687 10086
rect 743 10030 811 10086
rect 867 10030 935 10086
rect 991 10030 1059 10086
rect 1115 10030 1183 10086
rect 1239 10030 1307 10086
rect 1363 10030 1431 10086
rect 1487 10030 1555 10086
rect 1611 10030 1679 10086
rect 1735 10030 1803 10086
rect 1859 10030 1927 10086
rect 1983 10030 2051 10086
rect 2107 10030 2117 10086
rect 305 9962 2117 10030
rect 305 9906 315 9962
rect 371 9906 439 9962
rect 495 9906 563 9962
rect 619 9906 687 9962
rect 743 9906 811 9962
rect 867 9906 935 9962
rect 991 9906 1059 9962
rect 1115 9906 1183 9962
rect 1239 9906 1307 9962
rect 1363 9906 1431 9962
rect 1487 9906 1555 9962
rect 1611 9906 1679 9962
rect 1735 9906 1803 9962
rect 1859 9906 1927 9962
rect 1983 9906 2051 9962
rect 2107 9906 2117 9962
rect 305 9838 2117 9906
rect 305 9782 315 9838
rect 371 9782 439 9838
rect 495 9782 563 9838
rect 619 9782 687 9838
rect 743 9782 811 9838
rect 867 9782 935 9838
rect 991 9782 1059 9838
rect 1115 9782 1183 9838
rect 1239 9782 1307 9838
rect 1363 9782 1431 9838
rect 1487 9782 1555 9838
rect 1611 9782 1679 9838
rect 1735 9782 1803 9838
rect 1859 9782 1927 9838
rect 1983 9782 2051 9838
rect 2107 9782 2117 9838
rect 305 9714 2117 9782
rect 305 9658 315 9714
rect 371 9658 439 9714
rect 495 9658 563 9714
rect 619 9658 687 9714
rect 743 9658 811 9714
rect 867 9658 935 9714
rect 991 9658 1059 9714
rect 1115 9658 1183 9714
rect 1239 9658 1307 9714
rect 1363 9658 1431 9714
rect 1487 9658 1555 9714
rect 1611 9658 1679 9714
rect 1735 9658 1803 9714
rect 1859 9658 1927 9714
rect 1983 9658 2051 9714
rect 2107 9658 2117 9714
rect 305 9590 2117 9658
rect 305 9534 315 9590
rect 371 9534 439 9590
rect 495 9534 563 9590
rect 619 9534 687 9590
rect 743 9534 811 9590
rect 867 9534 935 9590
rect 991 9534 1059 9590
rect 1115 9534 1183 9590
rect 1239 9534 1307 9590
rect 1363 9534 1431 9590
rect 1487 9534 1555 9590
rect 1611 9534 1679 9590
rect 1735 9534 1803 9590
rect 1859 9534 1927 9590
rect 1983 9534 2051 9590
rect 2107 9534 2117 9590
rect 305 9466 2117 9534
rect 305 9410 315 9466
rect 371 9410 439 9466
rect 495 9410 563 9466
rect 619 9410 687 9466
rect 743 9410 811 9466
rect 867 9410 935 9466
rect 991 9410 1059 9466
rect 1115 9410 1183 9466
rect 1239 9410 1307 9466
rect 1363 9410 1431 9466
rect 1487 9410 1555 9466
rect 1611 9410 1679 9466
rect 1735 9410 1803 9466
rect 1859 9410 1927 9466
rect 1983 9410 2051 9466
rect 2107 9410 2117 9466
rect 305 9342 2117 9410
rect 305 9286 315 9342
rect 371 9286 439 9342
rect 495 9286 563 9342
rect 619 9286 687 9342
rect 743 9286 811 9342
rect 867 9286 935 9342
rect 991 9286 1059 9342
rect 1115 9286 1183 9342
rect 1239 9286 1307 9342
rect 1363 9286 1431 9342
rect 1487 9286 1555 9342
rect 1611 9286 1679 9342
rect 1735 9286 1803 9342
rect 1859 9286 1927 9342
rect 1983 9286 2051 9342
rect 2107 9286 2117 9342
rect 305 9218 2117 9286
rect 305 9162 315 9218
rect 371 9162 439 9218
rect 495 9162 563 9218
rect 619 9162 687 9218
rect 743 9162 811 9218
rect 867 9162 935 9218
rect 991 9162 1059 9218
rect 1115 9162 1183 9218
rect 1239 9162 1307 9218
rect 1363 9162 1431 9218
rect 1487 9162 1555 9218
rect 1611 9162 1679 9218
rect 1735 9162 1803 9218
rect 1859 9162 1927 9218
rect 1983 9162 2051 9218
rect 2107 9162 2117 9218
rect 305 9094 2117 9162
rect 305 9038 315 9094
rect 371 9038 439 9094
rect 495 9038 563 9094
rect 619 9038 687 9094
rect 743 9038 811 9094
rect 867 9038 935 9094
rect 991 9038 1059 9094
rect 1115 9038 1183 9094
rect 1239 9038 1307 9094
rect 1363 9038 1431 9094
rect 1487 9038 1555 9094
rect 1611 9038 1679 9094
rect 1735 9038 1803 9094
rect 1859 9038 1927 9094
rect 1983 9038 2051 9094
rect 2107 9038 2117 9094
rect 305 8970 2117 9038
rect 305 8914 315 8970
rect 371 8914 439 8970
rect 495 8914 563 8970
rect 619 8914 687 8970
rect 743 8914 811 8970
rect 867 8914 935 8970
rect 991 8914 1059 8970
rect 1115 8914 1183 8970
rect 1239 8914 1307 8970
rect 1363 8914 1431 8970
rect 1487 8914 1555 8970
rect 1611 8914 1679 8970
rect 1735 8914 1803 8970
rect 1859 8914 1927 8970
rect 1983 8914 2051 8970
rect 2107 8914 2117 8970
rect 305 8846 2117 8914
rect 305 8790 315 8846
rect 371 8790 439 8846
rect 495 8790 563 8846
rect 619 8790 687 8846
rect 743 8790 811 8846
rect 867 8790 935 8846
rect 991 8790 1059 8846
rect 1115 8790 1183 8846
rect 1239 8790 1307 8846
rect 1363 8790 1431 8846
rect 1487 8790 1555 8846
rect 1611 8790 1679 8846
rect 1735 8790 1803 8846
rect 1859 8790 1927 8846
rect 1983 8790 2051 8846
rect 2107 8790 2117 8846
rect 305 8722 2117 8790
rect 305 8666 315 8722
rect 371 8666 439 8722
rect 495 8666 563 8722
rect 619 8666 687 8722
rect 743 8666 811 8722
rect 867 8666 935 8722
rect 991 8666 1059 8722
rect 1115 8666 1183 8722
rect 1239 8666 1307 8722
rect 1363 8666 1431 8722
rect 1487 8666 1555 8722
rect 1611 8666 1679 8722
rect 1735 8666 1803 8722
rect 1859 8666 1927 8722
rect 1983 8666 2051 8722
rect 2107 8666 2117 8722
rect 305 8598 2117 8666
rect 305 8542 315 8598
rect 371 8542 439 8598
rect 495 8542 563 8598
rect 619 8542 687 8598
rect 743 8542 811 8598
rect 867 8542 935 8598
rect 991 8542 1059 8598
rect 1115 8542 1183 8598
rect 1239 8542 1307 8598
rect 1363 8542 1431 8598
rect 1487 8542 1555 8598
rect 1611 8542 1679 8598
rect 1735 8542 1803 8598
rect 1859 8542 1927 8598
rect 1983 8542 2051 8598
rect 2107 8542 2117 8598
rect 305 8474 2117 8542
rect 305 8418 315 8474
rect 371 8418 439 8474
rect 495 8418 563 8474
rect 619 8418 687 8474
rect 743 8418 811 8474
rect 867 8418 935 8474
rect 991 8418 1059 8474
rect 1115 8418 1183 8474
rect 1239 8418 1307 8474
rect 1363 8418 1431 8474
rect 1487 8418 1555 8474
rect 1611 8418 1679 8474
rect 1735 8418 1803 8474
rect 1859 8418 1927 8474
rect 1983 8418 2051 8474
rect 2107 8418 2117 8474
rect 305 8350 2117 8418
rect 305 8294 315 8350
rect 371 8294 439 8350
rect 495 8294 563 8350
rect 619 8294 687 8350
rect 743 8294 811 8350
rect 867 8294 935 8350
rect 991 8294 1059 8350
rect 1115 8294 1183 8350
rect 1239 8294 1307 8350
rect 1363 8294 1431 8350
rect 1487 8294 1555 8350
rect 1611 8294 1679 8350
rect 1735 8294 1803 8350
rect 1859 8294 1927 8350
rect 1983 8294 2051 8350
rect 2107 8294 2117 8350
rect 305 8226 2117 8294
rect 305 8170 315 8226
rect 371 8170 439 8226
rect 495 8170 563 8226
rect 619 8170 687 8226
rect 743 8170 811 8226
rect 867 8170 935 8226
rect 991 8170 1059 8226
rect 1115 8170 1183 8226
rect 1239 8170 1307 8226
rect 1363 8170 1431 8226
rect 1487 8170 1555 8226
rect 1611 8170 1679 8226
rect 1735 8170 1803 8226
rect 1859 8170 1927 8226
rect 1983 8170 2051 8226
rect 2107 8170 2117 8226
rect 305 8102 2117 8170
rect 305 8046 315 8102
rect 371 8046 439 8102
rect 495 8046 563 8102
rect 619 8046 687 8102
rect 743 8046 811 8102
rect 867 8046 935 8102
rect 991 8046 1059 8102
rect 1115 8046 1183 8102
rect 1239 8046 1307 8102
rect 1363 8046 1431 8102
rect 1487 8046 1555 8102
rect 1611 8046 1679 8102
rect 1735 8046 1803 8102
rect 1859 8046 1927 8102
rect 1983 8046 2051 8102
rect 2107 8046 2117 8102
rect 305 8036 2117 8046
rect 2798 10954 4734 10964
rect 2798 10898 2808 10954
rect 2864 10898 2932 10954
rect 2988 10898 3056 10954
rect 3112 10898 3180 10954
rect 3236 10898 3304 10954
rect 3360 10898 3428 10954
rect 3484 10898 3552 10954
rect 3608 10898 3676 10954
rect 3732 10898 3800 10954
rect 3856 10898 3924 10954
rect 3980 10898 4048 10954
rect 4104 10898 4172 10954
rect 4228 10898 4296 10954
rect 4352 10898 4420 10954
rect 4476 10898 4544 10954
rect 4600 10898 4668 10954
rect 4724 10898 4734 10954
rect 2798 10830 4734 10898
rect 2798 10774 2808 10830
rect 2864 10774 2932 10830
rect 2988 10774 3056 10830
rect 3112 10774 3180 10830
rect 3236 10774 3304 10830
rect 3360 10774 3428 10830
rect 3484 10774 3552 10830
rect 3608 10774 3676 10830
rect 3732 10774 3800 10830
rect 3856 10774 3924 10830
rect 3980 10774 4048 10830
rect 4104 10774 4172 10830
rect 4228 10774 4296 10830
rect 4352 10774 4420 10830
rect 4476 10774 4544 10830
rect 4600 10774 4668 10830
rect 4724 10774 4734 10830
rect 2798 10706 4734 10774
rect 2798 10650 2808 10706
rect 2864 10650 2932 10706
rect 2988 10650 3056 10706
rect 3112 10650 3180 10706
rect 3236 10650 3304 10706
rect 3360 10650 3428 10706
rect 3484 10650 3552 10706
rect 3608 10650 3676 10706
rect 3732 10650 3800 10706
rect 3856 10650 3924 10706
rect 3980 10650 4048 10706
rect 4104 10650 4172 10706
rect 4228 10650 4296 10706
rect 4352 10650 4420 10706
rect 4476 10650 4544 10706
rect 4600 10650 4668 10706
rect 4724 10650 4734 10706
rect 2798 10582 4734 10650
rect 2798 10526 2808 10582
rect 2864 10526 2932 10582
rect 2988 10526 3056 10582
rect 3112 10526 3180 10582
rect 3236 10526 3304 10582
rect 3360 10526 3428 10582
rect 3484 10526 3552 10582
rect 3608 10526 3676 10582
rect 3732 10526 3800 10582
rect 3856 10526 3924 10582
rect 3980 10526 4048 10582
rect 4104 10526 4172 10582
rect 4228 10526 4296 10582
rect 4352 10526 4420 10582
rect 4476 10526 4544 10582
rect 4600 10526 4668 10582
rect 4724 10526 4734 10582
rect 2798 10458 4734 10526
rect 2798 10402 2808 10458
rect 2864 10402 2932 10458
rect 2988 10402 3056 10458
rect 3112 10402 3180 10458
rect 3236 10402 3304 10458
rect 3360 10402 3428 10458
rect 3484 10402 3552 10458
rect 3608 10402 3676 10458
rect 3732 10402 3800 10458
rect 3856 10402 3924 10458
rect 3980 10402 4048 10458
rect 4104 10402 4172 10458
rect 4228 10402 4296 10458
rect 4352 10402 4420 10458
rect 4476 10402 4544 10458
rect 4600 10402 4668 10458
rect 4724 10402 4734 10458
rect 2798 10334 4734 10402
rect 2798 10278 2808 10334
rect 2864 10278 2932 10334
rect 2988 10278 3056 10334
rect 3112 10278 3180 10334
rect 3236 10278 3304 10334
rect 3360 10278 3428 10334
rect 3484 10278 3552 10334
rect 3608 10278 3676 10334
rect 3732 10278 3800 10334
rect 3856 10278 3924 10334
rect 3980 10278 4048 10334
rect 4104 10278 4172 10334
rect 4228 10278 4296 10334
rect 4352 10278 4420 10334
rect 4476 10278 4544 10334
rect 4600 10278 4668 10334
rect 4724 10278 4734 10334
rect 2798 10210 4734 10278
rect 2798 10154 2808 10210
rect 2864 10154 2932 10210
rect 2988 10154 3056 10210
rect 3112 10154 3180 10210
rect 3236 10154 3304 10210
rect 3360 10154 3428 10210
rect 3484 10154 3552 10210
rect 3608 10154 3676 10210
rect 3732 10154 3800 10210
rect 3856 10154 3924 10210
rect 3980 10154 4048 10210
rect 4104 10154 4172 10210
rect 4228 10154 4296 10210
rect 4352 10154 4420 10210
rect 4476 10154 4544 10210
rect 4600 10154 4668 10210
rect 4724 10154 4734 10210
rect 2798 10086 4734 10154
rect 2798 10030 2808 10086
rect 2864 10030 2932 10086
rect 2988 10030 3056 10086
rect 3112 10030 3180 10086
rect 3236 10030 3304 10086
rect 3360 10030 3428 10086
rect 3484 10030 3552 10086
rect 3608 10030 3676 10086
rect 3732 10030 3800 10086
rect 3856 10030 3924 10086
rect 3980 10030 4048 10086
rect 4104 10030 4172 10086
rect 4228 10030 4296 10086
rect 4352 10030 4420 10086
rect 4476 10030 4544 10086
rect 4600 10030 4668 10086
rect 4724 10030 4734 10086
rect 2798 9962 4734 10030
rect 2798 9906 2808 9962
rect 2864 9906 2932 9962
rect 2988 9906 3056 9962
rect 3112 9906 3180 9962
rect 3236 9906 3304 9962
rect 3360 9906 3428 9962
rect 3484 9906 3552 9962
rect 3608 9906 3676 9962
rect 3732 9906 3800 9962
rect 3856 9906 3924 9962
rect 3980 9906 4048 9962
rect 4104 9906 4172 9962
rect 4228 9906 4296 9962
rect 4352 9906 4420 9962
rect 4476 9906 4544 9962
rect 4600 9906 4668 9962
rect 4724 9906 4734 9962
rect 2798 9838 4734 9906
rect 2798 9782 2808 9838
rect 2864 9782 2932 9838
rect 2988 9782 3056 9838
rect 3112 9782 3180 9838
rect 3236 9782 3304 9838
rect 3360 9782 3428 9838
rect 3484 9782 3552 9838
rect 3608 9782 3676 9838
rect 3732 9782 3800 9838
rect 3856 9782 3924 9838
rect 3980 9782 4048 9838
rect 4104 9782 4172 9838
rect 4228 9782 4296 9838
rect 4352 9782 4420 9838
rect 4476 9782 4544 9838
rect 4600 9782 4668 9838
rect 4724 9782 4734 9838
rect 2798 9714 4734 9782
rect 2798 9658 2808 9714
rect 2864 9658 2932 9714
rect 2988 9658 3056 9714
rect 3112 9658 3180 9714
rect 3236 9658 3304 9714
rect 3360 9658 3428 9714
rect 3484 9658 3552 9714
rect 3608 9658 3676 9714
rect 3732 9658 3800 9714
rect 3856 9658 3924 9714
rect 3980 9658 4048 9714
rect 4104 9658 4172 9714
rect 4228 9658 4296 9714
rect 4352 9658 4420 9714
rect 4476 9658 4544 9714
rect 4600 9658 4668 9714
rect 4724 9658 4734 9714
rect 2798 9590 4734 9658
rect 2798 9534 2808 9590
rect 2864 9534 2932 9590
rect 2988 9534 3056 9590
rect 3112 9534 3180 9590
rect 3236 9534 3304 9590
rect 3360 9534 3428 9590
rect 3484 9534 3552 9590
rect 3608 9534 3676 9590
rect 3732 9534 3800 9590
rect 3856 9534 3924 9590
rect 3980 9534 4048 9590
rect 4104 9534 4172 9590
rect 4228 9534 4296 9590
rect 4352 9534 4420 9590
rect 4476 9534 4544 9590
rect 4600 9534 4668 9590
rect 4724 9534 4734 9590
rect 2798 9466 4734 9534
rect 2798 9410 2808 9466
rect 2864 9410 2932 9466
rect 2988 9410 3056 9466
rect 3112 9410 3180 9466
rect 3236 9410 3304 9466
rect 3360 9410 3428 9466
rect 3484 9410 3552 9466
rect 3608 9410 3676 9466
rect 3732 9410 3800 9466
rect 3856 9410 3924 9466
rect 3980 9410 4048 9466
rect 4104 9410 4172 9466
rect 4228 9410 4296 9466
rect 4352 9410 4420 9466
rect 4476 9410 4544 9466
rect 4600 9410 4668 9466
rect 4724 9410 4734 9466
rect 2798 9342 4734 9410
rect 2798 9286 2808 9342
rect 2864 9286 2932 9342
rect 2988 9286 3056 9342
rect 3112 9286 3180 9342
rect 3236 9286 3304 9342
rect 3360 9286 3428 9342
rect 3484 9286 3552 9342
rect 3608 9286 3676 9342
rect 3732 9286 3800 9342
rect 3856 9286 3924 9342
rect 3980 9286 4048 9342
rect 4104 9286 4172 9342
rect 4228 9286 4296 9342
rect 4352 9286 4420 9342
rect 4476 9286 4544 9342
rect 4600 9286 4668 9342
rect 4724 9286 4734 9342
rect 2798 9218 4734 9286
rect 2798 9162 2808 9218
rect 2864 9162 2932 9218
rect 2988 9162 3056 9218
rect 3112 9162 3180 9218
rect 3236 9162 3304 9218
rect 3360 9162 3428 9218
rect 3484 9162 3552 9218
rect 3608 9162 3676 9218
rect 3732 9162 3800 9218
rect 3856 9162 3924 9218
rect 3980 9162 4048 9218
rect 4104 9162 4172 9218
rect 4228 9162 4296 9218
rect 4352 9162 4420 9218
rect 4476 9162 4544 9218
rect 4600 9162 4668 9218
rect 4724 9162 4734 9218
rect 2798 9094 4734 9162
rect 2798 9038 2808 9094
rect 2864 9038 2932 9094
rect 2988 9038 3056 9094
rect 3112 9038 3180 9094
rect 3236 9038 3304 9094
rect 3360 9038 3428 9094
rect 3484 9038 3552 9094
rect 3608 9038 3676 9094
rect 3732 9038 3800 9094
rect 3856 9038 3924 9094
rect 3980 9038 4048 9094
rect 4104 9038 4172 9094
rect 4228 9038 4296 9094
rect 4352 9038 4420 9094
rect 4476 9038 4544 9094
rect 4600 9038 4668 9094
rect 4724 9038 4734 9094
rect 2798 8970 4734 9038
rect 2798 8914 2808 8970
rect 2864 8914 2932 8970
rect 2988 8914 3056 8970
rect 3112 8914 3180 8970
rect 3236 8914 3304 8970
rect 3360 8914 3428 8970
rect 3484 8914 3552 8970
rect 3608 8914 3676 8970
rect 3732 8914 3800 8970
rect 3856 8914 3924 8970
rect 3980 8914 4048 8970
rect 4104 8914 4172 8970
rect 4228 8914 4296 8970
rect 4352 8914 4420 8970
rect 4476 8914 4544 8970
rect 4600 8914 4668 8970
rect 4724 8914 4734 8970
rect 2798 8846 4734 8914
rect 2798 8790 2808 8846
rect 2864 8790 2932 8846
rect 2988 8790 3056 8846
rect 3112 8790 3180 8846
rect 3236 8790 3304 8846
rect 3360 8790 3428 8846
rect 3484 8790 3552 8846
rect 3608 8790 3676 8846
rect 3732 8790 3800 8846
rect 3856 8790 3924 8846
rect 3980 8790 4048 8846
rect 4104 8790 4172 8846
rect 4228 8790 4296 8846
rect 4352 8790 4420 8846
rect 4476 8790 4544 8846
rect 4600 8790 4668 8846
rect 4724 8790 4734 8846
rect 2798 8722 4734 8790
rect 2798 8666 2808 8722
rect 2864 8666 2932 8722
rect 2988 8666 3056 8722
rect 3112 8666 3180 8722
rect 3236 8666 3304 8722
rect 3360 8666 3428 8722
rect 3484 8666 3552 8722
rect 3608 8666 3676 8722
rect 3732 8666 3800 8722
rect 3856 8666 3924 8722
rect 3980 8666 4048 8722
rect 4104 8666 4172 8722
rect 4228 8666 4296 8722
rect 4352 8666 4420 8722
rect 4476 8666 4544 8722
rect 4600 8666 4668 8722
rect 4724 8666 4734 8722
rect 2798 8598 4734 8666
rect 2798 8542 2808 8598
rect 2864 8542 2932 8598
rect 2988 8542 3056 8598
rect 3112 8542 3180 8598
rect 3236 8542 3304 8598
rect 3360 8542 3428 8598
rect 3484 8542 3552 8598
rect 3608 8542 3676 8598
rect 3732 8542 3800 8598
rect 3856 8542 3924 8598
rect 3980 8542 4048 8598
rect 4104 8542 4172 8598
rect 4228 8542 4296 8598
rect 4352 8542 4420 8598
rect 4476 8542 4544 8598
rect 4600 8542 4668 8598
rect 4724 8542 4734 8598
rect 2798 8474 4734 8542
rect 2798 8418 2808 8474
rect 2864 8418 2932 8474
rect 2988 8418 3056 8474
rect 3112 8418 3180 8474
rect 3236 8418 3304 8474
rect 3360 8418 3428 8474
rect 3484 8418 3552 8474
rect 3608 8418 3676 8474
rect 3732 8418 3800 8474
rect 3856 8418 3924 8474
rect 3980 8418 4048 8474
rect 4104 8418 4172 8474
rect 4228 8418 4296 8474
rect 4352 8418 4420 8474
rect 4476 8418 4544 8474
rect 4600 8418 4668 8474
rect 4724 8418 4734 8474
rect 2798 8350 4734 8418
rect 2798 8294 2808 8350
rect 2864 8294 2932 8350
rect 2988 8294 3056 8350
rect 3112 8294 3180 8350
rect 3236 8294 3304 8350
rect 3360 8294 3428 8350
rect 3484 8294 3552 8350
rect 3608 8294 3676 8350
rect 3732 8294 3800 8350
rect 3856 8294 3924 8350
rect 3980 8294 4048 8350
rect 4104 8294 4172 8350
rect 4228 8294 4296 8350
rect 4352 8294 4420 8350
rect 4476 8294 4544 8350
rect 4600 8294 4668 8350
rect 4724 8294 4734 8350
rect 2798 8226 4734 8294
rect 2798 8170 2808 8226
rect 2864 8170 2932 8226
rect 2988 8170 3056 8226
rect 3112 8170 3180 8226
rect 3236 8170 3304 8226
rect 3360 8170 3428 8226
rect 3484 8170 3552 8226
rect 3608 8170 3676 8226
rect 3732 8170 3800 8226
rect 3856 8170 3924 8226
rect 3980 8170 4048 8226
rect 4104 8170 4172 8226
rect 4228 8170 4296 8226
rect 4352 8170 4420 8226
rect 4476 8170 4544 8226
rect 4600 8170 4668 8226
rect 4724 8170 4734 8226
rect 2798 8102 4734 8170
rect 2798 8046 2808 8102
rect 2864 8046 2932 8102
rect 2988 8046 3056 8102
rect 3112 8046 3180 8102
rect 3236 8046 3304 8102
rect 3360 8046 3428 8102
rect 3484 8046 3552 8102
rect 3608 8046 3676 8102
rect 3732 8046 3800 8102
rect 3856 8046 3924 8102
rect 3980 8046 4048 8102
rect 4104 8046 4172 8102
rect 4228 8046 4296 8102
rect 4352 8046 4420 8102
rect 4476 8046 4544 8102
rect 4600 8046 4668 8102
rect 4724 8046 4734 8102
rect 2798 8036 4734 8046
rect 5168 10954 7104 10964
rect 5168 10898 5178 10954
rect 5234 10898 5302 10954
rect 5358 10898 5426 10954
rect 5482 10898 5550 10954
rect 5606 10898 5674 10954
rect 5730 10898 5798 10954
rect 5854 10898 5922 10954
rect 5978 10898 6046 10954
rect 6102 10898 6170 10954
rect 6226 10898 6294 10954
rect 6350 10898 6418 10954
rect 6474 10898 6542 10954
rect 6598 10898 6666 10954
rect 6722 10898 6790 10954
rect 6846 10898 6914 10954
rect 6970 10898 7038 10954
rect 7094 10898 7104 10954
rect 5168 10830 7104 10898
rect 5168 10774 5178 10830
rect 5234 10774 5302 10830
rect 5358 10774 5426 10830
rect 5482 10774 5550 10830
rect 5606 10774 5674 10830
rect 5730 10774 5798 10830
rect 5854 10774 5922 10830
rect 5978 10774 6046 10830
rect 6102 10774 6170 10830
rect 6226 10774 6294 10830
rect 6350 10774 6418 10830
rect 6474 10774 6542 10830
rect 6598 10774 6666 10830
rect 6722 10774 6790 10830
rect 6846 10774 6914 10830
rect 6970 10774 7038 10830
rect 7094 10774 7104 10830
rect 5168 10706 7104 10774
rect 5168 10650 5178 10706
rect 5234 10650 5302 10706
rect 5358 10650 5426 10706
rect 5482 10650 5550 10706
rect 5606 10650 5674 10706
rect 5730 10650 5798 10706
rect 5854 10650 5922 10706
rect 5978 10650 6046 10706
rect 6102 10650 6170 10706
rect 6226 10650 6294 10706
rect 6350 10650 6418 10706
rect 6474 10650 6542 10706
rect 6598 10650 6666 10706
rect 6722 10650 6790 10706
rect 6846 10650 6914 10706
rect 6970 10650 7038 10706
rect 7094 10650 7104 10706
rect 5168 10582 7104 10650
rect 5168 10526 5178 10582
rect 5234 10526 5302 10582
rect 5358 10526 5426 10582
rect 5482 10526 5550 10582
rect 5606 10526 5674 10582
rect 5730 10526 5798 10582
rect 5854 10526 5922 10582
rect 5978 10526 6046 10582
rect 6102 10526 6170 10582
rect 6226 10526 6294 10582
rect 6350 10526 6418 10582
rect 6474 10526 6542 10582
rect 6598 10526 6666 10582
rect 6722 10526 6790 10582
rect 6846 10526 6914 10582
rect 6970 10526 7038 10582
rect 7094 10526 7104 10582
rect 5168 10458 7104 10526
rect 5168 10402 5178 10458
rect 5234 10402 5302 10458
rect 5358 10402 5426 10458
rect 5482 10402 5550 10458
rect 5606 10402 5674 10458
rect 5730 10402 5798 10458
rect 5854 10402 5922 10458
rect 5978 10402 6046 10458
rect 6102 10402 6170 10458
rect 6226 10402 6294 10458
rect 6350 10402 6418 10458
rect 6474 10402 6542 10458
rect 6598 10402 6666 10458
rect 6722 10402 6790 10458
rect 6846 10402 6914 10458
rect 6970 10402 7038 10458
rect 7094 10402 7104 10458
rect 5168 10334 7104 10402
rect 5168 10278 5178 10334
rect 5234 10278 5302 10334
rect 5358 10278 5426 10334
rect 5482 10278 5550 10334
rect 5606 10278 5674 10334
rect 5730 10278 5798 10334
rect 5854 10278 5922 10334
rect 5978 10278 6046 10334
rect 6102 10278 6170 10334
rect 6226 10278 6294 10334
rect 6350 10278 6418 10334
rect 6474 10278 6542 10334
rect 6598 10278 6666 10334
rect 6722 10278 6790 10334
rect 6846 10278 6914 10334
rect 6970 10278 7038 10334
rect 7094 10278 7104 10334
rect 5168 10210 7104 10278
rect 5168 10154 5178 10210
rect 5234 10154 5302 10210
rect 5358 10154 5426 10210
rect 5482 10154 5550 10210
rect 5606 10154 5674 10210
rect 5730 10154 5798 10210
rect 5854 10154 5922 10210
rect 5978 10154 6046 10210
rect 6102 10154 6170 10210
rect 6226 10154 6294 10210
rect 6350 10154 6418 10210
rect 6474 10154 6542 10210
rect 6598 10154 6666 10210
rect 6722 10154 6790 10210
rect 6846 10154 6914 10210
rect 6970 10154 7038 10210
rect 7094 10154 7104 10210
rect 5168 10086 7104 10154
rect 5168 10030 5178 10086
rect 5234 10030 5302 10086
rect 5358 10030 5426 10086
rect 5482 10030 5550 10086
rect 5606 10030 5674 10086
rect 5730 10030 5798 10086
rect 5854 10030 5922 10086
rect 5978 10030 6046 10086
rect 6102 10030 6170 10086
rect 6226 10030 6294 10086
rect 6350 10030 6418 10086
rect 6474 10030 6542 10086
rect 6598 10030 6666 10086
rect 6722 10030 6790 10086
rect 6846 10030 6914 10086
rect 6970 10030 7038 10086
rect 7094 10030 7104 10086
rect 5168 9962 7104 10030
rect 5168 9906 5178 9962
rect 5234 9906 5302 9962
rect 5358 9906 5426 9962
rect 5482 9906 5550 9962
rect 5606 9906 5674 9962
rect 5730 9906 5798 9962
rect 5854 9906 5922 9962
rect 5978 9906 6046 9962
rect 6102 9906 6170 9962
rect 6226 9906 6294 9962
rect 6350 9906 6418 9962
rect 6474 9906 6542 9962
rect 6598 9906 6666 9962
rect 6722 9906 6790 9962
rect 6846 9906 6914 9962
rect 6970 9906 7038 9962
rect 7094 9906 7104 9962
rect 5168 9838 7104 9906
rect 5168 9782 5178 9838
rect 5234 9782 5302 9838
rect 5358 9782 5426 9838
rect 5482 9782 5550 9838
rect 5606 9782 5674 9838
rect 5730 9782 5798 9838
rect 5854 9782 5922 9838
rect 5978 9782 6046 9838
rect 6102 9782 6170 9838
rect 6226 9782 6294 9838
rect 6350 9782 6418 9838
rect 6474 9782 6542 9838
rect 6598 9782 6666 9838
rect 6722 9782 6790 9838
rect 6846 9782 6914 9838
rect 6970 9782 7038 9838
rect 7094 9782 7104 9838
rect 5168 9714 7104 9782
rect 5168 9658 5178 9714
rect 5234 9658 5302 9714
rect 5358 9658 5426 9714
rect 5482 9658 5550 9714
rect 5606 9658 5674 9714
rect 5730 9658 5798 9714
rect 5854 9658 5922 9714
rect 5978 9658 6046 9714
rect 6102 9658 6170 9714
rect 6226 9658 6294 9714
rect 6350 9658 6418 9714
rect 6474 9658 6542 9714
rect 6598 9658 6666 9714
rect 6722 9658 6790 9714
rect 6846 9658 6914 9714
rect 6970 9658 7038 9714
rect 7094 9658 7104 9714
rect 5168 9590 7104 9658
rect 5168 9534 5178 9590
rect 5234 9534 5302 9590
rect 5358 9534 5426 9590
rect 5482 9534 5550 9590
rect 5606 9534 5674 9590
rect 5730 9534 5798 9590
rect 5854 9534 5922 9590
rect 5978 9534 6046 9590
rect 6102 9534 6170 9590
rect 6226 9534 6294 9590
rect 6350 9534 6418 9590
rect 6474 9534 6542 9590
rect 6598 9534 6666 9590
rect 6722 9534 6790 9590
rect 6846 9534 6914 9590
rect 6970 9534 7038 9590
rect 7094 9534 7104 9590
rect 5168 9466 7104 9534
rect 5168 9410 5178 9466
rect 5234 9410 5302 9466
rect 5358 9410 5426 9466
rect 5482 9410 5550 9466
rect 5606 9410 5674 9466
rect 5730 9410 5798 9466
rect 5854 9410 5922 9466
rect 5978 9410 6046 9466
rect 6102 9410 6170 9466
rect 6226 9410 6294 9466
rect 6350 9410 6418 9466
rect 6474 9410 6542 9466
rect 6598 9410 6666 9466
rect 6722 9410 6790 9466
rect 6846 9410 6914 9466
rect 6970 9410 7038 9466
rect 7094 9410 7104 9466
rect 5168 9342 7104 9410
rect 5168 9286 5178 9342
rect 5234 9286 5302 9342
rect 5358 9286 5426 9342
rect 5482 9286 5550 9342
rect 5606 9286 5674 9342
rect 5730 9286 5798 9342
rect 5854 9286 5922 9342
rect 5978 9286 6046 9342
rect 6102 9286 6170 9342
rect 6226 9286 6294 9342
rect 6350 9286 6418 9342
rect 6474 9286 6542 9342
rect 6598 9286 6666 9342
rect 6722 9286 6790 9342
rect 6846 9286 6914 9342
rect 6970 9286 7038 9342
rect 7094 9286 7104 9342
rect 5168 9218 7104 9286
rect 5168 9162 5178 9218
rect 5234 9162 5302 9218
rect 5358 9162 5426 9218
rect 5482 9162 5550 9218
rect 5606 9162 5674 9218
rect 5730 9162 5798 9218
rect 5854 9162 5922 9218
rect 5978 9162 6046 9218
rect 6102 9162 6170 9218
rect 6226 9162 6294 9218
rect 6350 9162 6418 9218
rect 6474 9162 6542 9218
rect 6598 9162 6666 9218
rect 6722 9162 6790 9218
rect 6846 9162 6914 9218
rect 6970 9162 7038 9218
rect 7094 9162 7104 9218
rect 5168 9094 7104 9162
rect 5168 9038 5178 9094
rect 5234 9038 5302 9094
rect 5358 9038 5426 9094
rect 5482 9038 5550 9094
rect 5606 9038 5674 9094
rect 5730 9038 5798 9094
rect 5854 9038 5922 9094
rect 5978 9038 6046 9094
rect 6102 9038 6170 9094
rect 6226 9038 6294 9094
rect 6350 9038 6418 9094
rect 6474 9038 6542 9094
rect 6598 9038 6666 9094
rect 6722 9038 6790 9094
rect 6846 9038 6914 9094
rect 6970 9038 7038 9094
rect 7094 9038 7104 9094
rect 5168 8970 7104 9038
rect 5168 8914 5178 8970
rect 5234 8914 5302 8970
rect 5358 8914 5426 8970
rect 5482 8914 5550 8970
rect 5606 8914 5674 8970
rect 5730 8914 5798 8970
rect 5854 8914 5922 8970
rect 5978 8914 6046 8970
rect 6102 8914 6170 8970
rect 6226 8914 6294 8970
rect 6350 8914 6418 8970
rect 6474 8914 6542 8970
rect 6598 8914 6666 8970
rect 6722 8914 6790 8970
rect 6846 8914 6914 8970
rect 6970 8914 7038 8970
rect 7094 8914 7104 8970
rect 5168 8846 7104 8914
rect 5168 8790 5178 8846
rect 5234 8790 5302 8846
rect 5358 8790 5426 8846
rect 5482 8790 5550 8846
rect 5606 8790 5674 8846
rect 5730 8790 5798 8846
rect 5854 8790 5922 8846
rect 5978 8790 6046 8846
rect 6102 8790 6170 8846
rect 6226 8790 6294 8846
rect 6350 8790 6418 8846
rect 6474 8790 6542 8846
rect 6598 8790 6666 8846
rect 6722 8790 6790 8846
rect 6846 8790 6914 8846
rect 6970 8790 7038 8846
rect 7094 8790 7104 8846
rect 5168 8722 7104 8790
rect 5168 8666 5178 8722
rect 5234 8666 5302 8722
rect 5358 8666 5426 8722
rect 5482 8666 5550 8722
rect 5606 8666 5674 8722
rect 5730 8666 5798 8722
rect 5854 8666 5922 8722
rect 5978 8666 6046 8722
rect 6102 8666 6170 8722
rect 6226 8666 6294 8722
rect 6350 8666 6418 8722
rect 6474 8666 6542 8722
rect 6598 8666 6666 8722
rect 6722 8666 6790 8722
rect 6846 8666 6914 8722
rect 6970 8666 7038 8722
rect 7094 8666 7104 8722
rect 5168 8598 7104 8666
rect 5168 8542 5178 8598
rect 5234 8542 5302 8598
rect 5358 8542 5426 8598
rect 5482 8542 5550 8598
rect 5606 8542 5674 8598
rect 5730 8542 5798 8598
rect 5854 8542 5922 8598
rect 5978 8542 6046 8598
rect 6102 8542 6170 8598
rect 6226 8542 6294 8598
rect 6350 8542 6418 8598
rect 6474 8542 6542 8598
rect 6598 8542 6666 8598
rect 6722 8542 6790 8598
rect 6846 8542 6914 8598
rect 6970 8542 7038 8598
rect 7094 8542 7104 8598
rect 5168 8474 7104 8542
rect 5168 8418 5178 8474
rect 5234 8418 5302 8474
rect 5358 8418 5426 8474
rect 5482 8418 5550 8474
rect 5606 8418 5674 8474
rect 5730 8418 5798 8474
rect 5854 8418 5922 8474
rect 5978 8418 6046 8474
rect 6102 8418 6170 8474
rect 6226 8418 6294 8474
rect 6350 8418 6418 8474
rect 6474 8418 6542 8474
rect 6598 8418 6666 8474
rect 6722 8418 6790 8474
rect 6846 8418 6914 8474
rect 6970 8418 7038 8474
rect 7094 8418 7104 8474
rect 5168 8350 7104 8418
rect 5168 8294 5178 8350
rect 5234 8294 5302 8350
rect 5358 8294 5426 8350
rect 5482 8294 5550 8350
rect 5606 8294 5674 8350
rect 5730 8294 5798 8350
rect 5854 8294 5922 8350
rect 5978 8294 6046 8350
rect 6102 8294 6170 8350
rect 6226 8294 6294 8350
rect 6350 8294 6418 8350
rect 6474 8294 6542 8350
rect 6598 8294 6666 8350
rect 6722 8294 6790 8350
rect 6846 8294 6914 8350
rect 6970 8294 7038 8350
rect 7094 8294 7104 8350
rect 5168 8226 7104 8294
rect 5168 8170 5178 8226
rect 5234 8170 5302 8226
rect 5358 8170 5426 8226
rect 5482 8170 5550 8226
rect 5606 8170 5674 8226
rect 5730 8170 5798 8226
rect 5854 8170 5922 8226
rect 5978 8170 6046 8226
rect 6102 8170 6170 8226
rect 6226 8170 6294 8226
rect 6350 8170 6418 8226
rect 6474 8170 6542 8226
rect 6598 8170 6666 8226
rect 6722 8170 6790 8226
rect 6846 8170 6914 8226
rect 6970 8170 7038 8226
rect 7094 8170 7104 8226
rect 5168 8102 7104 8170
rect 5168 8046 5178 8102
rect 5234 8046 5302 8102
rect 5358 8046 5426 8102
rect 5482 8046 5550 8102
rect 5606 8046 5674 8102
rect 5730 8046 5798 8102
rect 5854 8046 5922 8102
rect 5978 8046 6046 8102
rect 6102 8046 6170 8102
rect 6226 8046 6294 8102
rect 6350 8046 6418 8102
rect 6474 8046 6542 8102
rect 6598 8046 6666 8102
rect 6722 8046 6790 8102
rect 6846 8046 6914 8102
rect 6970 8046 7038 8102
rect 7094 8046 7104 8102
rect 5168 8036 7104 8046
rect 7874 10954 9810 10964
rect 7874 10898 7884 10954
rect 7940 10898 8008 10954
rect 8064 10898 8132 10954
rect 8188 10898 8256 10954
rect 8312 10898 8380 10954
rect 8436 10898 8504 10954
rect 8560 10898 8628 10954
rect 8684 10898 8752 10954
rect 8808 10898 8876 10954
rect 8932 10898 9000 10954
rect 9056 10898 9124 10954
rect 9180 10898 9248 10954
rect 9304 10898 9372 10954
rect 9428 10898 9496 10954
rect 9552 10898 9620 10954
rect 9676 10898 9744 10954
rect 9800 10898 9810 10954
rect 7874 10830 9810 10898
rect 7874 10774 7884 10830
rect 7940 10774 8008 10830
rect 8064 10774 8132 10830
rect 8188 10774 8256 10830
rect 8312 10774 8380 10830
rect 8436 10774 8504 10830
rect 8560 10774 8628 10830
rect 8684 10774 8752 10830
rect 8808 10774 8876 10830
rect 8932 10774 9000 10830
rect 9056 10774 9124 10830
rect 9180 10774 9248 10830
rect 9304 10774 9372 10830
rect 9428 10774 9496 10830
rect 9552 10774 9620 10830
rect 9676 10774 9744 10830
rect 9800 10774 9810 10830
rect 7874 10706 9810 10774
rect 7874 10650 7884 10706
rect 7940 10650 8008 10706
rect 8064 10650 8132 10706
rect 8188 10650 8256 10706
rect 8312 10650 8380 10706
rect 8436 10650 8504 10706
rect 8560 10650 8628 10706
rect 8684 10650 8752 10706
rect 8808 10650 8876 10706
rect 8932 10650 9000 10706
rect 9056 10650 9124 10706
rect 9180 10650 9248 10706
rect 9304 10650 9372 10706
rect 9428 10650 9496 10706
rect 9552 10650 9620 10706
rect 9676 10650 9744 10706
rect 9800 10650 9810 10706
rect 7874 10582 9810 10650
rect 7874 10526 7884 10582
rect 7940 10526 8008 10582
rect 8064 10526 8132 10582
rect 8188 10526 8256 10582
rect 8312 10526 8380 10582
rect 8436 10526 8504 10582
rect 8560 10526 8628 10582
rect 8684 10526 8752 10582
rect 8808 10526 8876 10582
rect 8932 10526 9000 10582
rect 9056 10526 9124 10582
rect 9180 10526 9248 10582
rect 9304 10526 9372 10582
rect 9428 10526 9496 10582
rect 9552 10526 9620 10582
rect 9676 10526 9744 10582
rect 9800 10526 9810 10582
rect 7874 10458 9810 10526
rect 7874 10402 7884 10458
rect 7940 10402 8008 10458
rect 8064 10402 8132 10458
rect 8188 10402 8256 10458
rect 8312 10402 8380 10458
rect 8436 10402 8504 10458
rect 8560 10402 8628 10458
rect 8684 10402 8752 10458
rect 8808 10402 8876 10458
rect 8932 10402 9000 10458
rect 9056 10402 9124 10458
rect 9180 10402 9248 10458
rect 9304 10402 9372 10458
rect 9428 10402 9496 10458
rect 9552 10402 9620 10458
rect 9676 10402 9744 10458
rect 9800 10402 9810 10458
rect 7874 10334 9810 10402
rect 7874 10278 7884 10334
rect 7940 10278 8008 10334
rect 8064 10278 8132 10334
rect 8188 10278 8256 10334
rect 8312 10278 8380 10334
rect 8436 10278 8504 10334
rect 8560 10278 8628 10334
rect 8684 10278 8752 10334
rect 8808 10278 8876 10334
rect 8932 10278 9000 10334
rect 9056 10278 9124 10334
rect 9180 10278 9248 10334
rect 9304 10278 9372 10334
rect 9428 10278 9496 10334
rect 9552 10278 9620 10334
rect 9676 10278 9744 10334
rect 9800 10278 9810 10334
rect 7874 10210 9810 10278
rect 7874 10154 7884 10210
rect 7940 10154 8008 10210
rect 8064 10154 8132 10210
rect 8188 10154 8256 10210
rect 8312 10154 8380 10210
rect 8436 10154 8504 10210
rect 8560 10154 8628 10210
rect 8684 10154 8752 10210
rect 8808 10154 8876 10210
rect 8932 10154 9000 10210
rect 9056 10154 9124 10210
rect 9180 10154 9248 10210
rect 9304 10154 9372 10210
rect 9428 10154 9496 10210
rect 9552 10154 9620 10210
rect 9676 10154 9744 10210
rect 9800 10154 9810 10210
rect 7874 10086 9810 10154
rect 7874 10030 7884 10086
rect 7940 10030 8008 10086
rect 8064 10030 8132 10086
rect 8188 10030 8256 10086
rect 8312 10030 8380 10086
rect 8436 10030 8504 10086
rect 8560 10030 8628 10086
rect 8684 10030 8752 10086
rect 8808 10030 8876 10086
rect 8932 10030 9000 10086
rect 9056 10030 9124 10086
rect 9180 10030 9248 10086
rect 9304 10030 9372 10086
rect 9428 10030 9496 10086
rect 9552 10030 9620 10086
rect 9676 10030 9744 10086
rect 9800 10030 9810 10086
rect 7874 9962 9810 10030
rect 7874 9906 7884 9962
rect 7940 9906 8008 9962
rect 8064 9906 8132 9962
rect 8188 9906 8256 9962
rect 8312 9906 8380 9962
rect 8436 9906 8504 9962
rect 8560 9906 8628 9962
rect 8684 9906 8752 9962
rect 8808 9906 8876 9962
rect 8932 9906 9000 9962
rect 9056 9906 9124 9962
rect 9180 9906 9248 9962
rect 9304 9906 9372 9962
rect 9428 9906 9496 9962
rect 9552 9906 9620 9962
rect 9676 9906 9744 9962
rect 9800 9906 9810 9962
rect 7874 9838 9810 9906
rect 7874 9782 7884 9838
rect 7940 9782 8008 9838
rect 8064 9782 8132 9838
rect 8188 9782 8256 9838
rect 8312 9782 8380 9838
rect 8436 9782 8504 9838
rect 8560 9782 8628 9838
rect 8684 9782 8752 9838
rect 8808 9782 8876 9838
rect 8932 9782 9000 9838
rect 9056 9782 9124 9838
rect 9180 9782 9248 9838
rect 9304 9782 9372 9838
rect 9428 9782 9496 9838
rect 9552 9782 9620 9838
rect 9676 9782 9744 9838
rect 9800 9782 9810 9838
rect 7874 9714 9810 9782
rect 7874 9658 7884 9714
rect 7940 9658 8008 9714
rect 8064 9658 8132 9714
rect 8188 9658 8256 9714
rect 8312 9658 8380 9714
rect 8436 9658 8504 9714
rect 8560 9658 8628 9714
rect 8684 9658 8752 9714
rect 8808 9658 8876 9714
rect 8932 9658 9000 9714
rect 9056 9658 9124 9714
rect 9180 9658 9248 9714
rect 9304 9658 9372 9714
rect 9428 9658 9496 9714
rect 9552 9658 9620 9714
rect 9676 9658 9744 9714
rect 9800 9658 9810 9714
rect 7874 9590 9810 9658
rect 7874 9534 7884 9590
rect 7940 9534 8008 9590
rect 8064 9534 8132 9590
rect 8188 9534 8256 9590
rect 8312 9534 8380 9590
rect 8436 9534 8504 9590
rect 8560 9534 8628 9590
rect 8684 9534 8752 9590
rect 8808 9534 8876 9590
rect 8932 9534 9000 9590
rect 9056 9534 9124 9590
rect 9180 9534 9248 9590
rect 9304 9534 9372 9590
rect 9428 9534 9496 9590
rect 9552 9534 9620 9590
rect 9676 9534 9744 9590
rect 9800 9534 9810 9590
rect 7874 9466 9810 9534
rect 7874 9410 7884 9466
rect 7940 9410 8008 9466
rect 8064 9410 8132 9466
rect 8188 9410 8256 9466
rect 8312 9410 8380 9466
rect 8436 9410 8504 9466
rect 8560 9410 8628 9466
rect 8684 9410 8752 9466
rect 8808 9410 8876 9466
rect 8932 9410 9000 9466
rect 9056 9410 9124 9466
rect 9180 9410 9248 9466
rect 9304 9410 9372 9466
rect 9428 9410 9496 9466
rect 9552 9410 9620 9466
rect 9676 9410 9744 9466
rect 9800 9410 9810 9466
rect 7874 9342 9810 9410
rect 7874 9286 7884 9342
rect 7940 9286 8008 9342
rect 8064 9286 8132 9342
rect 8188 9286 8256 9342
rect 8312 9286 8380 9342
rect 8436 9286 8504 9342
rect 8560 9286 8628 9342
rect 8684 9286 8752 9342
rect 8808 9286 8876 9342
rect 8932 9286 9000 9342
rect 9056 9286 9124 9342
rect 9180 9286 9248 9342
rect 9304 9286 9372 9342
rect 9428 9286 9496 9342
rect 9552 9286 9620 9342
rect 9676 9286 9744 9342
rect 9800 9286 9810 9342
rect 7874 9218 9810 9286
rect 7874 9162 7884 9218
rect 7940 9162 8008 9218
rect 8064 9162 8132 9218
rect 8188 9162 8256 9218
rect 8312 9162 8380 9218
rect 8436 9162 8504 9218
rect 8560 9162 8628 9218
rect 8684 9162 8752 9218
rect 8808 9162 8876 9218
rect 8932 9162 9000 9218
rect 9056 9162 9124 9218
rect 9180 9162 9248 9218
rect 9304 9162 9372 9218
rect 9428 9162 9496 9218
rect 9552 9162 9620 9218
rect 9676 9162 9744 9218
rect 9800 9162 9810 9218
rect 7874 9094 9810 9162
rect 7874 9038 7884 9094
rect 7940 9038 8008 9094
rect 8064 9038 8132 9094
rect 8188 9038 8256 9094
rect 8312 9038 8380 9094
rect 8436 9038 8504 9094
rect 8560 9038 8628 9094
rect 8684 9038 8752 9094
rect 8808 9038 8876 9094
rect 8932 9038 9000 9094
rect 9056 9038 9124 9094
rect 9180 9038 9248 9094
rect 9304 9038 9372 9094
rect 9428 9038 9496 9094
rect 9552 9038 9620 9094
rect 9676 9038 9744 9094
rect 9800 9038 9810 9094
rect 7874 8970 9810 9038
rect 7874 8914 7884 8970
rect 7940 8914 8008 8970
rect 8064 8914 8132 8970
rect 8188 8914 8256 8970
rect 8312 8914 8380 8970
rect 8436 8914 8504 8970
rect 8560 8914 8628 8970
rect 8684 8914 8752 8970
rect 8808 8914 8876 8970
rect 8932 8914 9000 8970
rect 9056 8914 9124 8970
rect 9180 8914 9248 8970
rect 9304 8914 9372 8970
rect 9428 8914 9496 8970
rect 9552 8914 9620 8970
rect 9676 8914 9744 8970
rect 9800 8914 9810 8970
rect 7874 8846 9810 8914
rect 7874 8790 7884 8846
rect 7940 8790 8008 8846
rect 8064 8790 8132 8846
rect 8188 8790 8256 8846
rect 8312 8790 8380 8846
rect 8436 8790 8504 8846
rect 8560 8790 8628 8846
rect 8684 8790 8752 8846
rect 8808 8790 8876 8846
rect 8932 8790 9000 8846
rect 9056 8790 9124 8846
rect 9180 8790 9248 8846
rect 9304 8790 9372 8846
rect 9428 8790 9496 8846
rect 9552 8790 9620 8846
rect 9676 8790 9744 8846
rect 9800 8790 9810 8846
rect 7874 8722 9810 8790
rect 7874 8666 7884 8722
rect 7940 8666 8008 8722
rect 8064 8666 8132 8722
rect 8188 8666 8256 8722
rect 8312 8666 8380 8722
rect 8436 8666 8504 8722
rect 8560 8666 8628 8722
rect 8684 8666 8752 8722
rect 8808 8666 8876 8722
rect 8932 8666 9000 8722
rect 9056 8666 9124 8722
rect 9180 8666 9248 8722
rect 9304 8666 9372 8722
rect 9428 8666 9496 8722
rect 9552 8666 9620 8722
rect 9676 8666 9744 8722
rect 9800 8666 9810 8722
rect 7874 8598 9810 8666
rect 7874 8542 7884 8598
rect 7940 8542 8008 8598
rect 8064 8542 8132 8598
rect 8188 8542 8256 8598
rect 8312 8542 8380 8598
rect 8436 8542 8504 8598
rect 8560 8542 8628 8598
rect 8684 8542 8752 8598
rect 8808 8542 8876 8598
rect 8932 8542 9000 8598
rect 9056 8542 9124 8598
rect 9180 8542 9248 8598
rect 9304 8542 9372 8598
rect 9428 8542 9496 8598
rect 9552 8542 9620 8598
rect 9676 8542 9744 8598
rect 9800 8542 9810 8598
rect 7874 8474 9810 8542
rect 7874 8418 7884 8474
rect 7940 8418 8008 8474
rect 8064 8418 8132 8474
rect 8188 8418 8256 8474
rect 8312 8418 8380 8474
rect 8436 8418 8504 8474
rect 8560 8418 8628 8474
rect 8684 8418 8752 8474
rect 8808 8418 8876 8474
rect 8932 8418 9000 8474
rect 9056 8418 9124 8474
rect 9180 8418 9248 8474
rect 9304 8418 9372 8474
rect 9428 8418 9496 8474
rect 9552 8418 9620 8474
rect 9676 8418 9744 8474
rect 9800 8418 9810 8474
rect 7874 8350 9810 8418
rect 7874 8294 7884 8350
rect 7940 8294 8008 8350
rect 8064 8294 8132 8350
rect 8188 8294 8256 8350
rect 8312 8294 8380 8350
rect 8436 8294 8504 8350
rect 8560 8294 8628 8350
rect 8684 8294 8752 8350
rect 8808 8294 8876 8350
rect 8932 8294 9000 8350
rect 9056 8294 9124 8350
rect 9180 8294 9248 8350
rect 9304 8294 9372 8350
rect 9428 8294 9496 8350
rect 9552 8294 9620 8350
rect 9676 8294 9744 8350
rect 9800 8294 9810 8350
rect 7874 8226 9810 8294
rect 7874 8170 7884 8226
rect 7940 8170 8008 8226
rect 8064 8170 8132 8226
rect 8188 8170 8256 8226
rect 8312 8170 8380 8226
rect 8436 8170 8504 8226
rect 8560 8170 8628 8226
rect 8684 8170 8752 8226
rect 8808 8170 8876 8226
rect 8932 8170 9000 8226
rect 9056 8170 9124 8226
rect 9180 8170 9248 8226
rect 9304 8170 9372 8226
rect 9428 8170 9496 8226
rect 9552 8170 9620 8226
rect 9676 8170 9744 8226
rect 9800 8170 9810 8226
rect 7874 8102 9810 8170
rect 7874 8046 7884 8102
rect 7940 8046 8008 8102
rect 8064 8046 8132 8102
rect 8188 8046 8256 8102
rect 8312 8046 8380 8102
rect 8436 8046 8504 8102
rect 8560 8046 8628 8102
rect 8684 8046 8752 8102
rect 8808 8046 8876 8102
rect 8932 8046 9000 8102
rect 9056 8046 9124 8102
rect 9180 8046 9248 8102
rect 9304 8046 9372 8102
rect 9428 8046 9496 8102
rect 9552 8046 9620 8102
rect 9676 8046 9744 8102
rect 9800 8046 9810 8102
rect 7874 8036 9810 8046
rect 10244 10954 12180 10964
rect 10244 10898 10254 10954
rect 10310 10898 10378 10954
rect 10434 10898 10502 10954
rect 10558 10898 10626 10954
rect 10682 10898 10750 10954
rect 10806 10898 10874 10954
rect 10930 10898 10998 10954
rect 11054 10898 11122 10954
rect 11178 10898 11246 10954
rect 11302 10898 11370 10954
rect 11426 10898 11494 10954
rect 11550 10898 11618 10954
rect 11674 10898 11742 10954
rect 11798 10898 11866 10954
rect 11922 10898 11990 10954
rect 12046 10898 12114 10954
rect 12170 10898 12180 10954
rect 10244 10830 12180 10898
rect 10244 10774 10254 10830
rect 10310 10774 10378 10830
rect 10434 10774 10502 10830
rect 10558 10774 10626 10830
rect 10682 10774 10750 10830
rect 10806 10774 10874 10830
rect 10930 10774 10998 10830
rect 11054 10774 11122 10830
rect 11178 10774 11246 10830
rect 11302 10774 11370 10830
rect 11426 10774 11494 10830
rect 11550 10774 11618 10830
rect 11674 10774 11742 10830
rect 11798 10774 11866 10830
rect 11922 10774 11990 10830
rect 12046 10774 12114 10830
rect 12170 10774 12180 10830
rect 10244 10706 12180 10774
rect 10244 10650 10254 10706
rect 10310 10650 10378 10706
rect 10434 10650 10502 10706
rect 10558 10650 10626 10706
rect 10682 10650 10750 10706
rect 10806 10650 10874 10706
rect 10930 10650 10998 10706
rect 11054 10650 11122 10706
rect 11178 10650 11246 10706
rect 11302 10650 11370 10706
rect 11426 10650 11494 10706
rect 11550 10650 11618 10706
rect 11674 10650 11742 10706
rect 11798 10650 11866 10706
rect 11922 10650 11990 10706
rect 12046 10650 12114 10706
rect 12170 10650 12180 10706
rect 10244 10582 12180 10650
rect 10244 10526 10254 10582
rect 10310 10526 10378 10582
rect 10434 10526 10502 10582
rect 10558 10526 10626 10582
rect 10682 10526 10750 10582
rect 10806 10526 10874 10582
rect 10930 10526 10998 10582
rect 11054 10526 11122 10582
rect 11178 10526 11246 10582
rect 11302 10526 11370 10582
rect 11426 10526 11494 10582
rect 11550 10526 11618 10582
rect 11674 10526 11742 10582
rect 11798 10526 11866 10582
rect 11922 10526 11990 10582
rect 12046 10526 12114 10582
rect 12170 10526 12180 10582
rect 10244 10458 12180 10526
rect 10244 10402 10254 10458
rect 10310 10402 10378 10458
rect 10434 10402 10502 10458
rect 10558 10402 10626 10458
rect 10682 10402 10750 10458
rect 10806 10402 10874 10458
rect 10930 10402 10998 10458
rect 11054 10402 11122 10458
rect 11178 10402 11246 10458
rect 11302 10402 11370 10458
rect 11426 10402 11494 10458
rect 11550 10402 11618 10458
rect 11674 10402 11742 10458
rect 11798 10402 11866 10458
rect 11922 10402 11990 10458
rect 12046 10402 12114 10458
rect 12170 10402 12180 10458
rect 10244 10334 12180 10402
rect 10244 10278 10254 10334
rect 10310 10278 10378 10334
rect 10434 10278 10502 10334
rect 10558 10278 10626 10334
rect 10682 10278 10750 10334
rect 10806 10278 10874 10334
rect 10930 10278 10998 10334
rect 11054 10278 11122 10334
rect 11178 10278 11246 10334
rect 11302 10278 11370 10334
rect 11426 10278 11494 10334
rect 11550 10278 11618 10334
rect 11674 10278 11742 10334
rect 11798 10278 11866 10334
rect 11922 10278 11990 10334
rect 12046 10278 12114 10334
rect 12170 10278 12180 10334
rect 10244 10210 12180 10278
rect 10244 10154 10254 10210
rect 10310 10154 10378 10210
rect 10434 10154 10502 10210
rect 10558 10154 10626 10210
rect 10682 10154 10750 10210
rect 10806 10154 10874 10210
rect 10930 10154 10998 10210
rect 11054 10154 11122 10210
rect 11178 10154 11246 10210
rect 11302 10154 11370 10210
rect 11426 10154 11494 10210
rect 11550 10154 11618 10210
rect 11674 10154 11742 10210
rect 11798 10154 11866 10210
rect 11922 10154 11990 10210
rect 12046 10154 12114 10210
rect 12170 10154 12180 10210
rect 10244 10086 12180 10154
rect 10244 10030 10254 10086
rect 10310 10030 10378 10086
rect 10434 10030 10502 10086
rect 10558 10030 10626 10086
rect 10682 10030 10750 10086
rect 10806 10030 10874 10086
rect 10930 10030 10998 10086
rect 11054 10030 11122 10086
rect 11178 10030 11246 10086
rect 11302 10030 11370 10086
rect 11426 10030 11494 10086
rect 11550 10030 11618 10086
rect 11674 10030 11742 10086
rect 11798 10030 11866 10086
rect 11922 10030 11990 10086
rect 12046 10030 12114 10086
rect 12170 10030 12180 10086
rect 10244 9962 12180 10030
rect 10244 9906 10254 9962
rect 10310 9906 10378 9962
rect 10434 9906 10502 9962
rect 10558 9906 10626 9962
rect 10682 9906 10750 9962
rect 10806 9906 10874 9962
rect 10930 9906 10998 9962
rect 11054 9906 11122 9962
rect 11178 9906 11246 9962
rect 11302 9906 11370 9962
rect 11426 9906 11494 9962
rect 11550 9906 11618 9962
rect 11674 9906 11742 9962
rect 11798 9906 11866 9962
rect 11922 9906 11990 9962
rect 12046 9906 12114 9962
rect 12170 9906 12180 9962
rect 10244 9838 12180 9906
rect 10244 9782 10254 9838
rect 10310 9782 10378 9838
rect 10434 9782 10502 9838
rect 10558 9782 10626 9838
rect 10682 9782 10750 9838
rect 10806 9782 10874 9838
rect 10930 9782 10998 9838
rect 11054 9782 11122 9838
rect 11178 9782 11246 9838
rect 11302 9782 11370 9838
rect 11426 9782 11494 9838
rect 11550 9782 11618 9838
rect 11674 9782 11742 9838
rect 11798 9782 11866 9838
rect 11922 9782 11990 9838
rect 12046 9782 12114 9838
rect 12170 9782 12180 9838
rect 10244 9714 12180 9782
rect 10244 9658 10254 9714
rect 10310 9658 10378 9714
rect 10434 9658 10502 9714
rect 10558 9658 10626 9714
rect 10682 9658 10750 9714
rect 10806 9658 10874 9714
rect 10930 9658 10998 9714
rect 11054 9658 11122 9714
rect 11178 9658 11246 9714
rect 11302 9658 11370 9714
rect 11426 9658 11494 9714
rect 11550 9658 11618 9714
rect 11674 9658 11742 9714
rect 11798 9658 11866 9714
rect 11922 9658 11990 9714
rect 12046 9658 12114 9714
rect 12170 9658 12180 9714
rect 10244 9590 12180 9658
rect 10244 9534 10254 9590
rect 10310 9534 10378 9590
rect 10434 9534 10502 9590
rect 10558 9534 10626 9590
rect 10682 9534 10750 9590
rect 10806 9534 10874 9590
rect 10930 9534 10998 9590
rect 11054 9534 11122 9590
rect 11178 9534 11246 9590
rect 11302 9534 11370 9590
rect 11426 9534 11494 9590
rect 11550 9534 11618 9590
rect 11674 9534 11742 9590
rect 11798 9534 11866 9590
rect 11922 9534 11990 9590
rect 12046 9534 12114 9590
rect 12170 9534 12180 9590
rect 10244 9466 12180 9534
rect 10244 9410 10254 9466
rect 10310 9410 10378 9466
rect 10434 9410 10502 9466
rect 10558 9410 10626 9466
rect 10682 9410 10750 9466
rect 10806 9410 10874 9466
rect 10930 9410 10998 9466
rect 11054 9410 11122 9466
rect 11178 9410 11246 9466
rect 11302 9410 11370 9466
rect 11426 9410 11494 9466
rect 11550 9410 11618 9466
rect 11674 9410 11742 9466
rect 11798 9410 11866 9466
rect 11922 9410 11990 9466
rect 12046 9410 12114 9466
rect 12170 9410 12180 9466
rect 10244 9342 12180 9410
rect 10244 9286 10254 9342
rect 10310 9286 10378 9342
rect 10434 9286 10502 9342
rect 10558 9286 10626 9342
rect 10682 9286 10750 9342
rect 10806 9286 10874 9342
rect 10930 9286 10998 9342
rect 11054 9286 11122 9342
rect 11178 9286 11246 9342
rect 11302 9286 11370 9342
rect 11426 9286 11494 9342
rect 11550 9286 11618 9342
rect 11674 9286 11742 9342
rect 11798 9286 11866 9342
rect 11922 9286 11990 9342
rect 12046 9286 12114 9342
rect 12170 9286 12180 9342
rect 10244 9218 12180 9286
rect 10244 9162 10254 9218
rect 10310 9162 10378 9218
rect 10434 9162 10502 9218
rect 10558 9162 10626 9218
rect 10682 9162 10750 9218
rect 10806 9162 10874 9218
rect 10930 9162 10998 9218
rect 11054 9162 11122 9218
rect 11178 9162 11246 9218
rect 11302 9162 11370 9218
rect 11426 9162 11494 9218
rect 11550 9162 11618 9218
rect 11674 9162 11742 9218
rect 11798 9162 11866 9218
rect 11922 9162 11990 9218
rect 12046 9162 12114 9218
rect 12170 9162 12180 9218
rect 10244 9094 12180 9162
rect 10244 9038 10254 9094
rect 10310 9038 10378 9094
rect 10434 9038 10502 9094
rect 10558 9038 10626 9094
rect 10682 9038 10750 9094
rect 10806 9038 10874 9094
rect 10930 9038 10998 9094
rect 11054 9038 11122 9094
rect 11178 9038 11246 9094
rect 11302 9038 11370 9094
rect 11426 9038 11494 9094
rect 11550 9038 11618 9094
rect 11674 9038 11742 9094
rect 11798 9038 11866 9094
rect 11922 9038 11990 9094
rect 12046 9038 12114 9094
rect 12170 9038 12180 9094
rect 10244 8970 12180 9038
rect 10244 8914 10254 8970
rect 10310 8914 10378 8970
rect 10434 8914 10502 8970
rect 10558 8914 10626 8970
rect 10682 8914 10750 8970
rect 10806 8914 10874 8970
rect 10930 8914 10998 8970
rect 11054 8914 11122 8970
rect 11178 8914 11246 8970
rect 11302 8914 11370 8970
rect 11426 8914 11494 8970
rect 11550 8914 11618 8970
rect 11674 8914 11742 8970
rect 11798 8914 11866 8970
rect 11922 8914 11990 8970
rect 12046 8914 12114 8970
rect 12170 8914 12180 8970
rect 10244 8846 12180 8914
rect 10244 8790 10254 8846
rect 10310 8790 10378 8846
rect 10434 8790 10502 8846
rect 10558 8790 10626 8846
rect 10682 8790 10750 8846
rect 10806 8790 10874 8846
rect 10930 8790 10998 8846
rect 11054 8790 11122 8846
rect 11178 8790 11246 8846
rect 11302 8790 11370 8846
rect 11426 8790 11494 8846
rect 11550 8790 11618 8846
rect 11674 8790 11742 8846
rect 11798 8790 11866 8846
rect 11922 8790 11990 8846
rect 12046 8790 12114 8846
rect 12170 8790 12180 8846
rect 10244 8722 12180 8790
rect 10244 8666 10254 8722
rect 10310 8666 10378 8722
rect 10434 8666 10502 8722
rect 10558 8666 10626 8722
rect 10682 8666 10750 8722
rect 10806 8666 10874 8722
rect 10930 8666 10998 8722
rect 11054 8666 11122 8722
rect 11178 8666 11246 8722
rect 11302 8666 11370 8722
rect 11426 8666 11494 8722
rect 11550 8666 11618 8722
rect 11674 8666 11742 8722
rect 11798 8666 11866 8722
rect 11922 8666 11990 8722
rect 12046 8666 12114 8722
rect 12170 8666 12180 8722
rect 10244 8598 12180 8666
rect 10244 8542 10254 8598
rect 10310 8542 10378 8598
rect 10434 8542 10502 8598
rect 10558 8542 10626 8598
rect 10682 8542 10750 8598
rect 10806 8542 10874 8598
rect 10930 8542 10998 8598
rect 11054 8542 11122 8598
rect 11178 8542 11246 8598
rect 11302 8542 11370 8598
rect 11426 8542 11494 8598
rect 11550 8542 11618 8598
rect 11674 8542 11742 8598
rect 11798 8542 11866 8598
rect 11922 8542 11990 8598
rect 12046 8542 12114 8598
rect 12170 8542 12180 8598
rect 10244 8474 12180 8542
rect 10244 8418 10254 8474
rect 10310 8418 10378 8474
rect 10434 8418 10502 8474
rect 10558 8418 10626 8474
rect 10682 8418 10750 8474
rect 10806 8418 10874 8474
rect 10930 8418 10998 8474
rect 11054 8418 11122 8474
rect 11178 8418 11246 8474
rect 11302 8418 11370 8474
rect 11426 8418 11494 8474
rect 11550 8418 11618 8474
rect 11674 8418 11742 8474
rect 11798 8418 11866 8474
rect 11922 8418 11990 8474
rect 12046 8418 12114 8474
rect 12170 8418 12180 8474
rect 10244 8350 12180 8418
rect 10244 8294 10254 8350
rect 10310 8294 10378 8350
rect 10434 8294 10502 8350
rect 10558 8294 10626 8350
rect 10682 8294 10750 8350
rect 10806 8294 10874 8350
rect 10930 8294 10998 8350
rect 11054 8294 11122 8350
rect 11178 8294 11246 8350
rect 11302 8294 11370 8350
rect 11426 8294 11494 8350
rect 11550 8294 11618 8350
rect 11674 8294 11742 8350
rect 11798 8294 11866 8350
rect 11922 8294 11990 8350
rect 12046 8294 12114 8350
rect 12170 8294 12180 8350
rect 10244 8226 12180 8294
rect 10244 8170 10254 8226
rect 10310 8170 10378 8226
rect 10434 8170 10502 8226
rect 10558 8170 10626 8226
rect 10682 8170 10750 8226
rect 10806 8170 10874 8226
rect 10930 8170 10998 8226
rect 11054 8170 11122 8226
rect 11178 8170 11246 8226
rect 11302 8170 11370 8226
rect 11426 8170 11494 8226
rect 11550 8170 11618 8226
rect 11674 8170 11742 8226
rect 11798 8170 11866 8226
rect 11922 8170 11990 8226
rect 12046 8170 12114 8226
rect 12170 8170 12180 8226
rect 10244 8102 12180 8170
rect 10244 8046 10254 8102
rect 10310 8046 10378 8102
rect 10434 8046 10502 8102
rect 10558 8046 10626 8102
rect 10682 8046 10750 8102
rect 10806 8046 10874 8102
rect 10930 8046 10998 8102
rect 11054 8046 11122 8102
rect 11178 8046 11246 8102
rect 11302 8046 11370 8102
rect 11426 8046 11494 8102
rect 11550 8046 11618 8102
rect 11674 8046 11742 8102
rect 11798 8046 11866 8102
rect 11922 8046 11990 8102
rect 12046 8046 12114 8102
rect 12170 8046 12180 8102
rect 10244 8036 12180 8046
rect 12861 10954 14673 10964
rect 12861 10898 12871 10954
rect 12927 10898 12995 10954
rect 13051 10898 13119 10954
rect 13175 10898 13243 10954
rect 13299 10898 13367 10954
rect 13423 10898 13491 10954
rect 13547 10898 13615 10954
rect 13671 10898 13739 10954
rect 13795 10898 13863 10954
rect 13919 10898 13987 10954
rect 14043 10898 14111 10954
rect 14167 10898 14235 10954
rect 14291 10898 14359 10954
rect 14415 10898 14483 10954
rect 14539 10898 14607 10954
rect 14663 10898 14673 10954
rect 12861 10830 14673 10898
rect 12861 10774 12871 10830
rect 12927 10774 12995 10830
rect 13051 10774 13119 10830
rect 13175 10774 13243 10830
rect 13299 10774 13367 10830
rect 13423 10774 13491 10830
rect 13547 10774 13615 10830
rect 13671 10774 13739 10830
rect 13795 10774 13863 10830
rect 13919 10774 13987 10830
rect 14043 10774 14111 10830
rect 14167 10774 14235 10830
rect 14291 10774 14359 10830
rect 14415 10774 14483 10830
rect 14539 10774 14607 10830
rect 14663 10774 14673 10830
rect 12861 10706 14673 10774
rect 12861 10650 12871 10706
rect 12927 10650 12995 10706
rect 13051 10650 13119 10706
rect 13175 10650 13243 10706
rect 13299 10650 13367 10706
rect 13423 10650 13491 10706
rect 13547 10650 13615 10706
rect 13671 10650 13739 10706
rect 13795 10650 13863 10706
rect 13919 10650 13987 10706
rect 14043 10650 14111 10706
rect 14167 10650 14235 10706
rect 14291 10650 14359 10706
rect 14415 10650 14483 10706
rect 14539 10650 14607 10706
rect 14663 10650 14673 10706
rect 12861 10582 14673 10650
rect 12861 10526 12871 10582
rect 12927 10526 12995 10582
rect 13051 10526 13119 10582
rect 13175 10526 13243 10582
rect 13299 10526 13367 10582
rect 13423 10526 13491 10582
rect 13547 10526 13615 10582
rect 13671 10526 13739 10582
rect 13795 10526 13863 10582
rect 13919 10526 13987 10582
rect 14043 10526 14111 10582
rect 14167 10526 14235 10582
rect 14291 10526 14359 10582
rect 14415 10526 14483 10582
rect 14539 10526 14607 10582
rect 14663 10526 14673 10582
rect 12861 10458 14673 10526
rect 12861 10402 12871 10458
rect 12927 10402 12995 10458
rect 13051 10402 13119 10458
rect 13175 10402 13243 10458
rect 13299 10402 13367 10458
rect 13423 10402 13491 10458
rect 13547 10402 13615 10458
rect 13671 10402 13739 10458
rect 13795 10402 13863 10458
rect 13919 10402 13987 10458
rect 14043 10402 14111 10458
rect 14167 10402 14235 10458
rect 14291 10402 14359 10458
rect 14415 10402 14483 10458
rect 14539 10402 14607 10458
rect 14663 10402 14673 10458
rect 12861 10334 14673 10402
rect 12861 10278 12871 10334
rect 12927 10278 12995 10334
rect 13051 10278 13119 10334
rect 13175 10278 13243 10334
rect 13299 10278 13367 10334
rect 13423 10278 13491 10334
rect 13547 10278 13615 10334
rect 13671 10278 13739 10334
rect 13795 10278 13863 10334
rect 13919 10278 13987 10334
rect 14043 10278 14111 10334
rect 14167 10278 14235 10334
rect 14291 10278 14359 10334
rect 14415 10278 14483 10334
rect 14539 10278 14607 10334
rect 14663 10278 14673 10334
rect 12861 10210 14673 10278
rect 12861 10154 12871 10210
rect 12927 10154 12995 10210
rect 13051 10154 13119 10210
rect 13175 10154 13243 10210
rect 13299 10154 13367 10210
rect 13423 10154 13491 10210
rect 13547 10154 13615 10210
rect 13671 10154 13739 10210
rect 13795 10154 13863 10210
rect 13919 10154 13987 10210
rect 14043 10154 14111 10210
rect 14167 10154 14235 10210
rect 14291 10154 14359 10210
rect 14415 10154 14483 10210
rect 14539 10154 14607 10210
rect 14663 10154 14673 10210
rect 12861 10086 14673 10154
rect 12861 10030 12871 10086
rect 12927 10030 12995 10086
rect 13051 10030 13119 10086
rect 13175 10030 13243 10086
rect 13299 10030 13367 10086
rect 13423 10030 13491 10086
rect 13547 10030 13615 10086
rect 13671 10030 13739 10086
rect 13795 10030 13863 10086
rect 13919 10030 13987 10086
rect 14043 10030 14111 10086
rect 14167 10030 14235 10086
rect 14291 10030 14359 10086
rect 14415 10030 14483 10086
rect 14539 10030 14607 10086
rect 14663 10030 14673 10086
rect 12861 9962 14673 10030
rect 12861 9906 12871 9962
rect 12927 9906 12995 9962
rect 13051 9906 13119 9962
rect 13175 9906 13243 9962
rect 13299 9906 13367 9962
rect 13423 9906 13491 9962
rect 13547 9906 13615 9962
rect 13671 9906 13739 9962
rect 13795 9906 13863 9962
rect 13919 9906 13987 9962
rect 14043 9906 14111 9962
rect 14167 9906 14235 9962
rect 14291 9906 14359 9962
rect 14415 9906 14483 9962
rect 14539 9906 14607 9962
rect 14663 9906 14673 9962
rect 12861 9838 14673 9906
rect 12861 9782 12871 9838
rect 12927 9782 12995 9838
rect 13051 9782 13119 9838
rect 13175 9782 13243 9838
rect 13299 9782 13367 9838
rect 13423 9782 13491 9838
rect 13547 9782 13615 9838
rect 13671 9782 13739 9838
rect 13795 9782 13863 9838
rect 13919 9782 13987 9838
rect 14043 9782 14111 9838
rect 14167 9782 14235 9838
rect 14291 9782 14359 9838
rect 14415 9782 14483 9838
rect 14539 9782 14607 9838
rect 14663 9782 14673 9838
rect 12861 9714 14673 9782
rect 12861 9658 12871 9714
rect 12927 9658 12995 9714
rect 13051 9658 13119 9714
rect 13175 9658 13243 9714
rect 13299 9658 13367 9714
rect 13423 9658 13491 9714
rect 13547 9658 13615 9714
rect 13671 9658 13739 9714
rect 13795 9658 13863 9714
rect 13919 9658 13987 9714
rect 14043 9658 14111 9714
rect 14167 9658 14235 9714
rect 14291 9658 14359 9714
rect 14415 9658 14483 9714
rect 14539 9658 14607 9714
rect 14663 9658 14673 9714
rect 12861 9590 14673 9658
rect 12861 9534 12871 9590
rect 12927 9534 12995 9590
rect 13051 9534 13119 9590
rect 13175 9534 13243 9590
rect 13299 9534 13367 9590
rect 13423 9534 13491 9590
rect 13547 9534 13615 9590
rect 13671 9534 13739 9590
rect 13795 9534 13863 9590
rect 13919 9534 13987 9590
rect 14043 9534 14111 9590
rect 14167 9534 14235 9590
rect 14291 9534 14359 9590
rect 14415 9534 14483 9590
rect 14539 9534 14607 9590
rect 14663 9534 14673 9590
rect 12861 9466 14673 9534
rect 12861 9410 12871 9466
rect 12927 9410 12995 9466
rect 13051 9410 13119 9466
rect 13175 9410 13243 9466
rect 13299 9410 13367 9466
rect 13423 9410 13491 9466
rect 13547 9410 13615 9466
rect 13671 9410 13739 9466
rect 13795 9410 13863 9466
rect 13919 9410 13987 9466
rect 14043 9410 14111 9466
rect 14167 9410 14235 9466
rect 14291 9410 14359 9466
rect 14415 9410 14483 9466
rect 14539 9410 14607 9466
rect 14663 9410 14673 9466
rect 12861 9342 14673 9410
rect 12861 9286 12871 9342
rect 12927 9286 12995 9342
rect 13051 9286 13119 9342
rect 13175 9286 13243 9342
rect 13299 9286 13367 9342
rect 13423 9286 13491 9342
rect 13547 9286 13615 9342
rect 13671 9286 13739 9342
rect 13795 9286 13863 9342
rect 13919 9286 13987 9342
rect 14043 9286 14111 9342
rect 14167 9286 14235 9342
rect 14291 9286 14359 9342
rect 14415 9286 14483 9342
rect 14539 9286 14607 9342
rect 14663 9286 14673 9342
rect 12861 9218 14673 9286
rect 12861 9162 12871 9218
rect 12927 9162 12995 9218
rect 13051 9162 13119 9218
rect 13175 9162 13243 9218
rect 13299 9162 13367 9218
rect 13423 9162 13491 9218
rect 13547 9162 13615 9218
rect 13671 9162 13739 9218
rect 13795 9162 13863 9218
rect 13919 9162 13987 9218
rect 14043 9162 14111 9218
rect 14167 9162 14235 9218
rect 14291 9162 14359 9218
rect 14415 9162 14483 9218
rect 14539 9162 14607 9218
rect 14663 9162 14673 9218
rect 12861 9094 14673 9162
rect 12861 9038 12871 9094
rect 12927 9038 12995 9094
rect 13051 9038 13119 9094
rect 13175 9038 13243 9094
rect 13299 9038 13367 9094
rect 13423 9038 13491 9094
rect 13547 9038 13615 9094
rect 13671 9038 13739 9094
rect 13795 9038 13863 9094
rect 13919 9038 13987 9094
rect 14043 9038 14111 9094
rect 14167 9038 14235 9094
rect 14291 9038 14359 9094
rect 14415 9038 14483 9094
rect 14539 9038 14607 9094
rect 14663 9038 14673 9094
rect 12861 8970 14673 9038
rect 12861 8914 12871 8970
rect 12927 8914 12995 8970
rect 13051 8914 13119 8970
rect 13175 8914 13243 8970
rect 13299 8914 13367 8970
rect 13423 8914 13491 8970
rect 13547 8914 13615 8970
rect 13671 8914 13739 8970
rect 13795 8914 13863 8970
rect 13919 8914 13987 8970
rect 14043 8914 14111 8970
rect 14167 8914 14235 8970
rect 14291 8914 14359 8970
rect 14415 8914 14483 8970
rect 14539 8914 14607 8970
rect 14663 8914 14673 8970
rect 12861 8846 14673 8914
rect 12861 8790 12871 8846
rect 12927 8790 12995 8846
rect 13051 8790 13119 8846
rect 13175 8790 13243 8846
rect 13299 8790 13367 8846
rect 13423 8790 13491 8846
rect 13547 8790 13615 8846
rect 13671 8790 13739 8846
rect 13795 8790 13863 8846
rect 13919 8790 13987 8846
rect 14043 8790 14111 8846
rect 14167 8790 14235 8846
rect 14291 8790 14359 8846
rect 14415 8790 14483 8846
rect 14539 8790 14607 8846
rect 14663 8790 14673 8846
rect 12861 8722 14673 8790
rect 12861 8666 12871 8722
rect 12927 8666 12995 8722
rect 13051 8666 13119 8722
rect 13175 8666 13243 8722
rect 13299 8666 13367 8722
rect 13423 8666 13491 8722
rect 13547 8666 13615 8722
rect 13671 8666 13739 8722
rect 13795 8666 13863 8722
rect 13919 8666 13987 8722
rect 14043 8666 14111 8722
rect 14167 8666 14235 8722
rect 14291 8666 14359 8722
rect 14415 8666 14483 8722
rect 14539 8666 14607 8722
rect 14663 8666 14673 8722
rect 12861 8598 14673 8666
rect 12861 8542 12871 8598
rect 12927 8542 12995 8598
rect 13051 8542 13119 8598
rect 13175 8542 13243 8598
rect 13299 8542 13367 8598
rect 13423 8542 13491 8598
rect 13547 8542 13615 8598
rect 13671 8542 13739 8598
rect 13795 8542 13863 8598
rect 13919 8542 13987 8598
rect 14043 8542 14111 8598
rect 14167 8542 14235 8598
rect 14291 8542 14359 8598
rect 14415 8542 14483 8598
rect 14539 8542 14607 8598
rect 14663 8542 14673 8598
rect 12861 8474 14673 8542
rect 12861 8418 12871 8474
rect 12927 8418 12995 8474
rect 13051 8418 13119 8474
rect 13175 8418 13243 8474
rect 13299 8418 13367 8474
rect 13423 8418 13491 8474
rect 13547 8418 13615 8474
rect 13671 8418 13739 8474
rect 13795 8418 13863 8474
rect 13919 8418 13987 8474
rect 14043 8418 14111 8474
rect 14167 8418 14235 8474
rect 14291 8418 14359 8474
rect 14415 8418 14483 8474
rect 14539 8418 14607 8474
rect 14663 8418 14673 8474
rect 12861 8350 14673 8418
rect 12861 8294 12871 8350
rect 12927 8294 12995 8350
rect 13051 8294 13119 8350
rect 13175 8294 13243 8350
rect 13299 8294 13367 8350
rect 13423 8294 13491 8350
rect 13547 8294 13615 8350
rect 13671 8294 13739 8350
rect 13795 8294 13863 8350
rect 13919 8294 13987 8350
rect 14043 8294 14111 8350
rect 14167 8294 14235 8350
rect 14291 8294 14359 8350
rect 14415 8294 14483 8350
rect 14539 8294 14607 8350
rect 14663 8294 14673 8350
rect 12861 8226 14673 8294
rect 12861 8170 12871 8226
rect 12927 8170 12995 8226
rect 13051 8170 13119 8226
rect 13175 8170 13243 8226
rect 13299 8170 13367 8226
rect 13423 8170 13491 8226
rect 13547 8170 13615 8226
rect 13671 8170 13739 8226
rect 13795 8170 13863 8226
rect 13919 8170 13987 8226
rect 14043 8170 14111 8226
rect 14167 8170 14235 8226
rect 14291 8170 14359 8226
rect 14415 8170 14483 8226
rect 14539 8170 14607 8226
rect 14663 8170 14673 8226
rect 12861 8102 14673 8170
rect 12861 8046 12871 8102
rect 12927 8046 12995 8102
rect 13051 8046 13119 8102
rect 13175 8046 13243 8102
rect 13299 8046 13367 8102
rect 13423 8046 13491 8102
rect 13547 8046 13615 8102
rect 13671 8046 13739 8102
rect 13795 8046 13863 8102
rect 13919 8046 13987 8102
rect 14043 8046 14111 8102
rect 14167 8046 14235 8102
rect 14291 8046 14359 8102
rect 14415 8046 14483 8102
rect 14539 8046 14607 8102
rect 14663 8046 14673 8102
rect 12861 8036 14673 8046
rect 10 8004 86 8014
rect 14892 8014 14902 10986
rect 14958 8014 14968 10986
rect 14892 8004 14968 8014
rect 10 7786 86 7796
rect 10 4814 20 7786
rect 76 4814 86 7786
rect 14892 7786 14968 7796
rect 305 7754 2117 7764
rect 305 7698 315 7754
rect 371 7698 439 7754
rect 495 7698 563 7754
rect 619 7698 687 7754
rect 743 7698 811 7754
rect 867 7698 935 7754
rect 991 7698 1059 7754
rect 1115 7698 1183 7754
rect 1239 7698 1307 7754
rect 1363 7698 1431 7754
rect 1487 7698 1555 7754
rect 1611 7698 1679 7754
rect 1735 7698 1803 7754
rect 1859 7698 1927 7754
rect 1983 7698 2051 7754
rect 2107 7698 2117 7754
rect 305 7630 2117 7698
rect 305 7574 315 7630
rect 371 7574 439 7630
rect 495 7574 563 7630
rect 619 7574 687 7630
rect 743 7574 811 7630
rect 867 7574 935 7630
rect 991 7574 1059 7630
rect 1115 7574 1183 7630
rect 1239 7574 1307 7630
rect 1363 7574 1431 7630
rect 1487 7574 1555 7630
rect 1611 7574 1679 7630
rect 1735 7574 1803 7630
rect 1859 7574 1927 7630
rect 1983 7574 2051 7630
rect 2107 7574 2117 7630
rect 305 7506 2117 7574
rect 305 7450 315 7506
rect 371 7450 439 7506
rect 495 7450 563 7506
rect 619 7450 687 7506
rect 743 7450 811 7506
rect 867 7450 935 7506
rect 991 7450 1059 7506
rect 1115 7450 1183 7506
rect 1239 7450 1307 7506
rect 1363 7450 1431 7506
rect 1487 7450 1555 7506
rect 1611 7450 1679 7506
rect 1735 7450 1803 7506
rect 1859 7450 1927 7506
rect 1983 7450 2051 7506
rect 2107 7450 2117 7506
rect 305 7382 2117 7450
rect 305 7326 315 7382
rect 371 7326 439 7382
rect 495 7326 563 7382
rect 619 7326 687 7382
rect 743 7326 811 7382
rect 867 7326 935 7382
rect 991 7326 1059 7382
rect 1115 7326 1183 7382
rect 1239 7326 1307 7382
rect 1363 7326 1431 7382
rect 1487 7326 1555 7382
rect 1611 7326 1679 7382
rect 1735 7326 1803 7382
rect 1859 7326 1927 7382
rect 1983 7326 2051 7382
rect 2107 7326 2117 7382
rect 305 7258 2117 7326
rect 305 7202 315 7258
rect 371 7202 439 7258
rect 495 7202 563 7258
rect 619 7202 687 7258
rect 743 7202 811 7258
rect 867 7202 935 7258
rect 991 7202 1059 7258
rect 1115 7202 1183 7258
rect 1239 7202 1307 7258
rect 1363 7202 1431 7258
rect 1487 7202 1555 7258
rect 1611 7202 1679 7258
rect 1735 7202 1803 7258
rect 1859 7202 1927 7258
rect 1983 7202 2051 7258
rect 2107 7202 2117 7258
rect 305 7134 2117 7202
rect 305 7078 315 7134
rect 371 7078 439 7134
rect 495 7078 563 7134
rect 619 7078 687 7134
rect 743 7078 811 7134
rect 867 7078 935 7134
rect 991 7078 1059 7134
rect 1115 7078 1183 7134
rect 1239 7078 1307 7134
rect 1363 7078 1431 7134
rect 1487 7078 1555 7134
rect 1611 7078 1679 7134
rect 1735 7078 1803 7134
rect 1859 7078 1927 7134
rect 1983 7078 2051 7134
rect 2107 7078 2117 7134
rect 305 7010 2117 7078
rect 305 6954 315 7010
rect 371 6954 439 7010
rect 495 6954 563 7010
rect 619 6954 687 7010
rect 743 6954 811 7010
rect 867 6954 935 7010
rect 991 6954 1059 7010
rect 1115 6954 1183 7010
rect 1239 6954 1307 7010
rect 1363 6954 1431 7010
rect 1487 6954 1555 7010
rect 1611 6954 1679 7010
rect 1735 6954 1803 7010
rect 1859 6954 1927 7010
rect 1983 6954 2051 7010
rect 2107 6954 2117 7010
rect 305 6886 2117 6954
rect 305 6830 315 6886
rect 371 6830 439 6886
rect 495 6830 563 6886
rect 619 6830 687 6886
rect 743 6830 811 6886
rect 867 6830 935 6886
rect 991 6830 1059 6886
rect 1115 6830 1183 6886
rect 1239 6830 1307 6886
rect 1363 6830 1431 6886
rect 1487 6830 1555 6886
rect 1611 6830 1679 6886
rect 1735 6830 1803 6886
rect 1859 6830 1927 6886
rect 1983 6830 2051 6886
rect 2107 6830 2117 6886
rect 305 6762 2117 6830
rect 305 6706 315 6762
rect 371 6706 439 6762
rect 495 6706 563 6762
rect 619 6706 687 6762
rect 743 6706 811 6762
rect 867 6706 935 6762
rect 991 6706 1059 6762
rect 1115 6706 1183 6762
rect 1239 6706 1307 6762
rect 1363 6706 1431 6762
rect 1487 6706 1555 6762
rect 1611 6706 1679 6762
rect 1735 6706 1803 6762
rect 1859 6706 1927 6762
rect 1983 6706 2051 6762
rect 2107 6706 2117 6762
rect 305 6638 2117 6706
rect 305 6582 315 6638
rect 371 6582 439 6638
rect 495 6582 563 6638
rect 619 6582 687 6638
rect 743 6582 811 6638
rect 867 6582 935 6638
rect 991 6582 1059 6638
rect 1115 6582 1183 6638
rect 1239 6582 1307 6638
rect 1363 6582 1431 6638
rect 1487 6582 1555 6638
rect 1611 6582 1679 6638
rect 1735 6582 1803 6638
rect 1859 6582 1927 6638
rect 1983 6582 2051 6638
rect 2107 6582 2117 6638
rect 305 6514 2117 6582
rect 305 6458 315 6514
rect 371 6458 439 6514
rect 495 6458 563 6514
rect 619 6458 687 6514
rect 743 6458 811 6514
rect 867 6458 935 6514
rect 991 6458 1059 6514
rect 1115 6458 1183 6514
rect 1239 6458 1307 6514
rect 1363 6458 1431 6514
rect 1487 6458 1555 6514
rect 1611 6458 1679 6514
rect 1735 6458 1803 6514
rect 1859 6458 1927 6514
rect 1983 6458 2051 6514
rect 2107 6458 2117 6514
rect 305 6390 2117 6458
rect 305 6334 315 6390
rect 371 6334 439 6390
rect 495 6334 563 6390
rect 619 6334 687 6390
rect 743 6334 811 6390
rect 867 6334 935 6390
rect 991 6334 1059 6390
rect 1115 6334 1183 6390
rect 1239 6334 1307 6390
rect 1363 6334 1431 6390
rect 1487 6334 1555 6390
rect 1611 6334 1679 6390
rect 1735 6334 1803 6390
rect 1859 6334 1927 6390
rect 1983 6334 2051 6390
rect 2107 6334 2117 6390
rect 305 6266 2117 6334
rect 305 6210 315 6266
rect 371 6210 439 6266
rect 495 6210 563 6266
rect 619 6210 687 6266
rect 743 6210 811 6266
rect 867 6210 935 6266
rect 991 6210 1059 6266
rect 1115 6210 1183 6266
rect 1239 6210 1307 6266
rect 1363 6210 1431 6266
rect 1487 6210 1555 6266
rect 1611 6210 1679 6266
rect 1735 6210 1803 6266
rect 1859 6210 1927 6266
rect 1983 6210 2051 6266
rect 2107 6210 2117 6266
rect 305 6142 2117 6210
rect 305 6086 315 6142
rect 371 6086 439 6142
rect 495 6086 563 6142
rect 619 6086 687 6142
rect 743 6086 811 6142
rect 867 6086 935 6142
rect 991 6086 1059 6142
rect 1115 6086 1183 6142
rect 1239 6086 1307 6142
rect 1363 6086 1431 6142
rect 1487 6086 1555 6142
rect 1611 6086 1679 6142
rect 1735 6086 1803 6142
rect 1859 6086 1927 6142
rect 1983 6086 2051 6142
rect 2107 6086 2117 6142
rect 305 6018 2117 6086
rect 305 5962 315 6018
rect 371 5962 439 6018
rect 495 5962 563 6018
rect 619 5962 687 6018
rect 743 5962 811 6018
rect 867 5962 935 6018
rect 991 5962 1059 6018
rect 1115 5962 1183 6018
rect 1239 5962 1307 6018
rect 1363 5962 1431 6018
rect 1487 5962 1555 6018
rect 1611 5962 1679 6018
rect 1735 5962 1803 6018
rect 1859 5962 1927 6018
rect 1983 5962 2051 6018
rect 2107 5962 2117 6018
rect 305 5894 2117 5962
rect 305 5838 315 5894
rect 371 5838 439 5894
rect 495 5838 563 5894
rect 619 5838 687 5894
rect 743 5838 811 5894
rect 867 5838 935 5894
rect 991 5838 1059 5894
rect 1115 5838 1183 5894
rect 1239 5838 1307 5894
rect 1363 5838 1431 5894
rect 1487 5838 1555 5894
rect 1611 5838 1679 5894
rect 1735 5838 1803 5894
rect 1859 5838 1927 5894
rect 1983 5838 2051 5894
rect 2107 5838 2117 5894
rect 305 5770 2117 5838
rect 305 5714 315 5770
rect 371 5714 439 5770
rect 495 5714 563 5770
rect 619 5714 687 5770
rect 743 5714 811 5770
rect 867 5714 935 5770
rect 991 5714 1059 5770
rect 1115 5714 1183 5770
rect 1239 5714 1307 5770
rect 1363 5714 1431 5770
rect 1487 5714 1555 5770
rect 1611 5714 1679 5770
rect 1735 5714 1803 5770
rect 1859 5714 1927 5770
rect 1983 5714 2051 5770
rect 2107 5714 2117 5770
rect 305 5646 2117 5714
rect 305 5590 315 5646
rect 371 5590 439 5646
rect 495 5590 563 5646
rect 619 5590 687 5646
rect 743 5590 811 5646
rect 867 5590 935 5646
rect 991 5590 1059 5646
rect 1115 5590 1183 5646
rect 1239 5590 1307 5646
rect 1363 5590 1431 5646
rect 1487 5590 1555 5646
rect 1611 5590 1679 5646
rect 1735 5590 1803 5646
rect 1859 5590 1927 5646
rect 1983 5590 2051 5646
rect 2107 5590 2117 5646
rect 305 5522 2117 5590
rect 305 5466 315 5522
rect 371 5466 439 5522
rect 495 5466 563 5522
rect 619 5466 687 5522
rect 743 5466 811 5522
rect 867 5466 935 5522
rect 991 5466 1059 5522
rect 1115 5466 1183 5522
rect 1239 5466 1307 5522
rect 1363 5466 1431 5522
rect 1487 5466 1555 5522
rect 1611 5466 1679 5522
rect 1735 5466 1803 5522
rect 1859 5466 1927 5522
rect 1983 5466 2051 5522
rect 2107 5466 2117 5522
rect 305 5398 2117 5466
rect 305 5342 315 5398
rect 371 5342 439 5398
rect 495 5342 563 5398
rect 619 5342 687 5398
rect 743 5342 811 5398
rect 867 5342 935 5398
rect 991 5342 1059 5398
rect 1115 5342 1183 5398
rect 1239 5342 1307 5398
rect 1363 5342 1431 5398
rect 1487 5342 1555 5398
rect 1611 5342 1679 5398
rect 1735 5342 1803 5398
rect 1859 5342 1927 5398
rect 1983 5342 2051 5398
rect 2107 5342 2117 5398
rect 305 5274 2117 5342
rect 305 5218 315 5274
rect 371 5218 439 5274
rect 495 5218 563 5274
rect 619 5218 687 5274
rect 743 5218 811 5274
rect 867 5218 935 5274
rect 991 5218 1059 5274
rect 1115 5218 1183 5274
rect 1239 5218 1307 5274
rect 1363 5218 1431 5274
rect 1487 5218 1555 5274
rect 1611 5218 1679 5274
rect 1735 5218 1803 5274
rect 1859 5218 1927 5274
rect 1983 5218 2051 5274
rect 2107 5218 2117 5274
rect 305 5150 2117 5218
rect 305 5094 315 5150
rect 371 5094 439 5150
rect 495 5094 563 5150
rect 619 5094 687 5150
rect 743 5094 811 5150
rect 867 5094 935 5150
rect 991 5094 1059 5150
rect 1115 5094 1183 5150
rect 1239 5094 1307 5150
rect 1363 5094 1431 5150
rect 1487 5094 1555 5150
rect 1611 5094 1679 5150
rect 1735 5094 1803 5150
rect 1859 5094 1927 5150
rect 1983 5094 2051 5150
rect 2107 5094 2117 5150
rect 305 5026 2117 5094
rect 305 4970 315 5026
rect 371 4970 439 5026
rect 495 4970 563 5026
rect 619 4970 687 5026
rect 743 4970 811 5026
rect 867 4970 935 5026
rect 991 4970 1059 5026
rect 1115 4970 1183 5026
rect 1239 4970 1307 5026
rect 1363 4970 1431 5026
rect 1487 4970 1555 5026
rect 1611 4970 1679 5026
rect 1735 4970 1803 5026
rect 1859 4970 1927 5026
rect 1983 4970 2051 5026
rect 2107 4970 2117 5026
rect 305 4902 2117 4970
rect 305 4846 315 4902
rect 371 4846 439 4902
rect 495 4846 563 4902
rect 619 4846 687 4902
rect 743 4846 811 4902
rect 867 4846 935 4902
rect 991 4846 1059 4902
rect 1115 4846 1183 4902
rect 1239 4846 1307 4902
rect 1363 4846 1431 4902
rect 1487 4846 1555 4902
rect 1611 4846 1679 4902
rect 1735 4846 1803 4902
rect 1859 4846 1927 4902
rect 1983 4846 2051 4902
rect 2107 4846 2117 4902
rect 305 4836 2117 4846
rect 2798 7754 4734 7764
rect 2798 7698 2808 7754
rect 2864 7698 2932 7754
rect 2988 7698 3056 7754
rect 3112 7698 3180 7754
rect 3236 7698 3304 7754
rect 3360 7698 3428 7754
rect 3484 7698 3552 7754
rect 3608 7698 3676 7754
rect 3732 7698 3800 7754
rect 3856 7698 3924 7754
rect 3980 7698 4048 7754
rect 4104 7698 4172 7754
rect 4228 7698 4296 7754
rect 4352 7698 4420 7754
rect 4476 7698 4544 7754
rect 4600 7698 4668 7754
rect 4724 7698 4734 7754
rect 2798 7630 4734 7698
rect 2798 7574 2808 7630
rect 2864 7574 2932 7630
rect 2988 7574 3056 7630
rect 3112 7574 3180 7630
rect 3236 7574 3304 7630
rect 3360 7574 3428 7630
rect 3484 7574 3552 7630
rect 3608 7574 3676 7630
rect 3732 7574 3800 7630
rect 3856 7574 3924 7630
rect 3980 7574 4048 7630
rect 4104 7574 4172 7630
rect 4228 7574 4296 7630
rect 4352 7574 4420 7630
rect 4476 7574 4544 7630
rect 4600 7574 4668 7630
rect 4724 7574 4734 7630
rect 2798 7506 4734 7574
rect 2798 7450 2808 7506
rect 2864 7450 2932 7506
rect 2988 7450 3056 7506
rect 3112 7450 3180 7506
rect 3236 7450 3304 7506
rect 3360 7450 3428 7506
rect 3484 7450 3552 7506
rect 3608 7450 3676 7506
rect 3732 7450 3800 7506
rect 3856 7450 3924 7506
rect 3980 7450 4048 7506
rect 4104 7450 4172 7506
rect 4228 7450 4296 7506
rect 4352 7450 4420 7506
rect 4476 7450 4544 7506
rect 4600 7450 4668 7506
rect 4724 7450 4734 7506
rect 2798 7382 4734 7450
rect 2798 7326 2808 7382
rect 2864 7326 2932 7382
rect 2988 7326 3056 7382
rect 3112 7326 3180 7382
rect 3236 7326 3304 7382
rect 3360 7326 3428 7382
rect 3484 7326 3552 7382
rect 3608 7326 3676 7382
rect 3732 7326 3800 7382
rect 3856 7326 3924 7382
rect 3980 7326 4048 7382
rect 4104 7326 4172 7382
rect 4228 7326 4296 7382
rect 4352 7326 4420 7382
rect 4476 7326 4544 7382
rect 4600 7326 4668 7382
rect 4724 7326 4734 7382
rect 2798 7258 4734 7326
rect 2798 7202 2808 7258
rect 2864 7202 2932 7258
rect 2988 7202 3056 7258
rect 3112 7202 3180 7258
rect 3236 7202 3304 7258
rect 3360 7202 3428 7258
rect 3484 7202 3552 7258
rect 3608 7202 3676 7258
rect 3732 7202 3800 7258
rect 3856 7202 3924 7258
rect 3980 7202 4048 7258
rect 4104 7202 4172 7258
rect 4228 7202 4296 7258
rect 4352 7202 4420 7258
rect 4476 7202 4544 7258
rect 4600 7202 4668 7258
rect 4724 7202 4734 7258
rect 2798 7134 4734 7202
rect 2798 7078 2808 7134
rect 2864 7078 2932 7134
rect 2988 7078 3056 7134
rect 3112 7078 3180 7134
rect 3236 7078 3304 7134
rect 3360 7078 3428 7134
rect 3484 7078 3552 7134
rect 3608 7078 3676 7134
rect 3732 7078 3800 7134
rect 3856 7078 3924 7134
rect 3980 7078 4048 7134
rect 4104 7078 4172 7134
rect 4228 7078 4296 7134
rect 4352 7078 4420 7134
rect 4476 7078 4544 7134
rect 4600 7078 4668 7134
rect 4724 7078 4734 7134
rect 2798 7010 4734 7078
rect 2798 6954 2808 7010
rect 2864 6954 2932 7010
rect 2988 6954 3056 7010
rect 3112 6954 3180 7010
rect 3236 6954 3304 7010
rect 3360 6954 3428 7010
rect 3484 6954 3552 7010
rect 3608 6954 3676 7010
rect 3732 6954 3800 7010
rect 3856 6954 3924 7010
rect 3980 6954 4048 7010
rect 4104 6954 4172 7010
rect 4228 6954 4296 7010
rect 4352 6954 4420 7010
rect 4476 6954 4544 7010
rect 4600 6954 4668 7010
rect 4724 6954 4734 7010
rect 2798 6886 4734 6954
rect 2798 6830 2808 6886
rect 2864 6830 2932 6886
rect 2988 6830 3056 6886
rect 3112 6830 3180 6886
rect 3236 6830 3304 6886
rect 3360 6830 3428 6886
rect 3484 6830 3552 6886
rect 3608 6830 3676 6886
rect 3732 6830 3800 6886
rect 3856 6830 3924 6886
rect 3980 6830 4048 6886
rect 4104 6830 4172 6886
rect 4228 6830 4296 6886
rect 4352 6830 4420 6886
rect 4476 6830 4544 6886
rect 4600 6830 4668 6886
rect 4724 6830 4734 6886
rect 2798 6762 4734 6830
rect 2798 6706 2808 6762
rect 2864 6706 2932 6762
rect 2988 6706 3056 6762
rect 3112 6706 3180 6762
rect 3236 6706 3304 6762
rect 3360 6706 3428 6762
rect 3484 6706 3552 6762
rect 3608 6706 3676 6762
rect 3732 6706 3800 6762
rect 3856 6706 3924 6762
rect 3980 6706 4048 6762
rect 4104 6706 4172 6762
rect 4228 6706 4296 6762
rect 4352 6706 4420 6762
rect 4476 6706 4544 6762
rect 4600 6706 4668 6762
rect 4724 6706 4734 6762
rect 2798 6638 4734 6706
rect 2798 6582 2808 6638
rect 2864 6582 2932 6638
rect 2988 6582 3056 6638
rect 3112 6582 3180 6638
rect 3236 6582 3304 6638
rect 3360 6582 3428 6638
rect 3484 6582 3552 6638
rect 3608 6582 3676 6638
rect 3732 6582 3800 6638
rect 3856 6582 3924 6638
rect 3980 6582 4048 6638
rect 4104 6582 4172 6638
rect 4228 6582 4296 6638
rect 4352 6582 4420 6638
rect 4476 6582 4544 6638
rect 4600 6582 4668 6638
rect 4724 6582 4734 6638
rect 2798 6514 4734 6582
rect 2798 6458 2808 6514
rect 2864 6458 2932 6514
rect 2988 6458 3056 6514
rect 3112 6458 3180 6514
rect 3236 6458 3304 6514
rect 3360 6458 3428 6514
rect 3484 6458 3552 6514
rect 3608 6458 3676 6514
rect 3732 6458 3800 6514
rect 3856 6458 3924 6514
rect 3980 6458 4048 6514
rect 4104 6458 4172 6514
rect 4228 6458 4296 6514
rect 4352 6458 4420 6514
rect 4476 6458 4544 6514
rect 4600 6458 4668 6514
rect 4724 6458 4734 6514
rect 2798 6390 4734 6458
rect 2798 6334 2808 6390
rect 2864 6334 2932 6390
rect 2988 6334 3056 6390
rect 3112 6334 3180 6390
rect 3236 6334 3304 6390
rect 3360 6334 3428 6390
rect 3484 6334 3552 6390
rect 3608 6334 3676 6390
rect 3732 6334 3800 6390
rect 3856 6334 3924 6390
rect 3980 6334 4048 6390
rect 4104 6334 4172 6390
rect 4228 6334 4296 6390
rect 4352 6334 4420 6390
rect 4476 6334 4544 6390
rect 4600 6334 4668 6390
rect 4724 6334 4734 6390
rect 2798 6266 4734 6334
rect 2798 6210 2808 6266
rect 2864 6210 2932 6266
rect 2988 6210 3056 6266
rect 3112 6210 3180 6266
rect 3236 6210 3304 6266
rect 3360 6210 3428 6266
rect 3484 6210 3552 6266
rect 3608 6210 3676 6266
rect 3732 6210 3800 6266
rect 3856 6210 3924 6266
rect 3980 6210 4048 6266
rect 4104 6210 4172 6266
rect 4228 6210 4296 6266
rect 4352 6210 4420 6266
rect 4476 6210 4544 6266
rect 4600 6210 4668 6266
rect 4724 6210 4734 6266
rect 2798 6142 4734 6210
rect 2798 6086 2808 6142
rect 2864 6086 2932 6142
rect 2988 6086 3056 6142
rect 3112 6086 3180 6142
rect 3236 6086 3304 6142
rect 3360 6086 3428 6142
rect 3484 6086 3552 6142
rect 3608 6086 3676 6142
rect 3732 6086 3800 6142
rect 3856 6086 3924 6142
rect 3980 6086 4048 6142
rect 4104 6086 4172 6142
rect 4228 6086 4296 6142
rect 4352 6086 4420 6142
rect 4476 6086 4544 6142
rect 4600 6086 4668 6142
rect 4724 6086 4734 6142
rect 2798 6018 4734 6086
rect 2798 5962 2808 6018
rect 2864 5962 2932 6018
rect 2988 5962 3056 6018
rect 3112 5962 3180 6018
rect 3236 5962 3304 6018
rect 3360 5962 3428 6018
rect 3484 5962 3552 6018
rect 3608 5962 3676 6018
rect 3732 5962 3800 6018
rect 3856 5962 3924 6018
rect 3980 5962 4048 6018
rect 4104 5962 4172 6018
rect 4228 5962 4296 6018
rect 4352 5962 4420 6018
rect 4476 5962 4544 6018
rect 4600 5962 4668 6018
rect 4724 5962 4734 6018
rect 2798 5894 4734 5962
rect 2798 5838 2808 5894
rect 2864 5838 2932 5894
rect 2988 5838 3056 5894
rect 3112 5838 3180 5894
rect 3236 5838 3304 5894
rect 3360 5838 3428 5894
rect 3484 5838 3552 5894
rect 3608 5838 3676 5894
rect 3732 5838 3800 5894
rect 3856 5838 3924 5894
rect 3980 5838 4048 5894
rect 4104 5838 4172 5894
rect 4228 5838 4296 5894
rect 4352 5838 4420 5894
rect 4476 5838 4544 5894
rect 4600 5838 4668 5894
rect 4724 5838 4734 5894
rect 2798 5770 4734 5838
rect 2798 5714 2808 5770
rect 2864 5714 2932 5770
rect 2988 5714 3056 5770
rect 3112 5714 3180 5770
rect 3236 5714 3304 5770
rect 3360 5714 3428 5770
rect 3484 5714 3552 5770
rect 3608 5714 3676 5770
rect 3732 5714 3800 5770
rect 3856 5714 3924 5770
rect 3980 5714 4048 5770
rect 4104 5714 4172 5770
rect 4228 5714 4296 5770
rect 4352 5714 4420 5770
rect 4476 5714 4544 5770
rect 4600 5714 4668 5770
rect 4724 5714 4734 5770
rect 2798 5646 4734 5714
rect 2798 5590 2808 5646
rect 2864 5590 2932 5646
rect 2988 5590 3056 5646
rect 3112 5590 3180 5646
rect 3236 5590 3304 5646
rect 3360 5590 3428 5646
rect 3484 5590 3552 5646
rect 3608 5590 3676 5646
rect 3732 5590 3800 5646
rect 3856 5590 3924 5646
rect 3980 5590 4048 5646
rect 4104 5590 4172 5646
rect 4228 5590 4296 5646
rect 4352 5590 4420 5646
rect 4476 5590 4544 5646
rect 4600 5590 4668 5646
rect 4724 5590 4734 5646
rect 2798 5522 4734 5590
rect 2798 5466 2808 5522
rect 2864 5466 2932 5522
rect 2988 5466 3056 5522
rect 3112 5466 3180 5522
rect 3236 5466 3304 5522
rect 3360 5466 3428 5522
rect 3484 5466 3552 5522
rect 3608 5466 3676 5522
rect 3732 5466 3800 5522
rect 3856 5466 3924 5522
rect 3980 5466 4048 5522
rect 4104 5466 4172 5522
rect 4228 5466 4296 5522
rect 4352 5466 4420 5522
rect 4476 5466 4544 5522
rect 4600 5466 4668 5522
rect 4724 5466 4734 5522
rect 2798 5398 4734 5466
rect 2798 5342 2808 5398
rect 2864 5342 2932 5398
rect 2988 5342 3056 5398
rect 3112 5342 3180 5398
rect 3236 5342 3304 5398
rect 3360 5342 3428 5398
rect 3484 5342 3552 5398
rect 3608 5342 3676 5398
rect 3732 5342 3800 5398
rect 3856 5342 3924 5398
rect 3980 5342 4048 5398
rect 4104 5342 4172 5398
rect 4228 5342 4296 5398
rect 4352 5342 4420 5398
rect 4476 5342 4544 5398
rect 4600 5342 4668 5398
rect 4724 5342 4734 5398
rect 2798 5274 4734 5342
rect 2798 5218 2808 5274
rect 2864 5218 2932 5274
rect 2988 5218 3056 5274
rect 3112 5218 3180 5274
rect 3236 5218 3304 5274
rect 3360 5218 3428 5274
rect 3484 5218 3552 5274
rect 3608 5218 3676 5274
rect 3732 5218 3800 5274
rect 3856 5218 3924 5274
rect 3980 5218 4048 5274
rect 4104 5218 4172 5274
rect 4228 5218 4296 5274
rect 4352 5218 4420 5274
rect 4476 5218 4544 5274
rect 4600 5218 4668 5274
rect 4724 5218 4734 5274
rect 2798 5150 4734 5218
rect 2798 5094 2808 5150
rect 2864 5094 2932 5150
rect 2988 5094 3056 5150
rect 3112 5094 3180 5150
rect 3236 5094 3304 5150
rect 3360 5094 3428 5150
rect 3484 5094 3552 5150
rect 3608 5094 3676 5150
rect 3732 5094 3800 5150
rect 3856 5094 3924 5150
rect 3980 5094 4048 5150
rect 4104 5094 4172 5150
rect 4228 5094 4296 5150
rect 4352 5094 4420 5150
rect 4476 5094 4544 5150
rect 4600 5094 4668 5150
rect 4724 5094 4734 5150
rect 2798 5026 4734 5094
rect 2798 4970 2808 5026
rect 2864 4970 2932 5026
rect 2988 4970 3056 5026
rect 3112 4970 3180 5026
rect 3236 4970 3304 5026
rect 3360 4970 3428 5026
rect 3484 4970 3552 5026
rect 3608 4970 3676 5026
rect 3732 4970 3800 5026
rect 3856 4970 3924 5026
rect 3980 4970 4048 5026
rect 4104 4970 4172 5026
rect 4228 4970 4296 5026
rect 4352 4970 4420 5026
rect 4476 4970 4544 5026
rect 4600 4970 4668 5026
rect 4724 4970 4734 5026
rect 2798 4902 4734 4970
rect 2798 4846 2808 4902
rect 2864 4846 2932 4902
rect 2988 4846 3056 4902
rect 3112 4846 3180 4902
rect 3236 4846 3304 4902
rect 3360 4846 3428 4902
rect 3484 4846 3552 4902
rect 3608 4846 3676 4902
rect 3732 4846 3800 4902
rect 3856 4846 3924 4902
rect 3980 4846 4048 4902
rect 4104 4846 4172 4902
rect 4228 4846 4296 4902
rect 4352 4846 4420 4902
rect 4476 4846 4544 4902
rect 4600 4846 4668 4902
rect 4724 4846 4734 4902
rect 2798 4836 4734 4846
rect 5168 7754 7104 7764
rect 5168 7698 5178 7754
rect 5234 7698 5302 7754
rect 5358 7698 5426 7754
rect 5482 7698 5550 7754
rect 5606 7698 5674 7754
rect 5730 7698 5798 7754
rect 5854 7698 5922 7754
rect 5978 7698 6046 7754
rect 6102 7698 6170 7754
rect 6226 7698 6294 7754
rect 6350 7698 6418 7754
rect 6474 7698 6542 7754
rect 6598 7698 6666 7754
rect 6722 7698 6790 7754
rect 6846 7698 6914 7754
rect 6970 7698 7038 7754
rect 7094 7698 7104 7754
rect 5168 7630 7104 7698
rect 5168 7574 5178 7630
rect 5234 7574 5302 7630
rect 5358 7574 5426 7630
rect 5482 7574 5550 7630
rect 5606 7574 5674 7630
rect 5730 7574 5798 7630
rect 5854 7574 5922 7630
rect 5978 7574 6046 7630
rect 6102 7574 6170 7630
rect 6226 7574 6294 7630
rect 6350 7574 6418 7630
rect 6474 7574 6542 7630
rect 6598 7574 6666 7630
rect 6722 7574 6790 7630
rect 6846 7574 6914 7630
rect 6970 7574 7038 7630
rect 7094 7574 7104 7630
rect 5168 7506 7104 7574
rect 5168 7450 5178 7506
rect 5234 7450 5302 7506
rect 5358 7450 5426 7506
rect 5482 7450 5550 7506
rect 5606 7450 5674 7506
rect 5730 7450 5798 7506
rect 5854 7450 5922 7506
rect 5978 7450 6046 7506
rect 6102 7450 6170 7506
rect 6226 7450 6294 7506
rect 6350 7450 6418 7506
rect 6474 7450 6542 7506
rect 6598 7450 6666 7506
rect 6722 7450 6790 7506
rect 6846 7450 6914 7506
rect 6970 7450 7038 7506
rect 7094 7450 7104 7506
rect 5168 7382 7104 7450
rect 5168 7326 5178 7382
rect 5234 7326 5302 7382
rect 5358 7326 5426 7382
rect 5482 7326 5550 7382
rect 5606 7326 5674 7382
rect 5730 7326 5798 7382
rect 5854 7326 5922 7382
rect 5978 7326 6046 7382
rect 6102 7326 6170 7382
rect 6226 7326 6294 7382
rect 6350 7326 6418 7382
rect 6474 7326 6542 7382
rect 6598 7326 6666 7382
rect 6722 7326 6790 7382
rect 6846 7326 6914 7382
rect 6970 7326 7038 7382
rect 7094 7326 7104 7382
rect 5168 7258 7104 7326
rect 5168 7202 5178 7258
rect 5234 7202 5302 7258
rect 5358 7202 5426 7258
rect 5482 7202 5550 7258
rect 5606 7202 5674 7258
rect 5730 7202 5798 7258
rect 5854 7202 5922 7258
rect 5978 7202 6046 7258
rect 6102 7202 6170 7258
rect 6226 7202 6294 7258
rect 6350 7202 6418 7258
rect 6474 7202 6542 7258
rect 6598 7202 6666 7258
rect 6722 7202 6790 7258
rect 6846 7202 6914 7258
rect 6970 7202 7038 7258
rect 7094 7202 7104 7258
rect 5168 7134 7104 7202
rect 5168 7078 5178 7134
rect 5234 7078 5302 7134
rect 5358 7078 5426 7134
rect 5482 7078 5550 7134
rect 5606 7078 5674 7134
rect 5730 7078 5798 7134
rect 5854 7078 5922 7134
rect 5978 7078 6046 7134
rect 6102 7078 6170 7134
rect 6226 7078 6294 7134
rect 6350 7078 6418 7134
rect 6474 7078 6542 7134
rect 6598 7078 6666 7134
rect 6722 7078 6790 7134
rect 6846 7078 6914 7134
rect 6970 7078 7038 7134
rect 7094 7078 7104 7134
rect 5168 7010 7104 7078
rect 5168 6954 5178 7010
rect 5234 6954 5302 7010
rect 5358 6954 5426 7010
rect 5482 6954 5550 7010
rect 5606 6954 5674 7010
rect 5730 6954 5798 7010
rect 5854 6954 5922 7010
rect 5978 6954 6046 7010
rect 6102 6954 6170 7010
rect 6226 6954 6294 7010
rect 6350 6954 6418 7010
rect 6474 6954 6542 7010
rect 6598 6954 6666 7010
rect 6722 6954 6790 7010
rect 6846 6954 6914 7010
rect 6970 6954 7038 7010
rect 7094 6954 7104 7010
rect 5168 6886 7104 6954
rect 5168 6830 5178 6886
rect 5234 6830 5302 6886
rect 5358 6830 5426 6886
rect 5482 6830 5550 6886
rect 5606 6830 5674 6886
rect 5730 6830 5798 6886
rect 5854 6830 5922 6886
rect 5978 6830 6046 6886
rect 6102 6830 6170 6886
rect 6226 6830 6294 6886
rect 6350 6830 6418 6886
rect 6474 6830 6542 6886
rect 6598 6830 6666 6886
rect 6722 6830 6790 6886
rect 6846 6830 6914 6886
rect 6970 6830 7038 6886
rect 7094 6830 7104 6886
rect 5168 6762 7104 6830
rect 5168 6706 5178 6762
rect 5234 6706 5302 6762
rect 5358 6706 5426 6762
rect 5482 6706 5550 6762
rect 5606 6706 5674 6762
rect 5730 6706 5798 6762
rect 5854 6706 5922 6762
rect 5978 6706 6046 6762
rect 6102 6706 6170 6762
rect 6226 6706 6294 6762
rect 6350 6706 6418 6762
rect 6474 6706 6542 6762
rect 6598 6706 6666 6762
rect 6722 6706 6790 6762
rect 6846 6706 6914 6762
rect 6970 6706 7038 6762
rect 7094 6706 7104 6762
rect 5168 6638 7104 6706
rect 5168 6582 5178 6638
rect 5234 6582 5302 6638
rect 5358 6582 5426 6638
rect 5482 6582 5550 6638
rect 5606 6582 5674 6638
rect 5730 6582 5798 6638
rect 5854 6582 5922 6638
rect 5978 6582 6046 6638
rect 6102 6582 6170 6638
rect 6226 6582 6294 6638
rect 6350 6582 6418 6638
rect 6474 6582 6542 6638
rect 6598 6582 6666 6638
rect 6722 6582 6790 6638
rect 6846 6582 6914 6638
rect 6970 6582 7038 6638
rect 7094 6582 7104 6638
rect 5168 6514 7104 6582
rect 5168 6458 5178 6514
rect 5234 6458 5302 6514
rect 5358 6458 5426 6514
rect 5482 6458 5550 6514
rect 5606 6458 5674 6514
rect 5730 6458 5798 6514
rect 5854 6458 5922 6514
rect 5978 6458 6046 6514
rect 6102 6458 6170 6514
rect 6226 6458 6294 6514
rect 6350 6458 6418 6514
rect 6474 6458 6542 6514
rect 6598 6458 6666 6514
rect 6722 6458 6790 6514
rect 6846 6458 6914 6514
rect 6970 6458 7038 6514
rect 7094 6458 7104 6514
rect 5168 6390 7104 6458
rect 5168 6334 5178 6390
rect 5234 6334 5302 6390
rect 5358 6334 5426 6390
rect 5482 6334 5550 6390
rect 5606 6334 5674 6390
rect 5730 6334 5798 6390
rect 5854 6334 5922 6390
rect 5978 6334 6046 6390
rect 6102 6334 6170 6390
rect 6226 6334 6294 6390
rect 6350 6334 6418 6390
rect 6474 6334 6542 6390
rect 6598 6334 6666 6390
rect 6722 6334 6790 6390
rect 6846 6334 6914 6390
rect 6970 6334 7038 6390
rect 7094 6334 7104 6390
rect 5168 6266 7104 6334
rect 5168 6210 5178 6266
rect 5234 6210 5302 6266
rect 5358 6210 5426 6266
rect 5482 6210 5550 6266
rect 5606 6210 5674 6266
rect 5730 6210 5798 6266
rect 5854 6210 5922 6266
rect 5978 6210 6046 6266
rect 6102 6210 6170 6266
rect 6226 6210 6294 6266
rect 6350 6210 6418 6266
rect 6474 6210 6542 6266
rect 6598 6210 6666 6266
rect 6722 6210 6790 6266
rect 6846 6210 6914 6266
rect 6970 6210 7038 6266
rect 7094 6210 7104 6266
rect 5168 6142 7104 6210
rect 5168 6086 5178 6142
rect 5234 6086 5302 6142
rect 5358 6086 5426 6142
rect 5482 6086 5550 6142
rect 5606 6086 5674 6142
rect 5730 6086 5798 6142
rect 5854 6086 5922 6142
rect 5978 6086 6046 6142
rect 6102 6086 6170 6142
rect 6226 6086 6294 6142
rect 6350 6086 6418 6142
rect 6474 6086 6542 6142
rect 6598 6086 6666 6142
rect 6722 6086 6790 6142
rect 6846 6086 6914 6142
rect 6970 6086 7038 6142
rect 7094 6086 7104 6142
rect 5168 6018 7104 6086
rect 5168 5962 5178 6018
rect 5234 5962 5302 6018
rect 5358 5962 5426 6018
rect 5482 5962 5550 6018
rect 5606 5962 5674 6018
rect 5730 5962 5798 6018
rect 5854 5962 5922 6018
rect 5978 5962 6046 6018
rect 6102 5962 6170 6018
rect 6226 5962 6294 6018
rect 6350 5962 6418 6018
rect 6474 5962 6542 6018
rect 6598 5962 6666 6018
rect 6722 5962 6790 6018
rect 6846 5962 6914 6018
rect 6970 5962 7038 6018
rect 7094 5962 7104 6018
rect 5168 5894 7104 5962
rect 5168 5838 5178 5894
rect 5234 5838 5302 5894
rect 5358 5838 5426 5894
rect 5482 5838 5550 5894
rect 5606 5838 5674 5894
rect 5730 5838 5798 5894
rect 5854 5838 5922 5894
rect 5978 5838 6046 5894
rect 6102 5838 6170 5894
rect 6226 5838 6294 5894
rect 6350 5838 6418 5894
rect 6474 5838 6542 5894
rect 6598 5838 6666 5894
rect 6722 5838 6790 5894
rect 6846 5838 6914 5894
rect 6970 5838 7038 5894
rect 7094 5838 7104 5894
rect 5168 5770 7104 5838
rect 5168 5714 5178 5770
rect 5234 5714 5302 5770
rect 5358 5714 5426 5770
rect 5482 5714 5550 5770
rect 5606 5714 5674 5770
rect 5730 5714 5798 5770
rect 5854 5714 5922 5770
rect 5978 5714 6046 5770
rect 6102 5714 6170 5770
rect 6226 5714 6294 5770
rect 6350 5714 6418 5770
rect 6474 5714 6542 5770
rect 6598 5714 6666 5770
rect 6722 5714 6790 5770
rect 6846 5714 6914 5770
rect 6970 5714 7038 5770
rect 7094 5714 7104 5770
rect 5168 5646 7104 5714
rect 5168 5590 5178 5646
rect 5234 5590 5302 5646
rect 5358 5590 5426 5646
rect 5482 5590 5550 5646
rect 5606 5590 5674 5646
rect 5730 5590 5798 5646
rect 5854 5590 5922 5646
rect 5978 5590 6046 5646
rect 6102 5590 6170 5646
rect 6226 5590 6294 5646
rect 6350 5590 6418 5646
rect 6474 5590 6542 5646
rect 6598 5590 6666 5646
rect 6722 5590 6790 5646
rect 6846 5590 6914 5646
rect 6970 5590 7038 5646
rect 7094 5590 7104 5646
rect 5168 5522 7104 5590
rect 5168 5466 5178 5522
rect 5234 5466 5302 5522
rect 5358 5466 5426 5522
rect 5482 5466 5550 5522
rect 5606 5466 5674 5522
rect 5730 5466 5798 5522
rect 5854 5466 5922 5522
rect 5978 5466 6046 5522
rect 6102 5466 6170 5522
rect 6226 5466 6294 5522
rect 6350 5466 6418 5522
rect 6474 5466 6542 5522
rect 6598 5466 6666 5522
rect 6722 5466 6790 5522
rect 6846 5466 6914 5522
rect 6970 5466 7038 5522
rect 7094 5466 7104 5522
rect 5168 5398 7104 5466
rect 5168 5342 5178 5398
rect 5234 5342 5302 5398
rect 5358 5342 5426 5398
rect 5482 5342 5550 5398
rect 5606 5342 5674 5398
rect 5730 5342 5798 5398
rect 5854 5342 5922 5398
rect 5978 5342 6046 5398
rect 6102 5342 6170 5398
rect 6226 5342 6294 5398
rect 6350 5342 6418 5398
rect 6474 5342 6542 5398
rect 6598 5342 6666 5398
rect 6722 5342 6790 5398
rect 6846 5342 6914 5398
rect 6970 5342 7038 5398
rect 7094 5342 7104 5398
rect 5168 5274 7104 5342
rect 5168 5218 5178 5274
rect 5234 5218 5302 5274
rect 5358 5218 5426 5274
rect 5482 5218 5550 5274
rect 5606 5218 5674 5274
rect 5730 5218 5798 5274
rect 5854 5218 5922 5274
rect 5978 5218 6046 5274
rect 6102 5218 6170 5274
rect 6226 5218 6294 5274
rect 6350 5218 6418 5274
rect 6474 5218 6542 5274
rect 6598 5218 6666 5274
rect 6722 5218 6790 5274
rect 6846 5218 6914 5274
rect 6970 5218 7038 5274
rect 7094 5218 7104 5274
rect 5168 5150 7104 5218
rect 5168 5094 5178 5150
rect 5234 5094 5302 5150
rect 5358 5094 5426 5150
rect 5482 5094 5550 5150
rect 5606 5094 5674 5150
rect 5730 5094 5798 5150
rect 5854 5094 5922 5150
rect 5978 5094 6046 5150
rect 6102 5094 6170 5150
rect 6226 5094 6294 5150
rect 6350 5094 6418 5150
rect 6474 5094 6542 5150
rect 6598 5094 6666 5150
rect 6722 5094 6790 5150
rect 6846 5094 6914 5150
rect 6970 5094 7038 5150
rect 7094 5094 7104 5150
rect 5168 5026 7104 5094
rect 5168 4970 5178 5026
rect 5234 4970 5302 5026
rect 5358 4970 5426 5026
rect 5482 4970 5550 5026
rect 5606 4970 5674 5026
rect 5730 4970 5798 5026
rect 5854 4970 5922 5026
rect 5978 4970 6046 5026
rect 6102 4970 6170 5026
rect 6226 4970 6294 5026
rect 6350 4970 6418 5026
rect 6474 4970 6542 5026
rect 6598 4970 6666 5026
rect 6722 4970 6790 5026
rect 6846 4970 6914 5026
rect 6970 4970 7038 5026
rect 7094 4970 7104 5026
rect 5168 4902 7104 4970
rect 5168 4846 5178 4902
rect 5234 4846 5302 4902
rect 5358 4846 5426 4902
rect 5482 4846 5550 4902
rect 5606 4846 5674 4902
rect 5730 4846 5798 4902
rect 5854 4846 5922 4902
rect 5978 4846 6046 4902
rect 6102 4846 6170 4902
rect 6226 4846 6294 4902
rect 6350 4846 6418 4902
rect 6474 4846 6542 4902
rect 6598 4846 6666 4902
rect 6722 4846 6790 4902
rect 6846 4846 6914 4902
rect 6970 4846 7038 4902
rect 7094 4846 7104 4902
rect 5168 4836 7104 4846
rect 7874 7754 9810 7764
rect 7874 7698 7884 7754
rect 7940 7698 8008 7754
rect 8064 7698 8132 7754
rect 8188 7698 8256 7754
rect 8312 7698 8380 7754
rect 8436 7698 8504 7754
rect 8560 7698 8628 7754
rect 8684 7698 8752 7754
rect 8808 7698 8876 7754
rect 8932 7698 9000 7754
rect 9056 7698 9124 7754
rect 9180 7698 9248 7754
rect 9304 7698 9372 7754
rect 9428 7698 9496 7754
rect 9552 7698 9620 7754
rect 9676 7698 9744 7754
rect 9800 7698 9810 7754
rect 7874 7630 9810 7698
rect 7874 7574 7884 7630
rect 7940 7574 8008 7630
rect 8064 7574 8132 7630
rect 8188 7574 8256 7630
rect 8312 7574 8380 7630
rect 8436 7574 8504 7630
rect 8560 7574 8628 7630
rect 8684 7574 8752 7630
rect 8808 7574 8876 7630
rect 8932 7574 9000 7630
rect 9056 7574 9124 7630
rect 9180 7574 9248 7630
rect 9304 7574 9372 7630
rect 9428 7574 9496 7630
rect 9552 7574 9620 7630
rect 9676 7574 9744 7630
rect 9800 7574 9810 7630
rect 7874 7506 9810 7574
rect 7874 7450 7884 7506
rect 7940 7450 8008 7506
rect 8064 7450 8132 7506
rect 8188 7450 8256 7506
rect 8312 7450 8380 7506
rect 8436 7450 8504 7506
rect 8560 7450 8628 7506
rect 8684 7450 8752 7506
rect 8808 7450 8876 7506
rect 8932 7450 9000 7506
rect 9056 7450 9124 7506
rect 9180 7450 9248 7506
rect 9304 7450 9372 7506
rect 9428 7450 9496 7506
rect 9552 7450 9620 7506
rect 9676 7450 9744 7506
rect 9800 7450 9810 7506
rect 7874 7382 9810 7450
rect 7874 7326 7884 7382
rect 7940 7326 8008 7382
rect 8064 7326 8132 7382
rect 8188 7326 8256 7382
rect 8312 7326 8380 7382
rect 8436 7326 8504 7382
rect 8560 7326 8628 7382
rect 8684 7326 8752 7382
rect 8808 7326 8876 7382
rect 8932 7326 9000 7382
rect 9056 7326 9124 7382
rect 9180 7326 9248 7382
rect 9304 7326 9372 7382
rect 9428 7326 9496 7382
rect 9552 7326 9620 7382
rect 9676 7326 9744 7382
rect 9800 7326 9810 7382
rect 7874 7258 9810 7326
rect 7874 7202 7884 7258
rect 7940 7202 8008 7258
rect 8064 7202 8132 7258
rect 8188 7202 8256 7258
rect 8312 7202 8380 7258
rect 8436 7202 8504 7258
rect 8560 7202 8628 7258
rect 8684 7202 8752 7258
rect 8808 7202 8876 7258
rect 8932 7202 9000 7258
rect 9056 7202 9124 7258
rect 9180 7202 9248 7258
rect 9304 7202 9372 7258
rect 9428 7202 9496 7258
rect 9552 7202 9620 7258
rect 9676 7202 9744 7258
rect 9800 7202 9810 7258
rect 7874 7134 9810 7202
rect 7874 7078 7884 7134
rect 7940 7078 8008 7134
rect 8064 7078 8132 7134
rect 8188 7078 8256 7134
rect 8312 7078 8380 7134
rect 8436 7078 8504 7134
rect 8560 7078 8628 7134
rect 8684 7078 8752 7134
rect 8808 7078 8876 7134
rect 8932 7078 9000 7134
rect 9056 7078 9124 7134
rect 9180 7078 9248 7134
rect 9304 7078 9372 7134
rect 9428 7078 9496 7134
rect 9552 7078 9620 7134
rect 9676 7078 9744 7134
rect 9800 7078 9810 7134
rect 7874 7010 9810 7078
rect 7874 6954 7884 7010
rect 7940 6954 8008 7010
rect 8064 6954 8132 7010
rect 8188 6954 8256 7010
rect 8312 6954 8380 7010
rect 8436 6954 8504 7010
rect 8560 6954 8628 7010
rect 8684 6954 8752 7010
rect 8808 6954 8876 7010
rect 8932 6954 9000 7010
rect 9056 6954 9124 7010
rect 9180 6954 9248 7010
rect 9304 6954 9372 7010
rect 9428 6954 9496 7010
rect 9552 6954 9620 7010
rect 9676 6954 9744 7010
rect 9800 6954 9810 7010
rect 7874 6886 9810 6954
rect 7874 6830 7884 6886
rect 7940 6830 8008 6886
rect 8064 6830 8132 6886
rect 8188 6830 8256 6886
rect 8312 6830 8380 6886
rect 8436 6830 8504 6886
rect 8560 6830 8628 6886
rect 8684 6830 8752 6886
rect 8808 6830 8876 6886
rect 8932 6830 9000 6886
rect 9056 6830 9124 6886
rect 9180 6830 9248 6886
rect 9304 6830 9372 6886
rect 9428 6830 9496 6886
rect 9552 6830 9620 6886
rect 9676 6830 9744 6886
rect 9800 6830 9810 6886
rect 7874 6762 9810 6830
rect 7874 6706 7884 6762
rect 7940 6706 8008 6762
rect 8064 6706 8132 6762
rect 8188 6706 8256 6762
rect 8312 6706 8380 6762
rect 8436 6706 8504 6762
rect 8560 6706 8628 6762
rect 8684 6706 8752 6762
rect 8808 6706 8876 6762
rect 8932 6706 9000 6762
rect 9056 6706 9124 6762
rect 9180 6706 9248 6762
rect 9304 6706 9372 6762
rect 9428 6706 9496 6762
rect 9552 6706 9620 6762
rect 9676 6706 9744 6762
rect 9800 6706 9810 6762
rect 7874 6638 9810 6706
rect 7874 6582 7884 6638
rect 7940 6582 8008 6638
rect 8064 6582 8132 6638
rect 8188 6582 8256 6638
rect 8312 6582 8380 6638
rect 8436 6582 8504 6638
rect 8560 6582 8628 6638
rect 8684 6582 8752 6638
rect 8808 6582 8876 6638
rect 8932 6582 9000 6638
rect 9056 6582 9124 6638
rect 9180 6582 9248 6638
rect 9304 6582 9372 6638
rect 9428 6582 9496 6638
rect 9552 6582 9620 6638
rect 9676 6582 9744 6638
rect 9800 6582 9810 6638
rect 7874 6514 9810 6582
rect 7874 6458 7884 6514
rect 7940 6458 8008 6514
rect 8064 6458 8132 6514
rect 8188 6458 8256 6514
rect 8312 6458 8380 6514
rect 8436 6458 8504 6514
rect 8560 6458 8628 6514
rect 8684 6458 8752 6514
rect 8808 6458 8876 6514
rect 8932 6458 9000 6514
rect 9056 6458 9124 6514
rect 9180 6458 9248 6514
rect 9304 6458 9372 6514
rect 9428 6458 9496 6514
rect 9552 6458 9620 6514
rect 9676 6458 9744 6514
rect 9800 6458 9810 6514
rect 7874 6390 9810 6458
rect 7874 6334 7884 6390
rect 7940 6334 8008 6390
rect 8064 6334 8132 6390
rect 8188 6334 8256 6390
rect 8312 6334 8380 6390
rect 8436 6334 8504 6390
rect 8560 6334 8628 6390
rect 8684 6334 8752 6390
rect 8808 6334 8876 6390
rect 8932 6334 9000 6390
rect 9056 6334 9124 6390
rect 9180 6334 9248 6390
rect 9304 6334 9372 6390
rect 9428 6334 9496 6390
rect 9552 6334 9620 6390
rect 9676 6334 9744 6390
rect 9800 6334 9810 6390
rect 7874 6266 9810 6334
rect 7874 6210 7884 6266
rect 7940 6210 8008 6266
rect 8064 6210 8132 6266
rect 8188 6210 8256 6266
rect 8312 6210 8380 6266
rect 8436 6210 8504 6266
rect 8560 6210 8628 6266
rect 8684 6210 8752 6266
rect 8808 6210 8876 6266
rect 8932 6210 9000 6266
rect 9056 6210 9124 6266
rect 9180 6210 9248 6266
rect 9304 6210 9372 6266
rect 9428 6210 9496 6266
rect 9552 6210 9620 6266
rect 9676 6210 9744 6266
rect 9800 6210 9810 6266
rect 7874 6142 9810 6210
rect 7874 6086 7884 6142
rect 7940 6086 8008 6142
rect 8064 6086 8132 6142
rect 8188 6086 8256 6142
rect 8312 6086 8380 6142
rect 8436 6086 8504 6142
rect 8560 6086 8628 6142
rect 8684 6086 8752 6142
rect 8808 6086 8876 6142
rect 8932 6086 9000 6142
rect 9056 6086 9124 6142
rect 9180 6086 9248 6142
rect 9304 6086 9372 6142
rect 9428 6086 9496 6142
rect 9552 6086 9620 6142
rect 9676 6086 9744 6142
rect 9800 6086 9810 6142
rect 7874 6018 9810 6086
rect 7874 5962 7884 6018
rect 7940 5962 8008 6018
rect 8064 5962 8132 6018
rect 8188 5962 8256 6018
rect 8312 5962 8380 6018
rect 8436 5962 8504 6018
rect 8560 5962 8628 6018
rect 8684 5962 8752 6018
rect 8808 5962 8876 6018
rect 8932 5962 9000 6018
rect 9056 5962 9124 6018
rect 9180 5962 9248 6018
rect 9304 5962 9372 6018
rect 9428 5962 9496 6018
rect 9552 5962 9620 6018
rect 9676 5962 9744 6018
rect 9800 5962 9810 6018
rect 7874 5894 9810 5962
rect 7874 5838 7884 5894
rect 7940 5838 8008 5894
rect 8064 5838 8132 5894
rect 8188 5838 8256 5894
rect 8312 5838 8380 5894
rect 8436 5838 8504 5894
rect 8560 5838 8628 5894
rect 8684 5838 8752 5894
rect 8808 5838 8876 5894
rect 8932 5838 9000 5894
rect 9056 5838 9124 5894
rect 9180 5838 9248 5894
rect 9304 5838 9372 5894
rect 9428 5838 9496 5894
rect 9552 5838 9620 5894
rect 9676 5838 9744 5894
rect 9800 5838 9810 5894
rect 7874 5770 9810 5838
rect 7874 5714 7884 5770
rect 7940 5714 8008 5770
rect 8064 5714 8132 5770
rect 8188 5714 8256 5770
rect 8312 5714 8380 5770
rect 8436 5714 8504 5770
rect 8560 5714 8628 5770
rect 8684 5714 8752 5770
rect 8808 5714 8876 5770
rect 8932 5714 9000 5770
rect 9056 5714 9124 5770
rect 9180 5714 9248 5770
rect 9304 5714 9372 5770
rect 9428 5714 9496 5770
rect 9552 5714 9620 5770
rect 9676 5714 9744 5770
rect 9800 5714 9810 5770
rect 7874 5646 9810 5714
rect 7874 5590 7884 5646
rect 7940 5590 8008 5646
rect 8064 5590 8132 5646
rect 8188 5590 8256 5646
rect 8312 5590 8380 5646
rect 8436 5590 8504 5646
rect 8560 5590 8628 5646
rect 8684 5590 8752 5646
rect 8808 5590 8876 5646
rect 8932 5590 9000 5646
rect 9056 5590 9124 5646
rect 9180 5590 9248 5646
rect 9304 5590 9372 5646
rect 9428 5590 9496 5646
rect 9552 5590 9620 5646
rect 9676 5590 9744 5646
rect 9800 5590 9810 5646
rect 7874 5522 9810 5590
rect 7874 5466 7884 5522
rect 7940 5466 8008 5522
rect 8064 5466 8132 5522
rect 8188 5466 8256 5522
rect 8312 5466 8380 5522
rect 8436 5466 8504 5522
rect 8560 5466 8628 5522
rect 8684 5466 8752 5522
rect 8808 5466 8876 5522
rect 8932 5466 9000 5522
rect 9056 5466 9124 5522
rect 9180 5466 9248 5522
rect 9304 5466 9372 5522
rect 9428 5466 9496 5522
rect 9552 5466 9620 5522
rect 9676 5466 9744 5522
rect 9800 5466 9810 5522
rect 7874 5398 9810 5466
rect 7874 5342 7884 5398
rect 7940 5342 8008 5398
rect 8064 5342 8132 5398
rect 8188 5342 8256 5398
rect 8312 5342 8380 5398
rect 8436 5342 8504 5398
rect 8560 5342 8628 5398
rect 8684 5342 8752 5398
rect 8808 5342 8876 5398
rect 8932 5342 9000 5398
rect 9056 5342 9124 5398
rect 9180 5342 9248 5398
rect 9304 5342 9372 5398
rect 9428 5342 9496 5398
rect 9552 5342 9620 5398
rect 9676 5342 9744 5398
rect 9800 5342 9810 5398
rect 7874 5274 9810 5342
rect 7874 5218 7884 5274
rect 7940 5218 8008 5274
rect 8064 5218 8132 5274
rect 8188 5218 8256 5274
rect 8312 5218 8380 5274
rect 8436 5218 8504 5274
rect 8560 5218 8628 5274
rect 8684 5218 8752 5274
rect 8808 5218 8876 5274
rect 8932 5218 9000 5274
rect 9056 5218 9124 5274
rect 9180 5218 9248 5274
rect 9304 5218 9372 5274
rect 9428 5218 9496 5274
rect 9552 5218 9620 5274
rect 9676 5218 9744 5274
rect 9800 5218 9810 5274
rect 7874 5150 9810 5218
rect 7874 5094 7884 5150
rect 7940 5094 8008 5150
rect 8064 5094 8132 5150
rect 8188 5094 8256 5150
rect 8312 5094 8380 5150
rect 8436 5094 8504 5150
rect 8560 5094 8628 5150
rect 8684 5094 8752 5150
rect 8808 5094 8876 5150
rect 8932 5094 9000 5150
rect 9056 5094 9124 5150
rect 9180 5094 9248 5150
rect 9304 5094 9372 5150
rect 9428 5094 9496 5150
rect 9552 5094 9620 5150
rect 9676 5094 9744 5150
rect 9800 5094 9810 5150
rect 7874 5026 9810 5094
rect 7874 4970 7884 5026
rect 7940 4970 8008 5026
rect 8064 4970 8132 5026
rect 8188 4970 8256 5026
rect 8312 4970 8380 5026
rect 8436 4970 8504 5026
rect 8560 4970 8628 5026
rect 8684 4970 8752 5026
rect 8808 4970 8876 5026
rect 8932 4970 9000 5026
rect 9056 4970 9124 5026
rect 9180 4970 9248 5026
rect 9304 4970 9372 5026
rect 9428 4970 9496 5026
rect 9552 4970 9620 5026
rect 9676 4970 9744 5026
rect 9800 4970 9810 5026
rect 7874 4902 9810 4970
rect 7874 4846 7884 4902
rect 7940 4846 8008 4902
rect 8064 4846 8132 4902
rect 8188 4846 8256 4902
rect 8312 4846 8380 4902
rect 8436 4846 8504 4902
rect 8560 4846 8628 4902
rect 8684 4846 8752 4902
rect 8808 4846 8876 4902
rect 8932 4846 9000 4902
rect 9056 4846 9124 4902
rect 9180 4846 9248 4902
rect 9304 4846 9372 4902
rect 9428 4846 9496 4902
rect 9552 4846 9620 4902
rect 9676 4846 9744 4902
rect 9800 4846 9810 4902
rect 7874 4836 9810 4846
rect 10244 7754 12180 7764
rect 10244 7698 10254 7754
rect 10310 7698 10378 7754
rect 10434 7698 10502 7754
rect 10558 7698 10626 7754
rect 10682 7698 10750 7754
rect 10806 7698 10874 7754
rect 10930 7698 10998 7754
rect 11054 7698 11122 7754
rect 11178 7698 11246 7754
rect 11302 7698 11370 7754
rect 11426 7698 11494 7754
rect 11550 7698 11618 7754
rect 11674 7698 11742 7754
rect 11798 7698 11866 7754
rect 11922 7698 11990 7754
rect 12046 7698 12114 7754
rect 12170 7698 12180 7754
rect 10244 7630 12180 7698
rect 10244 7574 10254 7630
rect 10310 7574 10378 7630
rect 10434 7574 10502 7630
rect 10558 7574 10626 7630
rect 10682 7574 10750 7630
rect 10806 7574 10874 7630
rect 10930 7574 10998 7630
rect 11054 7574 11122 7630
rect 11178 7574 11246 7630
rect 11302 7574 11370 7630
rect 11426 7574 11494 7630
rect 11550 7574 11618 7630
rect 11674 7574 11742 7630
rect 11798 7574 11866 7630
rect 11922 7574 11990 7630
rect 12046 7574 12114 7630
rect 12170 7574 12180 7630
rect 10244 7506 12180 7574
rect 10244 7450 10254 7506
rect 10310 7450 10378 7506
rect 10434 7450 10502 7506
rect 10558 7450 10626 7506
rect 10682 7450 10750 7506
rect 10806 7450 10874 7506
rect 10930 7450 10998 7506
rect 11054 7450 11122 7506
rect 11178 7450 11246 7506
rect 11302 7450 11370 7506
rect 11426 7450 11494 7506
rect 11550 7450 11618 7506
rect 11674 7450 11742 7506
rect 11798 7450 11866 7506
rect 11922 7450 11990 7506
rect 12046 7450 12114 7506
rect 12170 7450 12180 7506
rect 10244 7382 12180 7450
rect 10244 7326 10254 7382
rect 10310 7326 10378 7382
rect 10434 7326 10502 7382
rect 10558 7326 10626 7382
rect 10682 7326 10750 7382
rect 10806 7326 10874 7382
rect 10930 7326 10998 7382
rect 11054 7326 11122 7382
rect 11178 7326 11246 7382
rect 11302 7326 11370 7382
rect 11426 7326 11494 7382
rect 11550 7326 11618 7382
rect 11674 7326 11742 7382
rect 11798 7326 11866 7382
rect 11922 7326 11990 7382
rect 12046 7326 12114 7382
rect 12170 7326 12180 7382
rect 10244 7258 12180 7326
rect 10244 7202 10254 7258
rect 10310 7202 10378 7258
rect 10434 7202 10502 7258
rect 10558 7202 10626 7258
rect 10682 7202 10750 7258
rect 10806 7202 10874 7258
rect 10930 7202 10998 7258
rect 11054 7202 11122 7258
rect 11178 7202 11246 7258
rect 11302 7202 11370 7258
rect 11426 7202 11494 7258
rect 11550 7202 11618 7258
rect 11674 7202 11742 7258
rect 11798 7202 11866 7258
rect 11922 7202 11990 7258
rect 12046 7202 12114 7258
rect 12170 7202 12180 7258
rect 10244 7134 12180 7202
rect 10244 7078 10254 7134
rect 10310 7078 10378 7134
rect 10434 7078 10502 7134
rect 10558 7078 10626 7134
rect 10682 7078 10750 7134
rect 10806 7078 10874 7134
rect 10930 7078 10998 7134
rect 11054 7078 11122 7134
rect 11178 7078 11246 7134
rect 11302 7078 11370 7134
rect 11426 7078 11494 7134
rect 11550 7078 11618 7134
rect 11674 7078 11742 7134
rect 11798 7078 11866 7134
rect 11922 7078 11990 7134
rect 12046 7078 12114 7134
rect 12170 7078 12180 7134
rect 10244 7010 12180 7078
rect 10244 6954 10254 7010
rect 10310 6954 10378 7010
rect 10434 6954 10502 7010
rect 10558 6954 10626 7010
rect 10682 6954 10750 7010
rect 10806 6954 10874 7010
rect 10930 6954 10998 7010
rect 11054 6954 11122 7010
rect 11178 6954 11246 7010
rect 11302 6954 11370 7010
rect 11426 6954 11494 7010
rect 11550 6954 11618 7010
rect 11674 6954 11742 7010
rect 11798 6954 11866 7010
rect 11922 6954 11990 7010
rect 12046 6954 12114 7010
rect 12170 6954 12180 7010
rect 10244 6886 12180 6954
rect 10244 6830 10254 6886
rect 10310 6830 10378 6886
rect 10434 6830 10502 6886
rect 10558 6830 10626 6886
rect 10682 6830 10750 6886
rect 10806 6830 10874 6886
rect 10930 6830 10998 6886
rect 11054 6830 11122 6886
rect 11178 6830 11246 6886
rect 11302 6830 11370 6886
rect 11426 6830 11494 6886
rect 11550 6830 11618 6886
rect 11674 6830 11742 6886
rect 11798 6830 11866 6886
rect 11922 6830 11990 6886
rect 12046 6830 12114 6886
rect 12170 6830 12180 6886
rect 10244 6762 12180 6830
rect 10244 6706 10254 6762
rect 10310 6706 10378 6762
rect 10434 6706 10502 6762
rect 10558 6706 10626 6762
rect 10682 6706 10750 6762
rect 10806 6706 10874 6762
rect 10930 6706 10998 6762
rect 11054 6706 11122 6762
rect 11178 6706 11246 6762
rect 11302 6706 11370 6762
rect 11426 6706 11494 6762
rect 11550 6706 11618 6762
rect 11674 6706 11742 6762
rect 11798 6706 11866 6762
rect 11922 6706 11990 6762
rect 12046 6706 12114 6762
rect 12170 6706 12180 6762
rect 10244 6638 12180 6706
rect 10244 6582 10254 6638
rect 10310 6582 10378 6638
rect 10434 6582 10502 6638
rect 10558 6582 10626 6638
rect 10682 6582 10750 6638
rect 10806 6582 10874 6638
rect 10930 6582 10998 6638
rect 11054 6582 11122 6638
rect 11178 6582 11246 6638
rect 11302 6582 11370 6638
rect 11426 6582 11494 6638
rect 11550 6582 11618 6638
rect 11674 6582 11742 6638
rect 11798 6582 11866 6638
rect 11922 6582 11990 6638
rect 12046 6582 12114 6638
rect 12170 6582 12180 6638
rect 10244 6514 12180 6582
rect 10244 6458 10254 6514
rect 10310 6458 10378 6514
rect 10434 6458 10502 6514
rect 10558 6458 10626 6514
rect 10682 6458 10750 6514
rect 10806 6458 10874 6514
rect 10930 6458 10998 6514
rect 11054 6458 11122 6514
rect 11178 6458 11246 6514
rect 11302 6458 11370 6514
rect 11426 6458 11494 6514
rect 11550 6458 11618 6514
rect 11674 6458 11742 6514
rect 11798 6458 11866 6514
rect 11922 6458 11990 6514
rect 12046 6458 12114 6514
rect 12170 6458 12180 6514
rect 10244 6390 12180 6458
rect 10244 6334 10254 6390
rect 10310 6334 10378 6390
rect 10434 6334 10502 6390
rect 10558 6334 10626 6390
rect 10682 6334 10750 6390
rect 10806 6334 10874 6390
rect 10930 6334 10998 6390
rect 11054 6334 11122 6390
rect 11178 6334 11246 6390
rect 11302 6334 11370 6390
rect 11426 6334 11494 6390
rect 11550 6334 11618 6390
rect 11674 6334 11742 6390
rect 11798 6334 11866 6390
rect 11922 6334 11990 6390
rect 12046 6334 12114 6390
rect 12170 6334 12180 6390
rect 10244 6266 12180 6334
rect 10244 6210 10254 6266
rect 10310 6210 10378 6266
rect 10434 6210 10502 6266
rect 10558 6210 10626 6266
rect 10682 6210 10750 6266
rect 10806 6210 10874 6266
rect 10930 6210 10998 6266
rect 11054 6210 11122 6266
rect 11178 6210 11246 6266
rect 11302 6210 11370 6266
rect 11426 6210 11494 6266
rect 11550 6210 11618 6266
rect 11674 6210 11742 6266
rect 11798 6210 11866 6266
rect 11922 6210 11990 6266
rect 12046 6210 12114 6266
rect 12170 6210 12180 6266
rect 10244 6142 12180 6210
rect 10244 6086 10254 6142
rect 10310 6086 10378 6142
rect 10434 6086 10502 6142
rect 10558 6086 10626 6142
rect 10682 6086 10750 6142
rect 10806 6086 10874 6142
rect 10930 6086 10998 6142
rect 11054 6086 11122 6142
rect 11178 6086 11246 6142
rect 11302 6086 11370 6142
rect 11426 6086 11494 6142
rect 11550 6086 11618 6142
rect 11674 6086 11742 6142
rect 11798 6086 11866 6142
rect 11922 6086 11990 6142
rect 12046 6086 12114 6142
rect 12170 6086 12180 6142
rect 10244 6018 12180 6086
rect 10244 5962 10254 6018
rect 10310 5962 10378 6018
rect 10434 5962 10502 6018
rect 10558 5962 10626 6018
rect 10682 5962 10750 6018
rect 10806 5962 10874 6018
rect 10930 5962 10998 6018
rect 11054 5962 11122 6018
rect 11178 5962 11246 6018
rect 11302 5962 11370 6018
rect 11426 5962 11494 6018
rect 11550 5962 11618 6018
rect 11674 5962 11742 6018
rect 11798 5962 11866 6018
rect 11922 5962 11990 6018
rect 12046 5962 12114 6018
rect 12170 5962 12180 6018
rect 10244 5894 12180 5962
rect 10244 5838 10254 5894
rect 10310 5838 10378 5894
rect 10434 5838 10502 5894
rect 10558 5838 10626 5894
rect 10682 5838 10750 5894
rect 10806 5838 10874 5894
rect 10930 5838 10998 5894
rect 11054 5838 11122 5894
rect 11178 5838 11246 5894
rect 11302 5838 11370 5894
rect 11426 5838 11494 5894
rect 11550 5838 11618 5894
rect 11674 5838 11742 5894
rect 11798 5838 11866 5894
rect 11922 5838 11990 5894
rect 12046 5838 12114 5894
rect 12170 5838 12180 5894
rect 10244 5770 12180 5838
rect 10244 5714 10254 5770
rect 10310 5714 10378 5770
rect 10434 5714 10502 5770
rect 10558 5714 10626 5770
rect 10682 5714 10750 5770
rect 10806 5714 10874 5770
rect 10930 5714 10998 5770
rect 11054 5714 11122 5770
rect 11178 5714 11246 5770
rect 11302 5714 11370 5770
rect 11426 5714 11494 5770
rect 11550 5714 11618 5770
rect 11674 5714 11742 5770
rect 11798 5714 11866 5770
rect 11922 5714 11990 5770
rect 12046 5714 12114 5770
rect 12170 5714 12180 5770
rect 10244 5646 12180 5714
rect 10244 5590 10254 5646
rect 10310 5590 10378 5646
rect 10434 5590 10502 5646
rect 10558 5590 10626 5646
rect 10682 5590 10750 5646
rect 10806 5590 10874 5646
rect 10930 5590 10998 5646
rect 11054 5590 11122 5646
rect 11178 5590 11246 5646
rect 11302 5590 11370 5646
rect 11426 5590 11494 5646
rect 11550 5590 11618 5646
rect 11674 5590 11742 5646
rect 11798 5590 11866 5646
rect 11922 5590 11990 5646
rect 12046 5590 12114 5646
rect 12170 5590 12180 5646
rect 10244 5522 12180 5590
rect 10244 5466 10254 5522
rect 10310 5466 10378 5522
rect 10434 5466 10502 5522
rect 10558 5466 10626 5522
rect 10682 5466 10750 5522
rect 10806 5466 10874 5522
rect 10930 5466 10998 5522
rect 11054 5466 11122 5522
rect 11178 5466 11246 5522
rect 11302 5466 11370 5522
rect 11426 5466 11494 5522
rect 11550 5466 11618 5522
rect 11674 5466 11742 5522
rect 11798 5466 11866 5522
rect 11922 5466 11990 5522
rect 12046 5466 12114 5522
rect 12170 5466 12180 5522
rect 10244 5398 12180 5466
rect 10244 5342 10254 5398
rect 10310 5342 10378 5398
rect 10434 5342 10502 5398
rect 10558 5342 10626 5398
rect 10682 5342 10750 5398
rect 10806 5342 10874 5398
rect 10930 5342 10998 5398
rect 11054 5342 11122 5398
rect 11178 5342 11246 5398
rect 11302 5342 11370 5398
rect 11426 5342 11494 5398
rect 11550 5342 11618 5398
rect 11674 5342 11742 5398
rect 11798 5342 11866 5398
rect 11922 5342 11990 5398
rect 12046 5342 12114 5398
rect 12170 5342 12180 5398
rect 10244 5274 12180 5342
rect 10244 5218 10254 5274
rect 10310 5218 10378 5274
rect 10434 5218 10502 5274
rect 10558 5218 10626 5274
rect 10682 5218 10750 5274
rect 10806 5218 10874 5274
rect 10930 5218 10998 5274
rect 11054 5218 11122 5274
rect 11178 5218 11246 5274
rect 11302 5218 11370 5274
rect 11426 5218 11494 5274
rect 11550 5218 11618 5274
rect 11674 5218 11742 5274
rect 11798 5218 11866 5274
rect 11922 5218 11990 5274
rect 12046 5218 12114 5274
rect 12170 5218 12180 5274
rect 10244 5150 12180 5218
rect 10244 5094 10254 5150
rect 10310 5094 10378 5150
rect 10434 5094 10502 5150
rect 10558 5094 10626 5150
rect 10682 5094 10750 5150
rect 10806 5094 10874 5150
rect 10930 5094 10998 5150
rect 11054 5094 11122 5150
rect 11178 5094 11246 5150
rect 11302 5094 11370 5150
rect 11426 5094 11494 5150
rect 11550 5094 11618 5150
rect 11674 5094 11742 5150
rect 11798 5094 11866 5150
rect 11922 5094 11990 5150
rect 12046 5094 12114 5150
rect 12170 5094 12180 5150
rect 10244 5026 12180 5094
rect 10244 4970 10254 5026
rect 10310 4970 10378 5026
rect 10434 4970 10502 5026
rect 10558 4970 10626 5026
rect 10682 4970 10750 5026
rect 10806 4970 10874 5026
rect 10930 4970 10998 5026
rect 11054 4970 11122 5026
rect 11178 4970 11246 5026
rect 11302 4970 11370 5026
rect 11426 4970 11494 5026
rect 11550 4970 11618 5026
rect 11674 4970 11742 5026
rect 11798 4970 11866 5026
rect 11922 4970 11990 5026
rect 12046 4970 12114 5026
rect 12170 4970 12180 5026
rect 10244 4902 12180 4970
rect 10244 4846 10254 4902
rect 10310 4846 10378 4902
rect 10434 4846 10502 4902
rect 10558 4846 10626 4902
rect 10682 4846 10750 4902
rect 10806 4846 10874 4902
rect 10930 4846 10998 4902
rect 11054 4846 11122 4902
rect 11178 4846 11246 4902
rect 11302 4846 11370 4902
rect 11426 4846 11494 4902
rect 11550 4846 11618 4902
rect 11674 4846 11742 4902
rect 11798 4846 11866 4902
rect 11922 4846 11990 4902
rect 12046 4846 12114 4902
rect 12170 4846 12180 4902
rect 10244 4836 12180 4846
rect 12861 7754 14673 7764
rect 12861 7698 12871 7754
rect 12927 7698 12995 7754
rect 13051 7698 13119 7754
rect 13175 7698 13243 7754
rect 13299 7698 13367 7754
rect 13423 7698 13491 7754
rect 13547 7698 13615 7754
rect 13671 7698 13739 7754
rect 13795 7698 13863 7754
rect 13919 7698 13987 7754
rect 14043 7698 14111 7754
rect 14167 7698 14235 7754
rect 14291 7698 14359 7754
rect 14415 7698 14483 7754
rect 14539 7698 14607 7754
rect 14663 7698 14673 7754
rect 12861 7630 14673 7698
rect 12861 7574 12871 7630
rect 12927 7574 12995 7630
rect 13051 7574 13119 7630
rect 13175 7574 13243 7630
rect 13299 7574 13367 7630
rect 13423 7574 13491 7630
rect 13547 7574 13615 7630
rect 13671 7574 13739 7630
rect 13795 7574 13863 7630
rect 13919 7574 13987 7630
rect 14043 7574 14111 7630
rect 14167 7574 14235 7630
rect 14291 7574 14359 7630
rect 14415 7574 14483 7630
rect 14539 7574 14607 7630
rect 14663 7574 14673 7630
rect 12861 7506 14673 7574
rect 12861 7450 12871 7506
rect 12927 7450 12995 7506
rect 13051 7450 13119 7506
rect 13175 7450 13243 7506
rect 13299 7450 13367 7506
rect 13423 7450 13491 7506
rect 13547 7450 13615 7506
rect 13671 7450 13739 7506
rect 13795 7450 13863 7506
rect 13919 7450 13987 7506
rect 14043 7450 14111 7506
rect 14167 7450 14235 7506
rect 14291 7450 14359 7506
rect 14415 7450 14483 7506
rect 14539 7450 14607 7506
rect 14663 7450 14673 7506
rect 12861 7382 14673 7450
rect 12861 7326 12871 7382
rect 12927 7326 12995 7382
rect 13051 7326 13119 7382
rect 13175 7326 13243 7382
rect 13299 7326 13367 7382
rect 13423 7326 13491 7382
rect 13547 7326 13615 7382
rect 13671 7326 13739 7382
rect 13795 7326 13863 7382
rect 13919 7326 13987 7382
rect 14043 7326 14111 7382
rect 14167 7326 14235 7382
rect 14291 7326 14359 7382
rect 14415 7326 14483 7382
rect 14539 7326 14607 7382
rect 14663 7326 14673 7382
rect 12861 7258 14673 7326
rect 12861 7202 12871 7258
rect 12927 7202 12995 7258
rect 13051 7202 13119 7258
rect 13175 7202 13243 7258
rect 13299 7202 13367 7258
rect 13423 7202 13491 7258
rect 13547 7202 13615 7258
rect 13671 7202 13739 7258
rect 13795 7202 13863 7258
rect 13919 7202 13987 7258
rect 14043 7202 14111 7258
rect 14167 7202 14235 7258
rect 14291 7202 14359 7258
rect 14415 7202 14483 7258
rect 14539 7202 14607 7258
rect 14663 7202 14673 7258
rect 12861 7134 14673 7202
rect 12861 7078 12871 7134
rect 12927 7078 12995 7134
rect 13051 7078 13119 7134
rect 13175 7078 13243 7134
rect 13299 7078 13367 7134
rect 13423 7078 13491 7134
rect 13547 7078 13615 7134
rect 13671 7078 13739 7134
rect 13795 7078 13863 7134
rect 13919 7078 13987 7134
rect 14043 7078 14111 7134
rect 14167 7078 14235 7134
rect 14291 7078 14359 7134
rect 14415 7078 14483 7134
rect 14539 7078 14607 7134
rect 14663 7078 14673 7134
rect 12861 7010 14673 7078
rect 12861 6954 12871 7010
rect 12927 6954 12995 7010
rect 13051 6954 13119 7010
rect 13175 6954 13243 7010
rect 13299 6954 13367 7010
rect 13423 6954 13491 7010
rect 13547 6954 13615 7010
rect 13671 6954 13739 7010
rect 13795 6954 13863 7010
rect 13919 6954 13987 7010
rect 14043 6954 14111 7010
rect 14167 6954 14235 7010
rect 14291 6954 14359 7010
rect 14415 6954 14483 7010
rect 14539 6954 14607 7010
rect 14663 6954 14673 7010
rect 12861 6886 14673 6954
rect 12861 6830 12871 6886
rect 12927 6830 12995 6886
rect 13051 6830 13119 6886
rect 13175 6830 13243 6886
rect 13299 6830 13367 6886
rect 13423 6830 13491 6886
rect 13547 6830 13615 6886
rect 13671 6830 13739 6886
rect 13795 6830 13863 6886
rect 13919 6830 13987 6886
rect 14043 6830 14111 6886
rect 14167 6830 14235 6886
rect 14291 6830 14359 6886
rect 14415 6830 14483 6886
rect 14539 6830 14607 6886
rect 14663 6830 14673 6886
rect 12861 6762 14673 6830
rect 12861 6706 12871 6762
rect 12927 6706 12995 6762
rect 13051 6706 13119 6762
rect 13175 6706 13243 6762
rect 13299 6706 13367 6762
rect 13423 6706 13491 6762
rect 13547 6706 13615 6762
rect 13671 6706 13739 6762
rect 13795 6706 13863 6762
rect 13919 6706 13987 6762
rect 14043 6706 14111 6762
rect 14167 6706 14235 6762
rect 14291 6706 14359 6762
rect 14415 6706 14483 6762
rect 14539 6706 14607 6762
rect 14663 6706 14673 6762
rect 12861 6638 14673 6706
rect 12861 6582 12871 6638
rect 12927 6582 12995 6638
rect 13051 6582 13119 6638
rect 13175 6582 13243 6638
rect 13299 6582 13367 6638
rect 13423 6582 13491 6638
rect 13547 6582 13615 6638
rect 13671 6582 13739 6638
rect 13795 6582 13863 6638
rect 13919 6582 13987 6638
rect 14043 6582 14111 6638
rect 14167 6582 14235 6638
rect 14291 6582 14359 6638
rect 14415 6582 14483 6638
rect 14539 6582 14607 6638
rect 14663 6582 14673 6638
rect 12861 6514 14673 6582
rect 12861 6458 12871 6514
rect 12927 6458 12995 6514
rect 13051 6458 13119 6514
rect 13175 6458 13243 6514
rect 13299 6458 13367 6514
rect 13423 6458 13491 6514
rect 13547 6458 13615 6514
rect 13671 6458 13739 6514
rect 13795 6458 13863 6514
rect 13919 6458 13987 6514
rect 14043 6458 14111 6514
rect 14167 6458 14235 6514
rect 14291 6458 14359 6514
rect 14415 6458 14483 6514
rect 14539 6458 14607 6514
rect 14663 6458 14673 6514
rect 12861 6390 14673 6458
rect 12861 6334 12871 6390
rect 12927 6334 12995 6390
rect 13051 6334 13119 6390
rect 13175 6334 13243 6390
rect 13299 6334 13367 6390
rect 13423 6334 13491 6390
rect 13547 6334 13615 6390
rect 13671 6334 13739 6390
rect 13795 6334 13863 6390
rect 13919 6334 13987 6390
rect 14043 6334 14111 6390
rect 14167 6334 14235 6390
rect 14291 6334 14359 6390
rect 14415 6334 14483 6390
rect 14539 6334 14607 6390
rect 14663 6334 14673 6390
rect 12861 6266 14673 6334
rect 12861 6210 12871 6266
rect 12927 6210 12995 6266
rect 13051 6210 13119 6266
rect 13175 6210 13243 6266
rect 13299 6210 13367 6266
rect 13423 6210 13491 6266
rect 13547 6210 13615 6266
rect 13671 6210 13739 6266
rect 13795 6210 13863 6266
rect 13919 6210 13987 6266
rect 14043 6210 14111 6266
rect 14167 6210 14235 6266
rect 14291 6210 14359 6266
rect 14415 6210 14483 6266
rect 14539 6210 14607 6266
rect 14663 6210 14673 6266
rect 12861 6142 14673 6210
rect 12861 6086 12871 6142
rect 12927 6086 12995 6142
rect 13051 6086 13119 6142
rect 13175 6086 13243 6142
rect 13299 6086 13367 6142
rect 13423 6086 13491 6142
rect 13547 6086 13615 6142
rect 13671 6086 13739 6142
rect 13795 6086 13863 6142
rect 13919 6086 13987 6142
rect 14043 6086 14111 6142
rect 14167 6086 14235 6142
rect 14291 6086 14359 6142
rect 14415 6086 14483 6142
rect 14539 6086 14607 6142
rect 14663 6086 14673 6142
rect 12861 6018 14673 6086
rect 12861 5962 12871 6018
rect 12927 5962 12995 6018
rect 13051 5962 13119 6018
rect 13175 5962 13243 6018
rect 13299 5962 13367 6018
rect 13423 5962 13491 6018
rect 13547 5962 13615 6018
rect 13671 5962 13739 6018
rect 13795 5962 13863 6018
rect 13919 5962 13987 6018
rect 14043 5962 14111 6018
rect 14167 5962 14235 6018
rect 14291 5962 14359 6018
rect 14415 5962 14483 6018
rect 14539 5962 14607 6018
rect 14663 5962 14673 6018
rect 12861 5894 14673 5962
rect 12861 5838 12871 5894
rect 12927 5838 12995 5894
rect 13051 5838 13119 5894
rect 13175 5838 13243 5894
rect 13299 5838 13367 5894
rect 13423 5838 13491 5894
rect 13547 5838 13615 5894
rect 13671 5838 13739 5894
rect 13795 5838 13863 5894
rect 13919 5838 13987 5894
rect 14043 5838 14111 5894
rect 14167 5838 14235 5894
rect 14291 5838 14359 5894
rect 14415 5838 14483 5894
rect 14539 5838 14607 5894
rect 14663 5838 14673 5894
rect 12861 5770 14673 5838
rect 12861 5714 12871 5770
rect 12927 5714 12995 5770
rect 13051 5714 13119 5770
rect 13175 5714 13243 5770
rect 13299 5714 13367 5770
rect 13423 5714 13491 5770
rect 13547 5714 13615 5770
rect 13671 5714 13739 5770
rect 13795 5714 13863 5770
rect 13919 5714 13987 5770
rect 14043 5714 14111 5770
rect 14167 5714 14235 5770
rect 14291 5714 14359 5770
rect 14415 5714 14483 5770
rect 14539 5714 14607 5770
rect 14663 5714 14673 5770
rect 12861 5646 14673 5714
rect 12861 5590 12871 5646
rect 12927 5590 12995 5646
rect 13051 5590 13119 5646
rect 13175 5590 13243 5646
rect 13299 5590 13367 5646
rect 13423 5590 13491 5646
rect 13547 5590 13615 5646
rect 13671 5590 13739 5646
rect 13795 5590 13863 5646
rect 13919 5590 13987 5646
rect 14043 5590 14111 5646
rect 14167 5590 14235 5646
rect 14291 5590 14359 5646
rect 14415 5590 14483 5646
rect 14539 5590 14607 5646
rect 14663 5590 14673 5646
rect 12861 5522 14673 5590
rect 12861 5466 12871 5522
rect 12927 5466 12995 5522
rect 13051 5466 13119 5522
rect 13175 5466 13243 5522
rect 13299 5466 13367 5522
rect 13423 5466 13491 5522
rect 13547 5466 13615 5522
rect 13671 5466 13739 5522
rect 13795 5466 13863 5522
rect 13919 5466 13987 5522
rect 14043 5466 14111 5522
rect 14167 5466 14235 5522
rect 14291 5466 14359 5522
rect 14415 5466 14483 5522
rect 14539 5466 14607 5522
rect 14663 5466 14673 5522
rect 12861 5398 14673 5466
rect 12861 5342 12871 5398
rect 12927 5342 12995 5398
rect 13051 5342 13119 5398
rect 13175 5342 13243 5398
rect 13299 5342 13367 5398
rect 13423 5342 13491 5398
rect 13547 5342 13615 5398
rect 13671 5342 13739 5398
rect 13795 5342 13863 5398
rect 13919 5342 13987 5398
rect 14043 5342 14111 5398
rect 14167 5342 14235 5398
rect 14291 5342 14359 5398
rect 14415 5342 14483 5398
rect 14539 5342 14607 5398
rect 14663 5342 14673 5398
rect 12861 5274 14673 5342
rect 12861 5218 12871 5274
rect 12927 5218 12995 5274
rect 13051 5218 13119 5274
rect 13175 5218 13243 5274
rect 13299 5218 13367 5274
rect 13423 5218 13491 5274
rect 13547 5218 13615 5274
rect 13671 5218 13739 5274
rect 13795 5218 13863 5274
rect 13919 5218 13987 5274
rect 14043 5218 14111 5274
rect 14167 5218 14235 5274
rect 14291 5218 14359 5274
rect 14415 5218 14483 5274
rect 14539 5218 14607 5274
rect 14663 5218 14673 5274
rect 12861 5150 14673 5218
rect 12861 5094 12871 5150
rect 12927 5094 12995 5150
rect 13051 5094 13119 5150
rect 13175 5094 13243 5150
rect 13299 5094 13367 5150
rect 13423 5094 13491 5150
rect 13547 5094 13615 5150
rect 13671 5094 13739 5150
rect 13795 5094 13863 5150
rect 13919 5094 13987 5150
rect 14043 5094 14111 5150
rect 14167 5094 14235 5150
rect 14291 5094 14359 5150
rect 14415 5094 14483 5150
rect 14539 5094 14607 5150
rect 14663 5094 14673 5150
rect 12861 5026 14673 5094
rect 12861 4970 12871 5026
rect 12927 4970 12995 5026
rect 13051 4970 13119 5026
rect 13175 4970 13243 5026
rect 13299 4970 13367 5026
rect 13423 4970 13491 5026
rect 13547 4970 13615 5026
rect 13671 4970 13739 5026
rect 13795 4970 13863 5026
rect 13919 4970 13987 5026
rect 14043 4970 14111 5026
rect 14167 4970 14235 5026
rect 14291 4970 14359 5026
rect 14415 4970 14483 5026
rect 14539 4970 14607 5026
rect 14663 4970 14673 5026
rect 12861 4902 14673 4970
rect 12861 4846 12871 4902
rect 12927 4846 12995 4902
rect 13051 4846 13119 4902
rect 13175 4846 13243 4902
rect 13299 4846 13367 4902
rect 13423 4846 13491 4902
rect 13547 4846 13615 4902
rect 13671 4846 13739 4902
rect 13795 4846 13863 4902
rect 13919 4846 13987 4902
rect 14043 4846 14111 4902
rect 14167 4846 14235 4902
rect 14291 4846 14359 4902
rect 14415 4846 14483 4902
rect 14539 4846 14607 4902
rect 14663 4846 14673 4902
rect 12861 4836 14673 4846
rect 10 4804 86 4814
rect 14892 4814 14902 7786
rect 14958 4814 14968 7786
rect 14892 4804 14968 4814
rect 10 4586 86 4596
rect 10 1614 20 4586
rect 76 1614 86 4586
rect 14892 4586 14968 4596
rect 305 4554 2117 4564
rect 305 4498 315 4554
rect 371 4498 439 4554
rect 495 4498 563 4554
rect 619 4498 687 4554
rect 743 4498 811 4554
rect 867 4498 935 4554
rect 991 4498 1059 4554
rect 1115 4498 1183 4554
rect 1239 4498 1307 4554
rect 1363 4498 1431 4554
rect 1487 4498 1555 4554
rect 1611 4498 1679 4554
rect 1735 4498 1803 4554
rect 1859 4498 1927 4554
rect 1983 4498 2051 4554
rect 2107 4498 2117 4554
rect 305 4430 2117 4498
rect 305 4374 315 4430
rect 371 4374 439 4430
rect 495 4374 563 4430
rect 619 4374 687 4430
rect 743 4374 811 4430
rect 867 4374 935 4430
rect 991 4374 1059 4430
rect 1115 4374 1183 4430
rect 1239 4374 1307 4430
rect 1363 4374 1431 4430
rect 1487 4374 1555 4430
rect 1611 4374 1679 4430
rect 1735 4374 1803 4430
rect 1859 4374 1927 4430
rect 1983 4374 2051 4430
rect 2107 4374 2117 4430
rect 305 4306 2117 4374
rect 305 4250 315 4306
rect 371 4250 439 4306
rect 495 4250 563 4306
rect 619 4250 687 4306
rect 743 4250 811 4306
rect 867 4250 935 4306
rect 991 4250 1059 4306
rect 1115 4250 1183 4306
rect 1239 4250 1307 4306
rect 1363 4250 1431 4306
rect 1487 4250 1555 4306
rect 1611 4250 1679 4306
rect 1735 4250 1803 4306
rect 1859 4250 1927 4306
rect 1983 4250 2051 4306
rect 2107 4250 2117 4306
rect 305 4182 2117 4250
rect 305 4126 315 4182
rect 371 4126 439 4182
rect 495 4126 563 4182
rect 619 4126 687 4182
rect 743 4126 811 4182
rect 867 4126 935 4182
rect 991 4126 1059 4182
rect 1115 4126 1183 4182
rect 1239 4126 1307 4182
rect 1363 4126 1431 4182
rect 1487 4126 1555 4182
rect 1611 4126 1679 4182
rect 1735 4126 1803 4182
rect 1859 4126 1927 4182
rect 1983 4126 2051 4182
rect 2107 4126 2117 4182
rect 305 4058 2117 4126
rect 305 4002 315 4058
rect 371 4002 439 4058
rect 495 4002 563 4058
rect 619 4002 687 4058
rect 743 4002 811 4058
rect 867 4002 935 4058
rect 991 4002 1059 4058
rect 1115 4002 1183 4058
rect 1239 4002 1307 4058
rect 1363 4002 1431 4058
rect 1487 4002 1555 4058
rect 1611 4002 1679 4058
rect 1735 4002 1803 4058
rect 1859 4002 1927 4058
rect 1983 4002 2051 4058
rect 2107 4002 2117 4058
rect 305 3934 2117 4002
rect 305 3878 315 3934
rect 371 3878 439 3934
rect 495 3878 563 3934
rect 619 3878 687 3934
rect 743 3878 811 3934
rect 867 3878 935 3934
rect 991 3878 1059 3934
rect 1115 3878 1183 3934
rect 1239 3878 1307 3934
rect 1363 3878 1431 3934
rect 1487 3878 1555 3934
rect 1611 3878 1679 3934
rect 1735 3878 1803 3934
rect 1859 3878 1927 3934
rect 1983 3878 2051 3934
rect 2107 3878 2117 3934
rect 305 3810 2117 3878
rect 305 3754 315 3810
rect 371 3754 439 3810
rect 495 3754 563 3810
rect 619 3754 687 3810
rect 743 3754 811 3810
rect 867 3754 935 3810
rect 991 3754 1059 3810
rect 1115 3754 1183 3810
rect 1239 3754 1307 3810
rect 1363 3754 1431 3810
rect 1487 3754 1555 3810
rect 1611 3754 1679 3810
rect 1735 3754 1803 3810
rect 1859 3754 1927 3810
rect 1983 3754 2051 3810
rect 2107 3754 2117 3810
rect 305 3686 2117 3754
rect 305 3630 315 3686
rect 371 3630 439 3686
rect 495 3630 563 3686
rect 619 3630 687 3686
rect 743 3630 811 3686
rect 867 3630 935 3686
rect 991 3630 1059 3686
rect 1115 3630 1183 3686
rect 1239 3630 1307 3686
rect 1363 3630 1431 3686
rect 1487 3630 1555 3686
rect 1611 3630 1679 3686
rect 1735 3630 1803 3686
rect 1859 3630 1927 3686
rect 1983 3630 2051 3686
rect 2107 3630 2117 3686
rect 305 3562 2117 3630
rect 305 3506 315 3562
rect 371 3506 439 3562
rect 495 3506 563 3562
rect 619 3506 687 3562
rect 743 3506 811 3562
rect 867 3506 935 3562
rect 991 3506 1059 3562
rect 1115 3506 1183 3562
rect 1239 3506 1307 3562
rect 1363 3506 1431 3562
rect 1487 3506 1555 3562
rect 1611 3506 1679 3562
rect 1735 3506 1803 3562
rect 1859 3506 1927 3562
rect 1983 3506 2051 3562
rect 2107 3506 2117 3562
rect 305 3438 2117 3506
rect 305 3382 315 3438
rect 371 3382 439 3438
rect 495 3382 563 3438
rect 619 3382 687 3438
rect 743 3382 811 3438
rect 867 3382 935 3438
rect 991 3382 1059 3438
rect 1115 3382 1183 3438
rect 1239 3382 1307 3438
rect 1363 3382 1431 3438
rect 1487 3382 1555 3438
rect 1611 3382 1679 3438
rect 1735 3382 1803 3438
rect 1859 3382 1927 3438
rect 1983 3382 2051 3438
rect 2107 3382 2117 3438
rect 305 3314 2117 3382
rect 305 3258 315 3314
rect 371 3258 439 3314
rect 495 3258 563 3314
rect 619 3258 687 3314
rect 743 3258 811 3314
rect 867 3258 935 3314
rect 991 3258 1059 3314
rect 1115 3258 1183 3314
rect 1239 3258 1307 3314
rect 1363 3258 1431 3314
rect 1487 3258 1555 3314
rect 1611 3258 1679 3314
rect 1735 3258 1803 3314
rect 1859 3258 1927 3314
rect 1983 3258 2051 3314
rect 2107 3258 2117 3314
rect 305 3190 2117 3258
rect 305 3134 315 3190
rect 371 3134 439 3190
rect 495 3134 563 3190
rect 619 3134 687 3190
rect 743 3134 811 3190
rect 867 3134 935 3190
rect 991 3134 1059 3190
rect 1115 3134 1183 3190
rect 1239 3134 1307 3190
rect 1363 3134 1431 3190
rect 1487 3134 1555 3190
rect 1611 3134 1679 3190
rect 1735 3134 1803 3190
rect 1859 3134 1927 3190
rect 1983 3134 2051 3190
rect 2107 3134 2117 3190
rect 305 3066 2117 3134
rect 305 3010 315 3066
rect 371 3010 439 3066
rect 495 3010 563 3066
rect 619 3010 687 3066
rect 743 3010 811 3066
rect 867 3010 935 3066
rect 991 3010 1059 3066
rect 1115 3010 1183 3066
rect 1239 3010 1307 3066
rect 1363 3010 1431 3066
rect 1487 3010 1555 3066
rect 1611 3010 1679 3066
rect 1735 3010 1803 3066
rect 1859 3010 1927 3066
rect 1983 3010 2051 3066
rect 2107 3010 2117 3066
rect 305 2942 2117 3010
rect 305 2886 315 2942
rect 371 2886 439 2942
rect 495 2886 563 2942
rect 619 2886 687 2942
rect 743 2886 811 2942
rect 867 2886 935 2942
rect 991 2886 1059 2942
rect 1115 2886 1183 2942
rect 1239 2886 1307 2942
rect 1363 2886 1431 2942
rect 1487 2886 1555 2942
rect 1611 2886 1679 2942
rect 1735 2886 1803 2942
rect 1859 2886 1927 2942
rect 1983 2886 2051 2942
rect 2107 2886 2117 2942
rect 305 2818 2117 2886
rect 305 2762 315 2818
rect 371 2762 439 2818
rect 495 2762 563 2818
rect 619 2762 687 2818
rect 743 2762 811 2818
rect 867 2762 935 2818
rect 991 2762 1059 2818
rect 1115 2762 1183 2818
rect 1239 2762 1307 2818
rect 1363 2762 1431 2818
rect 1487 2762 1555 2818
rect 1611 2762 1679 2818
rect 1735 2762 1803 2818
rect 1859 2762 1927 2818
rect 1983 2762 2051 2818
rect 2107 2762 2117 2818
rect 305 2694 2117 2762
rect 305 2638 315 2694
rect 371 2638 439 2694
rect 495 2638 563 2694
rect 619 2638 687 2694
rect 743 2638 811 2694
rect 867 2638 935 2694
rect 991 2638 1059 2694
rect 1115 2638 1183 2694
rect 1239 2638 1307 2694
rect 1363 2638 1431 2694
rect 1487 2638 1555 2694
rect 1611 2638 1679 2694
rect 1735 2638 1803 2694
rect 1859 2638 1927 2694
rect 1983 2638 2051 2694
rect 2107 2638 2117 2694
rect 305 2570 2117 2638
rect 305 2514 315 2570
rect 371 2514 439 2570
rect 495 2514 563 2570
rect 619 2514 687 2570
rect 743 2514 811 2570
rect 867 2514 935 2570
rect 991 2514 1059 2570
rect 1115 2514 1183 2570
rect 1239 2514 1307 2570
rect 1363 2514 1431 2570
rect 1487 2514 1555 2570
rect 1611 2514 1679 2570
rect 1735 2514 1803 2570
rect 1859 2514 1927 2570
rect 1983 2514 2051 2570
rect 2107 2514 2117 2570
rect 305 2446 2117 2514
rect 305 2390 315 2446
rect 371 2390 439 2446
rect 495 2390 563 2446
rect 619 2390 687 2446
rect 743 2390 811 2446
rect 867 2390 935 2446
rect 991 2390 1059 2446
rect 1115 2390 1183 2446
rect 1239 2390 1307 2446
rect 1363 2390 1431 2446
rect 1487 2390 1555 2446
rect 1611 2390 1679 2446
rect 1735 2390 1803 2446
rect 1859 2390 1927 2446
rect 1983 2390 2051 2446
rect 2107 2390 2117 2446
rect 305 2322 2117 2390
rect 305 2266 315 2322
rect 371 2266 439 2322
rect 495 2266 563 2322
rect 619 2266 687 2322
rect 743 2266 811 2322
rect 867 2266 935 2322
rect 991 2266 1059 2322
rect 1115 2266 1183 2322
rect 1239 2266 1307 2322
rect 1363 2266 1431 2322
rect 1487 2266 1555 2322
rect 1611 2266 1679 2322
rect 1735 2266 1803 2322
rect 1859 2266 1927 2322
rect 1983 2266 2051 2322
rect 2107 2266 2117 2322
rect 305 2198 2117 2266
rect 305 2142 315 2198
rect 371 2142 439 2198
rect 495 2142 563 2198
rect 619 2142 687 2198
rect 743 2142 811 2198
rect 867 2142 935 2198
rect 991 2142 1059 2198
rect 1115 2142 1183 2198
rect 1239 2142 1307 2198
rect 1363 2142 1431 2198
rect 1487 2142 1555 2198
rect 1611 2142 1679 2198
rect 1735 2142 1803 2198
rect 1859 2142 1927 2198
rect 1983 2142 2051 2198
rect 2107 2142 2117 2198
rect 305 2074 2117 2142
rect 305 2018 315 2074
rect 371 2018 439 2074
rect 495 2018 563 2074
rect 619 2018 687 2074
rect 743 2018 811 2074
rect 867 2018 935 2074
rect 991 2018 1059 2074
rect 1115 2018 1183 2074
rect 1239 2018 1307 2074
rect 1363 2018 1431 2074
rect 1487 2018 1555 2074
rect 1611 2018 1679 2074
rect 1735 2018 1803 2074
rect 1859 2018 1927 2074
rect 1983 2018 2051 2074
rect 2107 2018 2117 2074
rect 305 1950 2117 2018
rect 305 1894 315 1950
rect 371 1894 439 1950
rect 495 1894 563 1950
rect 619 1894 687 1950
rect 743 1894 811 1950
rect 867 1894 935 1950
rect 991 1894 1059 1950
rect 1115 1894 1183 1950
rect 1239 1894 1307 1950
rect 1363 1894 1431 1950
rect 1487 1894 1555 1950
rect 1611 1894 1679 1950
rect 1735 1894 1803 1950
rect 1859 1894 1927 1950
rect 1983 1894 2051 1950
rect 2107 1894 2117 1950
rect 305 1826 2117 1894
rect 305 1770 315 1826
rect 371 1770 439 1826
rect 495 1770 563 1826
rect 619 1770 687 1826
rect 743 1770 811 1826
rect 867 1770 935 1826
rect 991 1770 1059 1826
rect 1115 1770 1183 1826
rect 1239 1770 1307 1826
rect 1363 1770 1431 1826
rect 1487 1770 1555 1826
rect 1611 1770 1679 1826
rect 1735 1770 1803 1826
rect 1859 1770 1927 1826
rect 1983 1770 2051 1826
rect 2107 1770 2117 1826
rect 305 1702 2117 1770
rect 305 1646 315 1702
rect 371 1646 439 1702
rect 495 1646 563 1702
rect 619 1646 687 1702
rect 743 1646 811 1702
rect 867 1646 935 1702
rect 991 1646 1059 1702
rect 1115 1646 1183 1702
rect 1239 1646 1307 1702
rect 1363 1646 1431 1702
rect 1487 1646 1555 1702
rect 1611 1646 1679 1702
rect 1735 1646 1803 1702
rect 1859 1646 1927 1702
rect 1983 1646 2051 1702
rect 2107 1646 2117 1702
rect 305 1636 2117 1646
rect 2798 4554 4734 4564
rect 2798 4498 2808 4554
rect 2864 4498 2932 4554
rect 2988 4498 3056 4554
rect 3112 4498 3180 4554
rect 3236 4498 3304 4554
rect 3360 4498 3428 4554
rect 3484 4498 3552 4554
rect 3608 4498 3676 4554
rect 3732 4498 3800 4554
rect 3856 4498 3924 4554
rect 3980 4498 4048 4554
rect 4104 4498 4172 4554
rect 4228 4498 4296 4554
rect 4352 4498 4420 4554
rect 4476 4498 4544 4554
rect 4600 4498 4668 4554
rect 4724 4498 4734 4554
rect 2798 4430 4734 4498
rect 2798 4374 2808 4430
rect 2864 4374 2932 4430
rect 2988 4374 3056 4430
rect 3112 4374 3180 4430
rect 3236 4374 3304 4430
rect 3360 4374 3428 4430
rect 3484 4374 3552 4430
rect 3608 4374 3676 4430
rect 3732 4374 3800 4430
rect 3856 4374 3924 4430
rect 3980 4374 4048 4430
rect 4104 4374 4172 4430
rect 4228 4374 4296 4430
rect 4352 4374 4420 4430
rect 4476 4374 4544 4430
rect 4600 4374 4668 4430
rect 4724 4374 4734 4430
rect 2798 4306 4734 4374
rect 2798 4250 2808 4306
rect 2864 4250 2932 4306
rect 2988 4250 3056 4306
rect 3112 4250 3180 4306
rect 3236 4250 3304 4306
rect 3360 4250 3428 4306
rect 3484 4250 3552 4306
rect 3608 4250 3676 4306
rect 3732 4250 3800 4306
rect 3856 4250 3924 4306
rect 3980 4250 4048 4306
rect 4104 4250 4172 4306
rect 4228 4250 4296 4306
rect 4352 4250 4420 4306
rect 4476 4250 4544 4306
rect 4600 4250 4668 4306
rect 4724 4250 4734 4306
rect 2798 4182 4734 4250
rect 2798 4126 2808 4182
rect 2864 4126 2932 4182
rect 2988 4126 3056 4182
rect 3112 4126 3180 4182
rect 3236 4126 3304 4182
rect 3360 4126 3428 4182
rect 3484 4126 3552 4182
rect 3608 4126 3676 4182
rect 3732 4126 3800 4182
rect 3856 4126 3924 4182
rect 3980 4126 4048 4182
rect 4104 4126 4172 4182
rect 4228 4126 4296 4182
rect 4352 4126 4420 4182
rect 4476 4126 4544 4182
rect 4600 4126 4668 4182
rect 4724 4126 4734 4182
rect 2798 4058 4734 4126
rect 2798 4002 2808 4058
rect 2864 4002 2932 4058
rect 2988 4002 3056 4058
rect 3112 4002 3180 4058
rect 3236 4002 3304 4058
rect 3360 4002 3428 4058
rect 3484 4002 3552 4058
rect 3608 4002 3676 4058
rect 3732 4002 3800 4058
rect 3856 4002 3924 4058
rect 3980 4002 4048 4058
rect 4104 4002 4172 4058
rect 4228 4002 4296 4058
rect 4352 4002 4420 4058
rect 4476 4002 4544 4058
rect 4600 4002 4668 4058
rect 4724 4002 4734 4058
rect 2798 3934 4734 4002
rect 2798 3878 2808 3934
rect 2864 3878 2932 3934
rect 2988 3878 3056 3934
rect 3112 3878 3180 3934
rect 3236 3878 3304 3934
rect 3360 3878 3428 3934
rect 3484 3878 3552 3934
rect 3608 3878 3676 3934
rect 3732 3878 3800 3934
rect 3856 3878 3924 3934
rect 3980 3878 4048 3934
rect 4104 3878 4172 3934
rect 4228 3878 4296 3934
rect 4352 3878 4420 3934
rect 4476 3878 4544 3934
rect 4600 3878 4668 3934
rect 4724 3878 4734 3934
rect 2798 3810 4734 3878
rect 2798 3754 2808 3810
rect 2864 3754 2932 3810
rect 2988 3754 3056 3810
rect 3112 3754 3180 3810
rect 3236 3754 3304 3810
rect 3360 3754 3428 3810
rect 3484 3754 3552 3810
rect 3608 3754 3676 3810
rect 3732 3754 3800 3810
rect 3856 3754 3924 3810
rect 3980 3754 4048 3810
rect 4104 3754 4172 3810
rect 4228 3754 4296 3810
rect 4352 3754 4420 3810
rect 4476 3754 4544 3810
rect 4600 3754 4668 3810
rect 4724 3754 4734 3810
rect 2798 3686 4734 3754
rect 2798 3630 2808 3686
rect 2864 3630 2932 3686
rect 2988 3630 3056 3686
rect 3112 3630 3180 3686
rect 3236 3630 3304 3686
rect 3360 3630 3428 3686
rect 3484 3630 3552 3686
rect 3608 3630 3676 3686
rect 3732 3630 3800 3686
rect 3856 3630 3924 3686
rect 3980 3630 4048 3686
rect 4104 3630 4172 3686
rect 4228 3630 4296 3686
rect 4352 3630 4420 3686
rect 4476 3630 4544 3686
rect 4600 3630 4668 3686
rect 4724 3630 4734 3686
rect 2798 3562 4734 3630
rect 2798 3506 2808 3562
rect 2864 3506 2932 3562
rect 2988 3506 3056 3562
rect 3112 3506 3180 3562
rect 3236 3506 3304 3562
rect 3360 3506 3428 3562
rect 3484 3506 3552 3562
rect 3608 3506 3676 3562
rect 3732 3506 3800 3562
rect 3856 3506 3924 3562
rect 3980 3506 4048 3562
rect 4104 3506 4172 3562
rect 4228 3506 4296 3562
rect 4352 3506 4420 3562
rect 4476 3506 4544 3562
rect 4600 3506 4668 3562
rect 4724 3506 4734 3562
rect 2798 3438 4734 3506
rect 2798 3382 2808 3438
rect 2864 3382 2932 3438
rect 2988 3382 3056 3438
rect 3112 3382 3180 3438
rect 3236 3382 3304 3438
rect 3360 3382 3428 3438
rect 3484 3382 3552 3438
rect 3608 3382 3676 3438
rect 3732 3382 3800 3438
rect 3856 3382 3924 3438
rect 3980 3382 4048 3438
rect 4104 3382 4172 3438
rect 4228 3382 4296 3438
rect 4352 3382 4420 3438
rect 4476 3382 4544 3438
rect 4600 3382 4668 3438
rect 4724 3382 4734 3438
rect 2798 3314 4734 3382
rect 2798 3258 2808 3314
rect 2864 3258 2932 3314
rect 2988 3258 3056 3314
rect 3112 3258 3180 3314
rect 3236 3258 3304 3314
rect 3360 3258 3428 3314
rect 3484 3258 3552 3314
rect 3608 3258 3676 3314
rect 3732 3258 3800 3314
rect 3856 3258 3924 3314
rect 3980 3258 4048 3314
rect 4104 3258 4172 3314
rect 4228 3258 4296 3314
rect 4352 3258 4420 3314
rect 4476 3258 4544 3314
rect 4600 3258 4668 3314
rect 4724 3258 4734 3314
rect 2798 3190 4734 3258
rect 2798 3134 2808 3190
rect 2864 3134 2932 3190
rect 2988 3134 3056 3190
rect 3112 3134 3180 3190
rect 3236 3134 3304 3190
rect 3360 3134 3428 3190
rect 3484 3134 3552 3190
rect 3608 3134 3676 3190
rect 3732 3134 3800 3190
rect 3856 3134 3924 3190
rect 3980 3134 4048 3190
rect 4104 3134 4172 3190
rect 4228 3134 4296 3190
rect 4352 3134 4420 3190
rect 4476 3134 4544 3190
rect 4600 3134 4668 3190
rect 4724 3134 4734 3190
rect 2798 3066 4734 3134
rect 2798 3010 2808 3066
rect 2864 3010 2932 3066
rect 2988 3010 3056 3066
rect 3112 3010 3180 3066
rect 3236 3010 3304 3066
rect 3360 3010 3428 3066
rect 3484 3010 3552 3066
rect 3608 3010 3676 3066
rect 3732 3010 3800 3066
rect 3856 3010 3924 3066
rect 3980 3010 4048 3066
rect 4104 3010 4172 3066
rect 4228 3010 4296 3066
rect 4352 3010 4420 3066
rect 4476 3010 4544 3066
rect 4600 3010 4668 3066
rect 4724 3010 4734 3066
rect 2798 2942 4734 3010
rect 2798 2886 2808 2942
rect 2864 2886 2932 2942
rect 2988 2886 3056 2942
rect 3112 2886 3180 2942
rect 3236 2886 3304 2942
rect 3360 2886 3428 2942
rect 3484 2886 3552 2942
rect 3608 2886 3676 2942
rect 3732 2886 3800 2942
rect 3856 2886 3924 2942
rect 3980 2886 4048 2942
rect 4104 2886 4172 2942
rect 4228 2886 4296 2942
rect 4352 2886 4420 2942
rect 4476 2886 4544 2942
rect 4600 2886 4668 2942
rect 4724 2886 4734 2942
rect 2798 2818 4734 2886
rect 2798 2762 2808 2818
rect 2864 2762 2932 2818
rect 2988 2762 3056 2818
rect 3112 2762 3180 2818
rect 3236 2762 3304 2818
rect 3360 2762 3428 2818
rect 3484 2762 3552 2818
rect 3608 2762 3676 2818
rect 3732 2762 3800 2818
rect 3856 2762 3924 2818
rect 3980 2762 4048 2818
rect 4104 2762 4172 2818
rect 4228 2762 4296 2818
rect 4352 2762 4420 2818
rect 4476 2762 4544 2818
rect 4600 2762 4668 2818
rect 4724 2762 4734 2818
rect 2798 2694 4734 2762
rect 2798 2638 2808 2694
rect 2864 2638 2932 2694
rect 2988 2638 3056 2694
rect 3112 2638 3180 2694
rect 3236 2638 3304 2694
rect 3360 2638 3428 2694
rect 3484 2638 3552 2694
rect 3608 2638 3676 2694
rect 3732 2638 3800 2694
rect 3856 2638 3924 2694
rect 3980 2638 4048 2694
rect 4104 2638 4172 2694
rect 4228 2638 4296 2694
rect 4352 2638 4420 2694
rect 4476 2638 4544 2694
rect 4600 2638 4668 2694
rect 4724 2638 4734 2694
rect 2798 2570 4734 2638
rect 2798 2514 2808 2570
rect 2864 2514 2932 2570
rect 2988 2514 3056 2570
rect 3112 2514 3180 2570
rect 3236 2514 3304 2570
rect 3360 2514 3428 2570
rect 3484 2514 3552 2570
rect 3608 2514 3676 2570
rect 3732 2514 3800 2570
rect 3856 2514 3924 2570
rect 3980 2514 4048 2570
rect 4104 2514 4172 2570
rect 4228 2514 4296 2570
rect 4352 2514 4420 2570
rect 4476 2514 4544 2570
rect 4600 2514 4668 2570
rect 4724 2514 4734 2570
rect 2798 2446 4734 2514
rect 2798 2390 2808 2446
rect 2864 2390 2932 2446
rect 2988 2390 3056 2446
rect 3112 2390 3180 2446
rect 3236 2390 3304 2446
rect 3360 2390 3428 2446
rect 3484 2390 3552 2446
rect 3608 2390 3676 2446
rect 3732 2390 3800 2446
rect 3856 2390 3924 2446
rect 3980 2390 4048 2446
rect 4104 2390 4172 2446
rect 4228 2390 4296 2446
rect 4352 2390 4420 2446
rect 4476 2390 4544 2446
rect 4600 2390 4668 2446
rect 4724 2390 4734 2446
rect 2798 2322 4734 2390
rect 2798 2266 2808 2322
rect 2864 2266 2932 2322
rect 2988 2266 3056 2322
rect 3112 2266 3180 2322
rect 3236 2266 3304 2322
rect 3360 2266 3428 2322
rect 3484 2266 3552 2322
rect 3608 2266 3676 2322
rect 3732 2266 3800 2322
rect 3856 2266 3924 2322
rect 3980 2266 4048 2322
rect 4104 2266 4172 2322
rect 4228 2266 4296 2322
rect 4352 2266 4420 2322
rect 4476 2266 4544 2322
rect 4600 2266 4668 2322
rect 4724 2266 4734 2322
rect 2798 2198 4734 2266
rect 2798 2142 2808 2198
rect 2864 2142 2932 2198
rect 2988 2142 3056 2198
rect 3112 2142 3180 2198
rect 3236 2142 3304 2198
rect 3360 2142 3428 2198
rect 3484 2142 3552 2198
rect 3608 2142 3676 2198
rect 3732 2142 3800 2198
rect 3856 2142 3924 2198
rect 3980 2142 4048 2198
rect 4104 2142 4172 2198
rect 4228 2142 4296 2198
rect 4352 2142 4420 2198
rect 4476 2142 4544 2198
rect 4600 2142 4668 2198
rect 4724 2142 4734 2198
rect 2798 2074 4734 2142
rect 2798 2018 2808 2074
rect 2864 2018 2932 2074
rect 2988 2018 3056 2074
rect 3112 2018 3180 2074
rect 3236 2018 3304 2074
rect 3360 2018 3428 2074
rect 3484 2018 3552 2074
rect 3608 2018 3676 2074
rect 3732 2018 3800 2074
rect 3856 2018 3924 2074
rect 3980 2018 4048 2074
rect 4104 2018 4172 2074
rect 4228 2018 4296 2074
rect 4352 2018 4420 2074
rect 4476 2018 4544 2074
rect 4600 2018 4668 2074
rect 4724 2018 4734 2074
rect 2798 1950 4734 2018
rect 2798 1894 2808 1950
rect 2864 1894 2932 1950
rect 2988 1894 3056 1950
rect 3112 1894 3180 1950
rect 3236 1894 3304 1950
rect 3360 1894 3428 1950
rect 3484 1894 3552 1950
rect 3608 1894 3676 1950
rect 3732 1894 3800 1950
rect 3856 1894 3924 1950
rect 3980 1894 4048 1950
rect 4104 1894 4172 1950
rect 4228 1894 4296 1950
rect 4352 1894 4420 1950
rect 4476 1894 4544 1950
rect 4600 1894 4668 1950
rect 4724 1894 4734 1950
rect 2798 1826 4734 1894
rect 2798 1770 2808 1826
rect 2864 1770 2932 1826
rect 2988 1770 3056 1826
rect 3112 1770 3180 1826
rect 3236 1770 3304 1826
rect 3360 1770 3428 1826
rect 3484 1770 3552 1826
rect 3608 1770 3676 1826
rect 3732 1770 3800 1826
rect 3856 1770 3924 1826
rect 3980 1770 4048 1826
rect 4104 1770 4172 1826
rect 4228 1770 4296 1826
rect 4352 1770 4420 1826
rect 4476 1770 4544 1826
rect 4600 1770 4668 1826
rect 4724 1770 4734 1826
rect 2798 1702 4734 1770
rect 2798 1646 2808 1702
rect 2864 1646 2932 1702
rect 2988 1646 3056 1702
rect 3112 1646 3180 1702
rect 3236 1646 3304 1702
rect 3360 1646 3428 1702
rect 3484 1646 3552 1702
rect 3608 1646 3676 1702
rect 3732 1646 3800 1702
rect 3856 1646 3924 1702
rect 3980 1646 4048 1702
rect 4104 1646 4172 1702
rect 4228 1646 4296 1702
rect 4352 1646 4420 1702
rect 4476 1646 4544 1702
rect 4600 1646 4668 1702
rect 4724 1646 4734 1702
rect 2798 1636 4734 1646
rect 5168 4554 7104 4564
rect 5168 4498 5178 4554
rect 5234 4498 5302 4554
rect 5358 4498 5426 4554
rect 5482 4498 5550 4554
rect 5606 4498 5674 4554
rect 5730 4498 5798 4554
rect 5854 4498 5922 4554
rect 5978 4498 6046 4554
rect 6102 4498 6170 4554
rect 6226 4498 6294 4554
rect 6350 4498 6418 4554
rect 6474 4498 6542 4554
rect 6598 4498 6666 4554
rect 6722 4498 6790 4554
rect 6846 4498 6914 4554
rect 6970 4498 7038 4554
rect 7094 4498 7104 4554
rect 5168 4430 7104 4498
rect 5168 4374 5178 4430
rect 5234 4374 5302 4430
rect 5358 4374 5426 4430
rect 5482 4374 5550 4430
rect 5606 4374 5674 4430
rect 5730 4374 5798 4430
rect 5854 4374 5922 4430
rect 5978 4374 6046 4430
rect 6102 4374 6170 4430
rect 6226 4374 6294 4430
rect 6350 4374 6418 4430
rect 6474 4374 6542 4430
rect 6598 4374 6666 4430
rect 6722 4374 6790 4430
rect 6846 4374 6914 4430
rect 6970 4374 7038 4430
rect 7094 4374 7104 4430
rect 5168 4306 7104 4374
rect 5168 4250 5178 4306
rect 5234 4250 5302 4306
rect 5358 4250 5426 4306
rect 5482 4250 5550 4306
rect 5606 4250 5674 4306
rect 5730 4250 5798 4306
rect 5854 4250 5922 4306
rect 5978 4250 6046 4306
rect 6102 4250 6170 4306
rect 6226 4250 6294 4306
rect 6350 4250 6418 4306
rect 6474 4250 6542 4306
rect 6598 4250 6666 4306
rect 6722 4250 6790 4306
rect 6846 4250 6914 4306
rect 6970 4250 7038 4306
rect 7094 4250 7104 4306
rect 5168 4182 7104 4250
rect 5168 4126 5178 4182
rect 5234 4126 5302 4182
rect 5358 4126 5426 4182
rect 5482 4126 5550 4182
rect 5606 4126 5674 4182
rect 5730 4126 5798 4182
rect 5854 4126 5922 4182
rect 5978 4126 6046 4182
rect 6102 4126 6170 4182
rect 6226 4126 6294 4182
rect 6350 4126 6418 4182
rect 6474 4126 6542 4182
rect 6598 4126 6666 4182
rect 6722 4126 6790 4182
rect 6846 4126 6914 4182
rect 6970 4126 7038 4182
rect 7094 4126 7104 4182
rect 5168 4058 7104 4126
rect 5168 4002 5178 4058
rect 5234 4002 5302 4058
rect 5358 4002 5426 4058
rect 5482 4002 5550 4058
rect 5606 4002 5674 4058
rect 5730 4002 5798 4058
rect 5854 4002 5922 4058
rect 5978 4002 6046 4058
rect 6102 4002 6170 4058
rect 6226 4002 6294 4058
rect 6350 4002 6418 4058
rect 6474 4002 6542 4058
rect 6598 4002 6666 4058
rect 6722 4002 6790 4058
rect 6846 4002 6914 4058
rect 6970 4002 7038 4058
rect 7094 4002 7104 4058
rect 5168 3934 7104 4002
rect 5168 3878 5178 3934
rect 5234 3878 5302 3934
rect 5358 3878 5426 3934
rect 5482 3878 5550 3934
rect 5606 3878 5674 3934
rect 5730 3878 5798 3934
rect 5854 3878 5922 3934
rect 5978 3878 6046 3934
rect 6102 3878 6170 3934
rect 6226 3878 6294 3934
rect 6350 3878 6418 3934
rect 6474 3878 6542 3934
rect 6598 3878 6666 3934
rect 6722 3878 6790 3934
rect 6846 3878 6914 3934
rect 6970 3878 7038 3934
rect 7094 3878 7104 3934
rect 5168 3810 7104 3878
rect 5168 3754 5178 3810
rect 5234 3754 5302 3810
rect 5358 3754 5426 3810
rect 5482 3754 5550 3810
rect 5606 3754 5674 3810
rect 5730 3754 5798 3810
rect 5854 3754 5922 3810
rect 5978 3754 6046 3810
rect 6102 3754 6170 3810
rect 6226 3754 6294 3810
rect 6350 3754 6418 3810
rect 6474 3754 6542 3810
rect 6598 3754 6666 3810
rect 6722 3754 6790 3810
rect 6846 3754 6914 3810
rect 6970 3754 7038 3810
rect 7094 3754 7104 3810
rect 5168 3686 7104 3754
rect 5168 3630 5178 3686
rect 5234 3630 5302 3686
rect 5358 3630 5426 3686
rect 5482 3630 5550 3686
rect 5606 3630 5674 3686
rect 5730 3630 5798 3686
rect 5854 3630 5922 3686
rect 5978 3630 6046 3686
rect 6102 3630 6170 3686
rect 6226 3630 6294 3686
rect 6350 3630 6418 3686
rect 6474 3630 6542 3686
rect 6598 3630 6666 3686
rect 6722 3630 6790 3686
rect 6846 3630 6914 3686
rect 6970 3630 7038 3686
rect 7094 3630 7104 3686
rect 5168 3562 7104 3630
rect 5168 3506 5178 3562
rect 5234 3506 5302 3562
rect 5358 3506 5426 3562
rect 5482 3506 5550 3562
rect 5606 3506 5674 3562
rect 5730 3506 5798 3562
rect 5854 3506 5922 3562
rect 5978 3506 6046 3562
rect 6102 3506 6170 3562
rect 6226 3506 6294 3562
rect 6350 3506 6418 3562
rect 6474 3506 6542 3562
rect 6598 3506 6666 3562
rect 6722 3506 6790 3562
rect 6846 3506 6914 3562
rect 6970 3506 7038 3562
rect 7094 3506 7104 3562
rect 5168 3438 7104 3506
rect 5168 3382 5178 3438
rect 5234 3382 5302 3438
rect 5358 3382 5426 3438
rect 5482 3382 5550 3438
rect 5606 3382 5674 3438
rect 5730 3382 5798 3438
rect 5854 3382 5922 3438
rect 5978 3382 6046 3438
rect 6102 3382 6170 3438
rect 6226 3382 6294 3438
rect 6350 3382 6418 3438
rect 6474 3382 6542 3438
rect 6598 3382 6666 3438
rect 6722 3382 6790 3438
rect 6846 3382 6914 3438
rect 6970 3382 7038 3438
rect 7094 3382 7104 3438
rect 5168 3314 7104 3382
rect 5168 3258 5178 3314
rect 5234 3258 5302 3314
rect 5358 3258 5426 3314
rect 5482 3258 5550 3314
rect 5606 3258 5674 3314
rect 5730 3258 5798 3314
rect 5854 3258 5922 3314
rect 5978 3258 6046 3314
rect 6102 3258 6170 3314
rect 6226 3258 6294 3314
rect 6350 3258 6418 3314
rect 6474 3258 6542 3314
rect 6598 3258 6666 3314
rect 6722 3258 6790 3314
rect 6846 3258 6914 3314
rect 6970 3258 7038 3314
rect 7094 3258 7104 3314
rect 5168 3190 7104 3258
rect 5168 3134 5178 3190
rect 5234 3134 5302 3190
rect 5358 3134 5426 3190
rect 5482 3134 5550 3190
rect 5606 3134 5674 3190
rect 5730 3134 5798 3190
rect 5854 3134 5922 3190
rect 5978 3134 6046 3190
rect 6102 3134 6170 3190
rect 6226 3134 6294 3190
rect 6350 3134 6418 3190
rect 6474 3134 6542 3190
rect 6598 3134 6666 3190
rect 6722 3134 6790 3190
rect 6846 3134 6914 3190
rect 6970 3134 7038 3190
rect 7094 3134 7104 3190
rect 5168 3066 7104 3134
rect 5168 3010 5178 3066
rect 5234 3010 5302 3066
rect 5358 3010 5426 3066
rect 5482 3010 5550 3066
rect 5606 3010 5674 3066
rect 5730 3010 5798 3066
rect 5854 3010 5922 3066
rect 5978 3010 6046 3066
rect 6102 3010 6170 3066
rect 6226 3010 6294 3066
rect 6350 3010 6418 3066
rect 6474 3010 6542 3066
rect 6598 3010 6666 3066
rect 6722 3010 6790 3066
rect 6846 3010 6914 3066
rect 6970 3010 7038 3066
rect 7094 3010 7104 3066
rect 5168 2942 7104 3010
rect 5168 2886 5178 2942
rect 5234 2886 5302 2942
rect 5358 2886 5426 2942
rect 5482 2886 5550 2942
rect 5606 2886 5674 2942
rect 5730 2886 5798 2942
rect 5854 2886 5922 2942
rect 5978 2886 6046 2942
rect 6102 2886 6170 2942
rect 6226 2886 6294 2942
rect 6350 2886 6418 2942
rect 6474 2886 6542 2942
rect 6598 2886 6666 2942
rect 6722 2886 6790 2942
rect 6846 2886 6914 2942
rect 6970 2886 7038 2942
rect 7094 2886 7104 2942
rect 5168 2818 7104 2886
rect 5168 2762 5178 2818
rect 5234 2762 5302 2818
rect 5358 2762 5426 2818
rect 5482 2762 5550 2818
rect 5606 2762 5674 2818
rect 5730 2762 5798 2818
rect 5854 2762 5922 2818
rect 5978 2762 6046 2818
rect 6102 2762 6170 2818
rect 6226 2762 6294 2818
rect 6350 2762 6418 2818
rect 6474 2762 6542 2818
rect 6598 2762 6666 2818
rect 6722 2762 6790 2818
rect 6846 2762 6914 2818
rect 6970 2762 7038 2818
rect 7094 2762 7104 2818
rect 5168 2694 7104 2762
rect 5168 2638 5178 2694
rect 5234 2638 5302 2694
rect 5358 2638 5426 2694
rect 5482 2638 5550 2694
rect 5606 2638 5674 2694
rect 5730 2638 5798 2694
rect 5854 2638 5922 2694
rect 5978 2638 6046 2694
rect 6102 2638 6170 2694
rect 6226 2638 6294 2694
rect 6350 2638 6418 2694
rect 6474 2638 6542 2694
rect 6598 2638 6666 2694
rect 6722 2638 6790 2694
rect 6846 2638 6914 2694
rect 6970 2638 7038 2694
rect 7094 2638 7104 2694
rect 5168 2570 7104 2638
rect 5168 2514 5178 2570
rect 5234 2514 5302 2570
rect 5358 2514 5426 2570
rect 5482 2514 5550 2570
rect 5606 2514 5674 2570
rect 5730 2514 5798 2570
rect 5854 2514 5922 2570
rect 5978 2514 6046 2570
rect 6102 2514 6170 2570
rect 6226 2514 6294 2570
rect 6350 2514 6418 2570
rect 6474 2514 6542 2570
rect 6598 2514 6666 2570
rect 6722 2514 6790 2570
rect 6846 2514 6914 2570
rect 6970 2514 7038 2570
rect 7094 2514 7104 2570
rect 5168 2446 7104 2514
rect 5168 2390 5178 2446
rect 5234 2390 5302 2446
rect 5358 2390 5426 2446
rect 5482 2390 5550 2446
rect 5606 2390 5674 2446
rect 5730 2390 5798 2446
rect 5854 2390 5922 2446
rect 5978 2390 6046 2446
rect 6102 2390 6170 2446
rect 6226 2390 6294 2446
rect 6350 2390 6418 2446
rect 6474 2390 6542 2446
rect 6598 2390 6666 2446
rect 6722 2390 6790 2446
rect 6846 2390 6914 2446
rect 6970 2390 7038 2446
rect 7094 2390 7104 2446
rect 5168 2322 7104 2390
rect 5168 2266 5178 2322
rect 5234 2266 5302 2322
rect 5358 2266 5426 2322
rect 5482 2266 5550 2322
rect 5606 2266 5674 2322
rect 5730 2266 5798 2322
rect 5854 2266 5922 2322
rect 5978 2266 6046 2322
rect 6102 2266 6170 2322
rect 6226 2266 6294 2322
rect 6350 2266 6418 2322
rect 6474 2266 6542 2322
rect 6598 2266 6666 2322
rect 6722 2266 6790 2322
rect 6846 2266 6914 2322
rect 6970 2266 7038 2322
rect 7094 2266 7104 2322
rect 5168 2198 7104 2266
rect 5168 2142 5178 2198
rect 5234 2142 5302 2198
rect 5358 2142 5426 2198
rect 5482 2142 5550 2198
rect 5606 2142 5674 2198
rect 5730 2142 5798 2198
rect 5854 2142 5922 2198
rect 5978 2142 6046 2198
rect 6102 2142 6170 2198
rect 6226 2142 6294 2198
rect 6350 2142 6418 2198
rect 6474 2142 6542 2198
rect 6598 2142 6666 2198
rect 6722 2142 6790 2198
rect 6846 2142 6914 2198
rect 6970 2142 7038 2198
rect 7094 2142 7104 2198
rect 5168 2074 7104 2142
rect 5168 2018 5178 2074
rect 5234 2018 5302 2074
rect 5358 2018 5426 2074
rect 5482 2018 5550 2074
rect 5606 2018 5674 2074
rect 5730 2018 5798 2074
rect 5854 2018 5922 2074
rect 5978 2018 6046 2074
rect 6102 2018 6170 2074
rect 6226 2018 6294 2074
rect 6350 2018 6418 2074
rect 6474 2018 6542 2074
rect 6598 2018 6666 2074
rect 6722 2018 6790 2074
rect 6846 2018 6914 2074
rect 6970 2018 7038 2074
rect 7094 2018 7104 2074
rect 5168 1950 7104 2018
rect 5168 1894 5178 1950
rect 5234 1894 5302 1950
rect 5358 1894 5426 1950
rect 5482 1894 5550 1950
rect 5606 1894 5674 1950
rect 5730 1894 5798 1950
rect 5854 1894 5922 1950
rect 5978 1894 6046 1950
rect 6102 1894 6170 1950
rect 6226 1894 6294 1950
rect 6350 1894 6418 1950
rect 6474 1894 6542 1950
rect 6598 1894 6666 1950
rect 6722 1894 6790 1950
rect 6846 1894 6914 1950
rect 6970 1894 7038 1950
rect 7094 1894 7104 1950
rect 5168 1826 7104 1894
rect 5168 1770 5178 1826
rect 5234 1770 5302 1826
rect 5358 1770 5426 1826
rect 5482 1770 5550 1826
rect 5606 1770 5674 1826
rect 5730 1770 5798 1826
rect 5854 1770 5922 1826
rect 5978 1770 6046 1826
rect 6102 1770 6170 1826
rect 6226 1770 6294 1826
rect 6350 1770 6418 1826
rect 6474 1770 6542 1826
rect 6598 1770 6666 1826
rect 6722 1770 6790 1826
rect 6846 1770 6914 1826
rect 6970 1770 7038 1826
rect 7094 1770 7104 1826
rect 5168 1702 7104 1770
rect 5168 1646 5178 1702
rect 5234 1646 5302 1702
rect 5358 1646 5426 1702
rect 5482 1646 5550 1702
rect 5606 1646 5674 1702
rect 5730 1646 5798 1702
rect 5854 1646 5922 1702
rect 5978 1646 6046 1702
rect 6102 1646 6170 1702
rect 6226 1646 6294 1702
rect 6350 1646 6418 1702
rect 6474 1646 6542 1702
rect 6598 1646 6666 1702
rect 6722 1646 6790 1702
rect 6846 1646 6914 1702
rect 6970 1646 7038 1702
rect 7094 1646 7104 1702
rect 5168 1636 7104 1646
rect 7874 4554 9810 4564
rect 7874 4498 7884 4554
rect 7940 4498 8008 4554
rect 8064 4498 8132 4554
rect 8188 4498 8256 4554
rect 8312 4498 8380 4554
rect 8436 4498 8504 4554
rect 8560 4498 8628 4554
rect 8684 4498 8752 4554
rect 8808 4498 8876 4554
rect 8932 4498 9000 4554
rect 9056 4498 9124 4554
rect 9180 4498 9248 4554
rect 9304 4498 9372 4554
rect 9428 4498 9496 4554
rect 9552 4498 9620 4554
rect 9676 4498 9744 4554
rect 9800 4498 9810 4554
rect 7874 4430 9810 4498
rect 7874 4374 7884 4430
rect 7940 4374 8008 4430
rect 8064 4374 8132 4430
rect 8188 4374 8256 4430
rect 8312 4374 8380 4430
rect 8436 4374 8504 4430
rect 8560 4374 8628 4430
rect 8684 4374 8752 4430
rect 8808 4374 8876 4430
rect 8932 4374 9000 4430
rect 9056 4374 9124 4430
rect 9180 4374 9248 4430
rect 9304 4374 9372 4430
rect 9428 4374 9496 4430
rect 9552 4374 9620 4430
rect 9676 4374 9744 4430
rect 9800 4374 9810 4430
rect 7874 4306 9810 4374
rect 7874 4250 7884 4306
rect 7940 4250 8008 4306
rect 8064 4250 8132 4306
rect 8188 4250 8256 4306
rect 8312 4250 8380 4306
rect 8436 4250 8504 4306
rect 8560 4250 8628 4306
rect 8684 4250 8752 4306
rect 8808 4250 8876 4306
rect 8932 4250 9000 4306
rect 9056 4250 9124 4306
rect 9180 4250 9248 4306
rect 9304 4250 9372 4306
rect 9428 4250 9496 4306
rect 9552 4250 9620 4306
rect 9676 4250 9744 4306
rect 9800 4250 9810 4306
rect 7874 4182 9810 4250
rect 7874 4126 7884 4182
rect 7940 4126 8008 4182
rect 8064 4126 8132 4182
rect 8188 4126 8256 4182
rect 8312 4126 8380 4182
rect 8436 4126 8504 4182
rect 8560 4126 8628 4182
rect 8684 4126 8752 4182
rect 8808 4126 8876 4182
rect 8932 4126 9000 4182
rect 9056 4126 9124 4182
rect 9180 4126 9248 4182
rect 9304 4126 9372 4182
rect 9428 4126 9496 4182
rect 9552 4126 9620 4182
rect 9676 4126 9744 4182
rect 9800 4126 9810 4182
rect 7874 4058 9810 4126
rect 7874 4002 7884 4058
rect 7940 4002 8008 4058
rect 8064 4002 8132 4058
rect 8188 4002 8256 4058
rect 8312 4002 8380 4058
rect 8436 4002 8504 4058
rect 8560 4002 8628 4058
rect 8684 4002 8752 4058
rect 8808 4002 8876 4058
rect 8932 4002 9000 4058
rect 9056 4002 9124 4058
rect 9180 4002 9248 4058
rect 9304 4002 9372 4058
rect 9428 4002 9496 4058
rect 9552 4002 9620 4058
rect 9676 4002 9744 4058
rect 9800 4002 9810 4058
rect 7874 3934 9810 4002
rect 7874 3878 7884 3934
rect 7940 3878 8008 3934
rect 8064 3878 8132 3934
rect 8188 3878 8256 3934
rect 8312 3878 8380 3934
rect 8436 3878 8504 3934
rect 8560 3878 8628 3934
rect 8684 3878 8752 3934
rect 8808 3878 8876 3934
rect 8932 3878 9000 3934
rect 9056 3878 9124 3934
rect 9180 3878 9248 3934
rect 9304 3878 9372 3934
rect 9428 3878 9496 3934
rect 9552 3878 9620 3934
rect 9676 3878 9744 3934
rect 9800 3878 9810 3934
rect 7874 3810 9810 3878
rect 7874 3754 7884 3810
rect 7940 3754 8008 3810
rect 8064 3754 8132 3810
rect 8188 3754 8256 3810
rect 8312 3754 8380 3810
rect 8436 3754 8504 3810
rect 8560 3754 8628 3810
rect 8684 3754 8752 3810
rect 8808 3754 8876 3810
rect 8932 3754 9000 3810
rect 9056 3754 9124 3810
rect 9180 3754 9248 3810
rect 9304 3754 9372 3810
rect 9428 3754 9496 3810
rect 9552 3754 9620 3810
rect 9676 3754 9744 3810
rect 9800 3754 9810 3810
rect 7874 3686 9810 3754
rect 7874 3630 7884 3686
rect 7940 3630 8008 3686
rect 8064 3630 8132 3686
rect 8188 3630 8256 3686
rect 8312 3630 8380 3686
rect 8436 3630 8504 3686
rect 8560 3630 8628 3686
rect 8684 3630 8752 3686
rect 8808 3630 8876 3686
rect 8932 3630 9000 3686
rect 9056 3630 9124 3686
rect 9180 3630 9248 3686
rect 9304 3630 9372 3686
rect 9428 3630 9496 3686
rect 9552 3630 9620 3686
rect 9676 3630 9744 3686
rect 9800 3630 9810 3686
rect 7874 3562 9810 3630
rect 7874 3506 7884 3562
rect 7940 3506 8008 3562
rect 8064 3506 8132 3562
rect 8188 3506 8256 3562
rect 8312 3506 8380 3562
rect 8436 3506 8504 3562
rect 8560 3506 8628 3562
rect 8684 3506 8752 3562
rect 8808 3506 8876 3562
rect 8932 3506 9000 3562
rect 9056 3506 9124 3562
rect 9180 3506 9248 3562
rect 9304 3506 9372 3562
rect 9428 3506 9496 3562
rect 9552 3506 9620 3562
rect 9676 3506 9744 3562
rect 9800 3506 9810 3562
rect 7874 3438 9810 3506
rect 7874 3382 7884 3438
rect 7940 3382 8008 3438
rect 8064 3382 8132 3438
rect 8188 3382 8256 3438
rect 8312 3382 8380 3438
rect 8436 3382 8504 3438
rect 8560 3382 8628 3438
rect 8684 3382 8752 3438
rect 8808 3382 8876 3438
rect 8932 3382 9000 3438
rect 9056 3382 9124 3438
rect 9180 3382 9248 3438
rect 9304 3382 9372 3438
rect 9428 3382 9496 3438
rect 9552 3382 9620 3438
rect 9676 3382 9744 3438
rect 9800 3382 9810 3438
rect 7874 3314 9810 3382
rect 7874 3258 7884 3314
rect 7940 3258 8008 3314
rect 8064 3258 8132 3314
rect 8188 3258 8256 3314
rect 8312 3258 8380 3314
rect 8436 3258 8504 3314
rect 8560 3258 8628 3314
rect 8684 3258 8752 3314
rect 8808 3258 8876 3314
rect 8932 3258 9000 3314
rect 9056 3258 9124 3314
rect 9180 3258 9248 3314
rect 9304 3258 9372 3314
rect 9428 3258 9496 3314
rect 9552 3258 9620 3314
rect 9676 3258 9744 3314
rect 9800 3258 9810 3314
rect 7874 3190 9810 3258
rect 7874 3134 7884 3190
rect 7940 3134 8008 3190
rect 8064 3134 8132 3190
rect 8188 3134 8256 3190
rect 8312 3134 8380 3190
rect 8436 3134 8504 3190
rect 8560 3134 8628 3190
rect 8684 3134 8752 3190
rect 8808 3134 8876 3190
rect 8932 3134 9000 3190
rect 9056 3134 9124 3190
rect 9180 3134 9248 3190
rect 9304 3134 9372 3190
rect 9428 3134 9496 3190
rect 9552 3134 9620 3190
rect 9676 3134 9744 3190
rect 9800 3134 9810 3190
rect 7874 3066 9810 3134
rect 7874 3010 7884 3066
rect 7940 3010 8008 3066
rect 8064 3010 8132 3066
rect 8188 3010 8256 3066
rect 8312 3010 8380 3066
rect 8436 3010 8504 3066
rect 8560 3010 8628 3066
rect 8684 3010 8752 3066
rect 8808 3010 8876 3066
rect 8932 3010 9000 3066
rect 9056 3010 9124 3066
rect 9180 3010 9248 3066
rect 9304 3010 9372 3066
rect 9428 3010 9496 3066
rect 9552 3010 9620 3066
rect 9676 3010 9744 3066
rect 9800 3010 9810 3066
rect 7874 2942 9810 3010
rect 7874 2886 7884 2942
rect 7940 2886 8008 2942
rect 8064 2886 8132 2942
rect 8188 2886 8256 2942
rect 8312 2886 8380 2942
rect 8436 2886 8504 2942
rect 8560 2886 8628 2942
rect 8684 2886 8752 2942
rect 8808 2886 8876 2942
rect 8932 2886 9000 2942
rect 9056 2886 9124 2942
rect 9180 2886 9248 2942
rect 9304 2886 9372 2942
rect 9428 2886 9496 2942
rect 9552 2886 9620 2942
rect 9676 2886 9744 2942
rect 9800 2886 9810 2942
rect 7874 2818 9810 2886
rect 7874 2762 7884 2818
rect 7940 2762 8008 2818
rect 8064 2762 8132 2818
rect 8188 2762 8256 2818
rect 8312 2762 8380 2818
rect 8436 2762 8504 2818
rect 8560 2762 8628 2818
rect 8684 2762 8752 2818
rect 8808 2762 8876 2818
rect 8932 2762 9000 2818
rect 9056 2762 9124 2818
rect 9180 2762 9248 2818
rect 9304 2762 9372 2818
rect 9428 2762 9496 2818
rect 9552 2762 9620 2818
rect 9676 2762 9744 2818
rect 9800 2762 9810 2818
rect 7874 2694 9810 2762
rect 7874 2638 7884 2694
rect 7940 2638 8008 2694
rect 8064 2638 8132 2694
rect 8188 2638 8256 2694
rect 8312 2638 8380 2694
rect 8436 2638 8504 2694
rect 8560 2638 8628 2694
rect 8684 2638 8752 2694
rect 8808 2638 8876 2694
rect 8932 2638 9000 2694
rect 9056 2638 9124 2694
rect 9180 2638 9248 2694
rect 9304 2638 9372 2694
rect 9428 2638 9496 2694
rect 9552 2638 9620 2694
rect 9676 2638 9744 2694
rect 9800 2638 9810 2694
rect 7874 2570 9810 2638
rect 7874 2514 7884 2570
rect 7940 2514 8008 2570
rect 8064 2514 8132 2570
rect 8188 2514 8256 2570
rect 8312 2514 8380 2570
rect 8436 2514 8504 2570
rect 8560 2514 8628 2570
rect 8684 2514 8752 2570
rect 8808 2514 8876 2570
rect 8932 2514 9000 2570
rect 9056 2514 9124 2570
rect 9180 2514 9248 2570
rect 9304 2514 9372 2570
rect 9428 2514 9496 2570
rect 9552 2514 9620 2570
rect 9676 2514 9744 2570
rect 9800 2514 9810 2570
rect 7874 2446 9810 2514
rect 7874 2390 7884 2446
rect 7940 2390 8008 2446
rect 8064 2390 8132 2446
rect 8188 2390 8256 2446
rect 8312 2390 8380 2446
rect 8436 2390 8504 2446
rect 8560 2390 8628 2446
rect 8684 2390 8752 2446
rect 8808 2390 8876 2446
rect 8932 2390 9000 2446
rect 9056 2390 9124 2446
rect 9180 2390 9248 2446
rect 9304 2390 9372 2446
rect 9428 2390 9496 2446
rect 9552 2390 9620 2446
rect 9676 2390 9744 2446
rect 9800 2390 9810 2446
rect 7874 2322 9810 2390
rect 7874 2266 7884 2322
rect 7940 2266 8008 2322
rect 8064 2266 8132 2322
rect 8188 2266 8256 2322
rect 8312 2266 8380 2322
rect 8436 2266 8504 2322
rect 8560 2266 8628 2322
rect 8684 2266 8752 2322
rect 8808 2266 8876 2322
rect 8932 2266 9000 2322
rect 9056 2266 9124 2322
rect 9180 2266 9248 2322
rect 9304 2266 9372 2322
rect 9428 2266 9496 2322
rect 9552 2266 9620 2322
rect 9676 2266 9744 2322
rect 9800 2266 9810 2322
rect 7874 2198 9810 2266
rect 7874 2142 7884 2198
rect 7940 2142 8008 2198
rect 8064 2142 8132 2198
rect 8188 2142 8256 2198
rect 8312 2142 8380 2198
rect 8436 2142 8504 2198
rect 8560 2142 8628 2198
rect 8684 2142 8752 2198
rect 8808 2142 8876 2198
rect 8932 2142 9000 2198
rect 9056 2142 9124 2198
rect 9180 2142 9248 2198
rect 9304 2142 9372 2198
rect 9428 2142 9496 2198
rect 9552 2142 9620 2198
rect 9676 2142 9744 2198
rect 9800 2142 9810 2198
rect 7874 2074 9810 2142
rect 7874 2018 7884 2074
rect 7940 2018 8008 2074
rect 8064 2018 8132 2074
rect 8188 2018 8256 2074
rect 8312 2018 8380 2074
rect 8436 2018 8504 2074
rect 8560 2018 8628 2074
rect 8684 2018 8752 2074
rect 8808 2018 8876 2074
rect 8932 2018 9000 2074
rect 9056 2018 9124 2074
rect 9180 2018 9248 2074
rect 9304 2018 9372 2074
rect 9428 2018 9496 2074
rect 9552 2018 9620 2074
rect 9676 2018 9744 2074
rect 9800 2018 9810 2074
rect 7874 1950 9810 2018
rect 7874 1894 7884 1950
rect 7940 1894 8008 1950
rect 8064 1894 8132 1950
rect 8188 1894 8256 1950
rect 8312 1894 8380 1950
rect 8436 1894 8504 1950
rect 8560 1894 8628 1950
rect 8684 1894 8752 1950
rect 8808 1894 8876 1950
rect 8932 1894 9000 1950
rect 9056 1894 9124 1950
rect 9180 1894 9248 1950
rect 9304 1894 9372 1950
rect 9428 1894 9496 1950
rect 9552 1894 9620 1950
rect 9676 1894 9744 1950
rect 9800 1894 9810 1950
rect 7874 1826 9810 1894
rect 7874 1770 7884 1826
rect 7940 1770 8008 1826
rect 8064 1770 8132 1826
rect 8188 1770 8256 1826
rect 8312 1770 8380 1826
rect 8436 1770 8504 1826
rect 8560 1770 8628 1826
rect 8684 1770 8752 1826
rect 8808 1770 8876 1826
rect 8932 1770 9000 1826
rect 9056 1770 9124 1826
rect 9180 1770 9248 1826
rect 9304 1770 9372 1826
rect 9428 1770 9496 1826
rect 9552 1770 9620 1826
rect 9676 1770 9744 1826
rect 9800 1770 9810 1826
rect 7874 1702 9810 1770
rect 7874 1646 7884 1702
rect 7940 1646 8008 1702
rect 8064 1646 8132 1702
rect 8188 1646 8256 1702
rect 8312 1646 8380 1702
rect 8436 1646 8504 1702
rect 8560 1646 8628 1702
rect 8684 1646 8752 1702
rect 8808 1646 8876 1702
rect 8932 1646 9000 1702
rect 9056 1646 9124 1702
rect 9180 1646 9248 1702
rect 9304 1646 9372 1702
rect 9428 1646 9496 1702
rect 9552 1646 9620 1702
rect 9676 1646 9744 1702
rect 9800 1646 9810 1702
rect 7874 1636 9810 1646
rect 10244 4554 12180 4564
rect 10244 4498 10254 4554
rect 10310 4498 10378 4554
rect 10434 4498 10502 4554
rect 10558 4498 10626 4554
rect 10682 4498 10750 4554
rect 10806 4498 10874 4554
rect 10930 4498 10998 4554
rect 11054 4498 11122 4554
rect 11178 4498 11246 4554
rect 11302 4498 11370 4554
rect 11426 4498 11494 4554
rect 11550 4498 11618 4554
rect 11674 4498 11742 4554
rect 11798 4498 11866 4554
rect 11922 4498 11990 4554
rect 12046 4498 12114 4554
rect 12170 4498 12180 4554
rect 10244 4430 12180 4498
rect 10244 4374 10254 4430
rect 10310 4374 10378 4430
rect 10434 4374 10502 4430
rect 10558 4374 10626 4430
rect 10682 4374 10750 4430
rect 10806 4374 10874 4430
rect 10930 4374 10998 4430
rect 11054 4374 11122 4430
rect 11178 4374 11246 4430
rect 11302 4374 11370 4430
rect 11426 4374 11494 4430
rect 11550 4374 11618 4430
rect 11674 4374 11742 4430
rect 11798 4374 11866 4430
rect 11922 4374 11990 4430
rect 12046 4374 12114 4430
rect 12170 4374 12180 4430
rect 10244 4306 12180 4374
rect 10244 4250 10254 4306
rect 10310 4250 10378 4306
rect 10434 4250 10502 4306
rect 10558 4250 10626 4306
rect 10682 4250 10750 4306
rect 10806 4250 10874 4306
rect 10930 4250 10998 4306
rect 11054 4250 11122 4306
rect 11178 4250 11246 4306
rect 11302 4250 11370 4306
rect 11426 4250 11494 4306
rect 11550 4250 11618 4306
rect 11674 4250 11742 4306
rect 11798 4250 11866 4306
rect 11922 4250 11990 4306
rect 12046 4250 12114 4306
rect 12170 4250 12180 4306
rect 10244 4182 12180 4250
rect 10244 4126 10254 4182
rect 10310 4126 10378 4182
rect 10434 4126 10502 4182
rect 10558 4126 10626 4182
rect 10682 4126 10750 4182
rect 10806 4126 10874 4182
rect 10930 4126 10998 4182
rect 11054 4126 11122 4182
rect 11178 4126 11246 4182
rect 11302 4126 11370 4182
rect 11426 4126 11494 4182
rect 11550 4126 11618 4182
rect 11674 4126 11742 4182
rect 11798 4126 11866 4182
rect 11922 4126 11990 4182
rect 12046 4126 12114 4182
rect 12170 4126 12180 4182
rect 10244 4058 12180 4126
rect 10244 4002 10254 4058
rect 10310 4002 10378 4058
rect 10434 4002 10502 4058
rect 10558 4002 10626 4058
rect 10682 4002 10750 4058
rect 10806 4002 10874 4058
rect 10930 4002 10998 4058
rect 11054 4002 11122 4058
rect 11178 4002 11246 4058
rect 11302 4002 11370 4058
rect 11426 4002 11494 4058
rect 11550 4002 11618 4058
rect 11674 4002 11742 4058
rect 11798 4002 11866 4058
rect 11922 4002 11990 4058
rect 12046 4002 12114 4058
rect 12170 4002 12180 4058
rect 10244 3934 12180 4002
rect 10244 3878 10254 3934
rect 10310 3878 10378 3934
rect 10434 3878 10502 3934
rect 10558 3878 10626 3934
rect 10682 3878 10750 3934
rect 10806 3878 10874 3934
rect 10930 3878 10998 3934
rect 11054 3878 11122 3934
rect 11178 3878 11246 3934
rect 11302 3878 11370 3934
rect 11426 3878 11494 3934
rect 11550 3878 11618 3934
rect 11674 3878 11742 3934
rect 11798 3878 11866 3934
rect 11922 3878 11990 3934
rect 12046 3878 12114 3934
rect 12170 3878 12180 3934
rect 10244 3810 12180 3878
rect 10244 3754 10254 3810
rect 10310 3754 10378 3810
rect 10434 3754 10502 3810
rect 10558 3754 10626 3810
rect 10682 3754 10750 3810
rect 10806 3754 10874 3810
rect 10930 3754 10998 3810
rect 11054 3754 11122 3810
rect 11178 3754 11246 3810
rect 11302 3754 11370 3810
rect 11426 3754 11494 3810
rect 11550 3754 11618 3810
rect 11674 3754 11742 3810
rect 11798 3754 11866 3810
rect 11922 3754 11990 3810
rect 12046 3754 12114 3810
rect 12170 3754 12180 3810
rect 10244 3686 12180 3754
rect 10244 3630 10254 3686
rect 10310 3630 10378 3686
rect 10434 3630 10502 3686
rect 10558 3630 10626 3686
rect 10682 3630 10750 3686
rect 10806 3630 10874 3686
rect 10930 3630 10998 3686
rect 11054 3630 11122 3686
rect 11178 3630 11246 3686
rect 11302 3630 11370 3686
rect 11426 3630 11494 3686
rect 11550 3630 11618 3686
rect 11674 3630 11742 3686
rect 11798 3630 11866 3686
rect 11922 3630 11990 3686
rect 12046 3630 12114 3686
rect 12170 3630 12180 3686
rect 10244 3562 12180 3630
rect 10244 3506 10254 3562
rect 10310 3506 10378 3562
rect 10434 3506 10502 3562
rect 10558 3506 10626 3562
rect 10682 3506 10750 3562
rect 10806 3506 10874 3562
rect 10930 3506 10998 3562
rect 11054 3506 11122 3562
rect 11178 3506 11246 3562
rect 11302 3506 11370 3562
rect 11426 3506 11494 3562
rect 11550 3506 11618 3562
rect 11674 3506 11742 3562
rect 11798 3506 11866 3562
rect 11922 3506 11990 3562
rect 12046 3506 12114 3562
rect 12170 3506 12180 3562
rect 10244 3438 12180 3506
rect 10244 3382 10254 3438
rect 10310 3382 10378 3438
rect 10434 3382 10502 3438
rect 10558 3382 10626 3438
rect 10682 3382 10750 3438
rect 10806 3382 10874 3438
rect 10930 3382 10998 3438
rect 11054 3382 11122 3438
rect 11178 3382 11246 3438
rect 11302 3382 11370 3438
rect 11426 3382 11494 3438
rect 11550 3382 11618 3438
rect 11674 3382 11742 3438
rect 11798 3382 11866 3438
rect 11922 3382 11990 3438
rect 12046 3382 12114 3438
rect 12170 3382 12180 3438
rect 10244 3314 12180 3382
rect 10244 3258 10254 3314
rect 10310 3258 10378 3314
rect 10434 3258 10502 3314
rect 10558 3258 10626 3314
rect 10682 3258 10750 3314
rect 10806 3258 10874 3314
rect 10930 3258 10998 3314
rect 11054 3258 11122 3314
rect 11178 3258 11246 3314
rect 11302 3258 11370 3314
rect 11426 3258 11494 3314
rect 11550 3258 11618 3314
rect 11674 3258 11742 3314
rect 11798 3258 11866 3314
rect 11922 3258 11990 3314
rect 12046 3258 12114 3314
rect 12170 3258 12180 3314
rect 10244 3190 12180 3258
rect 10244 3134 10254 3190
rect 10310 3134 10378 3190
rect 10434 3134 10502 3190
rect 10558 3134 10626 3190
rect 10682 3134 10750 3190
rect 10806 3134 10874 3190
rect 10930 3134 10998 3190
rect 11054 3134 11122 3190
rect 11178 3134 11246 3190
rect 11302 3134 11370 3190
rect 11426 3134 11494 3190
rect 11550 3134 11618 3190
rect 11674 3134 11742 3190
rect 11798 3134 11866 3190
rect 11922 3134 11990 3190
rect 12046 3134 12114 3190
rect 12170 3134 12180 3190
rect 10244 3066 12180 3134
rect 10244 3010 10254 3066
rect 10310 3010 10378 3066
rect 10434 3010 10502 3066
rect 10558 3010 10626 3066
rect 10682 3010 10750 3066
rect 10806 3010 10874 3066
rect 10930 3010 10998 3066
rect 11054 3010 11122 3066
rect 11178 3010 11246 3066
rect 11302 3010 11370 3066
rect 11426 3010 11494 3066
rect 11550 3010 11618 3066
rect 11674 3010 11742 3066
rect 11798 3010 11866 3066
rect 11922 3010 11990 3066
rect 12046 3010 12114 3066
rect 12170 3010 12180 3066
rect 10244 2942 12180 3010
rect 10244 2886 10254 2942
rect 10310 2886 10378 2942
rect 10434 2886 10502 2942
rect 10558 2886 10626 2942
rect 10682 2886 10750 2942
rect 10806 2886 10874 2942
rect 10930 2886 10998 2942
rect 11054 2886 11122 2942
rect 11178 2886 11246 2942
rect 11302 2886 11370 2942
rect 11426 2886 11494 2942
rect 11550 2886 11618 2942
rect 11674 2886 11742 2942
rect 11798 2886 11866 2942
rect 11922 2886 11990 2942
rect 12046 2886 12114 2942
rect 12170 2886 12180 2942
rect 10244 2818 12180 2886
rect 10244 2762 10254 2818
rect 10310 2762 10378 2818
rect 10434 2762 10502 2818
rect 10558 2762 10626 2818
rect 10682 2762 10750 2818
rect 10806 2762 10874 2818
rect 10930 2762 10998 2818
rect 11054 2762 11122 2818
rect 11178 2762 11246 2818
rect 11302 2762 11370 2818
rect 11426 2762 11494 2818
rect 11550 2762 11618 2818
rect 11674 2762 11742 2818
rect 11798 2762 11866 2818
rect 11922 2762 11990 2818
rect 12046 2762 12114 2818
rect 12170 2762 12180 2818
rect 10244 2694 12180 2762
rect 10244 2638 10254 2694
rect 10310 2638 10378 2694
rect 10434 2638 10502 2694
rect 10558 2638 10626 2694
rect 10682 2638 10750 2694
rect 10806 2638 10874 2694
rect 10930 2638 10998 2694
rect 11054 2638 11122 2694
rect 11178 2638 11246 2694
rect 11302 2638 11370 2694
rect 11426 2638 11494 2694
rect 11550 2638 11618 2694
rect 11674 2638 11742 2694
rect 11798 2638 11866 2694
rect 11922 2638 11990 2694
rect 12046 2638 12114 2694
rect 12170 2638 12180 2694
rect 10244 2570 12180 2638
rect 10244 2514 10254 2570
rect 10310 2514 10378 2570
rect 10434 2514 10502 2570
rect 10558 2514 10626 2570
rect 10682 2514 10750 2570
rect 10806 2514 10874 2570
rect 10930 2514 10998 2570
rect 11054 2514 11122 2570
rect 11178 2514 11246 2570
rect 11302 2514 11370 2570
rect 11426 2514 11494 2570
rect 11550 2514 11618 2570
rect 11674 2514 11742 2570
rect 11798 2514 11866 2570
rect 11922 2514 11990 2570
rect 12046 2514 12114 2570
rect 12170 2514 12180 2570
rect 10244 2446 12180 2514
rect 10244 2390 10254 2446
rect 10310 2390 10378 2446
rect 10434 2390 10502 2446
rect 10558 2390 10626 2446
rect 10682 2390 10750 2446
rect 10806 2390 10874 2446
rect 10930 2390 10998 2446
rect 11054 2390 11122 2446
rect 11178 2390 11246 2446
rect 11302 2390 11370 2446
rect 11426 2390 11494 2446
rect 11550 2390 11618 2446
rect 11674 2390 11742 2446
rect 11798 2390 11866 2446
rect 11922 2390 11990 2446
rect 12046 2390 12114 2446
rect 12170 2390 12180 2446
rect 10244 2322 12180 2390
rect 10244 2266 10254 2322
rect 10310 2266 10378 2322
rect 10434 2266 10502 2322
rect 10558 2266 10626 2322
rect 10682 2266 10750 2322
rect 10806 2266 10874 2322
rect 10930 2266 10998 2322
rect 11054 2266 11122 2322
rect 11178 2266 11246 2322
rect 11302 2266 11370 2322
rect 11426 2266 11494 2322
rect 11550 2266 11618 2322
rect 11674 2266 11742 2322
rect 11798 2266 11866 2322
rect 11922 2266 11990 2322
rect 12046 2266 12114 2322
rect 12170 2266 12180 2322
rect 10244 2198 12180 2266
rect 10244 2142 10254 2198
rect 10310 2142 10378 2198
rect 10434 2142 10502 2198
rect 10558 2142 10626 2198
rect 10682 2142 10750 2198
rect 10806 2142 10874 2198
rect 10930 2142 10998 2198
rect 11054 2142 11122 2198
rect 11178 2142 11246 2198
rect 11302 2142 11370 2198
rect 11426 2142 11494 2198
rect 11550 2142 11618 2198
rect 11674 2142 11742 2198
rect 11798 2142 11866 2198
rect 11922 2142 11990 2198
rect 12046 2142 12114 2198
rect 12170 2142 12180 2198
rect 10244 2074 12180 2142
rect 10244 2018 10254 2074
rect 10310 2018 10378 2074
rect 10434 2018 10502 2074
rect 10558 2018 10626 2074
rect 10682 2018 10750 2074
rect 10806 2018 10874 2074
rect 10930 2018 10998 2074
rect 11054 2018 11122 2074
rect 11178 2018 11246 2074
rect 11302 2018 11370 2074
rect 11426 2018 11494 2074
rect 11550 2018 11618 2074
rect 11674 2018 11742 2074
rect 11798 2018 11866 2074
rect 11922 2018 11990 2074
rect 12046 2018 12114 2074
rect 12170 2018 12180 2074
rect 10244 1950 12180 2018
rect 10244 1894 10254 1950
rect 10310 1894 10378 1950
rect 10434 1894 10502 1950
rect 10558 1894 10626 1950
rect 10682 1894 10750 1950
rect 10806 1894 10874 1950
rect 10930 1894 10998 1950
rect 11054 1894 11122 1950
rect 11178 1894 11246 1950
rect 11302 1894 11370 1950
rect 11426 1894 11494 1950
rect 11550 1894 11618 1950
rect 11674 1894 11742 1950
rect 11798 1894 11866 1950
rect 11922 1894 11990 1950
rect 12046 1894 12114 1950
rect 12170 1894 12180 1950
rect 10244 1826 12180 1894
rect 10244 1770 10254 1826
rect 10310 1770 10378 1826
rect 10434 1770 10502 1826
rect 10558 1770 10626 1826
rect 10682 1770 10750 1826
rect 10806 1770 10874 1826
rect 10930 1770 10998 1826
rect 11054 1770 11122 1826
rect 11178 1770 11246 1826
rect 11302 1770 11370 1826
rect 11426 1770 11494 1826
rect 11550 1770 11618 1826
rect 11674 1770 11742 1826
rect 11798 1770 11866 1826
rect 11922 1770 11990 1826
rect 12046 1770 12114 1826
rect 12170 1770 12180 1826
rect 10244 1702 12180 1770
rect 10244 1646 10254 1702
rect 10310 1646 10378 1702
rect 10434 1646 10502 1702
rect 10558 1646 10626 1702
rect 10682 1646 10750 1702
rect 10806 1646 10874 1702
rect 10930 1646 10998 1702
rect 11054 1646 11122 1702
rect 11178 1646 11246 1702
rect 11302 1646 11370 1702
rect 11426 1646 11494 1702
rect 11550 1646 11618 1702
rect 11674 1646 11742 1702
rect 11798 1646 11866 1702
rect 11922 1646 11990 1702
rect 12046 1646 12114 1702
rect 12170 1646 12180 1702
rect 10244 1636 12180 1646
rect 12861 4554 14673 4564
rect 12861 4498 12871 4554
rect 12927 4498 12995 4554
rect 13051 4498 13119 4554
rect 13175 4498 13243 4554
rect 13299 4498 13367 4554
rect 13423 4498 13491 4554
rect 13547 4498 13615 4554
rect 13671 4498 13739 4554
rect 13795 4498 13863 4554
rect 13919 4498 13987 4554
rect 14043 4498 14111 4554
rect 14167 4498 14235 4554
rect 14291 4498 14359 4554
rect 14415 4498 14483 4554
rect 14539 4498 14607 4554
rect 14663 4498 14673 4554
rect 12861 4430 14673 4498
rect 12861 4374 12871 4430
rect 12927 4374 12995 4430
rect 13051 4374 13119 4430
rect 13175 4374 13243 4430
rect 13299 4374 13367 4430
rect 13423 4374 13491 4430
rect 13547 4374 13615 4430
rect 13671 4374 13739 4430
rect 13795 4374 13863 4430
rect 13919 4374 13987 4430
rect 14043 4374 14111 4430
rect 14167 4374 14235 4430
rect 14291 4374 14359 4430
rect 14415 4374 14483 4430
rect 14539 4374 14607 4430
rect 14663 4374 14673 4430
rect 12861 4306 14673 4374
rect 12861 4250 12871 4306
rect 12927 4250 12995 4306
rect 13051 4250 13119 4306
rect 13175 4250 13243 4306
rect 13299 4250 13367 4306
rect 13423 4250 13491 4306
rect 13547 4250 13615 4306
rect 13671 4250 13739 4306
rect 13795 4250 13863 4306
rect 13919 4250 13987 4306
rect 14043 4250 14111 4306
rect 14167 4250 14235 4306
rect 14291 4250 14359 4306
rect 14415 4250 14483 4306
rect 14539 4250 14607 4306
rect 14663 4250 14673 4306
rect 12861 4182 14673 4250
rect 12861 4126 12871 4182
rect 12927 4126 12995 4182
rect 13051 4126 13119 4182
rect 13175 4126 13243 4182
rect 13299 4126 13367 4182
rect 13423 4126 13491 4182
rect 13547 4126 13615 4182
rect 13671 4126 13739 4182
rect 13795 4126 13863 4182
rect 13919 4126 13987 4182
rect 14043 4126 14111 4182
rect 14167 4126 14235 4182
rect 14291 4126 14359 4182
rect 14415 4126 14483 4182
rect 14539 4126 14607 4182
rect 14663 4126 14673 4182
rect 12861 4058 14673 4126
rect 12861 4002 12871 4058
rect 12927 4002 12995 4058
rect 13051 4002 13119 4058
rect 13175 4002 13243 4058
rect 13299 4002 13367 4058
rect 13423 4002 13491 4058
rect 13547 4002 13615 4058
rect 13671 4002 13739 4058
rect 13795 4002 13863 4058
rect 13919 4002 13987 4058
rect 14043 4002 14111 4058
rect 14167 4002 14235 4058
rect 14291 4002 14359 4058
rect 14415 4002 14483 4058
rect 14539 4002 14607 4058
rect 14663 4002 14673 4058
rect 12861 3934 14673 4002
rect 12861 3878 12871 3934
rect 12927 3878 12995 3934
rect 13051 3878 13119 3934
rect 13175 3878 13243 3934
rect 13299 3878 13367 3934
rect 13423 3878 13491 3934
rect 13547 3878 13615 3934
rect 13671 3878 13739 3934
rect 13795 3878 13863 3934
rect 13919 3878 13987 3934
rect 14043 3878 14111 3934
rect 14167 3878 14235 3934
rect 14291 3878 14359 3934
rect 14415 3878 14483 3934
rect 14539 3878 14607 3934
rect 14663 3878 14673 3934
rect 12861 3810 14673 3878
rect 12861 3754 12871 3810
rect 12927 3754 12995 3810
rect 13051 3754 13119 3810
rect 13175 3754 13243 3810
rect 13299 3754 13367 3810
rect 13423 3754 13491 3810
rect 13547 3754 13615 3810
rect 13671 3754 13739 3810
rect 13795 3754 13863 3810
rect 13919 3754 13987 3810
rect 14043 3754 14111 3810
rect 14167 3754 14235 3810
rect 14291 3754 14359 3810
rect 14415 3754 14483 3810
rect 14539 3754 14607 3810
rect 14663 3754 14673 3810
rect 12861 3686 14673 3754
rect 12861 3630 12871 3686
rect 12927 3630 12995 3686
rect 13051 3630 13119 3686
rect 13175 3630 13243 3686
rect 13299 3630 13367 3686
rect 13423 3630 13491 3686
rect 13547 3630 13615 3686
rect 13671 3630 13739 3686
rect 13795 3630 13863 3686
rect 13919 3630 13987 3686
rect 14043 3630 14111 3686
rect 14167 3630 14235 3686
rect 14291 3630 14359 3686
rect 14415 3630 14483 3686
rect 14539 3630 14607 3686
rect 14663 3630 14673 3686
rect 12861 3562 14673 3630
rect 12861 3506 12871 3562
rect 12927 3506 12995 3562
rect 13051 3506 13119 3562
rect 13175 3506 13243 3562
rect 13299 3506 13367 3562
rect 13423 3506 13491 3562
rect 13547 3506 13615 3562
rect 13671 3506 13739 3562
rect 13795 3506 13863 3562
rect 13919 3506 13987 3562
rect 14043 3506 14111 3562
rect 14167 3506 14235 3562
rect 14291 3506 14359 3562
rect 14415 3506 14483 3562
rect 14539 3506 14607 3562
rect 14663 3506 14673 3562
rect 12861 3438 14673 3506
rect 12861 3382 12871 3438
rect 12927 3382 12995 3438
rect 13051 3382 13119 3438
rect 13175 3382 13243 3438
rect 13299 3382 13367 3438
rect 13423 3382 13491 3438
rect 13547 3382 13615 3438
rect 13671 3382 13739 3438
rect 13795 3382 13863 3438
rect 13919 3382 13987 3438
rect 14043 3382 14111 3438
rect 14167 3382 14235 3438
rect 14291 3382 14359 3438
rect 14415 3382 14483 3438
rect 14539 3382 14607 3438
rect 14663 3382 14673 3438
rect 12861 3314 14673 3382
rect 12861 3258 12871 3314
rect 12927 3258 12995 3314
rect 13051 3258 13119 3314
rect 13175 3258 13243 3314
rect 13299 3258 13367 3314
rect 13423 3258 13491 3314
rect 13547 3258 13615 3314
rect 13671 3258 13739 3314
rect 13795 3258 13863 3314
rect 13919 3258 13987 3314
rect 14043 3258 14111 3314
rect 14167 3258 14235 3314
rect 14291 3258 14359 3314
rect 14415 3258 14483 3314
rect 14539 3258 14607 3314
rect 14663 3258 14673 3314
rect 12861 3190 14673 3258
rect 12861 3134 12871 3190
rect 12927 3134 12995 3190
rect 13051 3134 13119 3190
rect 13175 3134 13243 3190
rect 13299 3134 13367 3190
rect 13423 3134 13491 3190
rect 13547 3134 13615 3190
rect 13671 3134 13739 3190
rect 13795 3134 13863 3190
rect 13919 3134 13987 3190
rect 14043 3134 14111 3190
rect 14167 3134 14235 3190
rect 14291 3134 14359 3190
rect 14415 3134 14483 3190
rect 14539 3134 14607 3190
rect 14663 3134 14673 3190
rect 12861 3066 14673 3134
rect 12861 3010 12871 3066
rect 12927 3010 12995 3066
rect 13051 3010 13119 3066
rect 13175 3010 13243 3066
rect 13299 3010 13367 3066
rect 13423 3010 13491 3066
rect 13547 3010 13615 3066
rect 13671 3010 13739 3066
rect 13795 3010 13863 3066
rect 13919 3010 13987 3066
rect 14043 3010 14111 3066
rect 14167 3010 14235 3066
rect 14291 3010 14359 3066
rect 14415 3010 14483 3066
rect 14539 3010 14607 3066
rect 14663 3010 14673 3066
rect 12861 2942 14673 3010
rect 12861 2886 12871 2942
rect 12927 2886 12995 2942
rect 13051 2886 13119 2942
rect 13175 2886 13243 2942
rect 13299 2886 13367 2942
rect 13423 2886 13491 2942
rect 13547 2886 13615 2942
rect 13671 2886 13739 2942
rect 13795 2886 13863 2942
rect 13919 2886 13987 2942
rect 14043 2886 14111 2942
rect 14167 2886 14235 2942
rect 14291 2886 14359 2942
rect 14415 2886 14483 2942
rect 14539 2886 14607 2942
rect 14663 2886 14673 2942
rect 12861 2818 14673 2886
rect 12861 2762 12871 2818
rect 12927 2762 12995 2818
rect 13051 2762 13119 2818
rect 13175 2762 13243 2818
rect 13299 2762 13367 2818
rect 13423 2762 13491 2818
rect 13547 2762 13615 2818
rect 13671 2762 13739 2818
rect 13795 2762 13863 2818
rect 13919 2762 13987 2818
rect 14043 2762 14111 2818
rect 14167 2762 14235 2818
rect 14291 2762 14359 2818
rect 14415 2762 14483 2818
rect 14539 2762 14607 2818
rect 14663 2762 14673 2818
rect 12861 2694 14673 2762
rect 12861 2638 12871 2694
rect 12927 2638 12995 2694
rect 13051 2638 13119 2694
rect 13175 2638 13243 2694
rect 13299 2638 13367 2694
rect 13423 2638 13491 2694
rect 13547 2638 13615 2694
rect 13671 2638 13739 2694
rect 13795 2638 13863 2694
rect 13919 2638 13987 2694
rect 14043 2638 14111 2694
rect 14167 2638 14235 2694
rect 14291 2638 14359 2694
rect 14415 2638 14483 2694
rect 14539 2638 14607 2694
rect 14663 2638 14673 2694
rect 12861 2570 14673 2638
rect 12861 2514 12871 2570
rect 12927 2514 12995 2570
rect 13051 2514 13119 2570
rect 13175 2514 13243 2570
rect 13299 2514 13367 2570
rect 13423 2514 13491 2570
rect 13547 2514 13615 2570
rect 13671 2514 13739 2570
rect 13795 2514 13863 2570
rect 13919 2514 13987 2570
rect 14043 2514 14111 2570
rect 14167 2514 14235 2570
rect 14291 2514 14359 2570
rect 14415 2514 14483 2570
rect 14539 2514 14607 2570
rect 14663 2514 14673 2570
rect 12861 2446 14673 2514
rect 12861 2390 12871 2446
rect 12927 2390 12995 2446
rect 13051 2390 13119 2446
rect 13175 2390 13243 2446
rect 13299 2390 13367 2446
rect 13423 2390 13491 2446
rect 13547 2390 13615 2446
rect 13671 2390 13739 2446
rect 13795 2390 13863 2446
rect 13919 2390 13987 2446
rect 14043 2390 14111 2446
rect 14167 2390 14235 2446
rect 14291 2390 14359 2446
rect 14415 2390 14483 2446
rect 14539 2390 14607 2446
rect 14663 2390 14673 2446
rect 12861 2322 14673 2390
rect 12861 2266 12871 2322
rect 12927 2266 12995 2322
rect 13051 2266 13119 2322
rect 13175 2266 13243 2322
rect 13299 2266 13367 2322
rect 13423 2266 13491 2322
rect 13547 2266 13615 2322
rect 13671 2266 13739 2322
rect 13795 2266 13863 2322
rect 13919 2266 13987 2322
rect 14043 2266 14111 2322
rect 14167 2266 14235 2322
rect 14291 2266 14359 2322
rect 14415 2266 14483 2322
rect 14539 2266 14607 2322
rect 14663 2266 14673 2322
rect 12861 2198 14673 2266
rect 12861 2142 12871 2198
rect 12927 2142 12995 2198
rect 13051 2142 13119 2198
rect 13175 2142 13243 2198
rect 13299 2142 13367 2198
rect 13423 2142 13491 2198
rect 13547 2142 13615 2198
rect 13671 2142 13739 2198
rect 13795 2142 13863 2198
rect 13919 2142 13987 2198
rect 14043 2142 14111 2198
rect 14167 2142 14235 2198
rect 14291 2142 14359 2198
rect 14415 2142 14483 2198
rect 14539 2142 14607 2198
rect 14663 2142 14673 2198
rect 12861 2074 14673 2142
rect 12861 2018 12871 2074
rect 12927 2018 12995 2074
rect 13051 2018 13119 2074
rect 13175 2018 13243 2074
rect 13299 2018 13367 2074
rect 13423 2018 13491 2074
rect 13547 2018 13615 2074
rect 13671 2018 13739 2074
rect 13795 2018 13863 2074
rect 13919 2018 13987 2074
rect 14043 2018 14111 2074
rect 14167 2018 14235 2074
rect 14291 2018 14359 2074
rect 14415 2018 14483 2074
rect 14539 2018 14607 2074
rect 14663 2018 14673 2074
rect 12861 1950 14673 2018
rect 12861 1894 12871 1950
rect 12927 1894 12995 1950
rect 13051 1894 13119 1950
rect 13175 1894 13243 1950
rect 13299 1894 13367 1950
rect 13423 1894 13491 1950
rect 13547 1894 13615 1950
rect 13671 1894 13739 1950
rect 13795 1894 13863 1950
rect 13919 1894 13987 1950
rect 14043 1894 14111 1950
rect 14167 1894 14235 1950
rect 14291 1894 14359 1950
rect 14415 1894 14483 1950
rect 14539 1894 14607 1950
rect 14663 1894 14673 1950
rect 12861 1826 14673 1894
rect 12861 1770 12871 1826
rect 12927 1770 12995 1826
rect 13051 1770 13119 1826
rect 13175 1770 13243 1826
rect 13299 1770 13367 1826
rect 13423 1770 13491 1826
rect 13547 1770 13615 1826
rect 13671 1770 13739 1826
rect 13795 1770 13863 1826
rect 13919 1770 13987 1826
rect 14043 1770 14111 1826
rect 14167 1770 14235 1826
rect 14291 1770 14359 1826
rect 14415 1770 14483 1826
rect 14539 1770 14607 1826
rect 14663 1770 14673 1826
rect 12861 1702 14673 1770
rect 12861 1646 12871 1702
rect 12927 1646 12995 1702
rect 13051 1646 13119 1702
rect 13175 1646 13243 1702
rect 13299 1646 13367 1702
rect 13423 1646 13491 1702
rect 13547 1646 13615 1702
rect 13671 1646 13739 1702
rect 13795 1646 13863 1702
rect 13919 1646 13987 1702
rect 14043 1646 14111 1702
rect 14167 1646 14235 1702
rect 14291 1646 14359 1702
rect 14415 1646 14483 1702
rect 14539 1646 14607 1702
rect 14663 1646 14673 1702
rect 12861 1636 14673 1646
rect 10 1604 86 1614
rect 14892 1614 14902 4586
rect 14958 1614 14968 4586
rect 14892 1604 14968 1614
use M1_NWELL_CDNS_40661956134204  M1_NWELL_CDNS_40661956134204_0
timestamp 1669390400
transform 1 0 2735 0 1 50138
box 0 0 1 1
use M1_NWELL_CDNS_40661956134204  M1_NWELL_CDNS_40661956134204_1
timestamp 1669390400
transform 1 0 12243 0 1 50138
box 0 0 1 1
use M1_NWELL_CDNS_40661956134205  M1_NWELL_CDNS_40661956134205_0
timestamp 1669390400
transform 1 0 7489 0 1 47838
box 0 0 1 1
use M1_NWELL_CDNS_40661956134205  M1_NWELL_CDNS_40661956134205_1
timestamp 1669390400
transform 1 0 7489 0 1 52438
box 0 0 1 1
use M1_PSUB_CDNS_40661956134197  M1_PSUB_CDNS_40661956134197_0
timestamp 1669390400
transform 1 0 379 0 1 55155
box 0 0 1 1
use M1_PSUB_CDNS_40661956134197  M1_PSUB_CDNS_40661956134197_1
timestamp 1669390400
transform 1 0 14599 0 1 55155
box 0 0 1 1
use M1_PSUB_CDNS_40661956134198  M1_PSUB_CDNS_40661956134198_0
timestamp 1669390400
transform 1 0 7489 0 1 53228
box 0 0 1 1
use M1_PSUB_CDNS_40661956134198  M1_PSUB_CDNS_40661956134198_1
timestamp 1669390400
transform 1 0 7489 0 1 57082
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_0
timestamp 1669390400
transform 1 0 3293 0 1 51539
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_1
timestamp 1669390400
transform 1 0 3293 0 1 50605
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_2
timestamp 1669390400
transform 1 0 3293 0 1 49671
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_3
timestamp 1669390400
transform 1 0 3293 0 1 48737
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_4
timestamp 1669390400
transform -1 0 11685 0 1 50605
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_5
timestamp 1669390400
transform -1 0 11685 0 1 48737
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_6
timestamp 1669390400
transform -1 0 11685 0 1 49671
box 0 0 1 1
use M1_PSUB_CDNS_40661956134199  M1_PSUB_CDNS_40661956134199_7
timestamp 1669390400
transform -1 0 11685 0 1 51539
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_0
timestamp 1669390400
transform 1 0 7489 0 -1 51852
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_1
timestamp 1669390400
transform 1 0 7489 0 1 51226
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_2
timestamp 1669390400
transform 1 0 7489 0 1 50918
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_3
timestamp 1669390400
transform 1 0 7489 0 1 50292
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_4
timestamp 1669390400
transform 1 0 7489 0 1 49984
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_5
timestamp 1669390400
transform 1 0 7489 0 1 49358
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_6
timestamp 1669390400
transform 1 0 7489 0 1 49050
box 0 0 1 1
use M1_PSUB_CDNS_40661956134200  M1_PSUB_CDNS_40661956134200_7
timestamp 1669390400
transform 1 0 7489 0 1 48424
box 0 0 1 1
use M1_PSUB_CDNS_40661956134201  M1_PSUB_CDNS_40661956134201_0
timestamp 1669390400
transform 1 0 7489 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_40661956134201  M1_PSUB_CDNS_40661956134201_1
timestamp 1669390400
transform 1 0 7489 0 1 51072
box 0 0 1 1
use M1_PSUB_CDNS_40661956134201  M1_PSUB_CDNS_40661956134201_2
timestamp 1669390400
transform 1 0 7489 0 1 49204
box 0 0 1 1
use M1_PSUB_CDNS_40661956134202  M1_PSUB_CDNS_40661956134202_0
timestamp 1669390400
transform 1 0 7489 0 -1 52006
box 0 0 1 1
use M1_PSUB_CDNS_40661956134202  M1_PSUB_CDNS_40661956134202_1
timestamp 1669390400
transform 1 0 7489 0 1 48270
box 0 0 1 1
use M1_PSUB_CDNS_40661956134203  M1_PSUB_CDNS_40661956134203_0
timestamp 1669390400
transform 1 0 3139 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_40661956134203  M1_PSUB_CDNS_40661956134203_1
timestamp 1669390400
transform -1 0 11839 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_40661956134228  M1_PSUB_CDNS_40661956134228_0
timestamp 1669390400
transform -1 0 13496 0 1 34924
box 0 0 1 1
use M1_PSUB_CDNS_40661956134229  M1_PSUB_CDNS_40661956134229_0
timestamp 1669390400
transform -1 0 14487 0 1 21924
box 0 0 1 1
use M1_PSUB_CDNS_40661956134229  M1_PSUB_CDNS_40661956134229_1
timestamp 1669390400
transform 1 0 491 0 1 21924
box 0 0 1 1
use M1_PSUB_CDNS_40661956134230  M1_PSUB_CDNS_40661956134230_0
timestamp 1669390400
transform 1 0 1241 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_40661956134230  M1_PSUB_CDNS_40661956134230_1
timestamp 1669390400
transform -1 0 13737 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_0
timestamp 1669390400
transform 1 0 14930 0 1 13500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_1
timestamp 1669390400
transform 1 0 14930 0 1 27900
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_2
timestamp 1669390400
transform 1 0 48 0 1 13500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_3
timestamp 1669390400
transform 1 0 48 0 1 27900
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_4
timestamp 1669390400
transform 1 0 48 0 1 45500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_5
timestamp 1669390400
transform 1 0 48 0 1 48700
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_6
timestamp 1669390400
transform 1 0 48 0 1 51900
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_7
timestamp 1669390400
transform 1 0 48 0 1 53500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_8
timestamp 1669390400
transform 1 0 48 0 1 37500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_9
timestamp 1669390400
transform 1 0 14930 0 1 37500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_10
timestamp 1669390400
transform 1 0 14930 0 1 45500
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_11
timestamp 1669390400
transform 1 0 14930 0 1 48700
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_12
timestamp 1669390400
transform 1 0 14930 0 1 51900
box 0 0 1 1
use M2_M1_CDNS_40661956134115  M2_M1_CDNS_40661956134115_13
timestamp 1669390400
transform 1 0 14930 0 1 53500
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_0
timestamp 1669390400
transform 1 0 4951 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_1
timestamp 1669390400
transform 1 0 4951 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_2
timestamp 1669390400
transform 1 0 4951 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_3
timestamp 1669390400
transform 1 0 4951 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_4
timestamp 1669390400
transform 1 0 10027 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_5
timestamp 1669390400
transform 1 0 10027 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_6
timestamp 1669390400
transform 1 0 10027 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_40661956134126  M2_M1_CDNS_40661956134126_7
timestamp 1669390400
transform 1 0 10027 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_0
timestamp 1669390400
transform 1 0 8842 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_1
timestamp 1669390400
transform 1 0 13767 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_2
timestamp 1669390400
transform 1 0 11212 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_3
timestamp 1669390400
transform 1 0 3766 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_4
timestamp 1669390400
transform 1 0 1211 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_5
timestamp 1669390400
transform 1 0 6136 0 1 792
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_6
timestamp 1669390400
transform 1 0 6136 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_7
timestamp 1669390400
transform 1 0 3766 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_8
timestamp 1669390400
transform 1 0 1211 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_9
timestamp 1669390400
transform 1 0 13767 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_10
timestamp 1669390400
transform 1 0 11212 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134140  M2_M1_CDNS_40661956134140_11
timestamp 1669390400
transform 1 0 8842 0 1 57473
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_0
timestamp 1669390400
transform 1 0 3275 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134145  M2_M1_CDNS_40661956134145_1
timestamp 1669390400
transform -1 0 11703 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134152  M2_M1_CDNS_40661956134152_0
timestamp 1669390400
transform 1 0 3943 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_40661956134152  M2_M1_CDNS_40661956134152_1
timestamp 1669390400
transform 1 0 3943 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_40661956134152  M2_M1_CDNS_40661956134152_2
timestamp 1669390400
transform -1 0 11035 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_40661956134152  M2_M1_CDNS_40661956134152_3
timestamp 1669390400
transform -1 0 11035 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_40661956134206  M2_M1_CDNS_40661956134206_0
timestamp 1669390400
transform 1 0 4951 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_40661956134206  M2_M1_CDNS_40661956134206_1
timestamp 1669390400
transform 1 0 4951 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_40661956134206  M2_M1_CDNS_40661956134206_2
timestamp 1669390400
transform 1 0 10027 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_40661956134206  M2_M1_CDNS_40661956134206_3
timestamp 1669390400
transform 1 0 10027 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_40661956134207  M2_M1_CDNS_40661956134207_0
timestamp 1669390400
transform 1 0 7489 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_40661956134207  M2_M1_CDNS_40661956134207_1
timestamp 1669390400
transform 1 0 7489 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_40661956134218  M2_M1_CDNS_40661956134218_0
timestamp 1669390400
transform 1 0 2581 0 1 53595
box 0 0 1 1
use M2_M1_CDNS_40661956134218  M2_M1_CDNS_40661956134218_1
timestamp 1669390400
transform 1 0 2581 0 1 56715
box 0 0 1 1
use M2_M1_CDNS_40661956134218  M2_M1_CDNS_40661956134218_2
timestamp 1669390400
transform 1 0 12397 0 1 53595
box 0 0 1 1
use M2_M1_CDNS_40661956134218  M2_M1_CDNS_40661956134218_3
timestamp 1669390400
transform 1 0 12397 0 1 56715
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_0
timestamp 1669390400
transform -1 0 6136 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_1
timestamp 1669390400
transform 1 0 6136 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_2
timestamp 1669390400
transform 1 0 6136 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_3
timestamp 1669390400
transform 1 0 6136 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_4
timestamp 1669390400
transform -1 0 8842 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_5
timestamp 1669390400
transform 1 0 8842 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_6
timestamp 1669390400
transform 1 0 8842 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_40661956134247  M2_M1_CDNS_40661956134247_7
timestamp 1669390400
transform 1 0 8842 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_40661956134249  M2_M1_CDNS_40661956134249_0
timestamp 1669390400
transform -1 0 6136 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134249  M2_M1_CDNS_40661956134249_1
timestamp 1669390400
transform 1 0 3766 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134249  M2_M1_CDNS_40661956134249_2
timestamp 1669390400
transform -1 0 11212 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134249  M2_M1_CDNS_40661956134249_3
timestamp 1669390400
transform -1 0 8842 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134250  M2_M1_CDNS_40661956134250_0
timestamp 1669390400
transform 1 0 7489 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_40661956134250  M2_M1_CDNS_40661956134250_1
timestamp 1669390400
transform 1 0 7489 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_40661956134250  M2_M1_CDNS_40661956134250_2
timestamp 1669390400
transform 1 0 7489 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_40661956134250  M2_M1_CDNS_40661956134250_3
timestamp 1669390400
transform 1 0 7489 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_0
timestamp 1669390400
transform 1 0 3943 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_1
timestamp 1669390400
transform 1 0 3943 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_2
timestamp 1669390400
transform 1 0 3943 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_3
timestamp 1669390400
transform -1 0 11035 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_4
timestamp 1669390400
transform -1 0 11035 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134251  M2_M1_CDNS_40661956134251_5
timestamp 1669390400
transform -1 0 11035 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_40661956134252  M2_M1_CDNS_40661956134252_0
timestamp 1669390400
transform 1 0 1211 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134252  M2_M1_CDNS_40661956134252_1
timestamp 1669390400
transform -1 0 13767 0 1 57078
box 0 0 1 1
use M2_M1_CDNS_40661956134253  M2_M1_CDNS_40661956134253_0
timestamp 1669390400
transform 1 0 1489 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134253  M2_M1_CDNS_40661956134253_1
timestamp 1669390400
transform -1 0 13489 0 1 53349
box 0 0 1 1
use M2_M1_CDNS_40661956134254  M2_M1_CDNS_40661956134254_0
timestamp 1669390400
transform 1 0 4951 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_40661956134254  M2_M1_CDNS_40661956134254_1
timestamp 1669390400
transform 1 0 10027 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_40661956134255  M2_M1_CDNS_40661956134255_0
timestamp 1669390400
transform 1 0 6136 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_40661956134255  M2_M1_CDNS_40661956134255_1
timestamp 1669390400
transform 1 0 6136 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_40661956134255  M2_M1_CDNS_40661956134255_2
timestamp 1669390400
transform 1 0 8842 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_40661956134255  M2_M1_CDNS_40661956134255_3
timestamp 1669390400
transform 1 0 8842 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_40661956134256  M2_M1_CDNS_40661956134256_0
timestamp 1669390400
transform 1 0 2616 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134256  M2_M1_CDNS_40661956134256_1
timestamp 1669390400
transform 1 0 12362 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_0
timestamp 1669390400
transform 1 0 14930 0 1 9500
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_1
timestamp 1669390400
transform 1 0 14930 0 1 6300
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_2
timestamp 1669390400
transform 1 0 14930 0 1 3100
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_3
timestamp 1669390400
transform 1 0 48 0 1 3100
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_4
timestamp 1669390400
transform 1 0 48 0 1 9500
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_5
timestamp 1669390400
transform 1 0 48 0 1 6300
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_6
timestamp 1669390400
transform 1 0 48 0 1 35100
box 0 0 1 1
use M2_M1_CDNS_40661956134258  M2_M1_CDNS_40661956134258_7
timestamp 1669390400
transform 1 0 14930 0 1 35100
box 0 0 1 1
use M2_M1_CDNS_40661956134261  M2_M1_CDNS_40661956134261_0
timestamp 1669390400
transform 1 0 48 0 1 56639
box 0 0 1 1
use M2_M1_CDNS_40661956134261  M2_M1_CDNS_40661956134261_1
timestamp 1669390400
transform 1 0 14930 0 1 56639
box 0 0 1 1
use M2_M1_CDNS_40661956134263  M2_M1_CDNS_40661956134263_0
timestamp 1669390400
transform 1 0 4053 0 1 54943
box 0 0 1 1
use M2_M1_CDNS_40661956134263  M2_M1_CDNS_40661956134263_1
timestamp 1669390400
transform -1 0 10925 0 1 54943
box 0 0 1 1
use M2_M1_CDNS_40661956134264  M2_M1_CDNS_40661956134264_0
timestamp 1669390400
transform 1 0 581 0 1 54943
box 0 0 1 1
use M2_M1_CDNS_40661956134264  M2_M1_CDNS_40661956134264_1
timestamp 1669390400
transform -1 0 14397 0 1 54943
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_0
timestamp 1669390400
transform 1 0 14930 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_1
timestamp 1669390400
transform 1 0 14930 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_2
timestamp 1669390400
transform 1 0 48 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_3
timestamp 1669390400
transform 1 0 48 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_4
timestamp 1669390400
transform 1 0 48 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_5
timestamp 1669390400
transform 1 0 48 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_6
timestamp 1669390400
transform 1 0 48 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_7
timestamp 1669390400
transform 1 0 48 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_8
timestamp 1669390400
transform 1 0 48 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_9
timestamp 1669390400
transform 1 0 14930 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_10
timestamp 1669390400
transform 1 0 14930 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_11
timestamp 1669390400
transform 1 0 14930 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_12
timestamp 1669390400
transform 1 0 14930 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134114  M3_M2_CDNS_40661956134114_13
timestamp 1669390400
transform 1 0 14930 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_0
timestamp 1669390400
transform -1 0 13767 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_1
timestamp 1669390400
transform -1 0 13767 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_2
timestamp 1669390400
transform 1 0 1211 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_3
timestamp 1669390400
transform 1 0 1211 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_4
timestamp 1669390400
transform 1 0 1211 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_5
timestamp 1669390400
transform 1 0 1211 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_6
timestamp 1669390400
transform 1 0 1211 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_7
timestamp 1669390400
transform 1 0 1211 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_8
timestamp 1669390400
transform 1 0 1211 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_9
timestamp 1669390400
transform -1 0 13767 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_10
timestamp 1669390400
transform -1 0 13767 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_11
timestamp 1669390400
transform -1 0 13767 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_12
timestamp 1669390400
transform -1 0 13767 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134119  M3_M2_CDNS_40661956134119_13
timestamp 1669390400
transform -1 0 13767 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_0
timestamp 1669390400
transform -1 0 13767 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_1
timestamp 1669390400
transform -1 0 13767 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_2
timestamp 1669390400
transform -1 0 13767 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_3
timestamp 1669390400
transform 1 0 1211 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_4
timestamp 1669390400
transform 1 0 1211 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_5
timestamp 1669390400
transform 1 0 1211 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_6
timestamp 1669390400
transform 1 0 1211 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134156  M3_M2_CDNS_40661956134156_7
timestamp 1669390400
transform -1 0 13767 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134219  M3_M2_CDNS_40661956134219_0
timestamp 1669390400
transform 1 0 2330 0 1 50304
box 0 0 1 1
use M3_M2_CDNS_40661956134219  M3_M2_CDNS_40661956134219_1
timestamp 1669390400
transform 1 0 2330 0 1 39105
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_0
timestamp 1669390400
transform -1 0 8842 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_1
timestamp 1669390400
transform -1 0 8842 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_2
timestamp 1669390400
transform -1 0 11212 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_3
timestamp 1669390400
transform -1 0 11212 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_4
timestamp 1669390400
transform 1 0 6136 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_5
timestamp 1669390400
transform 1 0 3766 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_6
timestamp 1669390400
transform 1 0 3766 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_7
timestamp 1669390400
transform 1 0 6136 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_8
timestamp 1669390400
transform 1 0 3766 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_9
timestamp 1669390400
transform 1 0 6136 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_10
timestamp 1669390400
transform 1 0 6136 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_11
timestamp 1669390400
transform 1 0 6136 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_12
timestamp 1669390400
transform 1 0 6136 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_13
timestamp 1669390400
transform 1 0 6136 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_14
timestamp 1669390400
transform 1 0 3766 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_15
timestamp 1669390400
transform 1 0 3766 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_16
timestamp 1669390400
transform 1 0 3766 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_17
timestamp 1669390400
transform 1 0 3766 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_18
timestamp 1669390400
transform -1 0 8842 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_19
timestamp 1669390400
transform -1 0 8842 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_20
timestamp 1669390400
transform -1 0 8842 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_21
timestamp 1669390400
transform -1 0 8842 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_22
timestamp 1669390400
transform -1 0 8842 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_23
timestamp 1669390400
transform -1 0 11212 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_24
timestamp 1669390400
transform -1 0 11212 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_25
timestamp 1669390400
transform -1 0 11212 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_26
timestamp 1669390400
transform -1 0 11212 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661956134221  M3_M2_CDNS_40661956134221_27
timestamp 1669390400
transform -1 0 11212 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_0
timestamp 1669390400
transform -1 0 11212 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_1
timestamp 1669390400
transform -1 0 11212 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_2
timestamp 1669390400
transform -1 0 11212 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_3
timestamp 1669390400
transform -1 0 8842 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_4
timestamp 1669390400
transform -1 0 8842 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_5
timestamp 1669390400
transform -1 0 8842 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_6
timestamp 1669390400
transform 1 0 6136 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_7
timestamp 1669390400
transform 1 0 3766 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_8
timestamp 1669390400
transform 1 0 6136 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_9
timestamp 1669390400
transform 1 0 3766 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_10
timestamp 1669390400
transform 1 0 6136 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_11
timestamp 1669390400
transform 1 0 3766 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_12
timestamp 1669390400
transform 1 0 3766 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_13
timestamp 1669390400
transform 1 0 6136 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_14
timestamp 1669390400
transform -1 0 11212 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134222  M3_M2_CDNS_40661956134222_15
timestamp 1669390400
transform -1 0 8842 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_0
timestamp 1669390400
transform -1 0 10027 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_1
timestamp 1669390400
transform -1 0 12397 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_2
timestamp 1669390400
transform 1 0 4951 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_3
timestamp 1669390400
transform 1 0 2581 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_4
timestamp 1669390400
transform 1 0 2581 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_5
timestamp 1669390400
transform 1 0 4951 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_6
timestamp 1669390400
transform 1 0 4951 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_7
timestamp 1669390400
transform 1 0 2581 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_8
timestamp 1669390400
transform 1 0 2581 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_9
timestamp 1669390400
transform 1 0 4951 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_10
timestamp 1669390400
transform 1 0 2581 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_11
timestamp 1669390400
transform 1 0 2581 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_12
timestamp 1669390400
transform 1 0 4951 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_13
timestamp 1669390400
transform 1 0 4951 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_14
timestamp 1669390400
transform -1 0 12397 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_15
timestamp 1669390400
transform -1 0 12397 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_16
timestamp 1669390400
transform -1 0 12397 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_17
timestamp 1669390400
transform -1 0 12397 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_18
timestamp 1669390400
transform -1 0 10027 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_19
timestamp 1669390400
transform -1 0 10027 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_20
timestamp 1669390400
transform -1 0 10027 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_21
timestamp 1669390400
transform -1 0 10027 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_22
timestamp 1669390400
transform -1 0 10027 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_23
timestamp 1669390400
transform -1 0 12397 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_24
timestamp 1669390400
transform -1 0 12397 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_25
timestamp 1669390400
transform -1 0 10027 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_26
timestamp 1669390400
transform 1 0 2581 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661956134223  M3_M2_CDNS_40661956134223_27
timestamp 1669390400
transform 1 0 4951 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_0
timestamp 1669390400
transform 1 0 7489 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_1
timestamp 1669390400
transform 1 0 7489 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_2
timestamp 1669390400
transform 1 0 7489 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_3
timestamp 1669390400
transform 1 0 7489 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_4
timestamp 1669390400
transform 1 0 7489 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_5
timestamp 1669390400
transform 1 0 7489 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_40661956134225  M3_M2_CDNS_40661956134225_6
timestamp 1669390400
transform 1 0 7489 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_0
timestamp 1669390400
transform -1 0 12397 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_1
timestamp 1669390400
transform -1 0 12397 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_2
timestamp 1669390400
transform -1 0 12397 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_3
timestamp 1669390400
transform -1 0 12397 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_4
timestamp 1669390400
transform -1 0 10027 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_5
timestamp 1669390400
transform -1 0 10027 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_6
timestamp 1669390400
transform -1 0 10027 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_7
timestamp 1669390400
transform -1 0 10027 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_8
timestamp 1669390400
transform 1 0 2581 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_9
timestamp 1669390400
transform 1 0 4951 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_10
timestamp 1669390400
transform 1 0 2581 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_11
timestamp 1669390400
transform 1 0 4951 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_12
timestamp 1669390400
transform 1 0 4951 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_13
timestamp 1669390400
transform 1 0 2581 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_14
timestamp 1669390400
transform 1 0 2581 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_15
timestamp 1669390400
transform 1 0 4951 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_16
timestamp 1669390400
transform 1 0 2581 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_17
timestamp 1669390400
transform 1 0 4951 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_18
timestamp 1669390400
transform -1 0 10027 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661956134226  M3_M2_CDNS_40661956134226_19
timestamp 1669390400
transform -1 0 12397 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661956134227  M3_M2_CDNS_40661956134227_0
timestamp 1669390400
transform 1 0 7489 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661956134227  M3_M2_CDNS_40661956134227_1
timestamp 1669390400
transform 1 0 7489 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661956134227  M3_M2_CDNS_40661956134227_2
timestamp 1669390400
transform 1 0 7489 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661956134227  M3_M2_CDNS_40661956134227_3
timestamp 1669390400
transform 1 0 7489 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661956134227  M3_M2_CDNS_40661956134227_4
timestamp 1669390400
transform 1 0 7489 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661956134257  M3_M2_CDNS_40661956134257_0
timestamp 1669390400
transform 1 0 1211 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134257  M3_M2_CDNS_40661956134257_1
timestamp 1669390400
transform -1 0 13767 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_0
timestamp 1669390400
transform 1 0 14930 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_1
timestamp 1669390400
transform 1 0 14930 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_2
timestamp 1669390400
transform 1 0 14930 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_3
timestamp 1669390400
transform 1 0 48 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_4
timestamp 1669390400
transform 1 0 48 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_5
timestamp 1669390400
transform 1 0 48 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_6
timestamp 1669390400
transform 1 0 48 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134259  M3_M2_CDNS_40661956134259_7
timestamp 1669390400
transform 1 0 14930 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661956134260  M3_M2_CDNS_40661956134260_0
timestamp 1669390400
transform 1 0 48 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134260  M3_M2_CDNS_40661956134260_1
timestamp 1669390400
transform 1 0 14930 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134262  M3_M2_CDNS_40661956134262_0
timestamp 1669390400
transform 1 0 3766 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134262  M3_M2_CDNS_40661956134262_1
timestamp 1669390400
transform 1 0 6136 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134262  M3_M2_CDNS_40661956134262_2
timestamp 1669390400
transform -1 0 8842 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661956134262  M3_M2_CDNS_40661956134262_3
timestamp 1669390400
transform -1 0 11212 0 1 56639
box 0 0 1 1
use comp018green_esd_clamp_v5p0_DVSS  comp018green_esd_clamp_v5p0_DVSS_0
timestamp 1669390400
transform 1 0 1008 0 1 1090
box -747 -51 13709 46134
use nmoscap_6p0_CDNS_406619561348  nmoscap_6p0_CDNS_406619561348_0
timestamp 1669390400
transform 1 0 835 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619561348  nmoscap_6p0_CDNS_406619561348_1
timestamp 1669390400
transform 1 0 11143 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619561348  nmoscap_6p0_CDNS_406619561348_2
timestamp 1669390400
transform 1 0 4271 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619561348  nmoscap_6p0_CDNS_406619561348_3
timestamp 1669390400
transform 1 0 7707 0 1 53655
box 0 0 1 1
use np_6p0_CDNS_406619561349  np_6p0_CDNS_406619561349_0
timestamp 1669390400
transform 1 0 3489 0 1 51439
box 0 0 1 1
use np_6p0_CDNS_406619561349  np_6p0_CDNS_406619561349_1
timestamp 1669390400
transform 1 0 3489 0 1 50505
box 0 0 1 1
use np_6p0_CDNS_406619561349  np_6p0_CDNS_406619561349_2
timestamp 1669390400
transform 1 0 3489 0 1 49571
box 0 0 1 1
use np_6p0_CDNS_406619561349  np_6p0_CDNS_406619561349_3
timestamp 1669390400
transform 1 0 3489 0 1 48637
box 0 0 1 1
<< labels >>
rlabel metal3 s 705 6432 705 6432 4 DVSS
port 1 nsew
rlabel metal3 s 752 3261 752 3261 4 DVSS
port 1 nsew
rlabel metal3 s 774 9418 774 9418 4 DVSS
port 1 nsew
rlabel metal3 s 774 13611 774 13611 4 DVSS
port 1 nsew
rlabel metal3 s 774 11795 774 11795 4 DVDD
port 2 nsew
rlabel metal3 s 774 22234 774 22234 4 DVDD
port 2 nsew
rlabel metal3 s 774 19120 774 19120 4 DVDD
port 2 nsew
rlabel metal3 s 774 15905 774 15905 4 DVDD
port 2 nsew
rlabel metal3 s 774 27853 774 27853 4 DVSS
port 1 nsew
rlabel metal3 s 774 29488 774 29488 4 DVDD
port 2 nsew
rlabel metal3 s 774 25470 774 25470 4 DVDD
port 2 nsew
rlabel metal3 s 774 35106 774 35106 4 DVSS
port 1 nsew
rlabel metal3 s 774 31879 774 31879 4 DVDD
port 2 nsew
rlabel metal3 s 774 37534 774 37534 4 DVSS
port 1 nsew
rlabel metal3 s 774 38969 774 38969 4 VDD
port 3 nsew
rlabel metal3 s 774 45369 774 45369 4 DVSS
port 1 nsew
rlabel metal3 s 774 43934 774 43934 4 DVDD
port 2 nsew
rlabel metal3 s 774 42169 774 42169 4 DVDD
port 2 nsew
rlabel metal3 s 774 40734 774 40734 4 DVDD
port 2 nsew
rlabel metal3 s 774 51769 774 51769 4 DVSS
port 1 nsew
rlabel metal3 s 774 50334 774 50334 4 VDD
port 3 nsew
rlabel metal3 s 774 48569 774 48569 4 DVSS
port 1 nsew
rlabel metal3 s 774 53534 774 53534 4 DVSS
port 1 nsew
rlabel metal3 s 774 56560 774 56560 4 DVSS
port 1 nsew
rlabel metal3 s 774 54969 774 54969 4 DVDD
port 2 nsew
rlabel metal3 s 774 47134 774 47134 4 DVDD
port 2 nsew
<< properties >>
string GDS_END 4238378
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4210318
string path 344.175 29.750 344.175 0.000 
<< end >>
