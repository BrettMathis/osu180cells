magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 3740 1620
<< nmos >>
rect 190 190 250 360
rect 540 190 600 360
rect 710 190 770 360
rect 820 190 880 360
rect 1170 190 1230 360
rect 1330 190 1390 360
rect 1500 190 1560 360
rect 1610 190 1670 360
rect 1780 190 1840 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2170 190 2230 360
rect 2340 190 2400 360
rect 2690 190 2750 360
rect 2800 190 2860 360
rect 2970 190 3030 360
rect 3320 190 3380 360
rect 3490 190 3550 360
<< pmos >>
rect 190 1090 250 1430
rect 510 1090 570 1430
rect 680 1090 740 1430
rect 850 1090 910 1430
rect 1170 1090 1230 1430
rect 1330 1090 1390 1430
rect 1500 1090 1560 1430
rect 1610 1090 1670 1430
rect 1780 1090 1840 1430
rect 1890 1090 1950 1430
rect 2060 1090 2120 1430
rect 2170 1090 2230 1430
rect 2340 1090 2400 1430
rect 2660 1090 2720 1430
rect 2830 1090 2890 1430
rect 3000 1090 3060 1430
rect 3320 1090 3380 1430
rect 3490 1090 3550 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 350 360
rect 250 252 282 298
rect 328 252 350 298
rect 250 190 350 252
rect 440 298 540 360
rect 440 252 462 298
rect 508 252 540 298
rect 440 190 540 252
rect 600 298 710 360
rect 600 252 632 298
rect 678 252 710 298
rect 600 190 710 252
rect 770 190 820 360
rect 880 298 980 360
rect 880 252 912 298
rect 958 252 980 298
rect 880 190 980 252
rect 1070 298 1170 360
rect 1070 252 1092 298
rect 1138 252 1170 298
rect 1070 190 1170 252
rect 1230 190 1330 360
rect 1390 298 1500 360
rect 1390 252 1422 298
rect 1468 252 1500 298
rect 1390 190 1500 252
rect 1560 190 1610 360
rect 1670 258 1780 360
rect 1670 212 1702 258
rect 1748 212 1780 258
rect 1670 190 1780 212
rect 1840 190 1890 360
rect 1950 298 2060 360
rect 1950 252 1982 298
rect 2028 252 2060 298
rect 1950 190 2060 252
rect 2120 190 2170 360
rect 2230 298 2340 360
rect 2230 252 2262 298
rect 2308 252 2340 298
rect 2230 190 2340 252
rect 2400 298 2500 360
rect 2400 252 2432 298
rect 2478 252 2500 298
rect 2400 190 2500 252
rect 2590 298 2690 360
rect 2590 252 2612 298
rect 2658 252 2690 298
rect 2590 190 2690 252
rect 2750 190 2800 360
rect 2860 298 2970 360
rect 2860 252 2892 298
rect 2938 252 2970 298
rect 2860 190 2970 252
rect 3030 298 3130 360
rect 3030 252 3062 298
rect 3108 252 3130 298
rect 3030 190 3130 252
rect 3220 298 3320 360
rect 3220 252 3242 298
rect 3288 252 3320 298
rect 3220 190 3320 252
rect 3380 298 3490 360
rect 3380 252 3412 298
rect 3458 252 3490 298
rect 3380 190 3490 252
rect 3550 298 3650 360
rect 3550 252 3582 298
rect 3628 252 3650 298
rect 3550 190 3650 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 350 1430
rect 250 1143 282 1377
rect 328 1143 350 1377
rect 250 1090 350 1143
rect 410 1377 510 1430
rect 410 1143 432 1377
rect 478 1143 510 1377
rect 410 1090 510 1143
rect 570 1405 680 1430
rect 570 1265 602 1405
rect 648 1265 680 1405
rect 570 1090 680 1265
rect 740 1405 850 1430
rect 740 1265 772 1405
rect 818 1265 850 1405
rect 740 1090 850 1265
rect 910 1405 1010 1430
rect 910 1265 942 1405
rect 988 1265 1010 1405
rect 910 1090 1010 1265
rect 1070 1377 1170 1430
rect 1070 1143 1092 1377
rect 1138 1143 1170 1377
rect 1070 1090 1170 1143
rect 1230 1090 1330 1430
rect 1390 1377 1500 1430
rect 1390 1143 1422 1377
rect 1468 1143 1500 1377
rect 1390 1090 1500 1143
rect 1560 1090 1610 1430
rect 1670 1377 1780 1430
rect 1670 1143 1702 1377
rect 1748 1143 1780 1377
rect 1670 1090 1780 1143
rect 1840 1090 1890 1430
rect 1950 1405 2060 1430
rect 1950 1265 1982 1405
rect 2028 1265 2060 1405
rect 1950 1090 2060 1265
rect 2120 1090 2170 1430
rect 2230 1405 2340 1430
rect 2230 1265 2262 1405
rect 2308 1265 2340 1405
rect 2230 1090 2340 1265
rect 2400 1377 2500 1430
rect 2400 1143 2432 1377
rect 2478 1143 2500 1377
rect 2400 1090 2500 1143
rect 2560 1410 2660 1430
rect 2560 1270 2582 1410
rect 2628 1270 2660 1410
rect 2560 1090 2660 1270
rect 2720 1408 2830 1430
rect 2720 1362 2752 1408
rect 2798 1362 2830 1408
rect 2720 1090 2830 1362
rect 2890 1368 3000 1430
rect 2890 1322 2922 1368
rect 2968 1322 3000 1368
rect 2890 1090 3000 1322
rect 3060 1377 3160 1430
rect 3060 1143 3092 1377
rect 3138 1143 3160 1377
rect 3060 1090 3160 1143
rect 3220 1377 3320 1430
rect 3220 1143 3242 1377
rect 3288 1143 3320 1377
rect 3220 1090 3320 1143
rect 3380 1377 3490 1430
rect 3380 1143 3412 1377
rect 3458 1143 3490 1377
rect 3380 1090 3490 1143
rect 3550 1377 3650 1430
rect 3550 1143 3582 1377
rect 3628 1143 3650 1377
rect 3550 1090 3650 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 462 252 508 298
rect 632 252 678 298
rect 912 252 958 298
rect 1092 252 1138 298
rect 1422 252 1468 298
rect 1702 212 1748 258
rect 1982 252 2028 298
rect 2262 252 2308 298
rect 2432 252 2478 298
rect 2612 252 2658 298
rect 2892 252 2938 298
rect 3062 252 3108 298
rect 3242 252 3288 298
rect 3412 252 3458 298
rect 3582 252 3628 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 432 1143 478 1377
rect 602 1265 648 1405
rect 772 1265 818 1405
rect 942 1265 988 1405
rect 1092 1143 1138 1377
rect 1422 1143 1468 1377
rect 1702 1143 1748 1377
rect 1982 1265 2028 1405
rect 2262 1265 2308 1405
rect 2432 1143 2478 1377
rect 2582 1270 2628 1410
rect 2752 1362 2798 1408
rect 2922 1322 2968 1368
rect 3092 1143 3138 1377
rect 3242 1143 3288 1377
rect 3412 1143 3458 1377
rect 3582 1143 3628 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 340 98 430 120
rect 340 52 362 98
rect 408 52 430 98
rect 340 30 430 52
rect 580 98 670 120
rect 580 52 602 98
rect 648 52 670 98
rect 580 30 670 52
rect 820 98 910 120
rect 820 52 842 98
rect 888 52 910 98
rect 820 30 910 52
rect 1060 98 1150 120
rect 1060 52 1082 98
rect 1128 52 1150 98
rect 1060 30 1150 52
rect 1300 98 1390 120
rect 1300 52 1322 98
rect 1368 52 1390 98
rect 1300 30 1390 52
rect 1540 98 1630 120
rect 1540 52 1562 98
rect 1608 52 1630 98
rect 1540 30 1630 52
rect 1780 98 1870 120
rect 1780 52 1802 98
rect 1848 52 1870 98
rect 1780 30 1870 52
rect 2020 98 2110 120
rect 2020 52 2042 98
rect 2088 52 2110 98
rect 2020 30 2110 52
rect 2260 98 2350 120
rect 2260 52 2282 98
rect 2328 52 2350 98
rect 2260 30 2350 52
rect 2500 98 2590 120
rect 2500 52 2522 98
rect 2568 52 2590 98
rect 2500 30 2590 52
rect 2740 98 2830 120
rect 2740 52 2762 98
rect 2808 52 2830 98
rect 2740 30 2830 52
rect 2980 98 3070 120
rect 2980 52 3002 98
rect 3048 52 3070 98
rect 2980 30 3070 52
rect 3220 98 3310 120
rect 3220 52 3242 98
rect 3288 52 3310 98
rect 3220 30 3310 52
rect 3460 98 3550 120
rect 3460 52 3482 98
rect 3528 52 3550 98
rect 3460 30 3550 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 340 1568 430 1590
rect 340 1522 362 1568
rect 408 1522 430 1568
rect 340 1500 430 1522
rect 580 1568 670 1590
rect 580 1522 602 1568
rect 648 1522 670 1568
rect 580 1500 670 1522
rect 820 1568 910 1590
rect 820 1522 842 1568
rect 888 1522 910 1568
rect 820 1500 910 1522
rect 1060 1568 1150 1590
rect 1060 1522 1082 1568
rect 1128 1522 1150 1568
rect 1060 1500 1150 1522
rect 1300 1568 1390 1590
rect 1300 1522 1322 1568
rect 1368 1522 1390 1568
rect 1300 1500 1390 1522
rect 1540 1568 1630 1590
rect 1540 1522 1562 1568
rect 1608 1522 1630 1568
rect 1540 1500 1630 1522
rect 1780 1568 1870 1590
rect 1780 1522 1802 1568
rect 1848 1522 1870 1568
rect 1780 1500 1870 1522
rect 2020 1568 2110 1590
rect 2020 1522 2042 1568
rect 2088 1522 2110 1568
rect 2020 1500 2110 1522
rect 2260 1568 2350 1590
rect 2260 1522 2282 1568
rect 2328 1522 2350 1568
rect 2260 1500 2350 1522
rect 2500 1568 2590 1590
rect 2500 1522 2522 1568
rect 2568 1522 2590 1568
rect 2500 1500 2590 1522
rect 2740 1568 2830 1590
rect 2740 1522 2762 1568
rect 2808 1522 2830 1568
rect 2740 1500 2830 1522
rect 2980 1568 3070 1590
rect 2980 1522 3002 1568
rect 3048 1522 3070 1568
rect 2980 1500 3070 1522
rect 3220 1568 3310 1590
rect 3220 1522 3242 1568
rect 3288 1522 3310 1568
rect 3220 1500 3310 1522
rect 3460 1568 3550 1590
rect 3460 1522 3482 1568
rect 3528 1522 3550 1568
rect 3460 1500 3550 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 362 52 408 98
rect 602 52 648 98
rect 842 52 888 98
rect 1082 52 1128 98
rect 1322 52 1368 98
rect 1562 52 1608 98
rect 1802 52 1848 98
rect 2042 52 2088 98
rect 2282 52 2328 98
rect 2522 52 2568 98
rect 2762 52 2808 98
rect 3002 52 3048 98
rect 3242 52 3288 98
rect 3482 52 3528 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 362 1522 408 1568
rect 602 1522 648 1568
rect 842 1522 888 1568
rect 1082 1522 1128 1568
rect 1322 1522 1368 1568
rect 1562 1522 1608 1568
rect 1802 1522 1848 1568
rect 2042 1522 2088 1568
rect 2282 1522 2328 1568
rect 2522 1522 2568 1568
rect 2762 1522 2808 1568
rect 3002 1522 3048 1568
rect 3242 1522 3288 1568
rect 3482 1522 3528 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 510 1430 570 1480
rect 680 1430 740 1480
rect 850 1430 910 1480
rect 1170 1430 1230 1480
rect 1330 1430 1390 1480
rect 1500 1430 1560 1480
rect 1610 1430 1670 1480
rect 1780 1430 1840 1480
rect 1890 1430 1950 1480
rect 2060 1430 2120 1480
rect 2170 1430 2230 1480
rect 2340 1430 2400 1480
rect 2660 1430 2720 1480
rect 2830 1430 2890 1480
rect 3000 1430 3060 1480
rect 3320 1430 3380 1480
rect 3490 1430 3550 1480
rect 190 1040 250 1090
rect 120 1018 250 1040
rect 120 972 142 1018
rect 188 972 250 1018
rect 120 950 250 972
rect 190 360 250 950
rect 510 780 570 1090
rect 680 910 740 1090
rect 680 883 800 910
rect 680 837 707 883
rect 753 837 800 883
rect 680 810 800 837
rect 510 753 630 780
rect 510 707 557 753
rect 603 707 630 753
rect 510 680 630 707
rect 510 630 570 680
rect 510 590 600 630
rect 540 360 600 590
rect 680 450 740 810
rect 850 780 910 1090
rect 1170 780 1230 1090
rect 1330 910 1390 1090
rect 1330 883 1430 910
rect 1330 837 1357 883
rect 1403 837 1430 883
rect 1330 810 1430 837
rect 850 753 990 780
rect 850 707 907 753
rect 953 707 990 753
rect 850 680 990 707
rect 1170 753 1290 780
rect 1170 707 1217 753
rect 1263 707 1290 753
rect 1170 680 1290 707
rect 850 450 910 680
rect 680 410 770 450
rect 710 360 770 410
rect 820 410 910 450
rect 820 360 880 410
rect 1170 360 1230 680
rect 1500 640 1560 1090
rect 1610 1040 1670 1090
rect 1780 1040 1840 1090
rect 1610 1013 1840 1040
rect 1610 970 1647 1013
rect 1620 967 1647 970
rect 1693 970 1840 1013
rect 1693 967 1720 970
rect 1620 920 1720 967
rect 1890 640 1950 1090
rect 2060 910 2120 1090
rect 2020 883 2120 910
rect 2020 837 2047 883
rect 2093 837 2120 883
rect 2020 810 2120 837
rect 2170 780 2230 1090
rect 2340 910 2400 1090
rect 2340 883 2440 910
rect 2340 837 2367 883
rect 2413 837 2440 883
rect 2340 810 2440 837
rect 2160 753 2260 780
rect 2160 707 2187 753
rect 2233 707 2260 753
rect 2160 680 2260 707
rect 2020 640 2120 650
rect 1330 623 2120 640
rect 1330 580 2047 623
rect 1330 360 1390 580
rect 2020 577 2047 580
rect 2093 577 2120 623
rect 2020 550 2120 577
rect 1460 493 1560 520
rect 1620 500 1720 520
rect 1460 447 1487 493
rect 1533 447 1560 493
rect 1460 420 1560 447
rect 1500 360 1560 420
rect 1610 493 1840 500
rect 1610 447 1647 493
rect 1693 447 1840 493
rect 1610 420 1840 447
rect 1610 360 1670 420
rect 1780 360 1840 420
rect 1890 483 1990 510
rect 1890 437 1917 483
rect 1963 437 1990 483
rect 1890 410 1990 437
rect 1890 360 1950 410
rect 2060 360 2120 550
rect 2170 360 2230 680
rect 2340 360 2400 810
rect 2660 510 2720 1090
rect 2830 910 2890 1090
rect 2770 883 2890 910
rect 2770 837 2817 883
rect 2863 837 2890 883
rect 2770 810 2890 837
rect 2580 483 2720 510
rect 2580 437 2617 483
rect 2663 450 2720 483
rect 2830 450 2890 810
rect 3000 630 3060 1090
rect 3320 650 3380 1090
rect 3490 910 3550 1090
rect 3430 883 3550 910
rect 3430 837 3457 883
rect 3503 837 3550 883
rect 3430 810 3550 837
rect 2663 437 2750 450
rect 2580 410 2750 437
rect 2690 360 2750 410
rect 2800 410 2890 450
rect 2970 590 3060 630
rect 3260 623 3380 650
rect 2970 510 3030 590
rect 3260 577 3307 623
rect 3353 577 3380 623
rect 3260 550 3380 577
rect 2970 483 3090 510
rect 2970 437 3017 483
rect 3063 437 3090 483
rect 2970 410 3090 437
rect 2800 360 2860 410
rect 2970 360 3030 410
rect 3320 360 3380 550
rect 3490 360 3550 810
rect 190 140 250 190
rect 540 140 600 190
rect 710 140 770 190
rect 820 140 880 190
rect 1170 140 1230 190
rect 1330 140 1390 190
rect 1500 140 1560 190
rect 1610 140 1670 190
rect 1780 140 1840 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2170 140 2230 190
rect 2340 140 2400 190
rect 2690 140 2750 190
rect 2800 140 2860 190
rect 2970 140 3030 190
rect 3320 140 3380 190
rect 3490 140 3550 190
<< polycontact >>
rect 142 972 188 1018
rect 707 837 753 883
rect 557 707 603 753
rect 1357 837 1403 883
rect 907 707 953 753
rect 1217 707 1263 753
rect 1647 967 1693 1013
rect 2047 837 2093 883
rect 2367 837 2413 883
rect 2187 707 2233 753
rect 2047 577 2093 623
rect 1487 447 1533 493
rect 1647 447 1693 493
rect 1917 437 1963 483
rect 2817 837 2863 883
rect 2617 437 2663 483
rect 3457 837 3503 883
rect 3307 577 3353 623
rect 3017 437 3063 483
<< metal1 >>
rect 0 1590 3740 1620
rect -810 1568 3740 1590
rect -810 1522 112 1568
rect 158 1566 362 1568
rect 408 1566 602 1568
rect 648 1566 842 1568
rect 888 1566 1082 1568
rect 1128 1566 1322 1568
rect 1368 1566 1562 1568
rect 1608 1566 1802 1568
rect 1848 1566 2042 1568
rect 2088 1566 2282 1568
rect 2328 1566 2522 1568
rect 2568 1566 2762 1568
rect 2808 1566 3002 1568
rect 3048 1566 3242 1568
rect 3288 1566 3482 1568
rect -810 1514 114 1522
rect 166 1514 354 1566
rect 408 1522 594 1566
rect 648 1522 834 1566
rect 888 1522 1074 1566
rect 1128 1522 1314 1566
rect 1368 1522 1554 1566
rect 1608 1522 1794 1566
rect 1848 1522 2034 1566
rect 2088 1522 2274 1566
rect 2328 1522 2514 1566
rect 2568 1522 2754 1566
rect 2808 1522 2994 1566
rect 3048 1522 3234 1566
rect 3288 1522 3474 1566
rect 3528 1522 3740 1568
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1794 1522
rect 1846 1514 2034 1522
rect 2086 1514 2274 1522
rect 2326 1514 2514 1522
rect 2566 1514 2754 1522
rect 2806 1514 2994 1522
rect 3046 1514 3234 1522
rect 3286 1514 3474 1522
rect 3526 1514 3740 1522
rect -810 1500 3740 1514
rect -810 1470 2930 1500
rect -700 1060 -650 1470
rect -40 1210 10 1470
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1090 160 1143
rect 280 1377 330 1470
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 110 1018 210 1020
rect 110 1016 142 1018
rect -700 930 -600 990
rect 110 964 134 1016
rect 188 972 210 1018
rect 186 964 210 972
rect 110 960 210 964
rect -130 800 -30 860
rect 280 500 330 1143
rect 430 1377 480 1430
rect 430 1143 432 1377
rect 478 1143 480 1377
rect 430 730 480 1143
rect 600 1405 650 1430
rect 600 1265 602 1405
rect 648 1265 650 1405
rect 600 1190 650 1265
rect 770 1405 820 1470
rect 770 1265 772 1405
rect 818 1265 820 1405
rect 770 1240 820 1265
rect 890 1430 940 1470
rect 890 1405 990 1430
rect 890 1265 942 1405
rect 988 1265 990 1405
rect 890 1190 990 1265
rect 600 1140 990 1190
rect 1090 1377 1140 1470
rect 1450 1430 1500 1470
rect 1090 1143 1092 1377
rect 1138 1143 1140 1377
rect 890 1060 940 1140
rect 1090 1090 1140 1143
rect 1420 1377 1500 1430
rect 1420 1143 1422 1377
rect 1468 1210 1500 1377
rect 1700 1377 1750 1470
rect 1468 1143 1470 1210
rect 1420 1040 1470 1143
rect 1700 1143 1702 1377
rect 1748 1143 1750 1377
rect 1940 1430 1990 1470
rect 1940 1405 2030 1430
rect 1940 1310 1982 1405
rect 1980 1265 1982 1310
rect 2028 1265 2030 1405
rect 1980 1240 2030 1265
rect 2260 1405 2310 1470
rect 2600 1430 2650 1470
rect 2260 1265 2262 1405
rect 2308 1265 2310 1405
rect 2260 1240 2310 1265
rect 2430 1377 2480 1430
rect 1700 1090 1750 1143
rect 1800 1190 2030 1240
rect 1090 990 1470 1040
rect 1620 1013 1720 1020
rect 680 886 780 890
rect 680 860 704 886
rect 520 834 704 860
rect 756 834 780 886
rect 520 830 780 834
rect 1090 860 1140 990
rect 1620 967 1647 1013
rect 1693 967 1720 1013
rect 1620 960 1720 967
rect 1330 886 1560 890
rect 1330 883 1484 886
rect 520 800 750 830
rect 1090 800 1310 860
rect 1330 837 1357 883
rect 1403 837 1484 883
rect 1330 834 1484 837
rect 1536 860 1560 886
rect 1536 834 1630 860
rect 1330 830 1630 834
rect 1480 800 1630 830
rect 380 670 480 730
rect 530 756 630 760
rect 530 704 554 756
rect 606 704 630 756
rect 530 700 630 704
rect 430 550 480 670
rect 670 550 730 800
rect 1090 760 1160 800
rect 880 756 1160 760
rect 880 704 904 756
rect 956 704 1160 756
rect 880 700 1160 704
rect 1190 756 1290 760
rect 1190 704 1214 756
rect 1266 704 1290 756
rect 1190 700 1290 704
rect 430 500 730 550
rect 900 500 950 510
rect 1090 500 1160 700
rect 1480 500 1540 800
rect 1640 500 1700 960
rect 1800 740 1850 1190
rect 2430 1143 2432 1377
rect 2478 1143 2480 1377
rect 2580 1410 2650 1430
rect 2580 1270 2582 1410
rect 2628 1290 2650 1410
rect 2750 1408 2800 1470
rect 2750 1362 2752 1408
rect 2798 1400 2800 1408
rect 2798 1362 2820 1400
rect 2750 1340 2820 1362
rect 2770 1290 2820 1340
rect 2920 1368 2970 1430
rect 2920 1322 2922 1368
rect 2968 1322 2970 1368
rect 2920 1290 2970 1322
rect 2628 1270 2970 1290
rect 2580 1240 2970 1270
rect 3090 1377 3140 1430
rect 2150 1016 2250 1020
rect 2150 964 2174 1016
rect 2226 964 2250 1016
rect 2150 960 2250 964
rect 2430 1000 2480 1143
rect 2600 1060 2650 1240
rect 2610 1020 2670 1040
rect 2770 1020 2820 1240
rect 3090 1143 3092 1377
rect 3138 1143 3140 1377
rect 3090 1020 3140 1143
rect 3240 1377 3290 1430
rect 3240 1143 3242 1377
rect 3288 1143 3290 1377
rect 2610 1016 3170 1020
rect 1790 690 1850 740
rect 1910 886 2120 890
rect 1910 834 2044 886
rect 2096 834 2120 886
rect 1910 830 2120 834
rect 260 496 360 500
rect 260 444 284 496
rect 336 444 360 496
rect 260 440 360 444
rect 630 496 980 500
rect 630 444 904 496
rect 956 444 980 496
rect 1090 460 1290 500
rect 630 440 980 444
rect 1080 450 1290 460
rect 280 430 340 440
rect 110 330 160 360
rect -700 90 -650 330
rect -350 90 -300 330
rect 100 298 160 330
rect 100 252 112 298
rect 158 252 160 298
rect 100 120 160 252
rect 280 298 330 430
rect 630 410 750 440
rect 900 430 950 440
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 460 298 510 360
rect 460 252 462 298
rect 508 252 510 298
rect 460 120 510 252
rect 630 298 680 410
rect 1080 400 1180 450
rect 1210 360 1290 450
rect 1460 493 1560 500
rect 1460 447 1487 493
rect 1533 447 1560 493
rect 1460 440 1560 447
rect 1620 496 1720 500
rect 1620 444 1644 496
rect 1696 444 1720 496
rect 1620 440 1720 444
rect 1790 370 1840 690
rect 1910 490 1970 830
rect 1980 800 2080 830
rect 2170 760 2230 960
rect 2430 950 2540 1000
rect 2430 890 2480 950
rect 2340 886 2480 890
rect 2340 834 2364 886
rect 2416 860 2480 886
rect 2490 860 2540 950
rect 2610 964 2614 1016
rect 2666 964 3094 1016
rect 3146 964 3170 1016
rect 2610 960 3170 964
rect 2610 940 2670 960
rect 2770 930 2870 960
rect 2770 920 2860 930
rect 2770 890 2820 920
rect 2770 886 2890 890
rect 2416 834 2720 860
rect 2340 830 2720 834
rect 2430 800 2720 830
rect 2770 834 2814 886
rect 2866 834 2890 886
rect 2770 830 2890 834
rect 2490 760 2540 800
rect 2160 756 2260 760
rect 2160 704 2184 756
rect 2236 704 2260 756
rect 2160 700 2260 704
rect 2430 710 2540 760
rect 2020 626 2120 630
rect 2020 574 2044 626
rect 2096 574 2120 626
rect 2020 570 2120 574
rect 2430 626 2490 710
rect 2430 574 2434 626
rect 2486 574 2490 626
rect 2430 550 2490 574
rect 1890 483 1990 490
rect 1890 437 1917 483
rect 1963 437 1990 483
rect 1890 430 1990 437
rect 2430 430 2480 550
rect 2650 490 2700 800
rect 2590 486 2700 490
rect 2590 434 2614 486
rect 2666 434 2700 486
rect 2590 430 2700 434
rect 2430 380 2700 430
rect 1790 366 2060 370
rect 630 252 632 298
rect 678 252 680 298
rect 630 190 680 252
rect 910 298 960 360
rect 910 252 912 298
rect 958 252 960 298
rect 910 250 960 252
rect 890 120 960 250
rect 1090 298 1140 360
rect 1210 330 1470 360
rect 1210 310 1500 330
rect 1790 320 1984 366
rect 1090 252 1092 298
rect 1138 252 1140 298
rect 1090 120 1140 252
rect 1420 298 1500 310
rect 1420 252 1422 298
rect 1468 252 1500 298
rect 1420 190 1500 252
rect 1450 120 1500 190
rect 1700 258 1750 280
rect 1700 212 1702 258
rect 1748 212 1750 258
rect 1700 120 1750 212
rect 1800 120 1850 320
rect 1980 314 1984 320
rect 2036 314 2060 366
rect 2260 330 2310 360
rect 1980 310 2060 314
rect 1980 298 2030 310
rect 1980 252 1982 298
rect 2028 252 2030 298
rect 1980 190 2030 252
rect 2250 298 2310 330
rect 2250 252 2262 298
rect 2308 252 2310 298
rect 2250 120 2310 252
rect 2430 298 2480 380
rect 2610 330 2660 360
rect 2430 252 2432 298
rect 2478 252 2480 298
rect 2430 160 2480 252
rect 2600 298 2660 330
rect 2600 252 2612 298
rect 2658 252 2660 298
rect 2600 120 2660 252
rect 2770 160 2820 830
rect 3090 630 3140 960
rect 3240 890 3290 1143
rect 3410 1377 3460 1500
rect 3410 1143 3412 1377
rect 3458 1143 3460 1377
rect 3410 1090 3460 1143
rect 3580 1377 3630 1430
rect 3580 1143 3582 1377
rect 3628 1143 3630 1377
rect 3580 1030 3630 1143
rect 3580 1016 3680 1030
rect 3580 964 3604 1016
rect 3656 964 3680 1016
rect 3580 960 3680 964
rect 3580 950 3670 960
rect 3240 886 3530 890
rect 3240 834 3454 886
rect 3506 834 3530 886
rect 3240 830 3530 834
rect 2890 626 3380 630
rect 2890 574 3304 626
rect 3356 574 3380 626
rect 2890 570 3380 574
rect 2890 298 2940 570
rect 2990 486 3090 490
rect 2990 434 3014 486
rect 3066 434 3090 486
rect 3460 460 3510 830
rect 2990 430 3090 434
rect 3240 410 3510 460
rect 2890 252 2892 298
rect 2938 252 2940 298
rect 2890 190 2940 252
rect 3060 298 3110 360
rect 3060 252 3062 298
rect 3108 252 3110 298
rect 3060 120 3110 252
rect 3240 298 3290 410
rect 3240 252 3242 298
rect 3288 252 3290 298
rect 3240 190 3290 252
rect 3410 298 3460 360
rect 3410 252 3412 298
rect 3458 252 3460 298
rect 3410 120 3460 252
rect 3580 298 3630 950
rect 3580 252 3582 298
rect 3628 252 3630 298
rect 3580 190 3630 252
rect 0 106 3740 120
rect 0 98 114 106
rect 0 90 112 98
rect -810 52 112 90
rect 166 54 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 2566 98 2754 106
rect 2806 98 2994 106
rect 3046 98 3234 106
rect 3286 98 3474 106
rect 3526 98 3740 106
rect 408 54 594 98
rect 648 54 834 98
rect 888 54 1074 98
rect 1128 54 1314 98
rect 1368 54 1554 98
rect 1608 54 1794 98
rect 1848 54 2034 98
rect 2088 54 2274 98
rect 2328 54 2514 98
rect 2568 54 2754 98
rect 2808 54 2994 98
rect 3048 54 3234 98
rect 3288 54 3474 98
rect 158 52 362 54
rect 408 52 602 54
rect 648 52 842 54
rect 888 52 1082 54
rect 1128 52 1322 54
rect 1368 52 1562 54
rect 1608 52 1802 54
rect 1848 52 2042 54
rect 2088 52 2282 54
rect 2328 52 2522 54
rect 2568 52 2762 54
rect 2808 52 3002 54
rect 3048 52 3242 54
rect 3288 52 3482 54
rect 3528 52 3740 98
rect -810 0 3740 52
rect -810 -30 2930 0
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 114 1514 166 1522
rect 354 1522 362 1566
rect 362 1522 406 1566
rect 594 1522 602 1566
rect 602 1522 646 1566
rect 834 1522 842 1566
rect 842 1522 886 1566
rect 1074 1522 1082 1566
rect 1082 1522 1126 1566
rect 1314 1522 1322 1566
rect 1322 1522 1366 1566
rect 1554 1522 1562 1566
rect 1562 1522 1606 1566
rect 1794 1522 1802 1566
rect 1802 1522 1846 1566
rect 2034 1522 2042 1566
rect 2042 1522 2086 1566
rect 2274 1522 2282 1566
rect 2282 1522 2326 1566
rect 2514 1522 2522 1566
rect 2522 1522 2566 1566
rect 2754 1522 2762 1566
rect 2762 1522 2806 1566
rect 2994 1522 3002 1566
rect 3002 1522 3046 1566
rect 3234 1522 3242 1566
rect 3242 1522 3286 1566
rect 3474 1522 3482 1566
rect 3482 1522 3526 1566
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 1794 1514 1846 1522
rect 2034 1514 2086 1522
rect 2274 1514 2326 1522
rect 2514 1514 2566 1522
rect 2754 1514 2806 1522
rect 2994 1514 3046 1522
rect 3234 1514 3286 1522
rect 3474 1514 3526 1522
rect 134 972 142 1016
rect 142 972 186 1016
rect 134 964 186 972
rect 704 883 756 886
rect 704 837 707 883
rect 707 837 753 883
rect 753 837 756 883
rect 704 834 756 837
rect 1484 834 1536 886
rect 554 753 606 756
rect 554 707 557 753
rect 557 707 603 753
rect 603 707 606 753
rect 554 704 606 707
rect 904 753 956 756
rect 904 707 907 753
rect 907 707 953 753
rect 953 707 956 753
rect 904 704 956 707
rect 1214 753 1266 756
rect 1214 707 1217 753
rect 1217 707 1263 753
rect 1263 707 1266 753
rect 1214 704 1266 707
rect 2174 964 2226 1016
rect 2044 883 2096 886
rect 2044 837 2047 883
rect 2047 837 2093 883
rect 2093 837 2096 883
rect 2044 834 2096 837
rect 284 444 336 496
rect 904 444 956 496
rect 1644 493 1696 496
rect 1644 447 1647 493
rect 1647 447 1693 493
rect 1693 447 1696 493
rect 1644 444 1696 447
rect 2364 883 2416 886
rect 2364 837 2367 883
rect 2367 837 2413 883
rect 2413 837 2416 883
rect 2614 964 2666 1016
rect 3094 964 3146 1016
rect 2364 834 2416 837
rect 2814 883 2866 886
rect 2814 837 2817 883
rect 2817 837 2863 883
rect 2863 837 2866 883
rect 2814 834 2866 837
rect 2184 753 2236 756
rect 2184 707 2187 753
rect 2187 707 2233 753
rect 2233 707 2236 753
rect 2184 704 2236 707
rect 2044 623 2096 626
rect 2044 577 2047 623
rect 2047 577 2093 623
rect 2093 577 2096 623
rect 2044 574 2096 577
rect 2434 574 2486 626
rect 2614 483 2666 486
rect 2614 437 2617 483
rect 2617 437 2663 483
rect 2663 437 2666 483
rect 2614 434 2666 437
rect 1984 314 2036 366
rect 3604 964 3656 1016
rect 3454 883 3506 886
rect 3454 837 3457 883
rect 3457 837 3503 883
rect 3503 837 3506 883
rect 3454 834 3506 837
rect 3304 623 3356 626
rect 3304 577 3307 623
rect 3307 577 3353 623
rect 3353 577 3356 623
rect 3304 574 3356 577
rect 3014 483 3066 486
rect 3014 437 3017 483
rect 3017 437 3063 483
rect 3063 437 3066 483
rect 3014 434 3066 437
rect 114 98 166 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 2754 98 2806 106
rect 2994 98 3046 106
rect 3234 98 3286 106
rect 3474 98 3526 106
rect 354 54 362 98
rect 362 54 406 98
rect 594 54 602 98
rect 602 54 646 98
rect 834 54 842 98
rect 842 54 886 98
rect 1074 54 1082 98
rect 1082 54 1126 98
rect 1314 54 1322 98
rect 1322 54 1366 98
rect 1554 54 1562 98
rect 1562 54 1606 98
rect 1794 54 1802 98
rect 1802 54 1846 98
rect 2034 54 2042 98
rect 2042 54 2086 98
rect 2274 54 2282 98
rect 2282 54 2326 98
rect 2514 54 2522 98
rect 2522 54 2566 98
rect 2754 54 2762 98
rect 2762 54 2806 98
rect 2994 54 3002 98
rect 3002 54 3046 98
rect 3234 54 3242 98
rect 3242 54 3286 98
rect 3474 54 3482 98
rect 3482 54 3526 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect 1780 1570 1860 1580
rect 2020 1570 2100 1580
rect 2260 1570 2340 1580
rect 2500 1570 2580 1580
rect 2740 1570 2820 1580
rect 2980 1570 3060 1580
rect 3220 1570 3300 1580
rect 3460 1570 3540 1580
rect 90 1566 190 1570
rect 90 1550 114 1566
rect -710 1540 -630 1550
rect -470 1540 -390 1550
rect -230 1540 -150 1550
rect 10 1540 114 1550
rect -720 1480 -620 1540
rect -480 1480 -380 1540
rect -240 1480 -140 1540
rect 0 1514 114 1540
rect 166 1514 190 1566
rect 330 1566 430 1570
rect 330 1550 354 1566
rect 250 1540 354 1550
rect 0 1510 190 1514
rect 240 1514 354 1540
rect 406 1514 430 1566
rect 570 1566 670 1570
rect 570 1550 594 1566
rect 490 1540 594 1550
rect 240 1510 430 1514
rect 480 1514 594 1540
rect 646 1514 670 1566
rect 810 1566 910 1570
rect 810 1550 834 1566
rect 730 1540 834 1550
rect 480 1510 670 1514
rect 720 1514 834 1540
rect 886 1514 910 1566
rect 1050 1566 1150 1570
rect 1050 1550 1074 1566
rect 970 1540 1074 1550
rect 720 1510 910 1514
rect 960 1514 1074 1540
rect 1126 1514 1150 1566
rect 1290 1566 1390 1570
rect 1290 1550 1314 1566
rect 1210 1540 1314 1550
rect 960 1510 1150 1514
rect 1200 1514 1314 1540
rect 1366 1514 1390 1566
rect 1530 1566 1630 1570
rect 1530 1550 1554 1566
rect 1450 1540 1554 1550
rect 1200 1510 1390 1514
rect 1440 1514 1554 1540
rect 1606 1514 1630 1566
rect 1770 1566 1870 1570
rect 1770 1550 1794 1566
rect 1690 1540 1794 1550
rect 1440 1510 1630 1514
rect 1680 1514 1794 1540
rect 1846 1514 1870 1566
rect 2010 1566 2110 1570
rect 2010 1550 2034 1566
rect 1930 1540 2034 1550
rect 1680 1510 1870 1514
rect 1920 1514 2034 1540
rect 2086 1514 2110 1566
rect 2250 1566 2350 1570
rect 2250 1550 2274 1566
rect 2170 1540 2274 1550
rect 1920 1510 2110 1514
rect 2160 1514 2274 1540
rect 2326 1514 2350 1566
rect 2490 1566 2590 1570
rect 2490 1550 2514 1566
rect 2410 1540 2514 1550
rect 2160 1510 2350 1514
rect 2400 1514 2514 1540
rect 2566 1514 2590 1566
rect 2730 1566 2830 1570
rect 2730 1550 2754 1566
rect 2650 1540 2754 1550
rect 2400 1510 2590 1514
rect 2640 1514 2754 1540
rect 2806 1514 2830 1566
rect 2640 1510 2830 1514
rect 2970 1566 3070 1570
rect 2970 1514 2994 1566
rect 3046 1514 3070 1566
rect 2970 1510 3070 1514
rect 3210 1566 3310 1570
rect 3210 1514 3234 1566
rect 3286 1514 3310 1566
rect 3210 1510 3310 1514
rect 3450 1566 3550 1570
rect 3450 1514 3474 1566
rect 3526 1514 3550 1566
rect 3450 1510 3550 1514
rect 0 1500 180 1510
rect 240 1500 420 1510
rect 480 1500 660 1510
rect 720 1500 900 1510
rect 960 1500 1140 1510
rect 1200 1500 1380 1510
rect 1440 1500 1620 1510
rect 1680 1500 1860 1510
rect 1920 1500 2100 1510
rect 2160 1500 2340 1510
rect 2400 1500 2580 1510
rect 2640 1500 2820 1510
rect 2980 1500 3060 1510
rect 3220 1500 3300 1510
rect 3460 1500 3540 1510
rect 0 1480 100 1500
rect 240 1480 340 1500
rect 480 1480 580 1500
rect 720 1480 820 1500
rect 960 1480 1060 1500
rect 1200 1480 1300 1500
rect 1440 1480 1540 1500
rect 1680 1480 1780 1500
rect 1920 1480 2020 1500
rect 2160 1480 2260 1500
rect 2400 1480 2500 1500
rect 2640 1480 2740 1500
rect -710 1470 -630 1480
rect -470 1470 -390 1480
rect -230 1470 -150 1480
rect 10 1470 90 1480
rect 250 1470 330 1480
rect 490 1470 570 1480
rect 730 1470 810 1480
rect 970 1470 1050 1480
rect 1210 1470 1290 1480
rect 1450 1470 1530 1480
rect 1690 1470 1770 1480
rect 1930 1470 2010 1480
rect 2170 1470 2250 1480
rect 2410 1470 2490 1480
rect 2650 1470 2730 1480
rect 700 1120 2870 1150
rect -110 1090 2870 1120
rect -110 1060 2060 1090
rect -700 920 -600 1000
rect -110 870 -50 1060
rect 110 1016 210 1030
rect 110 964 134 1016
rect 186 964 210 1016
rect 110 950 210 964
rect 700 900 760 1060
rect 2000 900 2060 1060
rect 2160 1020 2240 1030
rect 2600 1020 2680 1030
rect 2150 1016 2690 1020
rect 2150 964 2174 1016
rect 2226 964 2614 1016
rect 2666 964 2690 1016
rect 2810 1000 2870 1090
rect 2780 990 2870 1000
rect 2150 960 2690 964
rect 2160 950 2240 960
rect 2600 950 2680 960
rect 2770 930 2870 990
rect 3070 1016 3170 1030
rect 3590 1020 3670 1030
rect 3070 964 3094 1016
rect 3146 964 3170 1016
rect 3070 950 3170 964
rect 3580 1016 3680 1020
rect 3580 964 3604 1016
rect 3656 964 3680 1016
rect 3580 960 3680 964
rect 3590 950 3670 960
rect 2780 920 2870 930
rect 2810 900 2870 920
rect 680 886 780 900
rect 680 870 704 886
rect -130 790 -30 870
rect 650 834 704 870
rect 756 860 780 886
rect 1460 890 1550 900
rect 2000 890 2120 900
rect 2350 890 2430 900
rect 1460 886 2440 890
rect 1210 860 1310 870
rect 1460 860 1484 886
rect 756 834 1484 860
rect 1536 834 2044 886
rect 2096 834 2364 886
rect 2416 834 2440 886
rect 2790 886 2890 900
rect 3440 890 3520 900
rect 2630 860 2710 870
rect 650 830 2440 834
rect 650 800 1630 830
rect 1980 820 2120 830
rect 2350 820 2430 830
rect 650 790 740 800
rect 1210 790 1310 800
rect 1540 790 1620 800
rect 1980 790 2080 820
rect 2620 800 2720 860
rect 2790 834 2814 886
rect 2866 834 2890 886
rect 2790 820 2890 834
rect 3430 886 3530 890
rect 3430 834 3454 886
rect 3506 834 3530 886
rect 3430 830 3530 834
rect 3440 820 3520 830
rect 2630 790 2710 800
rect 530 756 630 770
rect 380 660 480 740
rect 530 704 554 756
rect 606 704 630 756
rect 530 690 630 704
rect 880 756 980 770
rect 880 704 904 756
rect 956 704 980 756
rect 880 690 980 704
rect 1190 756 1290 770
rect 2170 760 2250 770
rect 1190 704 1214 756
rect 1266 704 1290 756
rect 1190 690 1290 704
rect 2160 756 2260 760
rect 2160 704 2184 756
rect 2236 704 2260 756
rect 2160 700 2260 704
rect 2170 690 2250 700
rect 260 500 360 510
rect 550 500 610 690
rect 2030 630 2110 640
rect 2420 630 2500 640
rect 3290 630 3370 640
rect 2020 626 2520 630
rect 2020 574 2044 626
rect 2096 574 2434 626
rect 2486 574 2520 626
rect 2020 570 2520 574
rect 3220 626 3380 630
rect 3220 574 3304 626
rect 3356 574 3380 626
rect 3220 570 3380 574
rect 2030 560 2110 570
rect 2420 560 2500 570
rect 3290 560 3370 570
rect 260 496 610 500
rect 260 444 284 496
rect 336 444 610 496
rect 260 440 610 444
rect 260 430 360 440
rect 550 240 610 440
rect 880 500 980 510
rect 1630 500 1710 510
rect 880 496 1720 500
rect 880 444 904 496
rect 956 444 1644 496
rect 1696 444 1720 496
rect 880 440 1720 444
rect 2590 486 2690 500
rect 880 430 980 440
rect 1630 430 1710 440
rect 2590 434 2614 486
rect 2666 434 2690 486
rect 2590 420 2690 434
rect 2970 486 3090 500
rect 2970 434 3014 486
rect 3066 434 3090 486
rect 2970 420 3090 434
rect 1970 370 2050 380
rect 2590 370 2670 420
rect 1960 366 2670 370
rect 1960 314 1984 366
rect 2036 314 2670 366
rect 1960 310 2670 314
rect 1970 300 2050 310
rect 2970 240 3030 420
rect 550 180 3030 240
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 2740 110 2820 120
rect 2980 110 3060 120
rect 3220 110 3300 120
rect 3460 110 3540 120
rect 90 106 190 110
rect 90 90 114 106
rect -710 80 -630 90
rect -470 80 -390 90
rect -230 80 -150 90
rect 10 80 114 90
rect -720 20 -620 80
rect -480 20 -380 80
rect -240 20 -140 80
rect 0 54 114 80
rect 166 54 190 106
rect 330 106 430 110
rect 330 90 354 106
rect 250 80 354 90
rect 0 50 190 54
rect 240 54 354 80
rect 406 54 430 106
rect 570 106 670 110
rect 570 90 594 106
rect 490 80 594 90
rect 240 50 430 54
rect 480 54 594 80
rect 646 54 670 106
rect 810 106 910 110
rect 810 90 834 106
rect 730 80 834 90
rect 480 50 670 54
rect 720 54 834 80
rect 886 54 910 106
rect 1050 106 1150 110
rect 1050 90 1074 106
rect 970 80 1074 90
rect 720 50 910 54
rect 960 54 1074 80
rect 1126 54 1150 106
rect 1290 106 1390 110
rect 1290 90 1314 106
rect 1210 80 1314 90
rect 960 50 1150 54
rect 1200 54 1314 80
rect 1366 54 1390 106
rect 1530 106 1630 110
rect 1530 90 1554 106
rect 1450 80 1554 90
rect 1200 50 1390 54
rect 1440 54 1554 80
rect 1606 54 1630 106
rect 1770 106 1870 110
rect 1770 90 1794 106
rect 1690 80 1794 90
rect 1440 50 1630 54
rect 1680 54 1794 80
rect 1846 54 1870 106
rect 2010 106 2110 110
rect 2010 90 2034 106
rect 1930 80 2034 90
rect 1680 50 1870 54
rect 1920 54 2034 80
rect 2086 54 2110 106
rect 2250 106 2350 110
rect 2250 90 2274 106
rect 2170 80 2274 90
rect 1920 50 2110 54
rect 2160 54 2274 80
rect 2326 54 2350 106
rect 2490 106 2590 110
rect 2490 90 2514 106
rect 2410 80 2514 90
rect 2160 50 2350 54
rect 2400 54 2514 80
rect 2566 54 2590 106
rect 2730 106 2830 110
rect 2730 90 2754 106
rect 2650 80 2754 90
rect 2400 50 2590 54
rect 2640 54 2754 80
rect 2806 54 2830 106
rect 2640 50 2830 54
rect 2970 106 3070 110
rect 2970 54 2994 106
rect 3046 54 3070 106
rect 2970 50 3070 54
rect 3210 106 3310 110
rect 3210 54 3234 106
rect 3286 54 3310 106
rect 3210 50 3310 54
rect 3450 106 3550 110
rect 3450 54 3474 106
rect 3526 54 3550 106
rect 3450 50 3550 54
rect 0 40 180 50
rect 240 40 420 50
rect 480 40 660 50
rect 720 40 900 50
rect 960 40 1140 50
rect 1200 40 1380 50
rect 1440 40 1620 50
rect 1680 40 1860 50
rect 1920 40 2100 50
rect 2160 40 2340 50
rect 2400 40 2580 50
rect 2640 40 2820 50
rect 2980 40 3060 50
rect 3220 40 3300 50
rect 3460 40 3540 50
rect 0 20 100 40
rect 240 20 340 40
rect 480 20 580 40
rect 720 20 820 40
rect 960 20 1060 40
rect 1200 20 1300 40
rect 1440 20 1540 40
rect 1680 20 1780 40
rect 1920 20 2020 40
rect 2160 20 2260 40
rect 2400 20 2500 40
rect 2640 20 2740 40
rect -710 10 -630 20
rect -470 10 -390 20
rect -230 10 -150 20
rect 10 10 90 20
rect 250 10 330 20
rect 490 10 570 20
rect 730 10 810 20
rect 970 10 1050 20
rect 1210 10 1290 20
rect 1450 10 1530 20
rect 1690 10 1770 20
rect 1930 10 2010 20
rect 2170 10 2250 20
rect 2410 10 2490 20
rect 2650 10 2730 20
<< labels >>
rlabel metal2 s -710 1470 -630 1550 4 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -710 10 -630 90 4 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 380 660 480 740 4 D
port 1 nsew signal input
rlabel metal2 s -110 790 -50 1120 4 SN
port 2 nsew signal output
rlabel metal2 s -700 920 -600 1000 4 RN
port 3 nsew signal input
rlabel metal2 s 2780 920 2860 1000 4 Q
port 4 nsew signal output
rlabel metal2 s 2630 790 2710 870 4 QN
port 5 nsew signal output
rlabel metal2 s 650 790 740 870 4 CLK
port 6 nsew clock input
rlabel metal2 s 1210 790 1310 870 1 CLK
port 6 nsew clock input
rlabel metal2 s 1540 790 1620 870 1 CLK
port 6 nsew clock input
rlabel metal2 s 650 800 1630 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 670 410 730 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 650 410 750 470 1 CLK
port 6 nsew clock input
rlabel metal1 s 520 800 750 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 1100 400 1160 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 1080 400 1180 460 1 CLK
port 6 nsew clock input
rlabel metal1 s 1100 800 1310 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 1530 800 1630 860 1 CLK
port 6 nsew clock input
rlabel metal1 s 380 670 480 730 1 D
port 1 nsew signal input
rlabel metal2 s 2770 930 2870 990 1 Q
port 4 nsew signal output
rlabel metal1 s 2770 160 2820 1400 1 Q
port 4 nsew signal output
rlabel metal1 s 2770 920 2860 1000 1 Q
port 4 nsew signal output
rlabel metal1 s 2770 930 2870 1000 1 Q
port 4 nsew signal output
rlabel metal2 s 2620 800 2720 860 1 QN
port 5 nsew signal output
rlabel metal1 s 2430 160 2480 430 1 QN
port 5 nsew signal output
rlabel metal1 s 2430 800 2480 1400 1 QN
port 5 nsew signal output
rlabel metal1 s 2430 380 2700 430 1 QN
port 5 nsew signal output
rlabel metal1 s 2650 380 2700 860 1 QN
port 5 nsew signal output
rlabel metal1 s 2430 800 2720 860 1 QN
port 5 nsew signal output
rlabel metal1 s -700 930 -600 990 3 RN
port 3 nsew signal input
rlabel metal2 s -130 790 -30 870 3 SN
port 2 nsew signal output
rlabel metal2 s 2000 790 2060 1120 1 SN
port 2 nsew signal output
rlabel metal2 s -110 1060 2060 1120 1 SN
port 2 nsew signal output
rlabel metal2 s 1980 790 2080 870 1 SN
port 2 nsew signal output
rlabel metal1 s -130 800 -30 860 3 SN
port 2 nsew signal output
rlabel metal1 s 1980 800 2080 860 1 SN
port 2 nsew signal output
rlabel metal2 s -720 1480 -620 1540 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -470 1470 -390 1550 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -480 1480 -380 1540 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -230 1470 -150 1550 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -240 1480 -140 1540 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 10 1470 90 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 0 1480 100 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 250 1470 330 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 240 1480 340 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 490 1470 570 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 480 1480 580 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 730 1470 810 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 720 1480 820 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 970 1470 1050 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 960 1480 1060 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1210 1470 1290 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1200 1480 1300 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1450 1470 1530 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1440 1480 1540 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1690 1470 1770 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1680 1480 1780 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1930 1470 2010 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 1920 1480 2020 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2170 1470 2250 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2160 1480 2260 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2410 1470 2490 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2400 1480 2500 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2650 1470 2730 1550 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s 2640 1480 2740 1540 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s -700 1060 -650 1590 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s -40 1210 10 1590 3 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 280 1060 330 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 890 1060 940 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 1450 1210 1500 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 1940 1310 1990 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s 2600 1060 2650 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal1 s -810 1470 2930 1590 1 VDD
port 14 nsew power bidirectional abutment
rlabel metal2 s -720 20 -620 80 3 VSS
port 15 nsew ground bidirectional
rlabel metal2 s -470 10 -390 90 3 VSS
port 15 nsew ground bidirectional
rlabel metal2 s -480 20 -380 80 3 VSS
port 15 nsew ground bidirectional
rlabel metal2 s -230 10 -150 90 3 VSS
port 15 nsew ground bidirectional
rlabel metal2 s -240 20 -140 80 3 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 10 10 90 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 0 20 100 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 250 10 330 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 240 20 340 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 490 10 570 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 480 20 580 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 730 10 810 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 720 20 820 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 970 10 1050 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 960 20 1060 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1210 10 1290 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1200 20 1300 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1450 10 1530 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1440 20 1540 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1690 10 1770 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1680 20 1780 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1930 10 2010 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 1920 20 2020 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2170 10 2250 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2160 20 2260 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2410 10 2490 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2400 20 2500 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2650 10 2730 90 1 VSS
port 15 nsew ground bidirectional
rlabel metal2 s 2640 20 2740 80 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s -700 -30 -650 330 3 VSS
port 15 nsew ground bidirectional
rlabel metal1 s -350 -30 -300 330 3 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 100 -30 150 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 280 -30 330 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 890 -30 940 250 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 1450 -30 1500 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 1800 -30 1850 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 2250 -30 2300 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s 2600 -30 2650 330 1 VSS
port 15 nsew ground bidirectional
rlabel metal1 s -810 -30 2930 90 1 VSS
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX -810 -30 2930 1590
string GDS_END 306764
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 268690
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
