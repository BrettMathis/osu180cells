magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 352 323
<< polysilicon >>
rect -31 182 89 254
rect -31 -74 89 -1
use pmos_5p04310590878119_256x8m81  pmos_5p04310590878119_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 302
<< properties >>
string GDS_END 360376
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 360062
<< end >>
