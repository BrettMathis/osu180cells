magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 1340 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 520 190 580 360
rect 750 190 810 360
rect 910 190 970 360
rect 1080 190 1140 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 520 700 580 1040
rect 750 700 810 1040
rect 910 700 970 1040
rect 1080 700 1140 1040
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 520 360
rect 580 258 750 360
rect 580 212 642 258
rect 688 212 750 258
rect 580 190 750 212
rect 810 190 910 360
rect 970 293 1080 360
rect 970 247 1002 293
rect 1048 247 1080 293
rect 970 190 1080 247
rect 1140 298 1240 360
rect 1140 252 1172 298
rect 1218 252 1240 298
rect 1140 190 1240 252
<< pdiff >>
rect 90 987 190 1040
rect 90 753 112 987
rect 158 753 190 987
rect 90 700 190 753
rect 250 1017 360 1040
rect 250 783 282 1017
rect 328 783 360 1017
rect 250 700 360 783
rect 420 700 520 1040
rect 580 1018 750 1040
rect 580 972 642 1018
rect 688 972 750 1018
rect 580 700 750 972
rect 810 700 910 1040
rect 970 1017 1080 1040
rect 970 783 1002 1017
rect 1048 783 1080 1017
rect 970 700 1080 783
rect 1140 987 1240 1040
rect 1140 753 1172 987
rect 1218 753 1240 987
rect 1140 700 1240 753
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 642 212 688 258
rect 1002 247 1048 293
rect 1172 252 1218 298
<< pdiffc >>
rect 112 753 158 987
rect 282 783 328 1017
rect 642 972 688 1018
rect 1002 783 1048 1017
rect 1172 753 1218 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 520 1040 580 1090
rect 750 1040 810 1090
rect 910 1040 970 1090
rect 1080 1040 1140 1090
rect 190 680 250 700
rect 360 680 420 700
rect 190 630 420 680
rect 520 680 580 700
rect 750 680 810 700
rect 520 658 620 680
rect 190 520 250 630
rect 520 612 547 658
rect 593 612 620 658
rect 520 590 620 612
rect 710 653 810 680
rect 710 607 737 653
rect 783 607 810 653
rect 910 680 970 700
rect 1080 680 1140 700
rect 910 630 1140 680
rect 710 580 810 607
rect 190 493 320 520
rect 190 447 247 493
rect 293 447 320 493
rect 190 420 320 447
rect 470 453 580 480
rect 190 380 420 420
rect 470 407 497 453
rect 543 407 580 453
rect 470 380 580 407
rect 190 360 250 380
rect 360 360 420 380
rect 520 360 580 380
rect 750 360 810 580
rect 870 558 970 580
rect 870 512 897 558
rect 943 512 970 558
rect 1080 520 1140 630
rect 870 490 970 512
rect 910 360 970 490
rect 1020 493 1140 520
rect 1020 447 1047 493
rect 1093 447 1140 493
rect 1020 420 1140 447
rect 1080 360 1140 420
rect 190 140 250 190
rect 360 140 420 190
rect 520 140 580 190
rect 750 140 810 190
rect 910 140 970 190
rect 1080 140 1140 190
<< polycontact >>
rect 547 612 593 658
rect 737 607 783 653
rect 247 447 293 493
rect 497 407 543 453
rect 897 512 943 558
rect 1047 447 1093 493
<< metal1 >>
rect 0 1178 1340 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1340 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1340 1176
rect 0 1110 1340 1124
rect 110 987 160 1040
rect 110 753 112 987
rect 158 753 160 987
rect 280 1017 330 1110
rect 280 783 282 1017
rect 328 783 330 1017
rect 640 1018 690 1040
rect 640 972 642 1018
rect 688 972 690 1018
rect 640 910 690 972
rect 630 890 690 910
rect 1000 1017 1050 1110
rect 610 886 710 890
rect 610 834 634 886
rect 686 834 710 886
rect 610 830 710 834
rect 280 760 330 783
rect 1000 783 1002 1017
rect 1048 783 1050 1017
rect 110 650 160 753
rect 540 730 940 780
rect 1000 760 1050 783
rect 1170 987 1220 1040
rect 540 660 600 730
rect 890 680 940 730
rect 1170 753 1172 987
rect 1218 753 1220 987
rect 1170 680 1220 753
rect 520 658 620 660
rect 110 600 470 650
rect 520 612 547 658
rect 593 612 620 658
rect 520 610 620 612
rect 730 653 790 680
rect 110 298 160 600
rect 410 560 470 600
rect 730 607 737 653
rect 783 607 790 653
rect 730 560 790 607
rect 890 620 1220 680
rect 890 570 950 620
rect 410 510 790 560
rect 870 558 970 570
rect 870 512 897 558
rect 943 512 970 558
rect 870 510 970 512
rect 220 496 320 500
rect 220 444 244 496
rect 296 444 320 496
rect 1020 496 1120 500
rect 1020 460 1044 496
rect 220 440 320 444
rect 470 453 1044 460
rect 470 407 497 453
rect 543 444 1044 453
rect 1096 444 1120 496
rect 543 440 1120 444
rect 543 407 1090 440
rect 470 400 1090 407
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 630 340 690 350
rect 280 252 282 298
rect 328 252 330 298
rect 610 336 710 340
rect 610 284 634 336
rect 686 284 710 336
rect 610 280 710 284
rect 1000 293 1050 350
rect 630 260 690 280
rect 280 120 330 252
rect 640 258 690 260
rect 640 212 642 258
rect 688 212 690 258
rect 640 190 690 212
rect 1000 247 1002 293
rect 1048 247 1050 293
rect 1000 120 1050 247
rect 1170 298 1220 620
rect 1170 252 1172 298
rect 1218 252 1220 298
rect 1170 190 1220 252
rect 0 106 1340 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1340 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1340 54
rect 0 0 1340 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 634 834 686 886
rect 244 493 296 496
rect 244 447 247 493
rect 247 447 293 493
rect 293 447 296 493
rect 244 444 296 447
rect 1044 493 1096 496
rect 1044 447 1047 493
rect 1047 447 1093 493
rect 1093 447 1096 493
rect 1044 444 1096 447
rect 634 284 686 336
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 630 900 690 910
rect 620 886 700 900
rect 620 834 634 886
rect 686 834 700 886
rect 620 820 700 834
rect 230 500 310 510
rect 220 496 320 500
rect 220 444 244 496
rect 296 444 320 496
rect 220 440 320 444
rect 230 430 310 440
rect 630 350 690 820
rect 1030 500 1110 510
rect 1020 496 1120 500
rect 1020 444 1044 496
rect 1096 444 1120 496
rect 1020 440 1120 444
rect 1030 430 1110 440
rect 610 336 710 350
rect 610 284 634 336
rect 686 284 710 336
rect 610 270 710 284
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 230 430 310 510 4 A
port 1 nsew signal input
rlabel metal2 s 630 270 690 910 4 Y
port 2 nsew signal output
rlabel metal2 s 1030 430 1110 510 4 B
port 3 nsew signal input
rlabel metal2 s 220 440 320 500 1 A
port 1 nsew signal input
rlabel metal1 s 220 440 320 500 1 A
port 1 nsew signal input
rlabel metal2 s 1020 440 1120 500 1 B
port 3 nsew signal input
rlabel metal1 s 470 400 1090 460 1 B
port 3 nsew signal input
rlabel metal1 s 1020 440 1120 500 1 B
port 3 nsew signal input
rlabel metal2 s 90 1120 190 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 280 760 330 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1000 760 1050 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1110 1340 1230 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 280 0 330 360 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 1000 0 1050 350 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 0 1340 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 620 820 700 900 1 Y
port 2 nsew signal output
rlabel metal2 s 610 270 710 350 1 Y
port 2 nsew signal output
rlabel metal1 s 630 830 690 910 1 Y
port 2 nsew signal output
rlabel metal1 s 640 830 690 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 610 830 710 890 1 Y
port 2 nsew signal output
rlabel metal1 s 640 190 690 350 1 Y
port 2 nsew signal output
rlabel metal1 s 630 260 690 350 1 Y
port 2 nsew signal output
rlabel metal1 s 610 280 710 340 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1340 1230
string GDS_END 467820
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 456294
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
