magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -71 65 71 71
rect -71 -65 -65 65
rect 65 -65 71 65
rect -71 -71 71 -65
<< via1 >>
rect -65 -65 65 65
<< metal2 >>
rect -71 65 71 71
rect -71 -65 -65 65
rect 65 -65 71 65
rect -71 -71 71 -65
<< properties >>
string GDS_END 400594
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 399886
<< end >>
