magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 464 5462 1094
rect -86 453 86 464
rect 4277 453 5462 464
<< pwell >>
rect 1836 456 3739 464
rect 1688 453 3739 456
rect -86 -86 5462 453
<< mvnmos >>
rect 124 156 244 274
rect 348 156 468 274
rect 516 156 636 274
rect 740 156 860 274
rect 908 156 1028 274
rect 1360 146 1480 304
rect 1584 146 1704 304
rect 1968 226 2088 344
rect 2192 226 2312 344
rect 2360 226 2480 344
rect 2560 226 2680 344
rect 2828 226 2948 344
rect 3032 226 3152 344
rect 3256 226 3376 344
rect 3480 226 3600 344
rect 3888 157 4008 275
rect 4056 157 4176 275
rect 4280 157 4400 275
rect 4540 69 4660 333
rect 4908 69 5028 333
rect 5132 69 5252 333
<< mvpmos >>
rect 154 652 254 852
rect 358 652 458 852
rect 506 652 606 852
rect 740 652 840 852
rect 888 652 988 852
rect 1320 608 1420 884
rect 1524 608 1624 884
rect 1872 588 1972 788
rect 2076 588 2176 788
rect 2280 588 2380 788
rect 2560 620 2660 820
rect 2908 705 3008 905
rect 3188 588 3288 788
rect 3392 588 3492 788
rect 3596 588 3696 788
rect 3954 652 4054 852
rect 4158 652 4258 852
rect 4408 573 4508 939
rect 4616 573 4716 939
rect 4900 573 5000 939
rect 5104 573 5204 939
<< mvndiff >>
rect 1272 291 1360 304
rect 36 215 124 274
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 274
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 274
rect 636 215 740 274
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 274
rect 1028 205 1160 274
rect 1028 156 1101 205
rect 1088 65 1101 156
rect 1147 65 1160 205
rect 1272 245 1285 291
rect 1331 245 1360 291
rect 1272 146 1360 245
rect 1480 205 1584 304
rect 1480 159 1509 205
rect 1555 159 1584 205
rect 1480 146 1584 159
rect 1704 291 1792 304
rect 1704 245 1733 291
rect 1779 245 1792 291
rect 1704 146 1792 245
rect 1880 285 1968 344
rect 1880 239 1893 285
rect 1939 239 1968 285
rect 1880 226 1968 239
rect 2088 331 2192 344
rect 2088 285 2117 331
rect 2163 285 2192 331
rect 2088 226 2192 285
rect 2312 226 2360 344
rect 2480 226 2560 344
rect 2680 285 2828 344
rect 2680 239 2709 285
rect 2755 239 2828 285
rect 2680 226 2828 239
rect 2948 226 3032 344
rect 3152 331 3256 344
rect 3152 285 3181 331
rect 3227 285 3256 331
rect 3152 226 3256 285
rect 3376 331 3480 344
rect 3376 285 3405 331
rect 3451 285 3480 331
rect 3376 226 3480 285
rect 3600 331 3688 344
rect 3600 285 3629 331
rect 3675 285 3688 331
rect 3600 226 3688 285
rect 4460 275 4540 333
rect 3800 262 3888 275
rect 1088 52 1160 65
rect 3800 216 3813 262
rect 3859 216 3888 262
rect 3800 157 3888 216
rect 4008 157 4056 275
rect 4176 216 4280 275
rect 4176 170 4205 216
rect 4251 170 4280 216
rect 4176 157 4280 170
rect 4400 157 4540 275
rect 4460 69 4540 157
rect 4660 320 4748 333
rect 4660 180 4689 320
rect 4735 180 4748 320
rect 4660 69 4748 180
rect 4820 309 4908 333
rect 4820 169 4833 309
rect 4879 169 4908 309
rect 4820 69 4908 169
rect 5028 309 5132 333
rect 5028 169 5057 309
rect 5103 169 5132 309
rect 5028 69 5132 169
rect 5252 309 5340 333
rect 5252 169 5281 309
rect 5327 169 5340 309
rect 5252 69 5340 169
<< mvpdiff >>
rect 66 805 154 852
rect 66 665 79 805
rect 125 665 154 805
rect 66 652 154 665
rect 254 805 358 852
rect 254 665 283 805
rect 329 665 358 805
rect 254 652 358 665
rect 458 652 506 852
rect 606 805 740 852
rect 606 665 665 805
rect 711 665 740 805
rect 606 652 740 665
rect 840 652 888 852
rect 988 839 1076 852
rect 988 699 1017 839
rect 1063 699 1076 839
rect 988 652 1076 699
rect 1232 676 1320 884
rect 1232 630 1245 676
rect 1291 630 1320 676
rect 1232 608 1320 630
rect 1420 871 1524 884
rect 1420 825 1449 871
rect 1495 825 1524 871
rect 1420 608 1524 825
rect 1624 676 1712 884
rect 2440 959 2512 972
rect 2440 913 2453 959
rect 2499 913 2512 959
rect 3068 959 3140 972
rect 2440 900 2512 913
rect 3068 913 3081 959
rect 3127 913 3140 959
rect 3068 905 3140 913
rect 2440 820 2500 900
rect 2440 788 2560 820
rect 1624 630 1653 676
rect 1699 630 1712 676
rect 1624 608 1712 630
rect 1784 768 1872 788
rect 1784 628 1797 768
rect 1843 628 1872 768
rect 1784 588 1872 628
rect 1972 775 2076 788
rect 1972 635 2001 775
rect 2047 635 2076 775
rect 1972 588 2076 635
rect 2176 711 2280 788
rect 2176 665 2205 711
rect 2251 665 2280 711
rect 2176 588 2280 665
rect 2380 620 2560 788
rect 2660 711 2748 820
rect 2660 665 2689 711
rect 2735 665 2748 711
rect 2820 764 2908 905
rect 2820 718 2833 764
rect 2879 718 2908 764
rect 2820 705 2908 718
rect 3008 900 3140 905
rect 3008 788 3128 900
rect 4320 917 4408 939
rect 4320 871 4333 917
rect 4379 871 4408 917
rect 4320 852 4408 871
rect 3866 839 3954 852
rect 3866 793 3879 839
rect 3925 793 3954 839
rect 3008 705 3188 788
rect 2660 620 2748 665
rect 2380 588 2460 620
rect 3108 588 3188 705
rect 3288 764 3392 788
rect 3288 624 3317 764
rect 3363 624 3392 764
rect 3288 588 3392 624
rect 3492 742 3596 788
rect 3492 602 3521 742
rect 3567 602 3596 742
rect 3492 588 3596 602
rect 3696 650 3784 788
rect 3866 652 3954 793
rect 4054 711 4158 852
rect 4054 665 4083 711
rect 4129 665 4158 711
rect 4054 652 4158 665
rect 4258 652 4408 852
rect 3696 604 3725 650
rect 3771 604 3784 650
rect 3696 588 3784 604
rect 4328 573 4408 652
rect 4508 711 4616 939
rect 4508 665 4537 711
rect 4583 665 4616 711
rect 4508 573 4616 665
rect 4716 805 4900 939
rect 4716 665 4745 805
rect 4791 665 4900 805
rect 4716 573 4900 665
rect 5000 805 5104 939
rect 5000 665 5029 805
rect 5075 665 5104 805
rect 5000 573 5104 665
rect 5204 805 5292 939
rect 5204 665 5233 805
rect 5279 665 5292 805
rect 5204 573 5292 665
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1101 65 1147 205
rect 1285 245 1331 291
rect 1509 159 1555 205
rect 1733 245 1779 291
rect 1893 239 1939 285
rect 2117 285 2163 331
rect 2709 239 2755 285
rect 3181 285 3227 331
rect 3405 285 3451 331
rect 3629 285 3675 331
rect 3813 216 3859 262
rect 4205 170 4251 216
rect 4689 180 4735 320
rect 4833 169 4879 309
rect 5057 169 5103 309
rect 5281 169 5327 309
<< mvpdiffc >>
rect 79 665 125 805
rect 283 665 329 805
rect 665 665 711 805
rect 1017 699 1063 839
rect 1245 630 1291 676
rect 1449 825 1495 871
rect 2453 913 2499 959
rect 3081 913 3127 959
rect 1653 630 1699 676
rect 1797 628 1843 768
rect 2001 635 2047 775
rect 2205 665 2251 711
rect 2689 665 2735 711
rect 2833 718 2879 764
rect 4333 871 4379 917
rect 3879 793 3925 839
rect 3317 624 3363 764
rect 3521 602 3567 742
rect 4083 665 4129 711
rect 3725 604 3771 650
rect 4537 665 4583 711
rect 4745 665 4791 805
rect 5029 665 5075 805
rect 5233 665 5279 805
<< polysilicon >>
rect 154 944 988 984
rect 154 852 254 944
rect 358 852 458 896
rect 506 852 606 896
rect 740 852 840 896
rect 888 852 988 944
rect 1524 944 2176 984
rect 1320 884 1420 928
rect 1524 884 1624 944
rect 154 608 254 652
rect 154 473 244 608
rect 124 460 244 473
rect 124 414 137 460
rect 183 414 244 460
rect 124 274 244 414
rect 358 458 458 652
rect 358 412 371 458
rect 417 412 458 458
rect 358 318 458 412
rect 506 460 606 652
rect 506 414 519 460
rect 565 414 606 460
rect 506 401 606 414
rect 740 458 840 652
rect 888 608 988 652
rect 2076 867 2176 944
rect 1872 788 1972 832
rect 2076 821 2117 867
rect 2163 821 2176 867
rect 2908 905 3008 949
rect 2076 788 2176 821
rect 2280 788 2380 832
rect 2560 820 2660 864
rect 1320 542 1420 608
rect 1524 564 1624 608
rect 3248 944 4054 984
rect 3248 832 3288 944
rect 3188 788 3288 832
rect 3392 867 3492 880
rect 3392 821 3405 867
rect 3451 821 3492 867
rect 3954 852 4054 944
rect 4408 939 4508 983
rect 4616 939 4716 983
rect 4900 939 5000 983
rect 5104 939 5204 983
rect 4158 852 4258 896
rect 3392 788 3492 821
rect 3596 788 3696 832
rect 2908 661 3008 705
rect 1320 496 1333 542
rect 1379 496 1420 542
rect 1320 483 1420 496
rect 740 412 753 458
rect 799 412 840 458
rect 740 318 840 412
rect 908 460 1028 473
rect 908 414 921 460
rect 967 414 1028 460
rect 348 274 468 318
rect 516 274 636 318
rect 740 274 860 318
rect 908 274 1028 414
rect 1360 348 1420 483
rect 1584 424 1624 564
rect 1872 502 1972 588
rect 2076 544 2176 588
rect 2280 544 2380 588
rect 1872 456 1885 502
rect 1931 476 1972 502
rect 2340 504 2380 544
rect 2340 491 2480 504
rect 1931 460 2292 476
rect 1931 456 2233 460
rect 1872 436 2233 456
rect 1584 411 1704 424
rect 1584 365 1597 411
rect 1643 365 1704 411
rect 2192 414 2233 436
rect 2279 414 2292 460
rect 2340 445 2401 491
rect 2447 445 2480 491
rect 2340 434 2480 445
rect 2192 388 2292 414
rect 1360 304 1480 348
rect 1584 304 1704 365
rect 1968 344 2088 388
rect 2192 344 2312 388
rect 2360 344 2480 434
rect 2560 388 2660 620
rect 2908 618 2948 661
rect 2828 605 2948 618
rect 2828 559 2861 605
rect 2907 559 2948 605
rect 2560 344 2680 388
rect 2828 344 2948 559
rect 3188 544 3288 588
rect 3188 499 3228 544
rect 3032 427 3228 499
rect 3392 528 3492 588
rect 3596 544 3696 588
rect 3392 457 3520 528
rect 3032 344 3152 427
rect 3480 388 3520 457
rect 3656 476 3696 544
rect 3656 460 3807 476
rect 3954 470 4054 652
rect 4158 471 4258 652
rect 4408 513 4508 573
rect 3656 414 3721 460
rect 3767 414 3807 460
rect 3656 404 3807 414
rect 3707 401 3807 404
rect 3888 460 4054 470
rect 3888 414 3962 460
rect 4008 414 4054 460
rect 3888 401 4054 414
rect 4136 460 4258 471
rect 4136 414 4183 460
rect 4229 414 4258 460
rect 4136 401 4258 414
rect 4328 460 4508 513
rect 4328 414 4341 460
rect 4387 441 4508 460
rect 4616 540 4716 573
rect 4616 494 4629 540
rect 4675 494 4716 540
rect 4900 529 5000 573
rect 4616 481 4716 494
rect 4908 513 5000 529
rect 5104 513 5204 573
rect 4387 414 4400 441
rect 3256 344 3376 388
rect 3480 344 3600 388
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 124 24 636 64
rect 3888 275 4008 401
rect 4136 319 4176 401
rect 4328 319 4400 414
rect 4616 377 4660 481
rect 4540 333 4660 377
rect 4908 460 5204 513
rect 4908 414 4921 460
rect 4967 441 5204 460
rect 4967 414 5028 441
rect 4908 333 5028 414
rect 5132 377 5204 441
rect 5132 333 5252 377
rect 4056 275 4176 319
rect 4280 275 4400 319
rect 1360 102 1480 146
rect 1584 64 1704 146
rect 1968 64 2088 226
rect 2192 182 2312 226
rect 2360 182 2480 226
rect 1584 24 2088 64
rect 2560 64 2680 226
rect 2828 182 2948 226
rect 3032 182 3152 226
rect 3256 193 3376 226
rect 3256 147 3269 193
rect 3315 147 3376 193
rect 3480 182 3600 226
rect 3256 134 3376 147
rect 3888 113 4008 157
rect 4056 113 4176 157
rect 4280 64 4400 157
rect 2560 24 4400 64
rect 4540 25 4660 69
rect 4908 25 5028 69
rect 5132 25 5252 69
<< polycontact >>
rect 137 414 183 460
rect 371 412 417 458
rect 519 414 565 460
rect 2117 821 2163 867
rect 3405 821 3451 867
rect 1333 496 1379 542
rect 753 412 799 458
rect 921 414 967 460
rect 1885 456 1931 502
rect 1597 365 1643 411
rect 2233 414 2279 460
rect 2401 445 2447 491
rect 2861 559 2907 605
rect 3721 414 3767 460
rect 3962 414 4008 460
rect 4183 414 4229 460
rect 4341 414 4387 460
rect 4629 494 4675 540
rect 4921 414 4967 460
rect 3269 147 3315 193
<< metal1 >>
rect 0 959 5376 1098
rect 0 918 2453 959
rect 79 805 125 816
rect 79 561 125 665
rect 283 805 329 918
rect 1017 839 1063 918
rect 283 654 329 665
rect 665 805 711 816
rect 1438 871 1506 918
rect 2442 913 2453 918
rect 2499 918 3081 959
rect 2499 913 2510 918
rect 3070 913 3081 918
rect 3127 918 5376 959
rect 3127 913 3138 918
rect 1438 825 1449 871
rect 1495 825 1506 871
rect 2106 821 2117 867
rect 2163 821 3405 867
rect 3451 821 3462 867
rect 3879 839 3925 918
rect 4333 917 4379 918
rect 4333 860 4379 871
rect 1017 688 1063 699
rect 1109 768 1843 779
rect 1109 733 1797 768
rect 665 642 711 665
rect 1109 642 1155 733
rect 665 596 1155 642
rect 1245 676 1518 687
rect 1291 630 1518 676
rect 1245 619 1518 630
rect 79 550 549 561
rect 79 515 967 550
rect 519 504 967 515
rect 30 414 137 460
rect 183 414 194 460
rect 30 354 194 414
rect 254 458 418 469
rect 254 412 371 458
rect 417 412 418 458
rect 254 354 418 412
rect 519 460 565 504
rect 921 460 967 504
rect 1262 496 1333 542
rect 1379 496 1426 542
rect 1262 466 1426 496
rect 519 308 565 414
rect 702 412 753 458
rect 799 412 866 458
rect 702 354 866 412
rect 921 403 967 414
rect 1472 422 1518 619
rect 1653 676 1699 687
rect 1653 513 1699 630
rect 1797 617 1843 628
rect 2001 775 2047 786
rect 3879 782 3925 793
rect 2833 764 3363 775
rect 2205 711 2735 722
rect 2251 665 2689 711
rect 2879 729 3317 764
rect 2879 718 3227 729
rect 2833 707 3227 718
rect 2205 654 2735 665
rect 2001 594 2047 635
rect 2861 605 2907 616
rect 2001 559 2861 594
rect 2001 548 2907 559
rect 1653 502 1931 513
rect 1653 467 1885 502
rect 1733 456 1885 467
rect 1733 445 1931 456
rect 1472 411 1643 422
rect 1472 400 1597 411
rect 1285 365 1597 400
rect 1285 354 1643 365
rect 49 262 565 308
rect 665 262 1239 308
rect 49 215 95 262
rect 665 215 711 262
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 665 158 711 169
rect 1101 205 1147 216
rect 0 65 1101 90
rect 1193 188 1239 262
rect 1285 291 1331 354
rect 1285 234 1331 245
rect 1377 262 1687 308
rect 1377 188 1423 262
rect 1193 142 1423 188
rect 1509 205 1555 216
rect 1509 90 1555 159
rect 1641 188 1687 262
rect 1733 291 1779 445
rect 2117 331 2163 548
rect 3181 502 3227 707
rect 3971 768 4675 814
rect 3317 613 3363 624
rect 3521 742 3843 753
rect 3567 736 3843 742
rect 3971 736 4017 768
rect 3567 707 4017 736
rect 3807 690 4017 707
rect 4080 711 4129 722
rect 4080 665 4083 711
rect 3521 594 3567 602
rect 2401 491 3227 502
rect 2233 460 2279 471
rect 2447 445 3227 491
rect 2401 434 3227 445
rect 2233 388 2279 414
rect 2233 342 3135 388
rect 1733 234 1779 245
rect 1893 285 1939 296
rect 2117 274 2163 285
rect 2709 285 2755 296
rect 1893 188 1939 239
rect 1641 142 1939 188
rect 2709 90 2755 239
rect 3089 204 3135 342
rect 3181 331 3227 434
rect 3181 274 3227 285
rect 3405 548 3567 594
rect 3725 650 3771 661
rect 3725 563 3771 604
rect 4080 654 4129 665
rect 4537 711 4583 722
rect 3405 331 3451 548
rect 3405 274 3451 285
rect 3629 517 3859 563
rect 3629 331 3675 517
rect 3629 274 3675 285
rect 3721 460 3767 471
rect 3721 204 3767 414
rect 3813 308 3859 517
rect 3950 460 4008 542
rect 3950 414 3962 460
rect 3950 354 4008 414
rect 4080 308 4126 654
rect 4286 471 4338 542
rect 4286 460 4387 471
rect 3813 262 4126 308
rect 4172 414 4183 460
rect 4229 414 4240 460
rect 4172 308 4240 414
rect 4286 414 4341 460
rect 4286 403 4387 414
rect 4286 354 4338 403
rect 4537 308 4583 665
rect 4629 540 4675 768
rect 4745 805 4791 918
rect 4745 654 4791 665
rect 5029 805 5075 816
rect 4629 483 4675 494
rect 5029 542 5075 665
rect 5233 805 5279 918
rect 5233 654 5279 665
rect 4921 460 4967 471
rect 4689 414 4921 439
rect 4689 393 4967 414
rect 4689 320 4735 393
rect 4172 262 4689 308
rect 3813 205 3859 216
rect 3089 193 3767 204
rect 3089 147 3269 193
rect 3315 147 3767 193
rect 3089 136 3767 147
rect 4194 170 4205 216
rect 4251 170 4262 216
rect 4194 90 4262 170
rect 4689 169 4735 180
rect 4833 309 4879 320
rect 4833 90 4879 169
rect 5029 309 5122 542
rect 5029 169 5057 309
rect 5103 169 5122 309
rect 5029 158 5122 169
rect 5281 309 5327 320
rect 5281 90 5327 169
rect 1147 65 5376 90
rect 0 -90 5376 65
<< labels >>
flabel metal1 s 1262 466 1426 542 0 FreeSans 200 0 0 0 CLK
port 6 nsew clock input
flabel metal1 s 702 354 866 458 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 5029 542 5075 816 0 FreeSans 200 0 0 0 Q
port 7 nsew default output
flabel metal1 s 4286 471 4338 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 30 354 194 460 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 3950 354 4008 542 0 FreeSans 200 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 254 354 418 469 0 FreeSans 200 0 0 0 SI
port 5 nsew default input
flabel metal1 s 0 918 5376 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 5281 296 5327 320 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 4286 403 4387 471 1 RN
port 2 nsew default input
rlabel metal1 s 4286 354 4338 403 1 RN
port 2 nsew default input
rlabel metal1 s 5029 158 5122 542 1 Q
port 7 nsew default output
rlabel metal1 s 5233 913 5279 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 913 4791 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4333 913 4379 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3879 913 3925 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3070 913 3138 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2442 913 2510 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1438 913 1506 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1017 913 1063 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 913 329 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5233 860 5279 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 860 4791 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4333 860 4379 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3879 860 3925 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1438 860 1506 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1017 860 1063 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 860 329 913 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5233 825 5279 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 825 4791 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3879 825 3925 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1438 825 1506 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1017 825 1063 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 825 329 860 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5233 782 5279 825 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 782 4791 825 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3879 782 3925 825 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1017 782 1063 825 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 782 329 825 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5233 688 5279 782 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 688 4791 782 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1017 688 1063 782 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 688 329 782 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5233 654 5279 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4745 654 4791 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 283 654 329 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4833 296 4879 320 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5281 216 5327 296 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 216 4879 296 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2709 216 2755 296 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5281 215 5327 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 215 4879 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4194 215 4262 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2709 215 2755 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1509 215 1555 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1101 215 1147 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5281 90 5327 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 90 4879 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4194 90 4262 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2709 90 2755 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1509 90 1555 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1101 90 1147 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5376 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5376 1008
string GDS_END 384052
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 371716
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
