magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 1800 1620
<< nmos >>
rect 200 190 260 360
rect 400 190 460 360
rect 540 190 600 360
rect 710 190 770 360
rect 850 190 910 360
rect 1050 190 1110 360
rect 1370 190 1430 360
rect 1540 190 1600 360
<< pmos >>
rect 200 1090 260 1430
rect 370 1090 430 1430
rect 540 1090 600 1430
rect 710 1090 770 1430
rect 880 1090 940 1430
rect 1050 1090 1110 1430
rect 1370 1090 1430 1430
rect 1540 1090 1600 1430
<< ndiff >>
rect 100 298 200 360
rect 100 252 122 298
rect 168 252 200 298
rect 100 190 200 252
rect 260 298 400 360
rect 260 252 307 298
rect 353 252 400 298
rect 260 190 400 252
rect 460 190 540 360
rect 600 298 710 360
rect 600 252 632 298
rect 678 252 710 298
rect 600 190 710 252
rect 770 190 850 360
rect 910 298 1050 360
rect 910 252 957 298
rect 1003 252 1050 298
rect 910 190 1050 252
rect 1110 298 1210 360
rect 1110 252 1142 298
rect 1188 252 1210 298
rect 1110 190 1210 252
rect 1270 298 1370 360
rect 1270 252 1292 298
rect 1338 252 1370 298
rect 1270 190 1370 252
rect 1430 298 1540 360
rect 1430 252 1462 298
rect 1508 252 1540 298
rect 1430 190 1540 252
rect 1600 298 1700 360
rect 1600 252 1632 298
rect 1678 252 1700 298
rect 1600 190 1700 252
<< pdiff >>
rect 100 1377 200 1430
rect 100 1143 122 1377
rect 168 1143 200 1377
rect 100 1090 200 1143
rect 260 1410 370 1430
rect 260 1270 292 1410
rect 338 1270 370 1410
rect 260 1090 370 1270
rect 430 1090 540 1430
rect 600 1377 710 1430
rect 600 1143 632 1377
rect 678 1143 710 1377
rect 600 1090 710 1143
rect 770 1090 880 1430
rect 940 1377 1050 1430
rect 940 1143 972 1377
rect 1018 1143 1050 1377
rect 940 1090 1050 1143
rect 1110 1377 1210 1430
rect 1110 1143 1142 1377
rect 1188 1143 1210 1377
rect 1110 1090 1210 1143
rect 1270 1377 1370 1430
rect 1270 1143 1292 1377
rect 1338 1143 1370 1377
rect 1270 1090 1370 1143
rect 1430 1377 1540 1430
rect 1430 1143 1462 1377
rect 1508 1143 1540 1377
rect 1430 1090 1540 1143
rect 1600 1377 1700 1430
rect 1600 1143 1632 1377
rect 1678 1143 1700 1377
rect 1600 1090 1700 1143
<< ndiffc >>
rect 122 252 168 298
rect 307 252 353 298
rect 632 252 678 298
rect 957 252 1003 298
rect 1142 252 1188 298
rect 1292 252 1338 298
rect 1462 252 1508 298
rect 1632 252 1678 298
<< pdiffc >>
rect 122 1143 168 1377
rect 292 1270 338 1410
rect 632 1143 678 1377
rect 972 1143 1018 1377
rect 1142 1143 1188 1377
rect 1292 1143 1338 1377
rect 1462 1143 1508 1377
rect 1632 1143 1678 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 340 98 430 120
rect 340 52 362 98
rect 408 52 430 98
rect 340 30 430 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1060 98 1150 120
rect 1060 52 1082 98
rect 1128 52 1150 98
rect 1060 30 1150 52
rect 1290 98 1390 120
rect 1290 52 1312 98
rect 1358 52 1390 98
rect 1290 30 1390 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 340 1568 430 1590
rect 340 1522 362 1568
rect 408 1522 430 1568
rect 340 1500 430 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1060 1568 1150 1590
rect 1060 1522 1082 1568
rect 1128 1522 1150 1568
rect 1060 1500 1150 1522
rect 1300 1568 1390 1590
rect 1300 1522 1322 1568
rect 1368 1522 1390 1568
rect 1300 1500 1390 1522
rect 1540 1568 1630 1590
rect 1540 1522 1562 1568
rect 1608 1522 1630 1568
rect 1540 1500 1630 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 362 52 408 98
rect 592 52 638 98
rect 832 52 878 98
rect 1082 52 1128 98
rect 1312 52 1358 98
rect 1552 52 1598 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 362 1522 408 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1082 1522 1128 1568
rect 1322 1522 1368 1568
rect 1562 1522 1608 1568
<< polysilicon >>
rect 200 1430 260 1480
rect 370 1430 430 1480
rect 540 1430 600 1480
rect 710 1430 770 1480
rect 880 1430 940 1480
rect 1050 1430 1110 1480
rect 1370 1430 1430 1480
rect 1540 1430 1600 1480
rect 200 910 260 1090
rect 370 910 430 1090
rect 540 1020 600 1090
rect 520 993 620 1020
rect 520 947 547 993
rect 593 947 620 993
rect 520 920 620 947
rect 710 910 770 1090
rect 200 883 320 910
rect 200 837 237 883
rect 283 837 320 883
rect 200 810 320 837
rect 370 883 470 910
rect 370 837 397 883
rect 443 837 470 883
rect 370 810 470 837
rect 690 883 790 910
rect 690 837 717 883
rect 763 837 790 883
rect 690 810 790 837
rect 200 360 260 810
rect 370 450 430 810
rect 710 700 770 810
rect 540 640 770 700
rect 880 780 940 1090
rect 1050 910 1110 1090
rect 1040 883 1140 910
rect 1040 837 1067 883
rect 1113 837 1140 883
rect 1040 810 1140 837
rect 880 753 1000 780
rect 880 707 927 753
rect 973 707 1000 753
rect 880 680 1000 707
rect 370 410 460 450
rect 400 360 460 410
rect 540 360 600 640
rect 690 563 790 590
rect 690 517 717 563
rect 763 517 790 563
rect 690 490 790 517
rect 710 360 770 490
rect 880 450 940 680
rect 850 410 940 450
rect 850 360 910 410
rect 1050 360 1110 810
rect 1370 780 1430 1090
rect 1540 910 1600 1090
rect 1480 883 1600 910
rect 1480 837 1507 883
rect 1553 837 1600 883
rect 1480 810 1600 837
rect 1350 758 1440 780
rect 1350 712 1372 758
rect 1418 712 1440 758
rect 1350 690 1440 712
rect 1370 360 1430 690
rect 1540 360 1600 810
rect 200 140 260 190
rect 400 140 460 190
rect 540 140 600 190
rect 710 140 770 190
rect 850 140 910 190
rect 1050 140 1110 190
rect 1370 140 1430 190
rect 1540 140 1600 190
<< polycontact >>
rect 547 947 593 993
rect 237 837 283 883
rect 397 837 443 883
rect 717 837 763 883
rect 1067 837 1113 883
rect 927 707 973 753
rect 717 517 763 563
rect 1507 837 1553 883
rect 1372 712 1418 758
<< metal1 >>
rect -1550 1568 1800 1620
rect -1550 1522 112 1568
rect 158 1566 362 1568
rect -1550 1514 114 1522
rect 166 1514 354 1566
rect 408 1522 592 1568
rect 638 1566 832 1568
rect 878 1566 1082 1568
rect 1128 1566 1322 1568
rect 1368 1566 1562 1568
rect 646 1522 832 1566
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1566
rect 1128 1522 1314 1566
rect 1368 1522 1554 1566
rect 1608 1522 1800 1568
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1800 1522
rect -1550 1500 1800 1514
rect -1260 1250 -1210 1500
rect -580 1090 -530 1500
rect -90 1090 -40 1500
rect 80 1377 170 1430
rect 80 1143 122 1377
rect 168 1143 170 1377
rect 290 1410 340 1500
rect 290 1270 292 1410
rect 338 1270 340 1410
rect 290 1250 340 1270
rect 630 1377 680 1430
rect 80 1020 170 1143
rect 630 1143 632 1377
rect 678 1143 680 1377
rect 630 1140 680 1143
rect 230 1090 680 1140
rect 970 1377 1020 1500
rect 970 1143 972 1377
rect 1018 1143 1020 1377
rect 970 1090 1020 1143
rect 1140 1377 1190 1430
rect 1140 1143 1142 1377
rect 1188 1143 1190 1377
rect 1140 1100 1190 1143
rect 1290 1377 1340 1430
rect 1290 1143 1292 1377
rect 1338 1143 1340 1377
rect 80 960 180 1020
rect -1180 830 -1080 890
rect -860 830 -760 890
rect -510 830 -410 890
rect 80 760 170 960
rect 230 890 280 1090
rect 1140 1050 1240 1100
rect 520 993 620 1000
rect 520 947 547 993
rect 593 947 620 993
rect 520 940 620 947
rect 220 883 310 890
rect 220 837 237 883
rect 283 837 310 883
rect 220 830 310 837
rect 370 886 470 890
rect 370 834 394 886
rect 446 834 470 886
rect 370 830 470 834
rect 70 756 170 760
rect 70 704 94 756
rect 146 704 170 756
rect 70 700 170 704
rect -1260 120 -1180 360
rect -610 120 -530 360
rect -90 120 -40 360
rect 80 298 170 700
rect 230 460 280 830
rect 540 570 600 940
rect 690 886 790 890
rect 690 834 714 886
rect 766 834 790 886
rect 690 830 790 834
rect 1040 886 1140 890
rect 1040 834 1064 886
rect 1116 834 1140 886
rect 1040 830 1140 834
rect 900 756 1000 760
rect 900 704 924 756
rect 976 704 1000 756
rect 900 700 1000 704
rect 1190 570 1240 1050
rect 1290 1060 1340 1143
rect 1460 1377 1510 1500
rect 1460 1143 1462 1377
rect 1508 1143 1510 1377
rect 1460 1090 1510 1143
rect 1630 1377 1680 1430
rect 1630 1143 1632 1377
rect 1678 1143 1680 1377
rect 1290 1020 1370 1060
rect 1630 1030 1680 1143
rect 1630 1020 1710 1030
rect 1290 1016 1390 1020
rect 1290 964 1314 1016
rect 1366 1010 1390 1016
rect 1630 1016 1730 1020
rect 1366 964 1560 1010
rect 1290 960 1560 964
rect 1290 950 1370 960
rect 1500 883 1560 960
rect 1500 837 1507 883
rect 1553 837 1560 883
rect 1350 758 1450 760
rect 1350 712 1372 758
rect 1418 756 1450 758
rect 1350 704 1374 712
rect 1426 704 1450 756
rect 1350 700 1450 704
rect 540 563 1240 570
rect 540 517 717 563
rect 763 517 1240 563
rect 540 510 1240 517
rect 230 410 680 460
rect 1190 440 1240 510
rect 1500 460 1560 837
rect 80 252 122 298
rect 168 252 170 298
rect 80 190 170 252
rect 290 298 370 360
rect 290 252 307 298
rect 353 252 370 298
rect 290 120 370 252
rect 630 298 680 410
rect 1140 390 1240 440
rect 1290 410 1560 460
rect 1630 964 1654 1016
rect 1706 964 1730 1016
rect 1630 960 1730 964
rect 1630 950 1710 960
rect 630 252 632 298
rect 678 252 680 298
rect 630 190 680 252
rect 940 298 1020 360
rect 940 252 957 298
rect 1003 252 1020 298
rect 940 120 1020 252
rect 1140 298 1190 390
rect 1140 252 1142 298
rect 1188 252 1190 298
rect 1140 190 1190 252
rect 1290 298 1340 410
rect 1290 252 1292 298
rect 1338 252 1340 298
rect 1290 190 1340 252
rect 1460 298 1510 360
rect 1460 252 1462 298
rect 1508 252 1510 298
rect 1460 120 1510 252
rect 1630 298 1680 950
rect 1630 252 1632 298
rect 1678 252 1680 298
rect 1630 190 1680 252
rect -1550 106 1800 120
rect -1550 98 114 106
rect -1550 52 112 98
rect 166 54 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 158 52 362 54
rect 408 52 592 98
rect 646 54 832 98
rect 886 54 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 638 52 832 54
rect 878 52 1082 54
rect 1128 52 1312 98
rect 1366 54 1552 98
rect 1606 54 1800 106
rect 1358 52 1552 54
rect 1598 52 1800 54
rect -1550 0 1800 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 114 1514 166 1522
rect 354 1522 362 1566
rect 362 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1522 1082 1566
rect 1082 1522 1126 1566
rect 1314 1522 1322 1566
rect 1322 1522 1366 1566
rect 1554 1522 1562 1566
rect 1562 1522 1606 1566
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 394 883 446 886
rect 394 837 397 883
rect 397 837 443 883
rect 443 837 446 883
rect 394 834 446 837
rect 94 704 146 756
rect 714 883 766 886
rect 714 837 717 883
rect 717 837 763 883
rect 763 837 766 883
rect 714 834 766 837
rect 1064 883 1116 886
rect 1064 837 1067 883
rect 1067 837 1113 883
rect 1113 837 1116 883
rect 1064 834 1116 837
rect 924 753 976 756
rect 924 707 927 753
rect 927 707 973 753
rect 973 707 976 753
rect 924 704 976 707
rect 1314 964 1366 1016
rect 1374 712 1418 756
rect 1418 712 1426 756
rect 1374 704 1426 712
rect 1654 964 1706 1016
rect 114 98 166 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 354 54 362 98
rect 362 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1074 54 1082 98
rect 1082 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
<< metal2 >>
rect -1450 1570 -1370 1580
rect -1210 1570 -1130 1580
rect -970 1570 -890 1580
rect -730 1570 -650 1580
rect -490 1570 -410 1580
rect -250 1570 -170 1580
rect -10 1570 70 1580
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect -1460 1510 -1360 1570
rect -1220 1510 -1120 1570
rect -980 1510 -880 1570
rect -740 1510 -640 1570
rect -500 1510 -400 1570
rect -260 1510 -160 1570
rect -20 1510 80 1570
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1510 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1510 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1510 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1510 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1510 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1510 1390 1514
rect 1530 1566 1630 1570
rect 1530 1514 1554 1566
rect 1606 1514 1630 1566
rect 1530 1510 1630 1514
rect -1450 1500 -1370 1510
rect -1210 1500 -1130 1510
rect -970 1500 -890 1510
rect -730 1500 -650 1510
rect -490 1500 -410 1510
rect -250 1500 -170 1510
rect -10 1500 70 1510
rect 100 1500 180 1510
rect 340 1500 420 1510
rect 580 1500 660 1510
rect 820 1500 900 1510
rect 1060 1500 1140 1510
rect 1300 1500 1380 1510
rect 1540 1500 1620 1510
rect 90 1020 170 1030
rect 1300 1020 1380 1030
rect 1640 1020 1720 1030
rect 80 960 180 1020
rect 1290 1016 1390 1020
rect 1290 964 1314 1016
rect 1366 964 1390 1016
rect 1290 960 1390 964
rect 1630 1016 1730 1020
rect 1630 964 1654 1016
rect 1706 964 1730 1016
rect 1630 960 1730 964
rect 90 950 170 960
rect 1300 950 1380 960
rect 1640 950 1720 960
rect -1180 820 -1080 900
rect -850 890 -770 900
rect -510 890 -410 900
rect -860 830 -410 890
rect -850 820 -770 830
rect -510 820 -410 830
rect 370 886 470 900
rect 700 890 780 900
rect 1040 890 1140 900
rect 370 834 394 886
rect 446 834 470 886
rect 370 820 470 834
rect 690 886 1140 890
rect 690 834 714 886
rect 766 834 1064 886
rect 1116 834 1140 886
rect 690 830 1140 834
rect 700 820 780 830
rect 1040 820 1140 830
rect 70 760 170 770
rect 910 760 990 770
rect 1350 760 1450 770
rect 70 756 1450 760
rect 70 704 94 756
rect 146 704 924 756
rect 976 704 1374 756
rect 1426 704 1450 756
rect 70 700 1450 704
rect 70 690 170 700
rect 910 690 990 700
rect 1350 690 1450 700
rect -1450 110 -1370 120
rect -1210 110 -1130 120
rect -970 110 -890 120
rect -730 110 -650 120
rect -490 110 -410 120
rect -250 110 -170 120
rect -10 110 70 120
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect -1460 50 -1360 110
rect -1220 50 -1120 110
rect -980 50 -880 110
rect -740 50 -640 110
rect -500 50 -400 110
rect -260 50 -160 110
rect -20 50 80 110
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect -1450 40 -1370 50
rect -1210 40 -1130 50
rect -970 40 -890 50
rect -730 40 -650 50
rect -490 40 -410 50
rect -250 40 -170 50
rect -10 40 70 50
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
<< labels >>
rlabel metal1 s -1260 1250 -1210 1620 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s -1260 0 -1180 360 4 VSS
port 9 nsew ground bidirectional
rlabel metal1 s -1180 830 -1080 890 4 D
port 1 nsew signal input
rlabel metal1 s -860 830 -760 890 4 CLK
port 2 nsew clock input
rlabel metal1 s 80 190 130 1430 4 Q
port 3 nsew signal output
rlabel metal1 s -510 830 -410 890 3 CLK
port 2 nsew clock input
rlabel metal2 s -850 820 -770 900 3 CLK
port 2 nsew clock input
rlabel metal2 s -860 830 -410 890 3 CLK
port 2 nsew clock input
rlabel metal2 s -510 820 -410 900 3 CLK
port 2 nsew clock input
rlabel metal2 s -1180 820 -1080 900 3 D
port 1 nsew signal input
rlabel metal1 s 80 950 160 1030 1 Q
port 3 nsew signal output
rlabel metal1 s 80 960 180 1020 1 Q
port 3 nsew signal output
rlabel metal2 s 90 950 170 1030 1 Q
port 3 nsew signal output
rlabel metal2 s 80 960 180 1020 1 Q
port 3 nsew signal output
rlabel metal1 s -580 1090 -530 1620 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s -90 1090 -40 1620 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s -1550 1500 250 1620 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -1450 1500 -1370 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -1460 1510 -1360 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -1210 1500 -1130 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -1220 1510 -1120 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -970 1500 -890 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -980 1510 -880 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -730 1500 -650 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -740 1510 -640 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -490 1500 -410 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -500 1510 -400 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -250 1500 -170 1580 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -260 1510 -160 1570 3 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -10 1500 70 1580 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s -20 1510 80 1570 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s -610 0 -530 360 3 VSS
port 9 nsew ground bidirectional
rlabel metal1 s -90 0 -40 360 3 VSS
port 9 nsew ground bidirectional
rlabel metal1 s -1550 0 250 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -1450 40 -1370 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -1460 50 -1360 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -1210 40 -1130 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -1220 50 -1120 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -970 40 -890 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -980 50 -880 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -730 40 -650 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -740 50 -640 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -490 40 -410 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -500 50 -400 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -250 40 -170 120 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -260 50 -160 110 3 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -10 40 70 120 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s -20 50 80 110 1 VSS
port 9 nsew ground bidirectional
<< properties >>
string FIXED_BBOX -1550 0 250 1620
string GDS_END 323918
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 306822
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
