magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal3 >>
rect 357 911 857 1215
use M2_M14310591302017_512x8m81  M2_M14310591302017_512x8m81_0
timestamp 1669390400
transform 1 0 607 0 1 993
box -236 -81 236 81
use M3_M24310591302016_512x8m81  M3_M24310591302016_512x8m81_0
timestamp 1669390400
transform 1 0 607 0 1 993
box -236 -81 236 81
<< properties >>
string GDS_END 2875778
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2875606
<< end >>
