magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 2662 1094
<< pwell >>
rect -86 -86 2662 453
<< mvnmos >>
rect 135 69 255 333
rect 359 69 479 333
rect 583 69 703 333
rect 1070 68 1190 332
rect 1372 68 1492 245
rect 1596 68 1716 245
rect 1856 68 1976 332
rect 2080 68 2200 332
rect 2304 68 2424 332
<< mvpmos >>
rect 145 573 245 933
rect 349 573 449 933
rect 654 573 754 933
rect 1080 573 1180 933
rect 1320 628 1420 925
rect 1524 628 1624 925
rect 1764 580 1864 940
rect 1968 580 2068 940
rect 2172 580 2272 940
<< mvndiff >>
rect 47 287 135 333
rect 47 147 60 287
rect 106 147 135 287
rect 47 69 135 147
rect 255 193 359 333
rect 255 147 284 193
rect 330 147 359 193
rect 255 69 359 147
rect 479 287 583 333
rect 479 147 508 287
rect 554 147 583 287
rect 479 69 583 147
rect 703 320 910 333
rect 703 274 851 320
rect 897 274 910 320
rect 703 69 910 274
rect 982 308 1070 332
rect 982 262 995 308
rect 1041 262 1070 308
rect 982 68 1070 262
rect 1190 245 1270 332
rect 1776 245 1856 332
rect 1190 124 1372 245
rect 1190 78 1258 124
rect 1304 78 1372 124
rect 1190 68 1372 78
rect 1492 227 1596 245
rect 1492 181 1521 227
rect 1567 181 1596 227
rect 1492 68 1596 181
rect 1716 221 1856 245
rect 1716 81 1745 221
rect 1791 81 1856 221
rect 1716 68 1856 81
rect 1976 309 2080 332
rect 1976 169 2005 309
rect 2051 169 2080 309
rect 1976 68 2080 169
rect 2200 193 2304 332
rect 2200 147 2229 193
rect 2275 147 2304 193
rect 2200 68 2304 147
rect 2424 319 2512 332
rect 2424 179 2453 319
rect 2499 179 2512 319
rect 2424 68 2512 179
rect 1250 65 1312 68
<< mvpdiff >>
rect 57 831 145 933
rect 57 691 70 831
rect 116 691 145 831
rect 57 573 145 691
rect 245 920 349 933
rect 245 780 274 920
rect 320 780 349 920
rect 245 573 349 780
rect 449 831 654 933
rect 449 691 579 831
rect 625 691 654 831
rect 449 573 654 691
rect 754 739 842 933
rect 754 599 783 739
rect 829 599 842 739
rect 754 573 842 599
rect 992 739 1080 933
rect 992 599 1005 739
rect 1051 599 1080 739
rect 992 573 1080 599
rect 1180 925 1260 933
rect 1684 925 1764 940
rect 1180 913 1320 925
rect 1180 867 1209 913
rect 1255 867 1320 913
rect 1180 628 1320 867
rect 1420 799 1524 925
rect 1420 659 1449 799
rect 1495 659 1524 799
rect 1420 628 1524 659
rect 1624 831 1764 925
rect 1624 691 1653 831
rect 1699 691 1764 831
rect 1624 628 1764 691
rect 1180 573 1260 628
rect 1684 580 1764 628
rect 1864 831 1968 940
rect 1864 691 1893 831
rect 1939 691 1968 831
rect 1864 580 1968 691
rect 2068 927 2172 940
rect 2068 787 2097 927
rect 2143 787 2172 927
rect 2068 580 2172 787
rect 2272 831 2360 940
rect 2272 691 2301 831
rect 2347 691 2360 831
rect 2272 580 2360 691
<< mvndiffc >>
rect 60 147 106 287
rect 284 147 330 193
rect 508 147 554 287
rect 851 274 897 320
rect 995 262 1041 308
rect 1258 78 1304 124
rect 1521 181 1567 227
rect 1745 81 1791 221
rect 2005 169 2051 309
rect 2229 147 2275 193
rect 2453 179 2499 319
<< mvpdiffc >>
rect 70 691 116 831
rect 274 780 320 920
rect 579 691 625 831
rect 783 599 829 739
rect 1005 599 1051 739
rect 1209 867 1255 913
rect 1449 659 1495 799
rect 1653 691 1699 831
rect 1893 691 1939 831
rect 2097 787 2143 927
rect 2301 691 2347 831
<< polysilicon >>
rect 145 933 245 977
rect 349 933 449 977
rect 654 933 754 977
rect 1080 933 1180 977
rect 1320 925 1420 969
rect 1524 925 1624 969
rect 1764 940 1864 984
rect 1968 940 2068 984
rect 2172 940 2272 984
rect 145 513 245 573
rect 349 513 449 573
rect 654 540 754 573
rect 145 473 567 513
rect 654 494 667 540
rect 713 494 754 540
rect 654 481 754 494
rect 145 425 255 473
rect 527 444 567 473
rect 135 412 255 425
rect 135 366 148 412
rect 194 366 255 412
rect 135 333 255 366
rect 359 412 479 425
rect 359 366 372 412
rect 418 366 479 412
rect 527 404 623 444
rect 1080 425 1180 573
rect 1320 452 1420 628
rect 359 333 479 366
rect 583 377 623 404
rect 1070 412 1180 425
rect 583 333 703 377
rect 1070 366 1083 412
rect 1129 376 1180 412
rect 1336 412 1420 452
rect 1129 366 1190 376
rect 1070 332 1190 366
rect 1336 366 1361 412
rect 1407 377 1420 412
rect 1524 584 1624 628
rect 1524 377 1623 584
rect 1764 547 1864 580
rect 1764 501 1791 547
rect 1837 520 1864 547
rect 1968 547 2068 580
rect 1968 520 1996 547
rect 1837 501 1996 520
rect 2042 520 2068 547
rect 2172 547 2272 580
rect 2172 520 2202 547
rect 2042 501 2202 520
rect 2248 501 2272 547
rect 1764 480 2272 501
rect 1856 412 2424 432
rect 1407 366 1716 377
rect 1336 353 1716 366
rect 135 25 255 69
rect 359 25 479 69
rect 583 25 703 69
rect 1372 305 1716 353
rect 1856 366 1889 412
rect 1935 392 2119 412
rect 1935 366 1976 392
rect 1856 332 1976 366
rect 2080 366 2119 392
rect 2165 392 2335 412
rect 2165 366 2200 392
rect 2080 332 2200 366
rect 2304 366 2335 392
rect 2381 366 2424 412
rect 2304 332 2424 366
rect 1372 245 1492 305
rect 1596 245 1716 305
rect 1070 24 1190 68
rect 1372 24 1492 68
rect 1596 24 1716 68
rect 1856 24 1976 68
rect 2080 24 2200 68
rect 2304 24 2424 68
<< polycontact >>
rect 667 494 713 540
rect 148 366 194 412
rect 372 366 418 412
rect 1083 366 1129 412
rect 1361 366 1407 412
rect 1791 501 1837 547
rect 1996 501 2042 547
rect 2202 501 2248 547
rect 1889 366 1935 412
rect 2119 366 2165 412
rect 2335 366 2381 412
<< metal1 >>
rect 0 927 2576 1098
rect 0 920 2097 927
rect 0 918 274 920
rect 70 831 116 842
rect 320 918 2097 920
rect 1209 913 1255 918
rect 1209 856 1255 867
rect 274 769 320 780
rect 579 831 1165 842
rect 70 634 116 691
rect 625 810 1165 831
rect 1653 831 1699 918
rect 625 799 1495 810
rect 625 796 1449 799
rect 579 680 625 691
rect 759 739 829 750
rect 70 588 713 634
rect 142 412 194 542
rect 667 540 713 588
rect 667 412 713 494
rect 142 366 148 412
rect 142 354 194 366
rect 240 366 372 412
rect 418 366 713 412
rect 759 599 783 739
rect 759 588 829 599
rect 240 308 286 366
rect 60 287 286 308
rect 759 298 805 588
rect 875 331 921 796
rect 1121 764 1449 796
rect 1005 739 1051 750
rect 1653 680 1699 691
rect 1893 831 1986 842
rect 1939 691 1986 831
rect 2143 918 2576 927
rect 2097 776 2143 787
rect 2301 831 2347 842
rect 1051 599 1396 634
rect 1005 588 1396 599
rect 1038 412 1129 542
rect 1038 366 1083 412
rect 1038 354 1129 366
rect 1350 412 1396 588
rect 1449 547 1495 659
rect 1893 639 1986 691
rect 2301 639 2347 691
rect 1893 593 2499 639
rect 1449 501 1791 547
rect 1837 501 1996 547
rect 2042 501 2202 547
rect 2248 501 2273 547
rect 1350 366 1361 412
rect 1407 366 1418 412
rect 106 262 286 287
rect 508 287 805 298
rect 60 136 106 147
rect 284 193 330 204
rect 284 90 330 147
rect 554 216 805 287
rect 851 320 921 331
rect 897 274 921 320
rect 1350 308 1418 366
rect 851 263 921 274
rect 984 262 995 308
rect 1041 262 1418 308
rect 1521 366 1889 412
rect 1935 366 2119 412
rect 2165 366 2335 412
rect 2381 366 2406 412
rect 1521 227 1567 366
rect 2453 320 2499 593
rect 2005 319 2499 320
rect 2005 309 2453 319
rect 554 181 1521 216
rect 554 170 1567 181
rect 1745 221 1791 232
rect 508 136 554 147
rect 1247 90 1258 124
rect 0 78 1258 90
rect 1304 90 1315 124
rect 1304 81 1745 90
rect 2051 274 2453 309
rect 2005 158 2051 169
rect 2229 193 2275 204
rect 2453 168 2499 179
rect 2229 90 2275 147
rect 1791 81 2576 90
rect 1304 78 2576 81
rect 0 -90 2576 78
<< labels >>
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1038 354 1129 542 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 2576 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1745 204 1791 232 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2301 639 2347 842 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
rlabel metal1 s 1893 639 1986 842 1 ZN
port 3 nsew default output
rlabel metal1 s 1893 593 2499 639 1 ZN
port 3 nsew default output
rlabel metal1 s 2453 320 2499 593 1 ZN
port 3 nsew default output
rlabel metal1 s 2005 274 2499 320 1 ZN
port 3 nsew default output
rlabel metal1 s 2453 168 2499 274 1 ZN
port 3 nsew default output
rlabel metal1 s 2005 168 2051 274 1 ZN
port 3 nsew default output
rlabel metal1 s 2005 158 2051 168 1 ZN
port 3 nsew default output
rlabel metal1 s 2097 856 2143 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1653 856 1699 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1209 856 1255 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 856 320 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2097 776 2143 856 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1653 776 1699 856 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 776 320 856 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1653 769 1699 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 769 320 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1653 680 1699 769 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2229 124 2275 204 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1745 124 1791 204 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 284 124 330 204 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2229 90 2275 124 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1745 90 1791 124 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1247 90 1315 124 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 284 90 330 124 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2576 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 1008
string GDS_END 918454
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 911698
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
