magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< obsv1 >>
rect 0 0 86372 46576
<< obsv2 >>
rect 0 0 86372 46576
<< metal3 >>
rect 1401 45776 2401 46576
rect 2626 45968 3626 46576
rect 4137 45776 5137 46576
rect 5362 45968 6362 46576
rect 6801 45776 7801 46576
rect 8026 45968 9026 46576
rect 9537 45776 10537 46576
rect 10762 45968 11762 46576
rect 12201 45776 13201 46576
rect 13426 45968 14426 46576
rect 14937 45776 15937 46576
rect 16162 45968 17162 46576
rect 17601 45776 18601 46576
rect 18826 45968 19826 46576
rect 20653 45776 21653 46576
rect 22258 45968 23258 46576
rect 23483 45776 24483 46576
rect 25158 45968 26158 46576
rect 26572 45776 27572 46576
rect 27877 45968 28877 46576
rect 29273 45968 30273 46576
rect 30710 45776 31710 46576
rect 32381 45968 33381 46576
rect 34024 45968 35024 46576
rect 35415 45776 36415 46576
rect 36948 45968 37948 46576
rect 38585 45776 39585 46576
rect 39882 45968 40882 46576
rect 41230 45776 42230 46576
rect 42430 45968 43430 46576
rect 43713 45968 44713 46576
rect 45069 45776 46069 46576
rect 46313 45776 47313 46576
rect 47538 45968 48538 46576
rect 48901 45776 49901 46576
rect 50465 45968 51465 46576
rect 52569 45776 53569 46576
rect 54262 45776 55262 46576
rect 55990 45968 56990 46576
rect 57547 45776 58547 46576
rect 58791 45968 59791 46576
rect 60977 45776 61977 46576
rect 62202 45968 63202 46576
rect 63713 45776 64713 46576
rect 64938 45968 65938 46576
rect 66377 45776 67377 46576
rect 67602 45968 68602 46576
rect 69113 45776 70113 46576
rect 70338 45968 71338 46576
rect 71777 45776 72777 46576
rect 73002 45968 74002 46576
rect 74513 45776 75513 46576
rect 75738 45968 76738 46576
rect 77177 45776 78177 46576
rect 78402 45968 79402 46576
rect 80229 45776 81229 46576
rect 81834 45968 82834 46576
rect 83059 45776 84059 46576
rect 84666 45776 85666 46576
rect 0 44776 86372 45776
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44328 27779 44376
rect 57051 44328 86372 44376
rect 0 44127 86372 44328
rect 0 44076 27779 44127
rect 30402 44126 54622 44127
rect 57051 44076 86372 44127
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 59421 42528 86372 42576
rect 0 42327 86372 42528
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 59421 42276 86372 42327
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 59421 40728 86372 40776
rect 0 40527 86372 40728
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 59421 40476 86372 40527
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 59421 38928 86372 38976
rect 0 38727 86372 38928
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 59421 38676 86372 38727
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 59421 37128 86372 37176
rect 0 36927 86372 37128
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 59421 36876 86372 36927
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 84666 35776 86372 36476
rect 0 35126 24920 35326
rect 0 35016 1014 35126
rect 60549 35298 60639 35370
rect 83360 35298 86372 35326
rect 60549 35158 86372 35298
rect 60549 35086 60639 35158
rect 83360 35126 86372 35158
rect 0 34962 25085 35016
rect 0 34536 27830 34962
rect 24942 34490 27830 34536
rect 85358 35016 86372 35126
rect 61311 34962 86372 35016
rect 60510 34536 86372 34962
rect 60510 34490 61754 34536
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 32318 27214 34124
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 32315 86372 34124
rect 57908 32199 58351 32315
rect 26772 31486 58351 32199
rect 26772 29714 58351 30105
rect 84666 29714 86372 32315
rect 0 29430 86372 29714
rect 0 26890 26070 28416
rect 26772 27382 58351 29430
rect 0 26435 27828 26890
rect 1271 26434 27828 26435
rect 1954 26433 2279 26434
rect 12754 26433 13079 26434
rect 58785 26890 86372 28416
rect 57295 26435 86372 26890
rect 61530 26434 84717 26435
rect 61530 26433 61855 26434
rect 72330 26433 72655 26434
rect 0 23380 1706 23938
rect 26770 23380 58348 24278
rect 84666 23380 86372 23938
rect 0 23370 86372 23380
rect 0 22938 27214 23370
rect 27387 22291 57677 23199
rect 57908 22938 86372 23370
rect 57908 22937 83763 22938
rect 27387 22282 27826 22291
rect 0 21827 27826 22282
rect 56078 22282 57677 22291
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 21827 86372 22282
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 19969 86372 20739
rect 0 18016 24250 19969
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 61807 16784 86372 17730
rect 24111 16597 27828 16598
rect 0 15015 27828 16597
rect 46982 15015 86372 16784
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14936 51760 14966
rect 0 14491 47683 14936
rect 0 14329 45977 14491
rect 0 14328 24250 14329
rect 24047 14178 27214 14179
rect 0 13461 27214 14178
rect 0 12846 1706 13461
rect 24047 12934 27214 13461
rect 27387 13760 45977 14329
rect 57295 14328 86372 14968
rect 57295 14327 83763 14328
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13245 49775 13760
rect 29478 13243 49775 13245
rect 41493 13078 49775 13243
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12606 34761 12846
rect 50228 13461 86372 13866
rect 50228 12846 58421 13461
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12606 86372 12846
rect 0 12046 86372 12606
rect 0 12036 24250 12046
rect 26772 12036 86372 12046
rect 26772 12035 84999 12036
rect 26772 11844 58351 12035
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 10176 27828 11491
rect 29478 11697 58351 11844
rect 29478 10756 41353 11697
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 34904 9972 41353 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 10740 86372 11491
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 8154 28729 9514
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 6982 27828 7595
rect 28178 7652 28729 8154
rect 41857 9502 51430 10420
rect 57295 10176 86372 10740
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 41857 9165 55482 9502
rect 29513 7900 41397 8582
rect 28178 7084 34622 7652
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 9012 55482 9165
rect 50922 7596 57736 9012
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 57909 8154 86372 9514
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7392 86372 7595
rect 34860 7088 86372 7392
rect 34860 6592 55482 7088
rect 34860 6573 41397 6592
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 0 5766 34622 6177
rect 23687 5629 27214 5630
rect 0 5175 27214 5629
rect 29458 5665 34622 5766
rect 50922 6199 55482 6592
rect 59309 6982 86372 7088
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 50922 5766 86372 6198
rect 50922 5605 55482 5766
rect 0 5174 24250 5175
rect 0 5173 3011 5174
rect 0 4515 1712 5173
rect 57909 5629 62429 5630
rect 57909 5175 86372 5629
rect 61802 5174 86372 5175
rect 83361 5173 86372 5174
rect 57909 4619 62429 4621
rect 23909 4515 62429 4619
rect 84660 4515 86372 5173
rect 0 4166 86372 4515
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3772 61215 3875
rect 0 3524 86372 3772
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 0 2854 1000 3420
rect 60886 3420 86372 3524
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
<< obsm3 >>
rect 0 45832 1345 46576
rect 2457 45912 2570 46576
rect 3682 45912 4081 46576
rect 2457 45832 4081 45912
rect 5193 45912 5306 46576
rect 6418 45912 6745 46576
rect 5193 45832 6745 45912
rect 7857 45912 7970 46576
rect 9082 45912 9481 46576
rect 7857 45832 9481 45912
rect 10593 45912 10706 46576
rect 11818 45912 12145 46576
rect 10593 45832 12145 45912
rect 13257 45912 13370 46576
rect 14482 45912 14881 46576
rect 13257 45832 14881 45912
rect 15993 45912 16106 46576
rect 17218 45912 17545 46576
rect 15993 45832 17545 45912
rect 18657 45912 18770 46576
rect 19882 45912 20597 46576
rect 18657 45832 20597 45912
rect 21709 45912 22202 46576
rect 23314 45912 23427 46576
rect 21709 45832 23427 45912
rect 24539 45912 25102 46576
rect 26214 45912 26516 46576
rect 24539 45832 26516 45912
rect 27628 45912 27821 46576
rect 28933 45912 29217 46576
rect 30329 45912 30654 46576
rect 27628 45832 30654 45912
rect 31766 45912 32325 46576
rect 33437 45912 33968 46576
rect 35080 45912 35359 46576
rect 31766 45832 35359 45912
rect 36471 45912 36892 46576
rect 38004 45912 38529 46576
rect 36471 45832 38529 45912
rect 39641 45912 39826 46576
rect 40938 45912 41174 46576
rect 39641 45832 41174 45912
rect 42286 45912 42374 46576
rect 43486 45912 43657 46576
rect 44769 45912 45013 46576
rect 42286 45832 45013 45912
rect 46125 45832 46257 46576
rect 47369 45912 47482 46576
rect 48594 45912 48845 46576
rect 47369 45832 48845 45912
rect 49957 45912 50409 46576
rect 51521 45912 52513 46576
rect 49957 45832 52513 45912
rect 53625 45832 54206 46576
rect 55318 45912 55934 46576
rect 57046 45912 57491 46576
rect 55318 45832 57491 45912
rect 58603 45912 58735 46576
rect 59847 45912 60921 46576
rect 58603 45832 60921 45912
rect 62033 45912 62146 46576
rect 63258 45912 63657 46576
rect 62033 45832 63657 45912
rect 64769 45912 64882 46576
rect 65994 45912 66321 46576
rect 64769 45832 66321 45912
rect 67433 45912 67546 46576
rect 68658 45912 69057 46576
rect 67433 45832 69057 45912
rect 70169 45912 70282 46576
rect 71394 45912 71721 46576
rect 70169 45832 71721 45912
rect 72833 45912 72946 46576
rect 74058 45912 74457 46576
rect 72833 45832 74457 45912
rect 75569 45912 75682 46576
rect 76794 45912 77121 46576
rect 75569 45832 77121 45912
rect 78233 45912 78346 46576
rect 79458 45912 80173 46576
rect 78233 45832 80173 45912
rect 81285 45912 81778 46576
rect 82890 45912 83003 46576
rect 81285 45832 83003 45912
rect 84115 45832 84610 46576
rect 85722 45832 86372 46576
rect 0 44632 86372 44720
rect 1070 44432 85302 44632
rect 27835 44384 56995 44432
rect 27835 44070 30346 44071
rect 54678 44070 56995 44071
rect 27835 44020 56995 44070
rect 1070 43820 85302 44020
rect 0 43732 86372 43820
rect 1762 42920 84610 43732
rect 0 42832 86372 42920
rect 1070 42632 85302 42832
rect 27328 42584 59365 42632
rect 27328 42270 30347 42271
rect 54678 42270 59365 42271
rect 27328 42220 59365 42270
rect 1070 42020 85302 42220
rect 0 41932 86372 42020
rect 1762 41120 84610 41932
rect 0 41032 86372 41120
rect 1070 40832 85302 41032
rect 27328 40784 59365 40832
rect 27328 40470 30347 40471
rect 54678 40470 59365 40471
rect 27328 40420 59365 40470
rect 1070 40220 85302 40420
rect 0 40132 86372 40220
rect 1762 39320 84610 40132
rect 0 39232 86372 39320
rect 1070 39032 85302 39232
rect 27328 38984 59365 39032
rect 27328 38670 30347 38671
rect 54678 38670 59365 38671
rect 27328 38620 59365 38670
rect 1070 38420 85302 38620
rect 0 38332 86372 38420
rect 1762 37520 84610 38332
rect 0 37432 86372 37520
rect 1070 37232 85302 37432
rect 27328 37184 59365 37232
rect 27328 36870 30347 36871
rect 54678 36870 59365 36871
rect 27328 36820 59365 36870
rect 1070 36620 85302 36820
rect 0 36532 86372 36620
rect 1762 35720 84610 36532
rect 0 35426 86372 35720
rect 0 35382 60493 35426
rect 24976 35072 60493 35382
rect 60695 35382 86372 35426
rect 60695 35354 83304 35382
rect 25141 35030 60493 35072
rect 60695 35072 83304 35102
rect 60695 35030 61255 35072
rect 25141 35018 61255 35030
rect 0 34434 24886 34480
rect 27886 34434 60454 35018
rect 61810 34434 86372 34480
rect 0 34182 86372 34434
rect 0 34181 2039 34182
rect 2244 34181 86372 34182
rect 25141 34180 61797 34181
rect 72439 34180 72597 34181
rect 27270 32262 57852 34180
rect 25141 32260 57852 32262
rect 3067 32259 57852 32260
rect 1762 32255 57852 32259
rect 1762 31430 26716 32255
rect 58407 31430 84610 32259
rect 1762 30161 84610 31430
rect 1762 29770 26716 30161
rect 58407 29770 84610 30161
rect 0 28472 26716 29374
rect 26126 27326 26716 28472
rect 58407 28472 86372 29374
rect 58407 27326 58729 28472
rect 26126 26946 58729 27326
rect 27884 26379 57239 26946
rect 0 26378 1215 26379
rect 27884 26378 61474 26379
rect 84773 26378 86372 26379
rect 0 26377 1898 26378
rect 2335 26377 12698 26378
rect 13135 26377 61474 26378
rect 61911 26377 72274 26378
rect 72711 26377 86372 26378
rect 0 24334 86372 26377
rect 0 23994 26714 24334
rect 1762 23436 26714 23994
rect 58404 23994 86372 24334
rect 58404 23436 84610 23994
rect 27270 23255 57852 23314
rect 27270 22882 27331 23255
rect 0 22338 27331 22882
rect 57733 22881 57852 23255
rect 83819 22881 86372 22882
rect 57733 22338 86372 22881
rect 1070 21770 23980 21771
rect 27882 21770 56022 22235
rect 83819 21770 85302 21771
rect 1070 21764 85302 21770
rect 1070 21763 44376 21764
rect 1070 21681 29465 21763
rect 1070 21226 29457 21681
rect 0 20795 29457 21226
rect 55701 21226 85302 21764
rect 55701 20795 86372 21226
rect 24306 17960 61751 19913
rect 0 17959 61769 17960
rect 83819 17959 86372 17960
rect 0 17786 86372 17959
rect 23734 16840 61751 17786
rect 23734 16654 46926 16840
rect 23734 16653 24055 16654
rect 27884 15071 46926 16654
rect 55701 14910 57239 14912
rect 51816 14880 57239 14910
rect 47739 14435 57239 14880
rect 24306 14272 27331 14273
rect 0 14235 27331 14272
rect 0 14234 23991 14235
rect 1762 12903 23991 13405
rect 27270 13189 27331 14235
rect 46033 14271 57239 14435
rect 83819 14271 86372 14272
rect 46033 14235 86372 14271
rect 46033 14234 83113 14235
rect 84277 14234 86372 14235
rect 46033 14233 61751 14234
rect 72485 14233 72551 14234
rect 46033 14073 61717 14233
rect 46033 13922 59770 14073
rect 46033 13816 50172 13922
rect 60082 13922 61717 14073
rect 27270 13187 29422 13189
rect 27270 13022 41437 13187
rect 49831 13022 50172 13816
rect 27270 12990 50172 13022
rect 1762 12902 23765 12903
rect 34817 12662 50172 12990
rect 58477 12902 59770 13405
rect 60082 12903 84610 13405
rect 60082 12902 83113 12903
rect 84277 12902 84610 12903
rect 24306 11980 26716 11990
rect 0 11788 26716 11980
rect 85055 11979 86372 11980
rect 0 11549 29422 11788
rect 3067 11547 23991 11549
rect 27884 10700 29422 11549
rect 58407 11641 86372 11979
rect 27884 10120 34848 10700
rect 0 10119 2173 10120
rect 0 10118 2193 10119
rect 24306 10118 34848 10120
rect 0 9916 34848 10118
rect 41409 11583 86372 11641
rect 41409 10684 42205 11583
rect 57792 11549 86372 11583
rect 57792 11547 61769 11549
rect 41409 10476 57239 10684
rect 41409 9916 41801 10476
rect 0 9572 41801 9916
rect 0 9571 23991 9572
rect 1070 9570 2170 9571
rect 24306 8097 28122 8098
rect 3067 8096 28122 8097
rect 0 7652 28122 8096
rect 3067 7651 23569 7652
rect 27884 7028 28122 7652
rect 28785 9109 41801 9572
rect 51486 10120 57239 10476
rect 51486 10119 61749 10120
rect 51486 10117 61769 10119
rect 84538 10117 86372 10120
rect 51486 9572 86372 10117
rect 51486 9558 57853 9572
rect 62334 9571 86372 9572
rect 72490 9570 72546 9571
rect 83290 9570 85302 9571
rect 28785 8638 50866 9109
rect 28785 7844 29457 8638
rect 28785 7708 34804 7844
rect 27884 6926 29481 7028
rect 1070 6925 2170 6926
rect 1070 6924 2193 6925
rect 24306 6924 29481 6926
rect 1070 6688 29481 6924
rect 34678 6688 34804 7708
rect 1070 6629 34804 6688
rect 41453 7448 50866 8638
rect 55538 9068 57853 9558
rect 57792 8098 57853 9068
rect 57792 8097 61746 8098
rect 57792 8096 61769 8097
rect 57792 7652 86372 8096
rect 62803 7651 83305 7652
rect 1070 6255 29402 6629
rect 3067 6254 23631 6255
rect 41453 6121 50866 6536
rect 0 5686 29402 5710
rect 0 5685 23631 5686
rect 27270 5609 29402 5686
rect 34678 5609 50866 6121
rect 27270 5549 50866 5609
rect 55538 6926 59253 7032
rect 55538 6925 61746 6926
rect 55538 6924 61769 6925
rect 84843 6924 85302 6926
rect 55538 6255 85302 6924
rect 62485 6254 83305 6255
rect 55538 5686 86372 5710
rect 55538 5549 57853 5686
rect 62485 5685 86372 5686
rect 27270 5119 57853 5549
rect 24306 5118 61746 5119
rect 3067 5117 83305 5118
rect 1768 4677 84604 5117
rect 1768 4675 57853 4677
rect 1768 4571 23853 4675
rect 62485 4571 84604 4677
rect 59379 4108 61732 4110
rect 24397 4004 61732 4108
rect 0 3932 86372 4004
rect 0 3931 27382 3932
rect 27834 3931 28708 3932
rect 28950 3931 41718 3932
rect 41960 3931 42243 3932
rect 42485 3931 46817 3932
rect 47059 3931 47265 3932
rect 47507 3931 47713 3932
rect 47955 3931 48161 3932
rect 48403 3931 57289 3932
rect 0 3828 23853 3931
rect 61271 3828 86372 3932
rect 24397 3365 60830 3468
rect 3067 3364 60830 3365
rect 1056 2910 85302 3364
rect 0 2288 86372 2446
rect 0 0 650 1176
rect 1762 0 1983 1176
rect 3095 0 3386 1176
rect 4498 988 5786 1176
rect 4498 0 4586 988
rect 5698 0 5786 988
rect 6898 0 6986 1176
rect 8098 0 8186 1176
rect 9298 988 10586 1176
rect 9298 0 9386 988
rect 10498 0 10586 988
rect 11698 0 12387 1176
rect 13499 0 14186 1176
rect 15298 988 16586 1176
rect 15298 0 15386 988
rect 16498 0 16586 988
rect 17698 0 17786 1176
rect 18898 0 18986 1176
rect 20098 988 21854 1176
rect 20098 0 20186 988
rect 21298 0 21854 988
rect 22966 0 23054 1176
rect 24166 0 24354 1176
rect 25466 0 25654 1176
rect 26766 0 26954 1176
rect 28066 0 28254 1176
rect 29366 0 29554 1176
rect 30666 988 35975 1176
rect 30666 0 31268 988
rect 32380 0 32966 988
rect 34078 0 34775 988
rect 35887 0 35975 988
rect 37087 988 39172 1176
rect 37087 0 37972 988
rect 39084 0 39172 988
rect 40284 988 42377 1176
rect 40284 0 41177 988
rect 42289 0 42377 988
rect 43489 988 44777 1176
rect 43489 0 43577 988
rect 44689 0 44777 988
rect 45889 988 47177 1176
rect 45889 0 45977 988
rect 47089 0 47177 988
rect 48289 0 48510 1176
rect 49622 0 49820 1176
rect 50932 988 54402 1176
rect 50932 0 51177 988
rect 52289 0 52422 988
rect 53534 0 54402 988
rect 55514 0 55702 1176
rect 56814 0 57002 1176
rect 58114 0 58302 1176
rect 59414 0 59602 1176
rect 60714 0 60902 1176
rect 62014 0 62239 1176
rect 63351 988 65362 1176
rect 63351 0 64162 988
rect 65274 0 65362 988
rect 66474 0 66562 1176
rect 67674 0 67762 1176
rect 68874 988 70162 1176
rect 68874 0 68962 988
rect 70074 0 70162 988
rect 71274 0 71961 1176
rect 73073 0 73762 1176
rect 74874 988 76162 1176
rect 74874 0 74962 988
rect 76074 0 76162 988
rect 77274 0 77362 1176
rect 78474 0 78562 1176
rect 79674 988 80962 1176
rect 79674 0 79762 988
rect 80874 0 80962 988
rect 82074 0 82363 1176
rect 83475 0 84610 1176
rect 85722 0 86372 1176
<< labels >>
rlabel metal2 s 34243 0 34467 200 6 A[0]
port 6 nsew signal input
rlabel metal2 s 32552 0 32776 200 6 A[1]
port 5 nsew signal input
rlabel metal2 s 30859 0 31083 200 6 A[2]
port 4 nsew signal input
rlabel metal2 s 56265 0 56489 200 6 A[3]
port 3 nsew signal input
rlabel metal2 s 55164 0 55388 200 6 A[4]
port 2 nsew signal input
rlabel metal2 s 54417 0 54641 200 6 A[5]
port 1 nsew signal input
rlabel metal2 s 50342 0 50566 200 6 CEN
port 7 nsew signal input
rlabel metal2 s 27936 0 28160 200 6 CLK
port 8 nsew signal input
rlabel metal2 s 1864 0 2088 200 6 D[0]
port 16 nsew signal input
rlabel metal2 s 12206 0 12430 200 6 D[1]
port 15 nsew signal input
rlabel metal2 s 13454 0 13678 200 6 D[2]
port 14 nsew signal input
rlabel metal2 s 23795 0 24019 200 6 D[3]
port 13 nsew signal input
rlabel metal2 s 61447 0 61671 200 6 D[4]
port 12 nsew signal input
rlabel metal2 s 71782 0 72006 200 6 D[5]
port 11 nsew signal input
rlabel metal2 s 73030 0 73254 200 6 D[6]
port 10 nsew signal input
rlabel metal2 s 83372 0 83596 200 6 D[7]
port 9 nsew signal input
rlabel metal2 s 40588 0 40812 200 6 GWEN
port 17 nsew signal input
rlabel metal2 s 3380 0 3604 200 6 Q[0]
port 25 nsew signal output
rlabel metal2 s 11533 0 11757 200 6 Q[1]
port 24 nsew signal output
rlabel metal2 s 14127 0 14351 200 6 Q[2]
port 23 nsew signal output
rlabel metal2 s 22279 0 22503 200 6 Q[3]
port 22 nsew signal output
rlabel metal2 s 62958 0 63182 200 6 Q[4]
port 21 nsew signal output
rlabel metal2 s 71109 0 71333 200 6 Q[5]
port 20 nsew signal output
rlabel metal2 s 73703 0 73927 200 6 Q[6]
port 19 nsew signal output
rlabel metal2 s 81855 0 82079 200 6 Q[7]
port 18 nsew signal output
rlabel metal2 s 2539 0 2763 200 6 WEN[0]
port 35 nsew signal input
rlabel metal2 s 12604 0 12828 200 6 WEN[1]
port 34 nsew signal input
rlabel metal2 s 13054 0 13278 200 6 WEN[2]
port 33 nsew signal input
rlabel metal2 s 23404 0 23628 200 6 WEN[3]
port 32 nsew signal input
rlabel metal2 s 62115 0 62339 200 6 WEN[4]
port 31 nsew signal input
rlabel metal2 s 72180 0 72404 200 6 WEN[5]
port 30 nsew signal input
rlabel metal2 s 72630 0 72854 200 6 WEN[6]
port 29 nsew signal input
rlabel metal2 s 82695 0 82919 200 6 WEN[7]
port 28 nsew signal input
rlabel metal3 s 0 42976 1706 43676 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 41176 1706 41876 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 39376 1706 40076 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 37576 1706 38276 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 35776 1706 36476 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 8152 1014 9515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 8152 3011 9514 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 2226 8154 28729 9515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 8153 24250 9514 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 28178 7084 28729 9516 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 24047 8154 28729 9516 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29537 6744 34622 7652 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 28178 7084 34622 7652 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 1401 44776 2401 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 4137 44776 5137 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 6801 44776 7801 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 9537 44776 10537 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 12201 44776 13201 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 14937 44776 15937 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 17601 44776 18601 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 20653 44776 21653 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23483 44776 24483 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26572 44776 27572 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 30710 44776 31710 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 35415 44776 36415 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 38585 44776 39585 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 41230 44776 42230 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 45069 44776 46069 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 46313 44776 47313 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 48901 44776 49901 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 52569 44776 53569 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 54262 44776 55262 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57547 44776 58547 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 60977 44776 61977 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 63713 44776 64713 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 66377 44776 67377 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 69113 44776 70113 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 71777 44776 72777 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 74513 44776 75513 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 77177 44776 78177 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 80229 44776 81229 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 83059 44776 84059 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 44776 85666 46576 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 44776 86372 45776 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 42976 86372 43676 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 41176 86372 41876 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 39376 86372 40076 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 37576 86372 38276 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 35776 86372 36476 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 29430 1706 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 2095 32315 2188 34126 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 32315 3011 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 32316 25085 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 32318 27214 34124 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26772 31486 58351 32199 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26772 27382 58351 30105 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57908 31486 58351 34124 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61853 32315 72383 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57908 32315 86372 34124 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 29430 86372 29714 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 29430 86372 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 72653 32315 86372 34125 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 22938 1706 23938 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 22938 27214 23380 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26770 23370 58348 24278 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57908 22937 83763 23380 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57908 22938 86372 23380 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 22938 86372 23938 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 18016 24250 20739 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29513 19969 55645 21625 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29521 19969 55645 21707 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 44432 19969 55645 21708 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61825 18015 83763 20739 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61807 18016 86372 20739 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 19969 86372 20739 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 12036 1706 14178 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23821 12046 34761 12847 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 13461 27214 14178 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 12036 24250 12846 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 24047 12046 27214 14179 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 24047 12046 34761 12934 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 34904 9972 41353 12606 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29478 10756 41353 12606 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29478 11697 58351 12606 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26772 11844 58351 12606 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 50228 12035 58421 13866 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 59826 12035 60026 14017 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 50228 13461 86372 13866 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61807 13461 72429 14178 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61773 13461 86372 14177 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 83169 12035 84221 12847 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 83169 13461 84221 14179 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 50228 12036 86372 12846 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 26772 12035 84999 12606 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 12036 86372 14178 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 72607 13461 86372 14178 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61802 8153 86372 9514 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 8154 62278 9516 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 8154 72434 9515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 72602 8152 83234 9515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61825 8152 86372 9514 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 85358 8152 86372 9515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 4060 1712 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 5173 3011 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 5174 24250 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 4060 24341 4515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 6 VDD
port 26 nsew power bidirectional
rlabel metal3 s 2626 45968 3626 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 4642 0 5642 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 5362 45968 6362 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 8026 45968 9026 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 9442 0 10442 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 10762 45968 11762 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 13426 45968 14426 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 15442 0 16442 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 16162 45968 17162 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 18826 45968 19826 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 20242 0 21242 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 22258 45968 23258 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 25158 45968 26158 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 1954 26433 2279 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 12754 26433 13079 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 26435 26070 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 1271 26434 27828 26890 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 10176 3011 11493 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2249 10174 24250 11491 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2229 10175 24250 11491 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24047 10176 27828 11493 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 34536 1014 35326 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 35126 24920 35326 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 34536 25085 35016 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24942 34490 27830 34962 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27877 45968 28877 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29273 45968 30273 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 31324 0 32324 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 32381 45968 33381 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 33022 0 34022 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34024 45968 35024 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34831 0 35831 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 36948 45968 37948 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 38028 0 39028 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 39882 45968 40882 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41233 0 42233 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 42430 45968 43430 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 43633 0 44633 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 43713 45968 44713 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 46033 0 47033 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 47538 45968 48538 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50465 45968 51465 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 51233 0 52233 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 52478 0 53478 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 55990 45968 56990 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 58791 45968 59791 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 62202 45968 63202 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 64218 0 65218 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 64938 45968 65938 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 67602 45968 68602 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 69018 0 70018 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 70338 45968 71338 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 73002 45968 74002 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 75018 0 76018 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 75738 45968 76738 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 78402 45968 79402 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 79818 0 80818 932 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 81834 45968 82834 46576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 44076 27779 44376 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30402 44126 54622 44328 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 44127 86372 44328 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57051 44076 86372 44376 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 42327 86372 42528 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 40527 86372 40728 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60549 35086 60639 35370 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60510 34490 61754 34962 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60549 35158 86372 35298 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61311 34536 86372 35016 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61530 26433 61855 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 72330 26433 72655 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61530 26434 84717 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 7088 57736 9012 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59309 6982 86372 7595 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 7088 62747 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 6 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 6 VSS
port 27 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 46576
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2322524
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2272312
<< end >>
