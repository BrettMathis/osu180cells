magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 1274
<< mvpmos >>
rect 0 0 120 1154
<< mvpdiff >>
rect -88 1141 0 1154
rect -88 1095 -75 1141
rect -29 1095 0 1141
rect -88 1033 0 1095
rect -88 987 -75 1033
rect -29 987 0 1033
rect -88 925 0 987
rect -88 879 -75 925
rect -29 879 0 925
rect -88 817 0 879
rect -88 771 -75 817
rect -29 771 0 817
rect -88 709 0 771
rect -88 663 -75 709
rect -29 663 0 709
rect -88 601 0 663
rect -88 555 -75 601
rect -29 555 0 601
rect -88 493 0 555
rect -88 447 -75 493
rect -29 447 0 493
rect -88 385 0 447
rect -88 339 -75 385
rect -29 339 0 385
rect -88 277 0 339
rect -88 231 -75 277
rect -29 231 0 277
rect -88 168 0 231
rect -88 122 -75 168
rect -29 122 0 168
rect -88 59 0 122
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1141 208 1154
rect 120 1095 149 1141
rect 195 1095 208 1141
rect 120 1033 208 1095
rect 120 987 149 1033
rect 195 987 208 1033
rect 120 925 208 987
rect 120 879 149 925
rect 195 879 208 925
rect 120 817 208 879
rect 120 771 149 817
rect 195 771 208 817
rect 120 709 208 771
rect 120 663 149 709
rect 195 663 208 709
rect 120 601 208 663
rect 120 555 149 601
rect 195 555 208 601
rect 120 493 208 555
rect 120 447 149 493
rect 195 447 208 493
rect 120 385 208 447
rect 120 339 149 385
rect 195 339 208 385
rect 120 277 208 339
rect 120 231 149 277
rect 195 231 208 277
rect 120 168 208 231
rect 120 122 149 168
rect 195 122 208 168
rect 120 59 208 122
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 1095 -29 1141
rect -75 987 -29 1033
rect -75 879 -29 925
rect -75 771 -29 817
rect -75 663 -29 709
rect -75 555 -29 601
rect -75 447 -29 493
rect -75 339 -29 385
rect -75 231 -29 277
rect -75 122 -29 168
rect -75 13 -29 59
rect 149 1095 195 1141
rect 149 987 195 1033
rect 149 879 195 925
rect 149 771 195 817
rect 149 663 195 709
rect 149 555 195 601
rect 149 447 195 493
rect 149 339 195 385
rect 149 231 195 277
rect 149 122 195 168
rect 149 13 195 59
<< polysilicon >>
rect 0 1154 120 1198
rect 0 -44 120 0
<< metal1 >>
rect -75 1141 -29 1154
rect -75 1033 -29 1095
rect -75 925 -29 987
rect -75 817 -29 879
rect -75 709 -29 771
rect -75 601 -29 663
rect -75 493 -29 555
rect -75 385 -29 447
rect -75 277 -29 339
rect -75 168 -29 231
rect -75 59 -29 122
rect -75 0 -29 13
rect 149 1141 195 1154
rect 149 1033 195 1095
rect 149 925 195 987
rect 149 817 195 879
rect 149 709 195 771
rect 149 601 195 663
rect 149 493 195 555
rect 149 385 195 447
rect 149 277 195 339
rect 149 168 195 231
rect 149 59 195 122
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 577 -52 577 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 577 172 577 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 31666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 29298
<< end >>
