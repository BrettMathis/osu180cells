* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__dffr_1 D RN Q QN CLK
X0 VDD a_41_109 a_145_109 VDD pmos_3p3 w=34 l=6
X1 a_173_109 a_41_109 VDD VDD pmos_3p3 w=34 l=6
X2 a_122_14 CLK VDD VDD pmos_3p3 w=34 l=6
X3 a_122_14 CLK VSS VSS nmos_3p3 w=17 l=6
X4 VDD a_205_68 a_201_109 VDD pmos_3p3 w=34 l=6
X5 a_62_98 CLK a_112_109 VDD pmos_3p3 w=34 l=6
X6 a_145_109 a_122_14 a_62_98 VDD pmos_3p3 w=34 l=6
X7 a_145_19 CLK a_62_98 VSS nmos_3p3 w=17 l=6
X8 a_25_19 RN VDD VDD pmos_3p3 w=34 l=6
X9 a_41_109 a_25_19 VSS VSS nmos_3p3 w=17 l=6
X10 a_62_98 a_122_14 a_112_19 VSS nmos_3p3 w=17 l=6
X11 a_112_109 D VDD VDD pmos_3p3 w=34 l=6
X12 a_205_68 a_184_19 VSS VSS nmos_3p3 w=17 l=6
X13 a_25_19 RN VSS VSS nmos_3p3 w=17 l=6
X14 VDD a_205_68 QN VDD pmos_3p3 w=34 l=6
X15 Q QN VDD VDD pmos_3p3 w=34 l=6
X16 a_201_19 a_122_14 a_184_19 VSS nmos_3p3 w=17 l=6
X17 VSS a_205_68 a_201_19 VSS nmos_3p3 w=17 l=6
X18 Q QN VSS VSS nmos_3p3 w=17 l=6
X19 a_205_68 a_25_19 a_273_109 VDD pmos_3p3 w=34 l=6
X20 a_273_109 a_184_19 VDD VDD pmos_3p3 w=34 l=6
X21 VSS a_205_68 QN VSS nmos_3p3 w=17 l=6
X22 VSS a_62_98 a_41_109 VSS nmos_3p3 w=17 l=6
X23 VDD a_62_98 a_57_109 VDD pmos_3p3 w=34 l=6
X24 a_112_19 D VSS VSS nmos_3p3 w=17 l=6
X25 VSS a_25_19 a_205_68 VSS nmos_3p3 w=17 l=6
X26 a_57_109 a_25_19 a_41_109 VDD pmos_3p3 w=34 l=6
X27 a_173_19 a_41_109 VSS VSS nmos_3p3 w=17 l=6
X28 a_201_109 CLK a_184_19 VDD pmos_3p3 w=34 l=6
X29 a_184_19 a_122_14 a_173_109 VDD pmos_3p3 w=34 l=6
X30 VSS a_41_109 a_145_19 VSS nmos_3p3 w=17 l=6
X31 a_184_19 CLK a_173_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
