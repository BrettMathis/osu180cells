magic
tech gf180mcuA
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect -236 75 236 81
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -81 236 -75
<< via1 >>
rect -230 49 -204 75
rect -168 49 -142 75
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect 142 49 168 75
rect 204 49 230 75
rect -230 -13 -204 13
rect -168 -13 -142 13
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect 142 -13 168 13
rect 204 -13 230 13
rect -230 -75 -204 -49
rect -168 -75 -142 -49
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect 142 -75 168 -49
rect 204 -75 230 -49
<< metal2 >>
rect -236 75 236 81
rect -236 49 -230 75
rect -204 49 -168 75
rect -142 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 142 75
rect 168 49 204 75
rect 230 49 236 75
rect -236 13 236 49
rect -236 -13 -230 13
rect -204 -13 -168 13
rect -142 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 142 13
rect 168 -13 204 13
rect 230 -13 236 13
rect -236 -49 236 -13
rect -236 -75 -230 -49
rect -204 -75 -168 -49
rect -142 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 142 -49
rect 168 -75 204 -49
rect 230 -75 236 -49
rect -236 -81 236 -75
<< properties >>
string GDS_END 833626
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 831958
<< end >>
