magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 228
rect 224 0 344 228
rect 448 0 568 228
rect 672 0 792 228
rect 896 0 1016 228
<< mvndiff >>
rect -88 215 0 228
rect -88 169 -75 215
rect -29 169 0 215
rect -88 59 0 169
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 215 224 228
rect 120 169 149 215
rect 195 169 224 215
rect 120 59 224 169
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 215 448 228
rect 344 169 373 215
rect 419 169 448 215
rect 344 59 448 169
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 215 672 228
rect 568 169 597 215
rect 643 169 672 215
rect 568 59 672 169
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 215 896 228
rect 792 169 821 215
rect 867 169 896 215
rect 792 59 896 169
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 215 1104 228
rect 1016 169 1045 215
rect 1091 169 1104 215
rect 1016 59 1104 169
rect 1016 13 1045 59
rect 1091 13 1104 59
rect 1016 0 1104 13
<< mvndiffc >>
rect -75 169 -29 215
rect -75 13 -29 59
rect 149 169 195 215
rect 149 13 195 59
rect 373 169 419 215
rect 373 13 419 59
rect 597 169 643 215
rect 597 13 643 59
rect 821 169 867 215
rect 821 13 867 59
rect 1045 169 1091 215
rect 1045 13 1091 59
<< polysilicon >>
rect 0 228 120 272
rect 224 228 344 272
rect 448 228 568 272
rect 672 228 792 272
rect 896 228 1016 272
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
<< metal1 >>
rect -75 215 -29 228
rect -75 59 -29 169
rect -75 0 -29 13
rect 149 215 195 228
rect 149 59 195 169
rect 149 0 195 13
rect 373 215 419 228
rect 373 59 419 169
rect 373 0 419 13
rect 597 215 643 228
rect 597 59 643 169
rect 597 0 643 13
rect 821 215 867 228
rect 821 59 867 169
rect 821 0 867 13
rect 1045 215 1091 228
rect 1045 59 1091 169
rect 1045 0 1091 13
<< labels >>
flabel metal1 s -52 114 -52 114 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 114 1068 114 0 FreeSans 200 0 0 0 D
flabel metal1 s 172 114 172 114 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 114 396 114 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 114 620 114 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 114 844 114 0 FreeSans 200 0 0 0 S
<< properties >>
string GDS_END 104628
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 101436
<< end >>
