magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 1240 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 470 190 530 360
rect 700 190 760 360
rect 810 190 870 360
rect 980 190 1040 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 470 1090 530 1430
rect 700 1090 760 1430
rect 810 1090 870 1430
rect 980 1090 1040 1430
<< ndiff >>
rect 560 360 660 370
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 470 360
rect 530 350 700 360
rect 530 210 592 350
rect 638 210 700 350
rect 530 190 700 210
rect 760 190 810 360
rect 870 298 980 360
rect 870 252 902 298
rect 948 252 980 298
rect 870 190 980 252
rect 1040 298 1140 360
rect 1040 252 1072 298
rect 1118 252 1140 298
rect 1040 190 1140 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1090 470 1430
rect 530 1377 700 1430
rect 530 1143 592 1377
rect 638 1143 700 1377
rect 530 1090 700 1143
rect 760 1090 810 1430
rect 870 1377 980 1430
rect 870 1143 902 1377
rect 948 1143 980 1377
rect 870 1090 980 1143
rect 1040 1377 1140 1430
rect 1040 1143 1072 1377
rect 1118 1143 1140 1377
rect 1040 1090 1140 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 592 210 638 350
rect 902 252 948 298
rect 1072 252 1118 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 592 1143 638 1377
rect 902 1143 948 1377
rect 1072 1143 1118 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 470 1430 530 1480
rect 700 1430 760 1480
rect 810 1430 870 1480
rect 980 1430 1040 1480
rect 190 520 250 1090
rect 360 780 420 1090
rect 310 753 420 780
rect 310 707 337 753
rect 383 707 420 753
rect 310 680 420 707
rect 470 910 530 1090
rect 470 883 610 910
rect 470 837 537 883
rect 583 837 610 883
rect 470 810 610 837
rect 190 493 350 520
rect 190 447 277 493
rect 323 470 350 493
rect 323 447 420 470
rect 190 410 420 447
rect 190 360 250 410
rect 360 360 420 410
rect 470 360 530 810
rect 700 780 760 1090
rect 810 1040 870 1090
rect 980 1040 1040 1090
rect 810 980 1040 1040
rect 690 753 810 780
rect 690 707 737 753
rect 783 707 810 753
rect 690 680 810 707
rect 980 520 1040 980
rect 580 500 680 520
rect 580 493 760 500
rect 580 447 607 493
rect 653 447 760 493
rect 870 493 1040 520
rect 870 470 897 493
rect 580 420 760 447
rect 700 360 760 420
rect 810 447 897 470
rect 943 447 1040 493
rect 810 420 1040 447
rect 810 360 870 420
rect 980 360 1040 420
rect 190 140 250 190
rect 360 140 420 190
rect 470 140 530 190
rect 700 140 760 190
rect 810 140 870 190
rect 980 140 1040 190
<< polycontact >>
rect 337 707 383 753
rect 537 837 583 883
rect 277 447 323 493
rect 737 707 783 753
rect 607 447 653 493
rect 897 447 943 493
<< metal1 >>
rect 0 1568 1240 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1240 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1240 1566
rect 0 1470 1240 1514
rect 110 1377 160 1430
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 760 160 1143
rect 280 1377 330 1470
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 590 1377 640 1430
rect 590 1170 592 1377
rect 280 1060 330 1143
rect 580 1146 592 1170
rect 580 1094 584 1146
rect 638 1143 640 1377
rect 636 1094 640 1143
rect 580 1030 640 1094
rect 900 1377 950 1470
rect 900 1143 902 1377
rect 948 1143 950 1377
rect 900 1060 950 1143
rect 1070 1377 1120 1430
rect 1070 1143 1072 1377
rect 1118 1143 1120 1377
rect 1070 890 1120 1143
rect 510 883 1120 890
rect 510 837 537 883
rect 583 837 1120 883
rect 510 830 1120 837
rect 110 753 660 760
rect 110 707 337 753
rect 383 707 660 753
rect 110 700 660 707
rect 110 298 160 700
rect 600 500 660 700
rect 710 756 810 760
rect 710 704 734 756
rect 786 704 810 756
rect 710 670 810 704
rect 250 496 350 500
rect 250 444 274 496
rect 326 444 350 496
rect 250 410 350 444
rect 580 493 680 500
rect 580 447 607 493
rect 653 447 680 493
rect 580 440 680 447
rect 870 496 970 500
rect 870 444 894 496
rect 946 444 970 496
rect 870 410 970 444
rect 580 366 640 390
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 580 314 584 366
rect 636 350 640 366
rect 580 250 592 314
rect 590 210 592 250
rect 638 210 640 350
rect 590 160 640 210
rect 900 298 950 360
rect 900 252 902 298
rect 948 252 950 298
rect 900 120 950 252
rect 1070 298 1120 830
rect 1070 252 1072 298
rect 1118 252 1120 298
rect 1070 190 1120 252
rect 0 106 1240 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1240 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1240 54
rect 0 -30 1240 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 584 1143 592 1146
rect 592 1143 636 1146
rect 584 1094 636 1143
rect 734 753 786 756
rect 734 707 737 753
rect 737 707 783 753
rect 783 707 786 753
rect 734 704 786 707
rect 274 493 326 496
rect 274 447 277 493
rect 277 447 323 493
rect 323 447 326 493
rect 274 444 326 447
rect 894 493 946 496
rect 894 447 897 493
rect 897 447 943 493
rect 943 447 946 493
rect 894 444 946 447
rect 584 350 636 366
rect 584 314 592 350
rect 592 314 636 350
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1480 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1480 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1480 1150 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 580 1470 660 1480
rect 820 1470 900 1480
rect 1060 1470 1140 1480
rect 580 1160 640 1190
rect 570 1146 650 1160
rect 570 1094 584 1146
rect 636 1094 650 1146
rect 570 1050 650 1094
rect 270 510 330 520
rect 260 496 340 510
rect 260 444 274 496
rect 326 444 340 496
rect 260 400 340 444
rect 270 240 330 400
rect 580 380 640 1050
rect 730 770 790 780
rect 720 756 800 770
rect 720 704 734 756
rect 786 704 800 756
rect 720 660 800 704
rect 560 366 660 380
rect 560 314 584 366
rect 636 314 660 366
rect 560 270 660 314
rect 730 240 790 660
rect 890 510 950 520
rect 880 500 960 510
rect 870 496 970 500
rect 870 444 894 496
rect 946 444 970 496
rect 870 410 970 444
rect 880 400 960 410
rect 890 390 950 400
rect 270 150 790 240
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 20 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 20 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 20 1150 54
rect 100 10 180 20
rect 340 10 420 20
rect 580 10 660 20
rect 820 10 900 20
rect 1060 10 1140 20
<< labels >>
rlabel metal2 s 100 1470 180 1550 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 100 10 180 90 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 270 150 330 490 4 A
port 1 nsew signal input
rlabel metal2 s 580 270 640 1160 4 Y
port 2 nsew signal output
rlabel metal2 s 890 390 950 490 4 B
port 3 nsew signal input
rlabel metal2 s 260 400 340 480 1 A
port 1 nsew signal input
rlabel metal2 s 270 150 790 210 1 A
port 1 nsew signal input
rlabel metal2 s 730 150 790 750 1 A
port 1 nsew signal input
rlabel metal2 s 720 660 800 740 1 A
port 1 nsew signal input
rlabel metal1 s 250 410 350 470 1 A
port 1 nsew signal input
rlabel metal1 s 710 670 810 730 1 A
port 1 nsew signal input
rlabel metal2 s 880 400 960 480 1 B
port 3 nsew signal input
rlabel metal2 s 870 410 970 470 1 B
port 3 nsew signal input
rlabel metal1 s 870 410 970 470 1 B
port 3 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 580 1470 660 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 570 1480 670 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 820 1470 900 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 810 1480 910 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1060 1470 1140 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 1050 1480 1150 1540 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 280 1060 330 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 900 1060 950 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1470 1240 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 580 10 660 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 20 670 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 820 10 900 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 810 20 910 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1060 10 1140 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 1050 20 1150 80 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 280 -30 330 330 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 900 -30 950 330 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 -30 1240 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 1050 650 1130 1 Y
port 2 nsew signal output
rlabel metal2 s 560 270 660 350 1 Y
port 2 nsew signal output
rlabel metal1 s 580 1030 640 1140 1 Y
port 2 nsew signal output
rlabel metal1 s 590 1030 640 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 590 160 640 360 1 Y
port 2 nsew signal output
rlabel metal1 s 580 250 640 360 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 1240 1590
string GDS_END 443480
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 431954
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
