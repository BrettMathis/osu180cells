magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -141 344 4676
<< polysilicon >>
rect -31 4535 89 4607
rect -31 -74 89 -1
use pmos_5p04310589983291_64x8m81  pmos_5p04310589983291_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 4656
<< properties >>
string GDS_END 650056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 649742
<< end >>
