magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal1 >>
rect 0 362 224 422
rect 0 -30 224 30
<< labels >>
rlabel metal1 s 0 362 224 422 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -30 224 30 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 392
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1127812
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1126780
<< end >>
