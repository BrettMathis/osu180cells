magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 1120 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
rect 870 1090 930 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 870 360
rect 760 252 792 298
rect 838 252 870 298
rect 760 190 870 252
rect 930 298 1030 360
rect 930 252 962 298
rect 1008 252 1030 298
rect 930 190 1030 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 870 1430
rect 760 1143 792 1377
rect 838 1143 870 1377
rect 760 1090 870 1143
rect 930 1377 1030 1430
rect 930 1143 962 1377
rect 1008 1143 1030 1377
rect 930 1090 1030 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
rect 962 252 1008 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
rect 962 1143 1008 1377
<< psubdiff >>
rect 90 98 190 120
rect 90 52 112 98
rect 158 52 190 98
rect 90 30 190 52
rect 330 98 430 120
rect 330 52 352 98
rect 398 52 430 98
rect 330 30 430 52
rect 570 98 670 120
rect 570 52 592 98
rect 638 52 670 98
rect 570 30 670 52
rect 810 98 910 120
rect 810 52 832 98
rect 878 52 910 98
rect 810 30 910 52
<< nsubdiff >>
rect 90 1568 190 1590
rect 90 1522 112 1568
rect 158 1522 190 1568
rect 90 1500 190 1522
rect 330 1568 430 1590
rect 330 1522 352 1568
rect 398 1522 430 1568
rect 330 1500 430 1522
rect 570 1568 670 1590
rect 570 1522 592 1568
rect 638 1522 670 1568
rect 570 1500 670 1522
rect 810 1568 910 1590
rect 810 1522 832 1568
rect 878 1522 910 1568
rect 810 1500 910 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 870 1430 930 1480
rect 190 910 250 1090
rect 360 1070 420 1090
rect 530 1070 590 1090
rect 700 1070 760 1090
rect 870 1070 930 1090
rect 360 1010 930 1070
rect 190 883 310 910
rect 190 837 237 883
rect 283 837 310 883
rect 190 810 310 837
rect 190 360 250 810
rect 360 670 420 1010
rect 300 633 420 670
rect 300 587 327 633
rect 373 587 420 633
rect 300 550 420 587
rect 360 440 420 550
rect 700 440 760 1010
rect 360 380 930 440
rect 360 360 420 380
rect 530 360 590 380
rect 700 360 760 380
rect 870 360 930 380
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
<< polycontact >>
rect 237 837 283 883
rect 327 587 373 633
<< metal1 >>
rect 0 1590 1120 1620
rect -170 1568 1120 1590
rect -170 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1120 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect -170 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1120 1566
rect -170 1500 1120 1514
rect -170 1470 950 1500
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 860 160 1143
rect 280 1377 330 1470
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 1000 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1030 500 1143
rect 620 1377 670 1470
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 1030 670 1143
rect 790 1377 840 1470
rect 790 1143 792 1377
rect 838 1143 840 1377
rect 790 1030 840 1143
rect 960 1377 1010 1500
rect 960 1143 962 1377
rect 1008 1143 1010 1377
rect 960 1090 1010 1143
rect 450 1026 870 1030
rect 450 1000 794 1026
rect 280 974 794 1000
rect 846 974 870 1026
rect 280 970 870 974
rect 280 940 700 970
rect 280 890 330 940
rect 40 800 160 860
rect 210 886 330 890
rect 210 834 234 886
rect 286 834 330 886
rect 210 830 330 834
rect 110 640 160 800
rect 280 640 330 830
rect 110 633 400 640
rect 110 587 327 633
rect 373 587 400 633
rect 110 580 400 587
rect 110 298 160 580
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 430 330 580
rect 450 460 500 940
rect 620 460 670 940
rect 790 460 840 970
rect 450 430 840 460
rect 280 410 840 430
rect 280 380 670 410
rect 280 298 330 380
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 450 298 500 380
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 380
rect 620 252 622 298
rect 668 252 670 298
rect 620 120 670 252
rect 790 298 840 410
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 960 298 1010 360
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 120 1010 252
rect 0 106 1120 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 0 90 112 98
rect -170 52 112 90
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1120 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1120 54
rect -170 0 1120 52
rect -170 -30 950 0
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 794 974 846 1026
rect 234 883 286 886
rect 234 837 237 883
rect 237 837 283 883
rect 283 837 286 883
rect 234 834 286 837
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 90 1566 190 1570
rect -70 1540 10 1550
rect -80 1480 20 1540
rect 90 1514 114 1566
rect 166 1550 190 1566
rect 330 1566 430 1570
rect 166 1540 250 1550
rect 166 1514 260 1540
rect 90 1510 260 1514
rect 330 1514 354 1566
rect 406 1550 430 1566
rect 570 1566 670 1570
rect 406 1540 490 1550
rect 406 1514 500 1540
rect 330 1510 500 1514
rect 570 1514 594 1566
rect 646 1550 670 1566
rect 810 1566 910 1570
rect 646 1540 730 1550
rect 646 1514 740 1540
rect 570 1510 740 1514
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1510 910 1514
rect 100 1500 260 1510
rect 340 1500 500 1510
rect 580 1500 740 1510
rect 820 1500 900 1510
rect 160 1480 260 1500
rect 400 1480 500 1500
rect 640 1480 740 1500
rect -70 1470 10 1480
rect 170 1470 250 1480
rect 410 1470 490 1480
rect 650 1470 730 1480
rect 770 1030 870 1040
rect 760 1026 870 1030
rect 600 1000 700 1010
rect 590 940 700 1000
rect 760 974 794 1026
rect 846 974 870 1026
rect 760 970 870 974
rect 770 960 870 970
rect 600 930 700 940
rect 220 890 300 900
rect 210 886 310 890
rect 50 860 130 870
rect 40 800 140 860
rect 210 834 234 886
rect 286 834 310 886
rect 210 830 310 834
rect 220 820 300 830
rect 50 790 130 800
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 90 106 190 110
rect -70 80 10 90
rect -80 20 20 80
rect 90 54 114 106
rect 166 90 190 106
rect 330 106 430 110
rect 166 80 250 90
rect 166 54 260 80
rect 90 50 260 54
rect 330 54 354 106
rect 406 90 430 106
rect 570 106 670 110
rect 406 80 490 90
rect 406 54 500 80
rect 330 50 500 54
rect 570 54 594 106
rect 646 90 670 106
rect 810 106 910 110
rect 646 80 730 90
rect 646 54 740 80
rect 570 50 740 54
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 100 40 260 50
rect 340 40 500 50
rect 580 40 740 50
rect 820 40 900 50
rect 160 20 260 40
rect 400 20 500 40
rect 640 20 740 40
rect -70 10 10 20
rect 170 10 250 20
rect 410 10 490 20
rect 650 10 730 20
<< labels >>
rlabel metal2 s -70 10 10 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s -70 1470 10 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 50 790 130 870 4 A
port 1 nsew signal input
rlabel metal2 s 590 940 700 1000 4 Y
port 2 nsew signal output
rlabel metal2 s 40 800 140 860 1 A
port 1 nsew signal input
rlabel metal1 s 40 800 140 860 1 A
port 1 nsew signal input
rlabel metal2 s -80 1480 20 1540 3 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 170 1470 250 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 160 1480 260 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 410 1470 490 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 400 1480 500 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 650 1470 730 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 640 1480 740 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 1060 840 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s -170 1470 950 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s -80 20 20 80 3 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 170 10 250 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 160 20 260 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 410 10 490 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 400 20 500 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 650 10 730 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 640 20 740 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 -30 840 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s -170 -30 950 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 600 930 700 1010 1 Y
port 2 nsew signal output
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 380 670 430 1 Y
port 2 nsew signal output
rlabel metal1 s 620 160 670 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 940 700 1000 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX -170 -30 950 1590
string GDS_END 74358
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 65430
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
