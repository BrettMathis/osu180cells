magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 341 89 414
rect 193 341 313 414
use pmos_5p04310590878166_256x8m81  pmos_5p04310590878166_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 462
<< properties >>
string GDS_END 374992
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 374614
<< end >>
