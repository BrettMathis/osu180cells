magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 3136 844
rect 273 610 319 724
rect 360 424 430 550
rect 165 360 430 424
rect 697 617 743 724
rect 273 60 319 163
rect 670 248 886 312
rect 677 60 723 165
rect 800 110 886 248
rect 1541 561 1610 724
rect 2045 506 2091 724
rect 1553 60 1599 179
rect 2248 424 2340 676
rect 2453 506 2499 724
rect 2656 424 2776 676
rect 2861 506 2907 724
rect 2248 360 2776 424
rect 2045 60 2091 211
rect 2248 106 2340 360
rect 2493 60 2539 211
rect 2656 106 2776 360
rect 2941 60 2987 211
rect 0 -60 3136 60
<< obsm1 >>
rect 38 278 115 678
rect 522 417 579 678
rect 1020 628 1301 674
rect 625 467 1020 513
rect 1151 417 1197 562
rect 522 371 1197 417
rect 38 232 472 278
rect 38 106 115 232
rect 522 106 590 371
rect 957 202 1003 371
rect 1255 295 1301 628
rect 1757 461 1803 645
rect 1424 415 1834 461
rect 1255 249 1716 295
rect 1255 152 1301 249
rect 1040 106 1301 152
rect 1766 106 1834 415
<< labels >>
rlabel metal1 s 670 248 886 312 6 D
port 1 nsew default input
rlabel metal1 s 800 110 886 248 6 D
port 1 nsew default input
rlabel metal1 s 360 424 430 550 6 E
port 2 nsew clock input
rlabel metal1 s 165 360 430 424 6 E
port 2 nsew clock input
rlabel metal1 s 2656 424 2776 676 6 Q
port 3 nsew default output
rlabel metal1 s 2248 424 2340 676 6 Q
port 3 nsew default output
rlabel metal1 s 2248 360 2776 424 6 Q
port 3 nsew default output
rlabel metal1 s 2656 106 2776 360 6 Q
port 3 nsew default output
rlabel metal1 s 2248 106 2340 360 6 Q
port 3 nsew default output
rlabel metal1 s 0 724 3136 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2861 617 2907 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2453 617 2499 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2045 617 2091 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 617 1610 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 697 617 743 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 617 319 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2861 610 2907 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2453 610 2499 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2045 610 2091 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 610 1610 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 610 319 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2861 561 2907 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2453 561 2499 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2045 561 2091 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1541 561 1610 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2861 506 2907 561 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2453 506 2499 561 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2045 506 2091 561 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2941 179 2987 211 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2493 179 2539 211 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2045 179 2091 211 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2941 165 2987 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2493 165 2539 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2045 165 2091 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 165 1599 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2941 163 2987 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2493 163 2539 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2045 163 2091 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 163 1599 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 163 723 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2941 60 2987 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2493 60 2539 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2045 60 2091 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 60 1599 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 60 723 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3136 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 586916
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 580658
<< end >>
