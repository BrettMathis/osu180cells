magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect 316 7520 475 7579
rect 316 7474 372 7520
rect 418 7474 475 7520
rect 316 7357 475 7474
rect 316 7311 372 7357
rect 418 7311 475 7357
rect 316 7193 475 7311
rect 316 7147 372 7193
rect 418 7147 475 7193
rect 316 7030 475 7147
rect 316 6984 372 7030
rect 418 6984 475 7030
rect 316 6925 475 6984
<< psubdiffcont >>
rect 372 7474 418 7520
rect 372 7311 418 7357
rect 372 7147 418 7193
rect 372 6984 418 7030
<< polysilicon >>
rect 751 6598 870 6639
rect 1265 6598 1384 6639
rect 465 6552 870 6598
rect 465 6506 539 6552
rect 585 6506 697 6552
rect 743 6506 870 6552
rect 465 6460 870 6506
rect 975 6552 1384 6598
rect 975 6506 1049 6552
rect 1095 6506 1207 6552
rect 1253 6506 1384 6552
rect 975 6460 1384 6506
rect 751 6419 870 6460
rect 1265 6419 1384 6460
<< polycontact >>
rect 539 6506 585 6552
rect 697 6506 743 6552
rect 1049 6506 1095 6552
rect 1207 6506 1253 6552
<< metal1 >>
rect 324 7777 756 7818
rect 324 7725 459 7777
rect 511 7725 666 7777
rect 718 7725 756 7777
rect 324 7670 756 7725
rect 325 7559 756 7670
rect 325 7520 459 7559
rect 325 7474 372 7520
rect 418 7507 459 7520
rect 511 7507 666 7559
rect 718 7507 756 7559
rect 418 7474 756 7507
rect 325 7357 756 7474
rect 325 7311 372 7357
rect 418 7341 756 7357
rect 418 7311 459 7341
rect 325 7289 459 7311
rect 511 7289 666 7341
rect 718 7289 756 7341
rect 325 7193 756 7289
rect 325 7147 372 7193
rect 418 7147 756 7193
rect 325 7123 756 7147
rect 325 7071 459 7123
rect 511 7071 666 7123
rect 718 7071 756 7123
rect 325 7030 756 7071
rect 1148 7777 1276 7817
rect 1148 7725 1186 7777
rect 1238 7725 1276 7777
rect 1148 7559 1276 7725
rect 1148 7507 1186 7559
rect 1238 7507 1276 7559
rect 1148 7341 1276 7507
rect 1148 7289 1186 7341
rect 1238 7289 1276 7341
rect 1148 7123 1276 7289
rect 1148 7071 1186 7123
rect 1238 7071 1276 7123
rect 1148 7031 1276 7071
rect 325 6984 372 7030
rect 418 6984 756 7030
rect 325 6678 756 6984
rect 421 6589 761 6596
rect 865 6589 980 6739
rect 421 6555 778 6589
rect 421 6503 459 6555
rect 511 6552 671 6555
rect 723 6552 778 6555
rect 511 6506 539 6552
rect 585 6506 671 6552
rect 743 6506 778 6552
rect 511 6503 671 6506
rect 723 6503 778 6506
rect 421 6469 778 6503
rect 865 6552 1288 6589
rect 865 6506 1049 6552
rect 1095 6506 1207 6552
rect 1253 6506 1288 6552
rect 865 6469 1288 6506
rect 421 6463 761 6469
rect 351 6344 756 6380
rect 350 6333 756 6344
rect 350 6292 769 6333
rect 865 6315 980 6469
rect 350 6240 679 6292
rect 731 6240 769 6292
rect 350 6075 769 6240
rect 350 6023 679 6075
rect 731 6023 769 6075
rect 350 5857 769 6023
rect 350 5805 679 5857
rect 731 5805 769 5857
rect 350 5639 769 5805
rect 350 5587 679 5639
rect 731 5587 769 5639
rect 350 5421 769 5587
rect 350 5369 679 5421
rect 731 5369 769 5421
rect 350 5204 769 5369
rect 350 5152 679 5204
rect 731 5152 769 5204
rect 350 5112 769 5152
rect 1155 6292 1283 6333
rect 1379 6315 1494 6739
rect 1155 6240 1193 6292
rect 1245 6240 1283 6292
rect 1155 6075 1283 6240
rect 1155 6023 1193 6075
rect 1245 6023 1283 6075
rect 1155 5857 1283 6023
rect 1155 5805 1193 5857
rect 1245 5805 1283 5857
rect 1155 5639 1283 5805
rect 1155 5587 1193 5639
rect 1245 5587 1283 5639
rect 1155 5421 1283 5587
rect 1155 5369 1193 5421
rect 1245 5369 1283 5421
rect 1155 5204 1283 5369
rect 1155 5152 1193 5204
rect 1245 5152 1283 5204
rect 1155 5112 1283 5152
rect 350 5111 763 5112
rect 1161 5111 1277 5112
rect 350 3776 756 5111
rect 351 3676 756 3776
rect 860 3987 984 4027
rect 860 3935 896 3987
rect 948 3935 984 3987
rect 860 3769 984 3935
rect 860 3717 896 3769
rect 948 3717 984 3769
rect 860 3677 984 3717
rect 1374 3987 1498 4027
rect 1374 3935 1410 3987
rect 1462 3935 1498 3987
rect 1374 3769 1498 3935
rect 1374 3717 1410 3769
rect 1462 3717 1498 3769
rect 1374 3677 1498 3717
rect -14 3481 1953 3574
rect -14 3279 1953 3372
rect -14 3078 1953 3170
rect -14 2876 1953 2968
rect -14 2674 1953 2767
rect -14 2472 1953 2565
rect 423 1624 547 1664
rect 423 1572 459 1624
rect 511 1572 547 1624
rect 423 1406 547 1572
rect 423 1354 459 1406
rect 511 1354 547 1406
rect 423 1314 547 1354
<< via1 >>
rect 459 7725 511 7777
rect 666 7725 718 7777
rect 459 7507 511 7559
rect 666 7507 718 7559
rect 459 7289 511 7341
rect 666 7289 718 7341
rect 459 7071 511 7123
rect 666 7071 718 7123
rect 1186 7725 1238 7777
rect 1186 7507 1238 7559
rect 1186 7289 1238 7341
rect 1186 7071 1238 7123
rect 459 6503 511 6555
rect 671 6552 723 6555
rect 671 6506 697 6552
rect 697 6506 723 6552
rect 671 6503 723 6506
rect 679 6240 731 6292
rect 679 6023 731 6075
rect 679 5805 731 5857
rect 679 5587 731 5639
rect 679 5369 731 5421
rect 679 5152 731 5204
rect 1193 6240 1245 6292
rect 1193 6023 1245 6075
rect 1193 5805 1245 5857
rect 1193 5587 1245 5639
rect 1193 5369 1245 5421
rect 1193 5152 1245 5204
rect 896 3935 948 3987
rect 896 3717 948 3769
rect 1410 3935 1462 3987
rect 1410 3717 1462 3769
rect 459 1572 511 1624
rect 459 1354 511 1406
<< metal2 >>
rect 421 7779 756 7818
rect 421 7723 457 7779
rect 513 7723 664 7779
rect 720 7723 756 7779
rect 421 7561 756 7723
rect 421 7505 457 7561
rect 513 7505 664 7561
rect 720 7505 756 7561
rect 421 7343 756 7505
rect 421 7287 457 7343
rect 513 7287 664 7343
rect 720 7287 756 7343
rect 421 7125 756 7287
rect 421 7069 457 7125
rect 513 7069 664 7125
rect 720 7069 756 7125
rect 421 7031 756 7069
rect 1148 7779 1276 7816
rect 1148 7723 1184 7779
rect 1240 7723 1276 7779
rect 1148 7561 1276 7723
rect 1148 7505 1184 7561
rect 1240 7505 1276 7561
rect 1148 7343 1276 7505
rect 1148 7287 1184 7343
rect 1240 7287 1276 7343
rect 1148 7125 1276 7287
rect 1148 7069 1184 7125
rect 1240 7069 1276 7125
rect 1148 7031 1276 7069
rect 421 6555 761 6596
rect 421 6503 459 6555
rect 511 6503 671 6555
rect 723 6503 761 6555
rect 421 6463 761 6503
rect 421 1624 550 6463
rect 641 6294 769 6333
rect 641 6238 677 6294
rect 733 6238 769 6294
rect 641 6077 769 6238
rect 641 6021 677 6077
rect 733 6021 769 6077
rect 641 5859 769 6021
rect 641 5803 677 5859
rect 733 5803 769 5859
rect 641 5641 769 5803
rect 641 5585 677 5641
rect 733 5585 769 5641
rect 641 5423 769 5585
rect 641 5367 677 5423
rect 733 5367 769 5423
rect 641 5206 769 5367
rect 641 5150 677 5206
rect 733 5150 769 5206
rect 641 5111 769 5150
rect 1155 6294 1283 6333
rect 1155 6238 1191 6294
rect 1247 6238 1283 6294
rect 1155 6077 1283 6238
rect 1155 6021 1191 6077
rect 1247 6021 1283 6077
rect 1155 5859 1283 6021
rect 1155 5803 1191 5859
rect 1247 5803 1283 5859
rect 1155 5641 1283 5803
rect 1155 5585 1191 5641
rect 1247 5585 1283 5641
rect 1155 5423 1283 5585
rect 1155 5367 1191 5423
rect 1247 5367 1283 5423
rect 1155 5206 1283 5367
rect 1155 5150 1191 5206
rect 1247 5150 1283 5206
rect 1155 5111 1283 5150
rect 1635 4233 1760 4272
rect 1635 4177 1670 4233
rect 1726 4177 1760 4233
rect 1635 4057 1760 4177
rect 860 3987 984 4027
rect 860 3935 896 3987
rect 948 3935 984 3987
rect 860 3769 984 3935
rect 1374 3987 1498 4027
rect 1374 3935 1410 3987
rect 1462 3935 1498 3987
rect 860 3717 896 3769
rect 948 3717 984 3769
rect 860 3677 984 3717
rect 1144 3757 1272 3796
rect 1144 3701 1180 3757
rect 1236 3701 1272 3757
rect 421 1572 459 1624
rect 511 1572 550 1624
rect 421 1406 550 1572
rect 421 1359 459 1406
rect 423 1354 459 1359
rect 511 1359 550 1406
rect 1144 3539 1272 3701
rect 1374 3769 1498 3935
rect 1374 3717 1410 3769
rect 1462 3717 1498 3769
rect 1374 3677 1498 3717
rect 1633 4015 1762 4057
rect 1633 3959 1670 4015
rect 1726 3959 1762 4015
rect 1144 3483 1180 3539
rect 1236 3483 1272 3539
rect 1144 1413 1272 3483
rect 1633 1615 1762 3959
rect 511 1354 547 1359
rect 423 1314 547 1354
rect 1144 1280 1762 1413
<< via2 >>
rect 457 7777 513 7779
rect 457 7725 459 7777
rect 459 7725 511 7777
rect 511 7725 513 7777
rect 457 7723 513 7725
rect 664 7777 720 7779
rect 664 7725 666 7777
rect 666 7725 718 7777
rect 718 7725 720 7777
rect 664 7723 720 7725
rect 457 7559 513 7561
rect 457 7507 459 7559
rect 459 7507 511 7559
rect 511 7507 513 7559
rect 457 7505 513 7507
rect 664 7559 720 7561
rect 664 7507 666 7559
rect 666 7507 718 7559
rect 718 7507 720 7559
rect 664 7505 720 7507
rect 457 7341 513 7343
rect 457 7289 459 7341
rect 459 7289 511 7341
rect 511 7289 513 7341
rect 457 7287 513 7289
rect 664 7341 720 7343
rect 664 7289 666 7341
rect 666 7289 718 7341
rect 718 7289 720 7341
rect 664 7287 720 7289
rect 457 7123 513 7125
rect 457 7071 459 7123
rect 459 7071 511 7123
rect 511 7071 513 7123
rect 457 7069 513 7071
rect 664 7123 720 7125
rect 664 7071 666 7123
rect 666 7071 718 7123
rect 718 7071 720 7123
rect 664 7069 720 7071
rect 1184 7777 1240 7779
rect 1184 7725 1186 7777
rect 1186 7725 1238 7777
rect 1238 7725 1240 7777
rect 1184 7723 1240 7725
rect 1184 7559 1240 7561
rect 1184 7507 1186 7559
rect 1186 7507 1238 7559
rect 1238 7507 1240 7559
rect 1184 7505 1240 7507
rect 1184 7341 1240 7343
rect 1184 7289 1186 7341
rect 1186 7289 1238 7341
rect 1238 7289 1240 7341
rect 1184 7287 1240 7289
rect 1184 7123 1240 7125
rect 1184 7071 1186 7123
rect 1186 7071 1238 7123
rect 1238 7071 1240 7123
rect 1184 7069 1240 7071
rect 677 6292 733 6294
rect 677 6240 679 6292
rect 679 6240 731 6292
rect 731 6240 733 6292
rect 677 6238 733 6240
rect 677 6075 733 6077
rect 677 6023 679 6075
rect 679 6023 731 6075
rect 731 6023 733 6075
rect 677 6021 733 6023
rect 677 5857 733 5859
rect 677 5805 679 5857
rect 679 5805 731 5857
rect 731 5805 733 5857
rect 677 5803 733 5805
rect 677 5639 733 5641
rect 677 5587 679 5639
rect 679 5587 731 5639
rect 731 5587 733 5639
rect 677 5585 733 5587
rect 677 5421 733 5423
rect 677 5369 679 5421
rect 679 5369 731 5421
rect 731 5369 733 5421
rect 677 5367 733 5369
rect 677 5204 733 5206
rect 677 5152 679 5204
rect 679 5152 731 5204
rect 731 5152 733 5204
rect 677 5150 733 5152
rect 1191 6292 1247 6294
rect 1191 6240 1193 6292
rect 1193 6240 1245 6292
rect 1245 6240 1247 6292
rect 1191 6238 1247 6240
rect 1191 6075 1247 6077
rect 1191 6023 1193 6075
rect 1193 6023 1245 6075
rect 1245 6023 1247 6075
rect 1191 6021 1247 6023
rect 1191 5857 1247 5859
rect 1191 5805 1193 5857
rect 1193 5805 1245 5857
rect 1245 5805 1247 5857
rect 1191 5803 1247 5805
rect 1191 5639 1247 5641
rect 1191 5587 1193 5639
rect 1193 5587 1245 5639
rect 1245 5587 1247 5639
rect 1191 5585 1247 5587
rect 1191 5421 1247 5423
rect 1191 5369 1193 5421
rect 1193 5369 1245 5421
rect 1245 5369 1247 5421
rect 1191 5367 1247 5369
rect 1191 5204 1247 5206
rect 1191 5152 1193 5204
rect 1193 5152 1245 5204
rect 1245 5152 1247 5204
rect 1191 5150 1247 5152
rect 1670 4177 1726 4233
rect 1180 3701 1236 3757
rect 1670 3959 1726 4015
rect 1180 3483 1236 3539
<< metal3 >>
rect 0 7779 1876 7883
rect 0 7723 457 7779
rect 513 7723 664 7779
rect 720 7723 1184 7779
rect 1240 7723 1876 7779
rect 0 7561 1876 7723
rect 0 7505 457 7561
rect 513 7505 664 7561
rect 720 7505 1184 7561
rect 1240 7505 1876 7561
rect 0 7343 1876 7505
rect 0 7287 457 7343
rect 513 7287 664 7343
rect 720 7287 1184 7343
rect 1240 7287 1876 7343
rect 0 7125 1876 7287
rect 0 7069 457 7125
rect 513 7069 664 7125
rect 720 7069 1184 7125
rect 1240 7069 1876 7125
rect 0 6975 1876 7069
rect 0 6294 1901 6636
rect 0 6238 677 6294
rect 733 6238 1191 6294
rect 1247 6238 1901 6294
rect 0 6077 1901 6238
rect 0 6021 677 6077
rect 733 6021 1191 6077
rect 1247 6021 1901 6077
rect 0 5859 1901 6021
rect 0 5803 677 5859
rect 733 5803 1191 5859
rect 1247 5803 1901 5859
rect 0 5641 1901 5803
rect 0 5585 677 5641
rect 733 5585 1191 5641
rect 1247 5585 1901 5641
rect 0 5423 1901 5585
rect 0 5367 677 5423
rect 733 5367 1191 5423
rect 1247 5367 1901 5423
rect 0 5206 1901 5367
rect 0 5150 677 5206
rect 733 5150 1191 5206
rect 1247 5150 1901 5206
rect 0 4458 1901 5150
rect 1635 4233 1761 4272
rect 1635 4177 1670 4233
rect 1726 4177 1761 4233
rect 1635 4163 1761 4177
rect 6 4030 1761 4163
rect 1635 4015 1761 4030
rect 1635 3959 1670 4015
rect 1726 3959 1761 4015
rect 1635 3920 1761 3959
rect 15 3757 1760 3796
rect 15 3701 1180 3757
rect 1236 3701 1760 3757
rect 15 3662 1760 3701
rect 1145 3539 1271 3662
rect 1145 3483 1180 3539
rect 1236 3483 1271 3539
rect 1145 3444 1271 3483
use M1_NWELL$$47822892_128x8m81  M1_NWELL$$47822892_128x8m81_0
timestamp 1669390400
transform 1 0 334 0 1 5060
box -221 -1452 221 1452
use M1_POLY2$$46559276_128x8m81_0  M1_POLY2$$46559276_128x8m81_0_0
timestamp 1669390400
transform 1 0 1151 0 1 6529
box 0 0 1 1
use M1_POLY2$$46559276_128x8m81_0  M1_POLY2$$46559276_128x8m81_0_1
timestamp 1669390400
transform 1 0 641 0 1 6529
box 0 0 1 1
use M1_PSUB$$47818796_128x8m81  M1_PSUB$$47818796_128x8m81_0
timestamp 1669390400
transform 1 0 395 0 1 7252
box 0 0 1 1
use M2_M1$$34864172_128x8m81  M2_M1$$34864172_128x8m81_0
timestamp 1669390400
transform 1 0 591 0 1 6529
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 1489
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1669390400
transform 1 0 922 0 1 3852
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1669390400
transform 1 0 1436 0 1 3852
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 5722
box 0 0 1 1
use M2_M1$$43377708_128x8m81  M2_M1$$43377708_128x8m81_1
timestamp 1669390400
transform 1 0 705 0 1 5722
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7424
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7424
box 0 0 1 1
use M2_M1$$43379756_128x8m81  M2_M1$$43379756_128x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7424
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_0
timestamp 1669390400
transform 1 0 1698 0 1 4096
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_1
timestamp 1669390400
transform 1 0 1208 0 1 3620
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7424
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7424
box 0 0 1 1
use M3_M2$$47333420_128x8m81  M3_M2$$47333420_128x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7424
box 0 0 1 1
use M3_M2$$47334444_128x8m81  M3_M2$$47334444_128x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 5722
box 0 0 1 1
use M3_M2$$47334444_128x8m81  M3_M2$$47334444_128x8m81_1
timestamp 1669390400
transform 1 0 705 0 1 5722
box 0 0 1 1
use alatch_128x8m81  alatch_128x8m81_0
timestamp 1669390400
transform 1 0 70 0 1 -632
box -90 -1 1692 2968
use nmos_1p2$$47514668_128x8m81  nmos_1p2$$47514668_128x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 6670
box -119 -73 177 980
use nmos_1p2$$47514668_128x8m81  nmos_1p2$$47514668_128x8m81_1
timestamp 1669390400
transform 1 0 782 0 1 6670
box -119 -73 177 980
use pmos_1p2$$46887980_128x8m81  pmos_1p2$$46887980_128x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 3668
box -286 -142 344 2862
use pmos_1p2$$46887980_128x8m81  pmos_1p2$$46887980_128x8m81_1
timestamp 1669390400
transform 1 0 782 0 1 3668
box -286 -142 344 2862
<< properties >>
string GDS_END 828400
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 825726
<< end >>
