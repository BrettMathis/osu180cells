magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 111 8 123
rect 0 0 8 12
<< labels >>
rlabel metal1 s 0 111 8 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 0 8 12 6 VSS
port 2 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 8 123
string GDS_END 353318
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 353042
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
