magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 454
<< mvndiff >>
rect -88 441 0 454
rect -88 395 -75 441
rect -29 395 0 441
rect -88 314 0 395
rect -88 268 -75 314
rect -29 268 0 314
rect -88 187 0 268
rect -88 141 -75 187
rect -29 141 0 187
rect -88 59 0 141
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 441 208 454
rect 120 395 149 441
rect 195 395 208 441
rect 120 314 208 395
rect 120 268 149 314
rect 195 268 208 314
rect 120 187 208 268
rect 120 141 149 187
rect 195 141 208 187
rect 120 59 208 141
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 395 -29 441
rect -75 268 -29 314
rect -75 141 -29 187
rect -75 13 -29 59
rect 149 395 195 441
rect 149 268 195 314
rect 149 141 195 187
rect 149 13 195 59
<< polysilicon >>
rect 0 454 120 498
rect 0 -44 120 0
<< metal1 >>
rect -75 441 -29 454
rect -75 314 -29 395
rect -75 187 -29 268
rect -75 59 -29 141
rect -75 0 -29 13
rect 149 441 195 454
rect 149 314 195 395
rect 149 187 195 268
rect 149 59 195 141
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 227 -52 227 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 227 172 227 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 10842
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 9434
<< end >>
