magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 4790 870
<< pwell >>
rect -86 -86 4790 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2812 68 2932 232
rect 3036 68 3156 232
rect 3260 68 3380 232
rect 3484 68 3604 232
rect 3708 68 3828 232
rect 3932 68 4052 232
rect 4156 68 4276 232
rect 4380 68 4500 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
rect 3708 472 3808 716
rect 3932 472 4032 716
rect 4156 472 4256 716
rect 4380 472 4480 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 244 192 348 232
rect 244 146 273 192
rect 319 146 348 192
rect 244 68 348 146
rect 468 127 572 232
rect 468 81 497 127
rect 543 81 572 127
rect 468 68 572 81
rect 692 192 796 232
rect 692 146 721 192
rect 767 146 796 192
rect 692 68 796 146
rect 916 127 1020 232
rect 916 81 945 127
rect 991 81 1020 127
rect 916 68 1020 81
rect 1140 192 1244 232
rect 1140 146 1169 192
rect 1215 146 1244 192
rect 1140 68 1244 146
rect 1364 127 1468 232
rect 1364 81 1393 127
rect 1439 81 1468 127
rect 1364 68 1468 81
rect 1588 192 1692 232
rect 1588 146 1617 192
rect 1663 146 1692 192
rect 1588 68 1692 146
rect 1812 127 1916 232
rect 1812 81 1841 127
rect 1887 81 1916 127
rect 1812 68 1916 81
rect 2036 192 2140 232
rect 2036 146 2065 192
rect 2111 146 2140 192
rect 2036 68 2140 146
rect 2260 127 2364 232
rect 2260 81 2289 127
rect 2335 81 2364 127
rect 2260 68 2364 81
rect 2484 192 2588 232
rect 2484 146 2513 192
rect 2559 146 2588 192
rect 2484 68 2588 146
rect 2708 127 2812 232
rect 2708 81 2737 127
rect 2783 81 2812 127
rect 2708 68 2812 81
rect 2932 192 3036 232
rect 2932 146 2961 192
rect 3007 146 3036 192
rect 2932 68 3036 146
rect 3156 127 3260 232
rect 3156 81 3185 127
rect 3231 81 3260 127
rect 3156 68 3260 81
rect 3380 192 3484 232
rect 3380 146 3409 192
rect 3455 146 3484 192
rect 3380 68 3484 146
rect 3604 127 3708 232
rect 3604 81 3633 127
rect 3679 81 3708 127
rect 3604 68 3708 81
rect 3828 192 3932 232
rect 3828 146 3857 192
rect 3903 146 3932 192
rect 3828 68 3932 146
rect 4052 127 4156 232
rect 4052 81 4081 127
rect 4127 81 4156 127
rect 4052 68 4156 81
rect 4276 192 4380 232
rect 4276 146 4305 192
rect 4351 146 4380 192
rect 4276 68 4380 146
rect 4500 192 4588 232
rect 4500 146 4529 192
rect 4575 146 4588 192
rect 4500 68 4588 146
<< mvpdiff >>
rect 36 687 124 716
rect 36 547 49 687
rect 95 547 124 687
rect 36 472 124 547
rect 224 664 348 716
rect 224 524 273 664
rect 319 524 348 664
rect 224 472 348 524
rect 448 703 572 716
rect 448 657 477 703
rect 523 657 572 703
rect 448 472 572 657
rect 672 664 796 716
rect 672 524 701 664
rect 747 524 796 664
rect 672 472 796 524
rect 896 703 1020 716
rect 896 657 925 703
rect 971 657 1020 703
rect 896 472 1020 657
rect 1120 664 1244 716
rect 1120 524 1149 664
rect 1195 524 1244 664
rect 1120 472 1244 524
rect 1344 703 1468 716
rect 1344 657 1373 703
rect 1419 657 1468 703
rect 1344 472 1468 657
rect 1568 664 1692 716
rect 1568 524 1597 664
rect 1643 524 1692 664
rect 1568 472 1692 524
rect 1792 703 1916 716
rect 1792 657 1821 703
rect 1867 657 1916 703
rect 1792 472 1916 657
rect 2016 664 2140 716
rect 2016 524 2045 664
rect 2091 524 2140 664
rect 2016 472 2140 524
rect 2240 703 2364 716
rect 2240 657 2269 703
rect 2315 657 2364 703
rect 2240 472 2364 657
rect 2464 664 2588 716
rect 2464 524 2493 664
rect 2539 524 2588 664
rect 2464 472 2588 524
rect 2688 703 2812 716
rect 2688 657 2717 703
rect 2763 657 2812 703
rect 2688 472 2812 657
rect 2912 664 3036 716
rect 2912 524 2941 664
rect 2987 524 3036 664
rect 2912 472 3036 524
rect 3136 703 3260 716
rect 3136 657 3165 703
rect 3211 657 3260 703
rect 3136 472 3260 657
rect 3360 664 3484 716
rect 3360 524 3389 664
rect 3435 524 3484 664
rect 3360 472 3484 524
rect 3584 703 3708 716
rect 3584 657 3613 703
rect 3659 657 3708 703
rect 3584 472 3708 657
rect 3808 664 3932 716
rect 3808 524 3837 664
rect 3883 524 3932 664
rect 3808 472 3932 524
rect 4032 703 4156 716
rect 4032 657 4061 703
rect 4107 657 4156 703
rect 4032 472 4156 657
rect 4256 664 4380 716
rect 4256 524 4285 664
rect 4331 524 4380 664
rect 4256 472 4380 524
rect 4480 687 4568 716
rect 4480 547 4509 687
rect 4555 547 4568 687
rect 4480 472 4568 547
<< mvndiffc >>
rect 49 146 95 192
rect 273 146 319 192
rect 497 81 543 127
rect 721 146 767 192
rect 945 81 991 127
rect 1169 146 1215 192
rect 1393 81 1439 127
rect 1617 146 1663 192
rect 1841 81 1887 127
rect 2065 146 2111 192
rect 2289 81 2335 127
rect 2513 146 2559 192
rect 2737 81 2783 127
rect 2961 146 3007 192
rect 3185 81 3231 127
rect 3409 146 3455 192
rect 3633 81 3679 127
rect 3857 146 3903 192
rect 4081 81 4127 127
rect 4305 146 4351 192
rect 4529 146 4575 192
<< mvpdiffc >>
rect 49 547 95 687
rect 273 524 319 664
rect 477 657 523 703
rect 701 524 747 664
rect 925 657 971 703
rect 1149 524 1195 664
rect 1373 657 1419 703
rect 1597 524 1643 664
rect 1821 657 1867 703
rect 2045 524 2091 664
rect 2269 657 2315 703
rect 2493 524 2539 664
rect 2717 657 2763 703
rect 2941 524 2987 664
rect 3165 657 3211 703
rect 3389 524 3435 664
rect 3613 657 3659 703
rect 3837 524 3883 664
rect 4061 657 4107 703
rect 4285 524 4331 664
rect 4509 547 4555 687
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 3708 716 3808 760
rect 3932 716 4032 760
rect 4156 716 4256 760
rect 4380 716 4480 760
rect 124 412 224 472
rect 348 412 448 472
rect 572 412 672 472
rect 796 412 896 472
rect 1020 412 1120 472
rect 1244 412 1344 472
rect 1468 412 1568 472
rect 1692 412 1792 472
rect 1916 412 2016 472
rect 2140 412 2240 472
rect 2364 412 2464 472
rect 2588 412 2688 472
rect 2812 412 2912 472
rect 3036 412 3136 472
rect 3260 412 3360 472
rect 3484 412 3584 472
rect 3708 412 3808 472
rect 3932 412 4032 472
rect 4156 412 4256 472
rect 4380 412 4480 472
rect 124 399 4480 412
rect 124 353 137 399
rect 1593 353 3008 399
rect 4464 353 4480 399
rect 124 340 4480 353
rect 124 232 244 340
rect 348 232 468 340
rect 572 232 692 340
rect 796 232 916 340
rect 1020 232 1140 340
rect 1244 232 1364 340
rect 1468 232 1588 340
rect 1692 232 1812 340
rect 1916 232 2036 340
rect 2140 232 2260 340
rect 2364 232 2484 340
rect 2588 232 2708 340
rect 2812 232 2932 340
rect 3036 232 3156 340
rect 3260 232 3380 340
rect 3484 232 3604 340
rect 3708 232 3828 340
rect 3932 232 4052 340
rect 4156 232 4276 340
rect 4380 288 4480 340
rect 4380 232 4500 288
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2812 24 2932 68
rect 3036 24 3156 68
rect 3260 24 3380 68
rect 3484 24 3604 68
rect 3708 24 3828 68
rect 3932 24 4052 68
rect 4156 24 4276 68
rect 4380 24 4500 68
<< polycontact >>
rect 137 353 1593 399
rect 3008 353 4464 399
<< metal1 >>
rect 0 724 4704 844
rect 49 687 95 724
rect 466 703 534 724
rect 49 528 95 547
rect 273 664 319 675
rect 466 657 477 703
rect 523 657 534 703
rect 914 703 982 724
rect 701 664 747 675
rect 319 524 701 611
rect 914 657 925 703
rect 971 657 982 703
rect 1362 703 1430 724
rect 1149 664 1195 675
rect 747 524 1149 611
rect 1362 657 1373 703
rect 1419 657 1430 703
rect 1810 703 1878 724
rect 1597 664 1643 675
rect 1195 524 1597 611
rect 1810 657 1821 703
rect 1867 657 1878 703
rect 2258 703 2326 724
rect 2045 664 2091 675
rect 1643 524 2045 611
rect 2258 657 2269 703
rect 2315 657 2326 703
rect 2706 703 2774 724
rect 2493 664 2539 675
rect 2091 524 2493 611
rect 2706 657 2717 703
rect 2763 657 2774 703
rect 3154 703 3222 724
rect 2941 664 2987 675
rect 2539 524 2941 611
rect 3154 657 3165 703
rect 3211 657 3222 703
rect 3602 703 3670 724
rect 3389 664 3435 675
rect 2987 524 3389 611
rect 3602 657 3613 703
rect 3659 657 3670 703
rect 4050 703 4118 724
rect 3837 664 3883 675
rect 3435 524 3837 611
rect 4050 657 4061 703
rect 4107 657 4118 703
rect 4509 687 4555 724
rect 4285 664 4331 675
rect 3883 524 4285 611
rect 4509 528 4555 547
rect 273 476 4331 524
rect 1679 463 2933 476
rect 122 399 1604 430
rect 122 353 137 399
rect 1593 353 1604 399
rect 2206 321 2386 463
rect 2997 399 4475 430
rect 2997 353 3008 399
rect 4464 353 4475 399
rect 1683 307 2954 321
rect 49 192 95 203
rect 262 192 4351 307
rect 262 146 273 192
rect 319 173 721 192
rect 319 146 330 173
rect 767 173 1169 192
rect 49 60 95 146
rect 721 135 767 146
rect 1215 173 1617 192
rect 1169 135 1215 146
rect 1663 173 2065 192
rect 1617 135 1663 146
rect 2111 173 2513 192
rect 2065 135 2111 146
rect 2559 173 2961 192
rect 2513 135 2559 146
rect 3007 173 3409 192
rect 2961 135 3007 146
rect 3455 173 3857 192
rect 3409 135 3455 146
rect 3903 173 4305 192
rect 3857 135 3903 146
rect 4305 135 4351 146
rect 4529 192 4575 203
rect 486 81 497 127
rect 543 81 554 127
rect 486 60 554 81
rect 934 81 945 127
rect 991 81 1002 127
rect 934 60 1002 81
rect 1382 81 1393 127
rect 1439 81 1450 127
rect 1382 60 1450 81
rect 1830 81 1841 127
rect 1887 81 1898 127
rect 1830 60 1898 81
rect 2278 81 2289 127
rect 2335 81 2346 127
rect 2278 60 2346 81
rect 2726 81 2737 127
rect 2783 81 2794 127
rect 2726 60 2794 81
rect 3174 81 3185 127
rect 3231 81 3242 127
rect 3174 60 3242 81
rect 3622 81 3633 127
rect 3679 81 3690 127
rect 3622 60 3690 81
rect 4070 81 4081 127
rect 4127 81 4138 127
rect 4070 60 4138 81
rect 4529 60 4575 146
rect 0 -60 4704 60
<< labels >>
flabel metal1 s 4529 127 4575 203 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 4285 611 4331 675 0 FreeSans 400 0 0 0 ZN
port 2 nsew default output
flabel metal1 s 122 353 1604 430 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 4704 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2997 353 4475 430 1 I
port 1 nsew default input
rlabel metal1 s 3837 611 3883 675 1 ZN
port 2 nsew default output
rlabel metal1 s 3389 611 3435 675 1 ZN
port 2 nsew default output
rlabel metal1 s 2941 611 2987 675 1 ZN
port 2 nsew default output
rlabel metal1 s 2493 611 2539 675 1 ZN
port 2 nsew default output
rlabel metal1 s 2045 611 2091 675 1 ZN
port 2 nsew default output
rlabel metal1 s 1597 611 1643 675 1 ZN
port 2 nsew default output
rlabel metal1 s 1149 611 1195 675 1 ZN
port 2 nsew default output
rlabel metal1 s 701 611 747 675 1 ZN
port 2 nsew default output
rlabel metal1 s 273 611 319 675 1 ZN
port 2 nsew default output
rlabel metal1 s 273 476 4331 611 1 ZN
port 2 nsew default output
rlabel metal1 s 1679 463 2933 476 1 ZN
port 2 nsew default output
rlabel metal1 s 2206 321 2386 463 1 ZN
port 2 nsew default output
rlabel metal1 s 1683 307 2954 321 1 ZN
port 2 nsew default output
rlabel metal1 s 262 173 4351 307 1 ZN
port 2 nsew default output
rlabel metal1 s 4305 146 4351 173 1 ZN
port 2 nsew default output
rlabel metal1 s 3857 146 3903 173 1 ZN
port 2 nsew default output
rlabel metal1 s 3409 146 3455 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2961 146 3007 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2513 146 2559 173 1 ZN
port 2 nsew default output
rlabel metal1 s 2065 146 2111 173 1 ZN
port 2 nsew default output
rlabel metal1 s 1617 146 1663 173 1 ZN
port 2 nsew default output
rlabel metal1 s 1169 146 1215 173 1 ZN
port 2 nsew default output
rlabel metal1 s 721 146 767 173 1 ZN
port 2 nsew default output
rlabel metal1 s 262 146 330 173 1 ZN
port 2 nsew default output
rlabel metal1 s 4305 135 4351 146 1 ZN
port 2 nsew default output
rlabel metal1 s 3857 135 3903 146 1 ZN
port 2 nsew default output
rlabel metal1 s 3409 135 3455 146 1 ZN
port 2 nsew default output
rlabel metal1 s 2961 135 3007 146 1 ZN
port 2 nsew default output
rlabel metal1 s 2513 135 2559 146 1 ZN
port 2 nsew default output
rlabel metal1 s 2065 135 2111 146 1 ZN
port 2 nsew default output
rlabel metal1 s 1617 135 1663 146 1 ZN
port 2 nsew default output
rlabel metal1 s 1169 135 1215 146 1 ZN
port 2 nsew default output
rlabel metal1 s 721 135 767 146 1 ZN
port 2 nsew default output
rlabel metal1 s 4509 657 4555 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4050 657 4118 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3602 657 3670 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3154 657 3222 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2706 657 2774 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2258 657 2326 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1810 657 1878 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1362 657 1430 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 914 657 982 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 466 657 534 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 528 4555 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 528 95 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 127 95 203 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 60 4575 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4704 60 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 784
string GDS_END 506656
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 496972
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
