magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 3136 844
rect 273 600 319 724
rect 698 424 809 559
rect 156 364 809 424
rect 402 248 540 318
rect 590 254 642 364
rect 1118 563 1186 724
rect 1526 563 1594 724
rect 1713 514 1759 724
rect 1008 360 1478 424
rect 2151 514 2197 724
rect 2372 468 2444 676
rect 2589 514 2635 724
rect 2793 468 2892 676
rect 2997 514 3043 724
rect 2372 422 3000 468
rect 273 60 319 223
rect 465 110 540 248
rect 1082 60 1150 213
rect 2934 278 3000 422
rect 2365 232 3000 278
rect 1693 60 1739 177
rect 2141 60 2187 177
rect 2365 109 2411 232
rect 2589 60 2635 177
rect 2813 109 2859 232
rect 3037 60 3083 177
rect 0 -60 3136 60
<< obsm1 >>
rect 38 516 115 676
rect 632 619 912 665
rect 38 470 632 516
rect 38 163 106 470
rect 864 314 912 619
rect 1333 516 1379 676
rect 962 470 1594 516
rect 1526 372 1594 470
rect 1917 468 1963 676
rect 1917 422 2179 468
rect 2133 372 2179 422
rect 1526 326 2072 372
rect 2133 326 2874 372
rect 864 268 1306 314
rect 864 212 912 268
rect 690 166 912 212
rect 1526 106 1594 326
rect 2133 278 2179 326
rect 1917 232 2179 278
rect 1917 109 1963 232
<< labels >>
rlabel metal1 s 402 248 540 318 6 D
port 1 nsew default input
rlabel metal1 s 465 110 540 248 6 D
port 1 nsew default input
rlabel metal1 s 698 424 809 559 6 E
port 2 nsew clock input
rlabel metal1 s 156 364 809 424 6 E
port 2 nsew clock input
rlabel metal1 s 590 254 642 364 6 E
port 2 nsew clock input
rlabel metal1 s 1008 360 1478 424 6 SETN
port 3 nsew default input
rlabel metal1 s 2793 468 2892 676 6 Q
port 4 nsew default output
rlabel metal1 s 2372 468 2444 676 6 Q
port 4 nsew default output
rlabel metal1 s 2372 422 3000 468 6 Q
port 4 nsew default output
rlabel metal1 s 2934 278 3000 422 6 Q
port 4 nsew default output
rlabel metal1 s 2365 232 3000 278 6 Q
port 4 nsew default output
rlabel metal1 s 2813 109 2859 232 6 Q
port 4 nsew default output
rlabel metal1 s 2365 109 2411 232 6 Q
port 4 nsew default output
rlabel metal1 s 0 724 3136 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2997 600 3043 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2589 600 2635 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2151 600 2197 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1713 600 1759 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 600 1594 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1118 600 1186 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 600 319 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2997 563 3043 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2589 563 2635 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2151 563 2197 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1713 563 1759 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 563 1594 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1118 563 1186 600 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2997 514 3043 563 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2589 514 2635 563 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2151 514 2197 563 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1713 514 1759 563 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 213 319 223 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1082 177 1150 213 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 177 319 213 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3037 60 3083 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2589 60 2635 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2141 60 2187 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1693 60 1739 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1082 60 1150 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 177 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3136 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 648044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 640586
<< end >>
