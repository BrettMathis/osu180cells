magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 960 1620
<< nmos >>
rect 190 190 250 360
rect 530 190 590 360
rect 700 190 760 360
<< pmos >>
rect 190 1090 250 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 350 360
rect 250 252 282 298
rect 328 252 350 298
rect 250 190 350 252
rect 430 298 530 360
rect 430 252 452 298
rect 498 252 530 298
rect 430 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 860 360
rect 760 252 792 298
rect 838 252 860 298
rect 760 190 860 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 350 1430
rect 250 1143 282 1377
rect 328 1143 350 1377
rect 250 1090 350 1143
rect 430 1377 530 1430
rect 430 1143 452 1377
rect 498 1143 530 1377
rect 430 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 860 1430
rect 760 1143 792 1377
rect 838 1143 860 1377
rect 760 1090 860 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
<< psubdiff >>
rect 90 98 190 120
rect 90 52 112 98
rect 158 52 190 98
rect 90 30 190 52
rect 330 98 430 120
rect 330 52 352 98
rect 398 52 430 98
rect 330 30 430 52
rect 570 98 670 120
rect 570 52 592 98
rect 638 52 670 98
rect 570 30 670 52
<< nsubdiff >>
rect 90 1568 190 1590
rect 90 1522 112 1568
rect 158 1522 190 1568
rect 90 1500 190 1522
rect 330 1568 430 1590
rect 330 1522 352 1568
rect 398 1522 430 1568
rect 330 1500 430 1522
rect 570 1568 670 1590
rect 570 1522 592 1568
rect 638 1522 670 1568
rect 570 1500 670 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 190 1060 250 1090
rect 530 1060 590 1090
rect 190 1010 590 1060
rect 190 650 250 1010
rect 300 890 400 920
rect 700 890 760 1090
rect 300 883 760 890
rect 300 837 327 883
rect 373 837 760 883
rect 300 830 760 837
rect 300 800 400 830
rect 120 630 250 650
rect 120 628 760 630
rect 120 582 142 628
rect 188 582 760 628
rect 120 580 760 582
rect 120 560 250 580
rect 190 360 250 560
rect 300 493 400 530
rect 300 447 327 493
rect 373 490 400 493
rect 373 447 590 490
rect 300 440 590 447
rect 300 410 400 440
rect 530 360 590 440
rect 700 360 760 580
rect 190 140 250 190
rect 530 140 590 190
rect 700 140 760 190
<< polycontact >>
rect 327 837 373 883
rect 142 582 188 628
rect 327 447 373 493
<< metal1 >>
rect 0 1590 960 1620
rect -20 1568 960 1590
rect -20 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 960 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect -20 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 960 1566
rect -20 1500 960 1514
rect -20 1470 940 1500
rect 90 1377 160 1470
rect 90 1143 112 1377
rect 158 1143 160 1377
rect 90 1090 160 1143
rect 280 1377 330 1430
rect 450 1400 500 1430
rect 620 1400 670 1430
rect 790 1400 840 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 90 1060 140 1090
rect 280 890 330 1143
rect 430 1377 500 1400
rect 430 1143 452 1377
rect 498 1143 500 1377
rect 280 883 400 890
rect 280 837 327 883
rect 373 837 400 883
rect 280 830 400 837
rect 110 628 210 630
rect 110 626 142 628
rect 110 600 134 626
rect 90 574 134 600
rect 188 582 210 628
rect 186 574 210 582
rect 90 570 210 574
rect 90 540 190 570
rect 280 500 330 830
rect 430 770 500 1143
rect 600 1377 670 1400
rect 600 1143 622 1377
rect 668 1143 670 1377
rect 600 1030 670 1143
rect 770 1377 840 1400
rect 770 1143 792 1377
rect 838 1143 840 1377
rect 600 1016 700 1030
rect 600 1000 624 1016
rect 580 964 624 1000
rect 676 964 700 1016
rect 580 950 700 964
rect 580 920 680 950
rect 430 756 570 770
rect 430 704 494 756
rect 546 704 570 756
rect 430 690 570 704
rect 430 660 550 690
rect 280 493 400 500
rect 280 447 327 493
rect 373 447 400 493
rect 280 440 400 447
rect 110 330 160 360
rect 90 298 160 330
rect 90 252 112 298
rect 158 252 160 298
rect 90 120 160 252
rect 280 298 330 440
rect 280 252 282 298
rect 328 252 330 298
rect 280 190 330 252
rect 430 298 500 660
rect 430 252 452 298
rect 498 252 500 298
rect 430 190 500 252
rect 600 298 670 920
rect 770 900 840 1143
rect 750 886 850 900
rect 750 870 774 886
rect 730 834 774 870
rect 826 834 850 886
rect 730 820 850 834
rect 730 790 840 820
rect 600 252 622 298
rect 668 252 670 298
rect 600 190 670 252
rect 770 298 840 790
rect 770 252 792 298
rect 838 252 840 298
rect 770 190 840 252
rect 430 160 480 190
rect 600 160 650 190
rect 770 160 820 190
rect 0 106 960 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 0 90 112 98
rect -20 52 112 90
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 960 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 960 54
rect -20 0 960 52
rect -20 -30 940 0
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 134 582 142 626
rect 142 582 186 626
rect 134 574 186 582
rect 624 964 676 1016
rect 494 704 546 756
rect 774 834 826 886
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 90 1566 190 1570
rect 90 1550 114 1566
rect 80 1540 114 1550
rect 70 1514 114 1540
rect 166 1514 190 1566
rect 330 1566 430 1570
rect 330 1550 354 1566
rect 320 1540 354 1550
rect 70 1510 190 1514
rect 310 1514 354 1540
rect 406 1514 430 1566
rect 570 1566 670 1570
rect 570 1550 594 1566
rect 560 1540 594 1550
rect 310 1510 430 1514
rect 550 1514 594 1540
rect 646 1514 670 1566
rect 550 1510 670 1514
rect 70 1500 180 1510
rect 310 1500 420 1510
rect 550 1500 660 1510
rect 70 1480 170 1500
rect 310 1480 410 1500
rect 550 1480 650 1500
rect 80 1470 160 1480
rect 320 1470 400 1480
rect 560 1470 640 1480
rect 600 1016 700 1030
rect 600 1000 624 1016
rect 580 964 624 1000
rect 676 964 700 1016
rect 580 950 700 964
rect 580 920 680 950
rect 750 886 850 900
rect 750 870 774 886
rect 730 834 774 870
rect 826 834 850 886
rect 730 820 850 834
rect 730 790 830 820
rect 470 756 570 770
rect 470 740 494 756
rect 450 704 494 740
rect 546 704 570 756
rect 450 690 570 704
rect 450 660 550 690
rect 110 626 210 640
rect 110 610 134 626
rect 90 574 134 610
rect 186 574 210 626
rect 90 560 210 574
rect 90 530 190 560
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 90 106 190 110
rect 90 90 114 106
rect 80 80 114 90
rect 70 54 114 80
rect 166 54 190 106
rect 330 106 430 110
rect 330 90 354 106
rect 320 80 354 90
rect 70 50 190 54
rect 310 54 354 80
rect 406 54 430 106
rect 570 106 670 110
rect 570 90 594 106
rect 560 80 594 90
rect 310 50 430 54
rect 550 54 594 80
rect 646 54 670 106
rect 550 50 670 54
rect 70 40 180 50
rect 310 40 420 50
rect 550 40 660 50
rect 70 20 170 40
rect 310 20 410 40
rect 550 20 650 40
rect 80 10 160 20
rect 320 10 400 20
rect 560 10 640 20
<< labels >>
rlabel metal2 s 80 10 160 90 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 80 1470 160 1550 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 920 680 1000 4 Y
port 1 nsew signal output
rlabel metal2 s 90 530 190 610 4 Sel
port 2 nsew signal output
rlabel metal2 s 450 660 550 740 4 A
port 3 nsew signal input
rlabel metal2 s 730 790 830 870 4 B
port 4 nsew signal input
rlabel metal1 s 430 160 480 1400 1 A
port 3 nsew signal input
rlabel metal1 s 430 660 550 740 1 A
port 3 nsew signal input
rlabel metal1 s 770 160 820 1400 1 B
port 4 nsew signal input
rlabel metal1 s 730 790 830 870 1 B
port 4 nsew signal input
rlabel metal1 s 90 540 190 600 1 Sel
port 2 nsew signal output
rlabel metal2 s 70 1480 170 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 320 1470 400 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 310 1480 410 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 560 1470 640 1550 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 550 1480 650 1540 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 90 1060 140 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s -20 1470 940 1590 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 70 20 170 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 320 10 400 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 310 20 410 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 560 10 640 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 550 20 650 80 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 90 -30 140 330 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s -20 -30 940 90 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 600 160 650 1400 1 Y
port 1 nsew signal output
rlabel metal1 s 580 920 680 1000 1 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX -20 -30 940 1590
string GDS_END 401092
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 392854
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
