* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addf_1 B CI CO S VDD VSS A
X0 a_680_156# B a_512_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X1 CO a_952_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 a_1992_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X3 VSS A a_1072_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X4 a_3048_156# B a_952_112# VSUBS nmos_6p0 w=0.38u l=0.6u
X5 VSS CI a_1072_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X6 a_2012_472# A VDD w_n86_352# pmos_6p0 w=0.7u l=0.5u
X7 a_1072_496# B VDD w_n86_352# pmos_6p0 w=0.66u l=0.5u
X8 a_512_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X9 a_124_46# CI a_680_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X10 a_3028_472# B a_952_112# w_n86_352# pmos_6p0 w=0.7u l=0.5u
X11 VDD CI a_1072_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X12 a_1072_156# B VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X13 a_680_496# B a_512_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X14 a_1072_156# a_952_112# a_124_46# VSUBS nmos_6p0 w=0.38u l=0.6u
X15 VSS A a_3048_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X16 VDD A a_1072_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X17 a_952_112# CI a_1992_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X18 VDD a_124_46# S w_n86_352# pmos_6p0 w=1.215u l=0.5u
X19 VDD A a_3028_472# w_n86_352# pmos_6p0 w=0.7u l=0.5u
X20 a_952_112# CI a_2012_472# w_n86_352# pmos_6p0 w=0.7u l=0.5u
X21 CO a_952_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X22 VDD B a_2012_472# w_n86_352# pmos_6p0 w=0.7u l=0.5u
X23 VSS a_124_46# S VSUBS nmos_6p0 w=0.71u l=0.6u
X24 a_1072_496# a_952_112# a_124_46# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X25 a_512_496# A VDD w_n86_352# pmos_6p0 w=0.66u l=0.5u
X26 VSS B a_1992_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X27 a_124_46# CI a_680_156# VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addf_2 VDD B CI CO S VSS A
X0 S a_132_24# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X1 a_912_156# B a_744_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_1284_492# a_1184_112# a_132_24# w_n86_352# pmos_6p0 w=0.68u l=0.5u
X3 a_1184_112# CI a_2248_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X4 CO a_1184_112# VDD w_n86_352# pmos_6p0 w=1.195u l=0.5u
X5 VDD a_1184_112# CO w_n86_352# pmos_6p0 w=1.195u l=0.5u
X6 a_1284_492# B VDD w_n86_352# pmos_6p0 w=0.68u l=0.5u
X7 VSS A a_3216_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X8 a_912_492# B a_744_492# w_n86_352# pmos_6p0 w=0.68u l=0.5u
X9 a_3216_472# B a_1184_112# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X10 VSS B a_2248_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X11 S a_132_24# VDD w_n86_352# pmos_6p0 w=1.12u l=0.5u
X12 VDD CI a_1284_492# w_n86_352# pmos_6p0 w=0.68u l=0.5u
X13 VSS CI a_1304_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X14 VDD A a_1284_492# w_n86_352# pmos_6p0 w=0.68u l=0.5u
X15 VDD A a_3216_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X16 VSS A a_1304_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X17 VDD B a_2248_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X18 a_3216_156# B a_1184_112# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 VDD a_132_24# S w_n86_352# pmos_6p0 w=1.12u l=0.5u
X20 a_744_492# A VDD w_n86_352# pmos_6p0 w=0.68u l=0.5u
X21 a_744_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X22 a_1304_156# a_1184_112# a_132_24# VSUBS nmos_6p0 w=0.38u l=0.6u
X23 a_2248_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X24 CO a_1184_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X25 a_2248_472# A VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X26 a_1184_112# CI a_2248_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X27 VSS a_132_24# S VSUBS nmos_6p0 w=0.815u l=0.6u
X28 a_1304_156# B VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X29 a_132_24# CI a_912_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X30 VSS a_1184_112# CO VSUBS nmos_6p0 w=0.815u l=0.6u
X31 a_132_24# CI a_912_492# w_n86_352# pmos_6p0 w=0.68u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addf_4 B CI CO S VDD VSS A
X0 a_1640_112# CI a_2748_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X1 VSS a_1640_112# CO VSUBS nmos_6p0 w=0.815u l=0.6u
X2 VSS a_1640_112# CO VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_1200_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X4 VDD a_140_24# S w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_140_24# CI a_1368_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X6 VDD a_1640_112# CO w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 S a_140_24# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X8 VSS A a_3696_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X9 VDD A a_1760_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X10 a_2728_156# A VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X11 CO a_1640_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_1368_496# B a_1200_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X13 VSS B a_2728_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X14 a_1760_156# a_1640_112# a_140_24# VSUBS nmos_6p0 w=0.38u l=0.6u
X15 CO a_1640_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X16 VDD A a_3676_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X17 a_2748_472# A VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X18 a_3696_156# B a_1640_112# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 a_3676_472# B a_1640_112# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X20 S a_140_24# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X21 CO a_1640_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X22 S a_140_24# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X23 VDD a_140_24# S w_n86_352# pmos_6p0 w=1.095u l=0.5u
X24 a_1760_496# a_1640_112# a_140_24# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X25 a_1200_496# A VDD w_n86_352# pmos_6p0 w=0.66u l=0.5u
X26 a_1760_496# B VDD w_n86_352# pmos_6p0 w=0.66u l=0.5u
X27 VDD a_1640_112# CO w_n86_352# pmos_6p0 w=1.215u l=0.5u
X28 a_140_24# CI a_1368_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X29 VDD CI a_1760_496# w_n86_352# pmos_6p0 w=0.66u l=0.5u
X30 S a_140_24# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X31 CO a_1640_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X32 VSS a_140_24# S VSUBS nmos_6p0 w=0.815u l=0.6u
X33 a_1640_112# CI a_2728_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X34 a_1760_156# B VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X35 VSS CI a_1760_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X36 VDD B a_2748_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X37 VSS a_140_24# S VSUBS nmos_6p0 w=0.815u l=0.6u
X38 a_1368_156# B a_1200_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X39 VSS A a_1760_156# VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addf_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addh_1 CO S VDD VSS A B
X0 VSS a_124_24# a_844_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X1 VDD B a_124_24# w_n86_352# pmos_6p0 w=0.635u l=0.5u
X2 S a_1052_148# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_1052_148# A a_1052_589# w_n86_352# pmos_6p0 w=0.635u l=0.5u
X4 a_844_148# A a_1052_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X5 S a_1052_148# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_1052_589# B VDD w_n86_352# pmos_6p0 w=0.635u l=0.5u
X7 a_124_24# B a_516_136# VSUBS nmos_6p0 w=0.48u l=0.6u
X8 a_516_136# A VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X9 VDD a_124_24# CO w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD a_124_24# a_1052_148# w_n86_352# pmos_6p0 w=0.635u l=0.5u
X11 VSS a_124_24# CO VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_124_24# A VDD w_n86_352# pmos_6p0 w=0.635u l=0.5u
X13 a_1052_148# B a_844_148# VSUBS nmos_6p0 w=0.42u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addh_2 CO S VDD VSS A B
X0 a_128_24# A VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X1 VDD B a_128_24# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 a_1064_69# A a_1272_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_128_24# B a_696_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X4 VDD a_128_24# CO w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 a_1272_520# B VDD w_n86_352# pmos_6p0 w=0.975u l=0.5u
X6 S a_1272_69# VDD w_n86_352# pmos_6p0 w=0.975u l=0.5u
X7 VDD a_128_24# a_1272_69# w_n86_352# pmos_6p0 w=0.975u l=0.5u
X8 CO a_128_24# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 a_696_69# A VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X10 CO a_128_24# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X11 a_1272_69# B a_1064_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X12 VSS a_128_24# a_1064_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X13 a_1272_69# A a_1272_520# w_n86_352# pmos_6p0 w=0.975u l=0.5u
X14 VSS a_128_24# CO VSUBS nmos_6p0 w=0.815u l=0.6u
X15 VSS a_1272_69# S VSUBS nmos_6p0 w=0.815u l=0.6u
X16 S a_1272_69# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X17 VDD a_1272_69# S w_n86_352# pmos_6p0 w=0.975u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__addh_4 B CO S VDD VSS A
X0 VSS A a_672_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VSS a_224_518# a_1126_156# VSUBS nmos_6p0 w=0.61u l=0.6u
X2 VDD a_1116_518# S w_n86_352# pmos_6p0 w=0.99u l=0.5u
X3 a_672_68# B a_224_518# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 CO a_224_518# VSS VSUBS nmos_6p0 w=1.05u l=0.6u
X5 S a_1116_518# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 S a_1116_518# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD B a_1330_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X8 a_1910_518# B VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X9 S a_1116_518# VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X10 a_1126_156# a_224_518# VSS VSUBS nmos_6p0 w=0.61u l=0.6u
X11 VSS a_224_518# CO VSUBS nmos_6p0 w=1.05u l=0.6u
X12 VSS a_1116_518# S VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD a_224_518# CO w_n86_352# pmos_6p0 w=0.99u l=0.5u
X14 a_224_518# B VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X15 a_1126_156# B a_1116_518# VSUBS nmos_6p0 w=0.61u l=0.6u
X16 a_1126_156# A a_1116_518# VSUBS nmos_6p0 w=0.61u l=0.6u
X17 VDD a_224_518# a_1116_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X18 a_244_68# A VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 VDD A a_224_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X20 CO a_224_518# VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X21 S a_1116_518# VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X22 a_1330_518# A a_1116_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X23 VDD a_224_518# CO w_n86_352# pmos_6p0 w=0.99u l=0.5u
X24 VDD B a_224_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X25 VSS a_224_518# CO VSUBS nmos_6p0 w=1.05u l=0.6u
X26 a_224_518# A VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X27 a_1116_518# a_224_518# VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X28 a_224_518# B a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X29 a_1116_518# B a_1126_156# VSUBS nmos_6p0 w=0.61u l=0.6u
X30 a_1116_518# A a_1126_156# VSUBS nmos_6p0 w=0.61u l=0.6u
X31 a_1116_518# A a_1910_518# w_n86_352# pmos_6p0 w=0.99u l=0.5u
X32 CO a_224_518# VSS VSUBS nmos_6p0 w=1.05u l=0.6u
X33 VDD a_1116_518# S w_n86_352# pmos_6p0 w=0.99u l=0.5u
X34 CO a_224_518# VDD w_n86_352# pmos_6p0 w=0.99u l=0.5u
X35 VSS a_1116_518# S VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__addh_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2
X0 a_244_159# A1 a_36_159# VSUBS nmos_6p0 w=0.365u l=0.6u
X1 a_36_159# A1 VDD w_n86_352# pmos_6p0 w=0.6u l=0.5u
X2 VDD A2 a_36_159# w_n86_352# pmos_6p0 w=0.6u l=0.5u
X3 Z a_36_159# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 Z a_36_159# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X5 VSS A2 a_244_159# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 VDD VSS Z A1 A2
X0 a_247_68# A1 a_39_68# VSUBS nmos_6p0 w=0.815u l=0.6u
X1 Z a_39_68# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 Z a_39_68# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X3 VDD a_39_68# Z w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 a_39_68# A1 VDD w_n86_352# pmos_6p0 w=1.07u l=0.5u
X5 VSS a_39_68# Z VSUBS nmos_6p0 w=0.815u l=0.6u
X6 VDD A2 a_39_68# w_n86_352# pmos_6p0 w=1.07u l=0.5u
X7 VSS A2 a_247_68# VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A2 VDD VSS Z A1
X0 VSS A2 a_659_69# VSUBS nmos_6p0 w=0.775u l=0.6u
X1 a_224_490# A1 VDD w_n86_352# pmos_6p0 w=1.125u l=0.5u
X2 Z a_224_490# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 VDD A2 a_224_490# w_n86_352# pmos_6p0 w=1.125u l=0.5u
X4 VDD a_224_490# Z w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 Z a_224_490# VSS VSUBS nmos_6p0 w=0.775u l=0.6u
X6 Z a_224_490# VSS VSUBS nmos_6p0 w=0.775u l=0.6u
X7 VSS a_224_490# Z VSUBS nmos_6p0 w=0.775u l=0.6u
X8 a_224_490# A1 a_244_69# VSUBS nmos_6p0 w=0.775u l=0.6u
X9 a_659_69# A1 a_224_490# VSUBS nmos_6p0 w=0.775u l=0.6u
X10 a_244_69# A2 VSS VSUBS nmos_6p0 w=0.775u l=0.6u
X11 a_224_490# A2 VDD w_n86_352# pmos_6p0 w=1.125u l=0.5u
X12 Z a_224_490# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X13 VSS a_224_490# Z VSUBS nmos_6p0 w=0.775u l=0.6u
X14 VDD A1 a_224_490# w_n86_352# pmos_6p0 w=1.125u l=0.5u
X15 VDD a_224_490# Z w_n86_352# pmos_6p0 w=1.215u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2
X0 VDD A1 a_36_148# w_n86_352# pmos_6p0 w=0.535u l=0.5u
X1 a_36_148# A2 VDD w_n86_352# pmos_6p0 w=0.535u l=0.5u
X2 VDD A3 a_36_148# w_n86_352# pmos_6p0 w=0.535u l=0.5u
X3 Z a_36_148# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 a_428_148# A2 a_244_148# VSUBS nmos_6p0 w=0.38u l=0.6u
X5 Z a_36_148# VSS VSUBS nmos_6p0 w=0.775u l=0.6u
X6 VSS A3 a_428_148# VSUBS nmos_6p0 w=0.38u l=0.6u
X7 a_244_148# A1 a_36_148# VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A3 VDD VSS Z A1 A2
X0 Z a_47_69# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X1 Z a_47_69# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 VDD A1 a_47_69# w_n86_352# pmos_6p0 w=0.985u l=0.5u
X3 a_47_69# A2 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X4 VDD a_47_69# Z w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 VSS a_47_69# Z VSUBS nmos_6p0 w=0.815u l=0.6u
X6 VSS A3 a_439_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X7 VDD A3 a_47_69# w_n86_352# pmos_6p0 w=0.985u l=0.5u
X8 a_255_69# A1 a_47_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X9 a_439_69# A2 a_255_69# VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A2 A3 VDD VSS Z A1
X0 a_224_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_224_472# Z VSUBS nmos_6p0 w=0.76u l=0.6u
X2 VSS a_224_472# Z VSUBS nmos_6p0 w=0.76u l=0.6u
X3 VDD A2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_260_69# A3 VSS VSUBS nmos_6p0 w=0.76u l=0.6u
X5 VSS A3 a_1040_69# VSUBS nmos_6p0 w=0.76u l=0.6u
X6 a_224_472# A1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_856_69# A1 a_224_472# VSUBS nmos_6p0 w=0.76u l=0.6u
X8 VDD A1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 Z a_224_472# VSS VSUBS nmos_6p0 w=0.76u l=0.6u
X10 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_224_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 Z a_224_472# VSS VSUBS nmos_6p0 w=0.76u l=0.6u
X13 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_224_472# A1 a_428_69# VSUBS nmos_6p0 w=0.76u l=0.6u
X15 VDD A3 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_428_69# A2 a_260_69# VSUBS nmos_6p0 w=0.76u l=0.6u
X17 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 a_1040_69# A2 a_856_69# VSUBS nmos_6p0 w=0.76u l=0.6u
X19 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and3_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A3 A4 VDD VSS Z A1 A2
X0 a_256_148# A1 a_48_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X1 a_48_148# A1 VDD w_n86_352# pmos_6p0 w=0.6u l=0.5u
X2 a_440_148# A2 a_256_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X3 Z a_48_148# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X4 VDD A2 a_48_148# w_n86_352# pmos_6p0 w=0.6u l=0.5u
X5 Z a_48_148# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_644_148# A3 a_440_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X7 a_48_148# A3 VDD w_n86_352# pmos_6p0 w=0.6u l=0.5u
X8 VSS A4 a_644_148# VSUBS nmos_6p0 w=0.42u l=0.6u
X9 VDD A4 a_48_148# w_n86_352# pmos_6p0 w=0.6u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A3 A4 VDD VSS Z A1 A2
X0 Z a_47_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_643_68# A3 a_439_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_255_68# A1 a_47_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_439_68# A2 a_255_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS a_47_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_47_68# A1 VDD w_n86_352# pmos_6p0 w=0.855u l=0.5u
X6 Z a_47_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD A2 a_47_68# w_n86_352# pmos_6p0 w=0.855u l=0.5u
X8 VSS A4 a_643_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_47_68# A3 VDD w_n86_352# pmos_6p0 w=0.855u l=0.5u
X10 VDD a_47_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VDD A4 a_47_68# w_n86_352# pmos_6p0 w=0.855u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A2 A3 A4 VDD VSS Z A1
X0 Z a_227_494# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_227_494# Z VSUBS nmos_6p0 w=0.645u l=0.6u
X2 VDD A1 a_227_494# w_n86_352# pmos_6p0 w=1.11u l=0.5u
X3 a_227_494# A1 VDD w_n86_352# pmos_6p0 w=1.11u l=0.5u
X4 VDD a_227_494# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_635_68# A2 a_431_68# VSUBS nmos_6p0 w=0.645u l=0.6u
X6 VDD A2 a_227_494# w_n86_352# pmos_6p0 w=1.11u l=0.5u
X7 a_247_68# A4 VSS VSUBS nmos_6p0 w=0.645u l=0.6u
X8 a_227_494# A3 VDD w_n86_352# pmos_6p0 w=1.11u l=0.5u
X9 VDD A4 a_227_494# w_n86_352# pmos_6p0 w=1.11u l=0.5u
X10 a_1451_68# A3 a_1247_68# VSUBS nmos_6p0 w=0.645u l=0.6u
X11 Z a_227_494# VSS VSUBS nmos_6p0 w=0.645u l=0.6u
X12 a_1247_68# A2 a_1063_68# VSUBS nmos_6p0 w=0.645u l=0.6u
X13 a_227_494# A1 a_635_68# VSUBS nmos_6p0 w=0.645u l=0.6u
X14 a_227_494# A4 VDD w_n86_352# pmos_6p0 w=1.11u l=0.5u
X15 Z a_227_494# VSS VSUBS nmos_6p0 w=0.645u l=0.6u
X16 VDD A3 a_227_494# w_n86_352# pmos_6p0 w=1.11u l=0.5u
X17 a_1063_68# A1 a_227_494# VSUBS nmos_6p0 w=0.645u l=0.6u
X18 Z a_227_494# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_431_68# A3 a_247_68# VSUBS nmos_6p0 w=0.645u l=0.6u
X20 VSS a_227_494# Z VSUBS nmos_6p0 w=0.645u l=0.6u
X21 a_227_494# A2 VDD w_n86_352# pmos_6p0 w=1.11u l=0.5u
X22 VDD a_227_494# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VSS A4 a_1451_68# VSUBS nmos_6p0 w=0.645u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__and4_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__antenna.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD
D0 VSUBS I np_6p0 pj=1.86u area=0.2052p
D1 I w_n86_352# pn_6p0 pj=1.86u area=0.2052p
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__antenna.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2
X0 VDD B a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X1 ZN A2 a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 a_36_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 VSS B ZN VSUBS nmos_6p0 w=0.51u l=0.6u
X4 ZN A1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_244_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2
X0 ZN A2 a_49_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X1 VSS B ZN VSUBS nmos_6p0 w=0.565u l=0.6u
X2 ZN A1 a_741_69# VSUBS nmos_6p0 w=0.775u l=0.6u
X3 a_1133_69# A1 ZN VSUBS nmos_6p0 w=0.775u l=0.6u
X4 VSS A2 a_1133_69# VSUBS nmos_6p0 w=0.775u l=0.6u
X5 VDD B a_49_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 ZN A1 a_49_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 a_741_69# A2 VSS VSUBS nmos_6p0 w=0.775u l=0.6u
X8 a_49_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 ZN B VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X10 a_49_472# A2 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X11 a_49_472# B VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A2 B VDD VSS ZN A1
X0 a_288_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_1072_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS B ZN VSUBS nmos_6p0 w=0.51u l=0.6u
X3 a_76_476# A1 ZN w_n86_352# pmos_6p0 w=1.2u l=0.5u
X4 ZN A1 a_288_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN A1 a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X6 a_76_476# A2 ZN w_n86_352# pmos_6p0 w=1.2u l=0.5u
X7 a_76_476# B VDD w_n86_352# pmos_6p0 w=1.2u l=0.5u
X8 ZN B VSS VSUBS nmos_6p0 w=0.51u l=0.6u
X9 a_680_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD B a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X11 VDD B a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X12 a_76_476# B VDD w_n86_352# pmos_6p0 w=1.2u l=0.5u
X13 ZN B VSS VSUBS nmos_6p0 w=0.51u l=0.6u
X14 ZN A2 a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X15 a_76_476# A1 ZN w_n86_352# pmos_6p0 w=1.2u l=0.5u
X16 a_1464_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 ZN A1 a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X18 VSS A2 a_1464_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_76_476# A2 ZN w_n86_352# pmos_6p0 w=1.2u l=0.5u
X20 VSS A2 a_680_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X21 ZN A2 a_76_476# w_n86_352# pmos_6p0 w=1.2u l=0.5u
X22 VSS B ZN VSUBS nmos_6p0 w=0.51u l=0.6u
X23 ZN A1 a_1072_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi21_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2
X0 a_665_69# A1 ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X1 VSS A2 a_665_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X2 ZN B1 a_257_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X3 VDD B2 a_49_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 a_49_472# B1 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 ZN A1 a_49_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 a_49_472# A2 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 a_257_69# B2 VSS VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 B1 B2 VDD VSS ZN A1 A2
X0 VSS B2 a_659_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X1 VDD B2 a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 ZN A1 a_1060_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_36_472# B1 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 a_1060_69# A2 VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X5 VDD B1 a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 VSS A2 a_1468_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X7 a_36_472# B2 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X8 ZN A2 a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 a_36_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X10 ZN B1 a_244_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X11 a_659_69# B1 ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_244_69# B2 VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X13 ZN A1 a_36_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X14 a_1468_69# A1 ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X15 a_36_472# A2 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A2 B1 B2 VDD VSS ZN A1
X0 VSS B2 a_1468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN A2 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_36_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VDD B2 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_36_497# B1 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_2356_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD B1 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 ZN B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_244_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_1468_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_36_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 ZN A1 a_2764_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_2764_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD B2 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 ZN A1 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 ZN A1 a_1948_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_652_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VSS B2 a_652_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VSS A2 a_3260_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_36_497# A2 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 a_3260_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_36_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X22 a_36_497# B1 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 ZN B1 a_1060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X24 ZN A1 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X25 a_1948_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X26 VSS A2 a_2356_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X27 a_1060_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X28 VDD B1 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X29 ZN A2 a_36_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X30 a_36_497# A2 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X31 a_36_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi22_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 B C VDD VSS ZN A1 A2
X0 ZN C VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X1 ZN A2 a_37_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 VSS B ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_37_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 VDD C a_653_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 a_245_90# A2 VSS VSUBS nmos_6p0 w=0.71u l=0.6u
X6 ZN A1 a_245_90# VSUBS nmos_6p0 w=0.71u l=0.6u
X7 a_653_472# B a_37_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2
X0 a_36_488# B a_1492_488# w_n86_352# pmos_6p0 w=1.14u l=0.5u
X1 a_636_68# A1 ZN VSUBS nmos_6p0 w=0.78u l=0.6u
X2 a_1492_488# C VDD w_n86_352# pmos_6p0 w=1.14u l=0.5u
X3 VSS A2 a_636_68# VSUBS nmos_6p0 w=0.78u l=0.6u
X4 VSS B ZN VSUBS nmos_6p0 w=0.515u l=0.6u
X5 VSS C ZN VSUBS nmos_6p0 w=0.515u l=0.6u
X6 a_244_68# A2 VSS VSUBS nmos_6p0 w=0.78u l=0.6u
X7 ZN A1 a_244_68# VSUBS nmos_6p0 w=0.78u l=0.6u
X8 ZN C VSS VSUBS nmos_6p0 w=0.515u l=0.6u
X9 VDD C a_1044_488# w_n86_352# pmos_6p0 w=1.14u l=0.5u
X10 ZN A1 a_36_488# w_n86_352# pmos_6p0 w=1.14u l=0.5u
X11 ZN B VSS VSUBS nmos_6p0 w=0.515u l=0.6u
X12 a_36_488# A2 ZN w_n86_352# pmos_6p0 w=1.14u l=0.5u
X13 ZN A2 a_36_488# w_n86_352# pmos_6p0 w=1.14u l=0.5u
X14 a_1044_488# B a_36_488# w_n86_352# pmos_6p0 w=1.14u l=0.5u
X15 a_36_488# A1 ZN w_n86_352# pmos_6p0 w=1.14u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1
X0 a_170_472# A2 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS B ZN VSUBS nmos_6p0 w=0.46u l=0.6u
X2 a_786_69# A1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X3 a_3662_472# C VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN A2 a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_170_472# B a_3662_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_1194_69# A2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X7 ZN A1 a_1194_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X8 VSS C ZN VSUBS nmos_6p0 w=0.46u l=0.6u
X9 a_170_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN B VSS VSUBS nmos_6p0 w=0.46u l=0.6u
X11 a_3126_472# B a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN A1 a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 ZN A1 a_358_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X14 ZN C VSS VSUBS nmos_6p0 w=0.46u l=0.6u
X15 VDD C a_3126_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 VSS A2 a_1602_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X17 VSS B ZN VSUBS nmos_6p0 w=0.46u l=0.6u
X18 a_1602_69# A1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X19 a_170_472# A2 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 a_2034_472# B a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_2590_472# C VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 a_358_69# A2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X23 VSS A2 a_786_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X24 a_170_472# B a_2590_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X25 VSS C ZN VSUBS nmos_6p0 w=0.46u l=0.6u
X26 ZN B VSS VSUBS nmos_6p0 w=0.46u l=0.6u
X27 ZN A2 a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 a_170_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 ZN C VSS VSUBS nmos_6p0 w=0.46u l=0.6u
X30 VDD C a_2034_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 ZN A1 a_170_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi211_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 B2 C VDD VSS ZN A1 A2 B1
X0 a_940_90# A2 VSS VSUBS nmos_6p0 w=0.71u l=0.6u
X1 VSS C ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X2 a_672_472# C a_56_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 VDD B2 a_56_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 ZN A1 a_940_90# VSUBS nmos_6p0 w=0.71u l=0.6u
X5 a_56_472# B1 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 a_672_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 ZN A2 a_672_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X8 a_244_90# B2 VSS VSUBS nmos_6p0 w=0.71u l=0.6u
X9 ZN B1 a_244_90# VSUBS nmos_6p0 w=0.71u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 B1 B2 VDD VSS ZN A1 A2 C
X0 a_244_492# C a_56_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X1 ZN A2 a_56_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X2 VDD B2 a_244_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X3 ZN A1 a_56_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X4 a_56_492# A1 ZN w_n86_352# pmos_6p0 w=1.12u l=0.5u
X5 a_56_492# A2 ZN w_n86_352# pmos_6p0 w=1.12u l=0.5u
X6 a_512_68# B2 VSS VSUBS nmos_6p0 w=0.715u l=0.6u
X7 ZN C VSS VSUBS nmos_6p0 w=0.575u l=0.6u
X8 a_244_492# B2 VDD w_n86_352# pmos_6p0 w=1.12u l=0.5u
X9 a_948_68# B1 ZN VSUBS nmos_6p0 w=0.715u l=0.6u
X10 VSS B2 a_948_68# VSUBS nmos_6p0 w=0.715u l=0.6u
X11 a_56_492# C a_244_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X12 VSS C ZN VSUBS nmos_6p0 w=0.405u l=0.6u
X13 VDD B1 a_244_492# w_n86_352# pmos_6p0 w=1.12u l=0.5u
X14 a_2267_68# A2 VSS VSUBS nmos_6p0 w=0.715u l=0.6u
X15 a_1875_68# A1 ZN VSUBS nmos_6p0 w=0.715u l=0.6u
X16 VSS A2 a_1875_68# VSUBS nmos_6p0 w=0.715u l=0.6u
X17 ZN A1 a_2267_68# VSUBS nmos_6p0 w=0.715u l=0.6u
X18 a_244_492# B1 VDD w_n86_352# pmos_6p0 w=1.12u l=0.5u
X19 ZN B1 a_512_68# VSUBS nmos_6p0 w=0.715u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A2 B1 B2 C VDD VSS ZN A1
X0 a_1478_69# B2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X1 VDD B1 a_234_508# w_n86_352# pmos_6p0 w=1.035u l=0.5u
X2 ZN A1 a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 ZN C VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X4 a_3320_69# A2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X5 ZN A1 a_3320_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X6 a_234_508# B1 VDD w_n86_352# pmos_6p0 w=1.035u l=0.5u
X7 ZN C VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X8 a_1822_472# C a_234_508# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 a_1822_472# A2 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X10 ZN B1 a_662_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X11 a_662_69# B2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X12 VSS C ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X13 a_1822_472# C a_234_508# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X14 ZN A2 a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X15 a_4136_69# A2 VSS VSUBS nmos_6p0 w=0.77u l=0.6u
X16 VSS B2 a_1070_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X17 VDD B2 a_234_508# w_n86_352# pmos_6p0 w=1.035u l=0.5u
X18 VSS A2 a_3728_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X19 a_234_508# C a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X20 a_1822_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X21 a_234_508# C a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X22 ZN A2 a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X23 a_1070_69# B1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X24 a_234_508# B2 VDD w_n86_352# pmos_6p0 w=1.035u l=0.5u
X25 ZN A1 a_1822_472# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X26 a_1822_472# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X27 VDD B1 a_234_508# w_n86_352# pmos_6p0 w=1.035u l=0.5u
X28 a_1822_472# A2 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X29 a_2912_69# A1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X30 VSS A2 a_2912_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X31 a_234_508# B1 VDD w_n86_352# pmos_6p0 w=1.035u l=0.5u
X32 a_3728_69# A1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X33 ZN A1 a_4136_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X34 a_244_69# B1 ZN VSUBS nmos_6p0 w=0.77u l=0.6u
X35 VSS C ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X36 VDD B2 a_234_508# w_n86_352# pmos_6p0 w=1.035u l=0.5u
X37 ZN B1 a_1478_69# VSUBS nmos_6p0 w=0.77u l=0.6u
X38 a_234_508# B2 VDD w_n86_352# pmos_6p0 w=1.035u l=0.5u
X39 VSS B2 a_244_69# VSUBS nmos_6p0 w=0.77u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi221_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 VSS VDD C2 C1 B2 B1 A2 A1 ZN
X0 VSS B2 a_744_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VDD C1 a_255_484# w_n86_352# pmos_6p0 w=1.16u l=0.5u
X2 ZN A2 a_619_484# w_n86_352# pmos_6p0 w=1.16u l=0.5u
X3 a_744_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_291_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_1235_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_619_484# A1 ZN w_n86_352# pmos_6p0 w=1.16u l=0.5u
X7 a_255_484# B1 a_619_484# w_n86_352# pmos_6p0 w=1.16u l=0.5u
X8 a_619_484# B2 a_255_484# w_n86_352# pmos_6p0 w=1.16u l=0.5u
X9 a_255_484# C2 VDD w_n86_352# pmos_6p0 w=1.16u l=0.5u
X10 ZN C1 a_291_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 ZN A1 a_1235_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 B2 B1 A2 A1 ZN VSS VDD C2 C1
X0 a_1191_68# B1 ZN VSUBS nmos_6p0 w=0.8u l=0.6u
X1 a_1619_68# B2 VSS VSUBS nmos_6p0 w=0.8u l=0.6u
X2 ZN A1 a_2438_68# VSUBS nmos_6p0 w=0.8u l=0.6u
X3 a_231_472# B1 a_1003_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_697_68# C2 VSS VSUBS nmos_6p0 w=0.8u l=0.6u
X5 a_1003_472# A2 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS C2 a_251_68# VSUBS nmos_6p0 w=0.8u l=0.6u
X7 ZN C1 a_697_68# VSUBS nmos_6p0 w=0.8u l=0.6u
X8 a_231_472# C1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_1003_472# B2 a_231_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN A2 a_1003_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN A1 a_1003_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 VSS B2 a_1191_68# VSUBS nmos_6p0 w=0.8u l=0.6u
X13 a_231_472# B2 a_1003_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_1003_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VDD C2 a_231_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_231_472# C2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 ZN B1 a_1619_68# VSUBS nmos_6p0 w=0.8u l=0.6u
X18 VDD C1 a_231_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_2438_68# A2 VSS VSUBS nmos_6p0 w=0.8u l=0.6u
X20 a_2030_68# A1 ZN VSUBS nmos_6p0 w=0.8u l=0.6u
X21 a_251_68# C1 ZN VSUBS nmos_6p0 w=0.8u l=0.6u
X22 a_1003_472# B1 a_231_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VSS A2 a_2030_68# VSUBS nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 ZN VSS VDD C2 C1 B2 B1 A2
X0 ZN C1 a_1468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_1812_472# A2 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 ZN B1 a_2428_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A2 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN A1 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS A2 a_4468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_224_472# C1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_1812_472# A2 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN B1 a_3244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_3244_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD C2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS B2 a_2836_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN A2 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_224_472# C2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 ZN A1 a_4876_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1812_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_2010_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VSS A2 a_3652_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VSS C2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_3652_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD C1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_244_68# C1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_1812_472# B2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 a_1468_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 a_2428_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_224_472# C1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X26 a_4468_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X27 a_224_472# B2 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 a_224_472# B1 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 a_4060_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X30 a_1812_472# B1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 a_652_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X32 ZN C1 a_652_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X33 VDD C2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X34 a_2836_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X35 a_224_472# B2 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X36 a_224_472# B1 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X37 VSS C2 a_1060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X38 a_224_472# C2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X39 VSS B2 a_2010_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X40 a_4876_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X41 a_1812_472# B1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X42 VDD C1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X43 a_1812_472# B2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X44 a_1060_68# C1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X45 ZN A1 a_4060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X46 ZN A1 a_1812_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X47 a_1812_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__aoi222_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD
X0 Z a_36_160# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 Z a_36_160# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VDD I a_36_160# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X3 VSS I a_36_160# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD
X0 VDD I a_36_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_36_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_36_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 Z a_36_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD
X0 VDD I a_36_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_36_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_36_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 Z a_36_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_36_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 Z a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 Z a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS
X0 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS
X0 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 Z I VDD VSS
X0 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X17 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X19 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X23 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X26 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X30 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X32 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X33 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X34 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X35 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 Z I VDD VSS
X0 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X10 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X19 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X26 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X27 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X29 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X31 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X32 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X33 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X34 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X35 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X36 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X37 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X38 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X39 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X40 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X41 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X42 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X43 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X44 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X45 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X46 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X47 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_20.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 VDD VSS Z I
X0 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X13 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X25 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X26 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X31 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X32 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X33 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X34 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X35 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X36 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X37 a_224_472# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X38 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X39 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X40 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X41 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X42 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X43 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X44 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X45 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X46 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X47 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X48 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X49 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X50 a_224_472# I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X51 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X52 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X53 VDD I a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X54 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X55 VDD a_224_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X56 VSS a_224_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X57 Z a_224_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X58 Z a_224_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X59 VSS I a_224_472# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__buf_20.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_1 EN VDD VSS Z I
X0 Z a_468_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 Z a_448_592# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_468_93# a_36_93# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X3 VDD EN a_36_93# w_n86_352# pmos_6p0 w=0.62u l=0.5u
X4 a_448_592# EN a_468_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 a_448_592# EN VDD w_n86_352# pmos_6p0 w=0.62u l=0.5u
X6 VSS EN a_36_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_468_93# a_36_93# a_448_592# w_n86_352# pmos_6p0 w=0.62u l=0.5u
X8 VSS I a_468_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 VDD I a_448_592# w_n86_352# pmos_6p0 w=0.62u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_2 I VDD VSS EN Z
X0 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X1 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X4 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X5 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_476_527# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD EN a_36_68# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X8 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X11 a_468_68# a_36_68# a_476_527# w_n86_352# pmos_6p0 w=0.945u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_3 EN VDD VSS Z I
X0 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X1 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X4 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X5 a_476_527# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD EN a_36_68# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X7 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS I a_468_68# VSUBS nmos_6p0 w=0.54u l=0.6u
X9 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.01u l=0.5u
X10 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X11 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.01u l=0.5u
X12 a_468_68# I VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X13 a_468_68# a_36_68# a_476_527# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X14 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_4 Z EN I VSS VDD
X0 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X1 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X3 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X4 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X5 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X6 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_476_527# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD EN a_36_68# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X9 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X10 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X13 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X14 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_468_68# a_36_68# a_476_527# w_n86_352# pmos_6p0 w=0.945u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_8 Z EN I VSS VDD
X0 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X2 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X4 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X7 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X8 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X10 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_476_527# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VDD EN a_36_68# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X13 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X14 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X15 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X19 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X20 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X21 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X22 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X23 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X25 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X26 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X27 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X28 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X29 a_468_68# a_36_68# a_476_527# w_n86_352# pmos_6p0 w=0.945u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_12 VDD VSS I Z EN
X0 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X2 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X3 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X5 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X6 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X7 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X9 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X11 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X12 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X16 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_476_527# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD EN a_36_68# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X19 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X20 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X24 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X25 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X26 VSS I a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X27 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X28 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X29 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X30 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X31 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X32 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X33 a_468_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X35 a_468_68# a_36_68# a_476_527# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X36 Z a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X37 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X38 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X39 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X40 VSS a_468_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X41 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_16 I VDD VSS Z EN
X0 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X1 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.15u l=0.5u
X3 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X4 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.15u l=0.5u
X6 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.15u l=0.5u
X8 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.15u l=0.5u
X9 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X10 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X12 a_468_69# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.15u l=0.5u
X15 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X17 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X18 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.15u l=0.5u
X20 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X21 VSS I a_468_69# VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD EN a_36_69# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X23 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X24 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_476_527# I VDD w_n86_352# pmos_6p0 w=1.15u l=0.5u
X26 VSS I a_468_69# VSUBS nmos_6p0 w=0.82u l=0.6u
X27 VSS I a_468_69# VSUBS nmos_6p0 w=0.82u l=0.6u
X28 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X29 a_468_69# a_36_69# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X30 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X31 a_476_527# EN VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X32 VDD I a_476_527# w_n86_352# pmos_6p0 w=1.175u l=0.5u
X33 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X34 VSS I a_468_69# VSUBS nmos_6p0 w=0.82u l=0.6u
X35 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X36 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X37 a_468_69# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X38 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X39 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X40 a_468_69# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X41 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X42 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X43 a_476_527# EN a_468_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X44 Z a_476_527# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X45 a_468_69# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X46 VSS EN a_36_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X47 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X48 a_468_69# a_36_69# a_476_527# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X49 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X50 VDD a_476_527# Z w_n86_352# pmos_6p0 w=1.175u l=0.5u
X51 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X52 Z a_468_69# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X53 VSS a_468_69# Z VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__bufz_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD
X0 Z a_36_113# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 Z a_36_113# VSS VSUBS nmos_6p0 w=0.495u l=0.6u
X2 VSS I a_36_113# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 VDD I a_36_113# w_n86_352# pmos_6p0 w=1.05u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I
X0 Z a_36_160# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_36_160# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X2 Z a_36_160# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X3 VDD I a_36_160# w_n86_352# pmos_6p0 w=1.02u l=0.5u
X4 VSS I a_36_160# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VDD a_36_160# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I
X0 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X1 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_224_552# I VSS VSUBS nmos_6p0 w=0.605u l=0.6u
X3 Z a_224_552# VSS VSUBS nmos_6p0 w=0.455u l=0.6u
X4 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X6 VSS a_224_552# Z VSUBS nmos_6p0 w=0.455u l=0.6u
X7 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VSS a_224_552# Z VSUBS nmos_6p0 w=0.455u l=0.6u
X9 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 Z a_224_552# VSS VSUBS nmos_6p0 w=0.455u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I
X0 Z a_224_552# VSS VSUBS nmos_6p0 w=0.455u l=0.6u
X1 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X2 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 Z a_224_552# VSS VSUBS nmos_6p0 w=0.455u l=0.6u
X4 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X6 a_224_552# I VSS VSUBS nmos_6p0 w=0.605u l=0.6u
X7 VSS a_224_552# Z VSUBS nmos_6p0 w=0.455u l=0.6u
X8 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VSS a_224_552# Z VSUBS nmos_6p0 w=0.455u l=0.6u
X10 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I
X0 Z a_224_552# VSS VSUBS nmos_6p0 w=0.43u l=0.6u
X1 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_224_552# I VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X3 VSS a_224_552# Z VSUBS nmos_6p0 w=0.43u l=0.6u
X4 Z a_224_552# VSS VSUBS nmos_6p0 w=0.43u l=0.6u
X5 VSS a_224_552# Z VSUBS nmos_6p0 w=0.43u l=0.6u
X6 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X8 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X9 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS I a_224_552# VSUBS nmos_6p0 w=0.405u l=0.6u
X12 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X13 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VSS a_224_552# Z VSUBS nmos_6p0 w=0.43u l=0.6u
X15 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 Z a_224_552# VSS VSUBS nmos_6p0 w=0.43u l=0.6u
X17 VSS a_224_552# Z VSUBS nmos_6p0 w=0.43u l=0.6u
X18 Z a_224_552# VSS VSUBS nmos_6p0 w=0.43u l=0.6u
X19 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X21 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 a_224_552# I VSS VSUBS nmos_6p0 w=0.405u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 VDD VSS Z I
X0 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X2 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X3 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X7 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X9 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
X10 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
X11 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X12 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X13 VSS I a_224_552# VSUBS nmos_6p0 w=0.365u l=0.6u
X14 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
X15 a_224_552# I VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X16 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VSS I a_224_552# VSUBS nmos_6p0 w=0.365u l=0.6u
X19 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X20 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
X22 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X24 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X25 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
X26 a_224_552# I VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X27 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X28 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X30 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 a_224_552# I VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X32 Z a_224_552# VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X33 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X34 VSS a_224_552# Z VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I
X0 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X2 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X3 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X7 a_224_552# I VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X8 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X9 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X10 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X12 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X13 VSS I a_224_552# VSUBS nmos_6p0 w=0.405u l=0.6u
X14 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X15 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X16 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X18 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X22 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X24 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X25 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X26 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X28 VSS I a_224_552# VSUBS nmos_6p0 w=0.405u l=0.6u
X29 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X30 a_224_552# I VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X31 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X32 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X33 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X34 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X35 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X36 VSS I a_224_552# VSUBS nmos_6p0 w=0.405u l=0.6u
X37 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X38 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X39 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X40 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
X41 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X42 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X43 a_224_552# I VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X44 Z a_224_552# VSS VSUBS nmos_6p0 w=0.485u l=0.6u
X45 VSS a_224_552# Z VSUBS nmos_6p0 w=0.485u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_20.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 VDD VSS Z I
X0 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X2 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X4 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS I a_224_552# VSUBS nmos_6p0 w=0.38u l=0.6u
X6 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X7 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X8 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_224_552# I VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X10 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X11 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X12 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X14 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X15 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X16 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X17 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X19 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X23 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X25 a_224_552# I VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X26 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X28 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X30 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X31 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X32 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X33 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X34 VSS I a_224_552# VSUBS nmos_6p0 w=0.38u l=0.6u
X35 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X36 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X37 a_224_552# I VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X38 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X39 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X40 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X41 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X42 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X43 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X44 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X45 VSS I a_224_552# VSUBS nmos_6p0 w=0.38u l=0.6u
X46 a_224_552# I VDD w_n86_352# pmos_6p0 w=0.82u l=0.5u
X47 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X48 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X49 VDD I a_224_552# w_n86_352# pmos_6p0 w=0.82u l=0.5u
X50 Z a_224_552# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X51 VSS I a_224_552# VSUBS nmos_6p0 w=0.38u l=0.6u
X52 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X53 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
X54 VDD a_224_552# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X55 Z a_224_552# VSS VSUBS nmos_6p0 w=0.47u l=0.6u
X56 a_224_552# I VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X57 VSS a_224_552# Z VSUBS nmos_6p0 w=0.47u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkbuf_20.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X2 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X3 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 VDD ZN I VSS
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X4 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 VDD VSS ZN I
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X3 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X5 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X6 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 VDD VSS ZN I
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X4 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X6 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X7 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X9 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X11 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X13 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 VDD VSS ZN I
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X2 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X3 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X5 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X8 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X11 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X12 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X13 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X15 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X19 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X20 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_16 VDD VSS ZN I
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X5 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X6 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X10 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X11 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X13 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X15 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X16 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X17 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X19 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X20 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X21 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X25 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X26 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X27 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X29 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_20.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 VDD VSS ZN I
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X3 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X6 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X7 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X9 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X12 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X14 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X15 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X16 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X18 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X20 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X21 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X24 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X25 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X26 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X28 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X32 ZN I VSS VSUBS nmos_6p0 w=0.48u l=0.6u
X33 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X34 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X35 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X36 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
X37 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X38 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X39 VSS I ZN VSUBS nmos_6p0 w=0.48u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__clkinv_20.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 CLKN VDD VSS D Q
X0 a_1301_500# a_474_472# a_1070_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X1 VDD a_2406_24# a_2238_185# w_n86_352# pmos_6p0 w=1.075u l=0.5u
X2 VDD CLKN a_62_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X3 VDD a_1358_112# a_1301_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X4 a_2406_24# a_1993_500# VDD w_n86_352# pmos_6p0 w=1.075u l=0.5u
X5 a_474_472# a_62_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X6 Q a_2406_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_1993_500# a_474_472# a_1358_112# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X8 a_862_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2238_185# a_62_124# a_1993_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X10 a_474_472# a_62_124# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X11 a_1358_112# a_1070_500# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_2406_24# a_1993_500# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X13 VSS a_1358_112# a_1310_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1310_156# a_62_124# a_1070_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_2238_185# a_474_472# a_1993_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 Q a_2406_24# VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X17 VSS a_2406_24# a_2238_185# VSUBS nmos_6p0 w=0.63u l=0.6u
X18 VSS CLKN a_62_124# VSUBS nmos_6p0 w=0.465u l=0.6u
X19 a_862_156# D VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X20 a_1358_112# a_1070_500# VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X21 a_1070_500# a_62_124# a_862_156# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X22 a_1070_500# a_474_472# a_862_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_1993_500# a_62_124# a_1358_112# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D Q VDD VSS CLKN
X0 Q a_2432_24# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 a_1301_500# a_474_472# a_1070_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X2 VDD a_2432_24# a_2238_185# w_n86_352# pmos_6p0 w=1.075u l=0.5u
X3 VDD CLKN a_62_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X4 VDD a_2432_24# Q w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 VDD a_1358_112# a_1301_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X6 a_2432_24# a_1993_500# VDD w_n86_352# pmos_6p0 w=1.075u l=0.5u
X7 a_474_472# a_62_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X8 Q a_2432_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_1993_500# a_474_472# a_1358_112# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X10 a_862_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_2238_185# a_62_124# a_1993_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X12 a_474_472# a_62_124# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X13 a_1358_112# a_1070_500# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VSS a_1358_112# a_1310_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_1310_156# a_62_124# a_1070_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2238_185# a_474_472# a_1993_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 VSS a_2432_24# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_2432_24# a_1993_500# VSS VSUBS nmos_6p0 w=0.945u l=0.6u
X19 VSS CLKN a_62_124# VSUBS nmos_6p0 w=0.465u l=0.6u
X20 a_862_156# D VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X21 a_1358_112# a_1070_500# VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X22 a_1070_500# a_62_124# a_862_156# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X23 a_1070_500# a_474_472# a_862_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X24 a_1993_500# a_62_124# a_1358_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 VSS a_2432_24# a_2238_185# VSUBS nmos_6p0 w=0.945u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_4 D Q VDD VSS CLKN
X0 a_1301_500# a_474_472# a_1070_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X1 VDD a_2432_24# a_2238_185# w_n86_352# pmos_6p0 w=1.075u l=0.5u
X2 VDD CLKN a_62_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X3 VDD a_1358_112# a_1301_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X4 a_2432_24# a_1993_500# VDD w_n86_352# pmos_6p0 w=1.075u l=0.5u
X5 a_474_472# a_62_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X6 VSS a_2432_24# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_1993_500# a_474_472# a_1358_112# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X8 a_862_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2238_185# a_62_124# a_1993_500# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X10 a_474_472# a_62_124# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X11 a_1358_112# a_1070_500# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VSS a_1358_112# a_1310_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 VDD a_2432_24# Q w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 Q a_2432_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1310_156# a_62_124# a_1070_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2238_185# a_474_472# a_1993_500# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 VDD a_2432_24# Q w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 a_2432_24# a_1993_500# VSS VSUBS nmos_6p0 w=0.945u l=0.6u
X19 Q a_2432_24# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 VSS CLKN a_62_124# VSUBS nmos_6p0 w=0.465u l=0.6u
X21 a_862_156# D VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X22 VSS a_2432_24# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_1358_112# a_1070_500# VDD w_n86_352# pmos_6p0 w=0.495u l=0.5u
X24 a_1070_500# a_62_124# a_862_156# w_n86_352# pmos_6p0 w=0.495u l=0.5u
X25 Q a_2432_24# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X26 a_1070_500# a_474_472# a_862_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 a_1993_500# a_62_124# a_1358_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 Q a_2432_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X29 VSS a_2432_24# a_2238_185# VSUBS nmos_6p0 w=0.945u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D VSS CLKN RN Q VDD
X0 a_3030_156# RN VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X1 a_2268_156# a_36_124# a_1356_112# VSUBS nmos_6p0 w=0.39u l=0.6u
X2 a_2268_156# a_448_472# a_1356_112# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X3 a_1476_156# a_1356_112# a_1304_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X4 a_1024_476# a_36_124# a_820_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X5 a_1356_112# a_1024_476# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X6 VDD a_2268_156# a_2682_301# w_n86_352# pmos_6p0 w=0.94u l=0.5u
X7 VSS a_2682_301# a_2563_527# VSUBS nmos_6p0 w=0.39u l=0.6u
X8 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.405u l=0.6u
X9 a_1228_476# a_448_472# a_1024_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X10 a_1228_476# RN VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
X11 a_1356_112# a_1024_476# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X12 a_1024_476# a_448_472# a_820_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X13 VDD a_2682_301# a_2563_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X14 a_2682_301# RN VDD w_n86_352# pmos_6p0 w=0.94u l=0.5u
X15 a_1304_156# a_36_124# a_1024_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X16 Q a_2682_301# VSS VSUBS nmos_6p0 w=0.795u l=0.6u
X17 VDD a_1356_112# a_1228_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X18 a_2563_527# a_448_472# a_2268_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X19 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X20 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X21 a_2563_527# a_36_124# a_2268_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X22 a_820_476# D VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X23 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X24 Q a_2682_301# VDD w_n86_352# pmos_6p0 w=1.175u l=0.5u
X25 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X26 a_2682_301# a_2268_156# a_3030_156# VSUBS nmos_6p0 w=0.4u l=0.6u
X27 a_820_476# D VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 D Q RN VDD VSS CLKN
X0 a_3030_156# RN VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X1 a_2268_156# a_36_124# a_1356_112# VSUBS nmos_6p0 w=0.39u l=0.6u
X2 a_2268_156# a_448_472# a_1356_112# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X3 a_1476_156# a_1356_112# a_1304_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X4 a_1024_476# a_36_124# a_820_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X5 a_1356_112# a_1024_476# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X6 VSS a_2682_301# a_2563_527# VSUBS nmos_6p0 w=0.39u l=0.6u
X7 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.405u l=0.6u
X8 a_1228_476# a_448_472# a_1024_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X9 a_1228_476# RN VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
X10 a_1356_112# a_1024_476# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X11 VDD a_2268_156# a_2682_301# w_n86_352# pmos_6p0 w=1.09u l=0.5u
X12 a_1024_476# a_448_472# a_820_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X13 VDD a_2682_301# a_2563_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X14 Q a_2682_301# VDD w_n86_352# pmos_6p0 w=1.185u l=0.5u
X15 a_1304_156# a_36_124# a_1024_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X16 Q a_2682_301# VSS VSUBS nmos_6p0 w=0.795u l=0.6u
X17 VDD a_1356_112# a_1228_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X18 a_2563_527# a_448_472# a_2268_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X19 a_2682_301# a_2268_156# a_3030_156# VSUBS nmos_6p0 w=0.825u l=0.6u
X20 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X21 VDD a_2682_301# Q w_n86_352# pmos_6p0 w=1.185u l=0.5u
X22 a_2682_301# RN VDD w_n86_352# pmos_6p0 w=1.09u l=0.5u
X23 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X24 VSS a_2682_301# Q VSUBS nmos_6p0 w=0.795u l=0.6u
X25 a_2563_527# a_36_124# a_2268_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X26 a_820_476# D VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X27 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X28 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X29 a_820_476# D VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 D Q RN VDD VSS CLKN
X0 a_3030_156# RN VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X1 a_2268_156# a_36_124# a_1356_112# VSUBS nmos_6p0 w=0.39u l=0.6u
X2 a_2268_156# a_448_472# a_1356_112# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X3 a_1476_156# a_1356_112# a_1304_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X4 a_1024_476# a_36_124# a_820_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X5 a_1356_112# a_1024_476# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X6 VSS a_2682_301# a_2563_527# VSUBS nmos_6p0 w=0.39u l=0.6u
X7 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.405u l=0.6u
X8 a_1228_476# a_448_472# a_1024_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X9 a_1228_476# RN VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
X10 a_1356_112# a_1024_476# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X11 VDD a_2268_156# a_2682_301# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 a_1024_476# a_448_472# a_820_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X13 Q a_2682_301# VSS VSUBS nmos_6p0 w=0.795u l=0.6u
X14 VDD a_2682_301# a_2563_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X15 Q a_2682_301# VDD w_n86_352# pmos_6p0 w=1.205u l=0.5u
X16 VDD a_2682_301# Q w_n86_352# pmos_6p0 w=1.205u l=0.5u
X17 a_1304_156# a_36_124# a_1024_476# VSUBS nmos_6p0 w=0.39u l=0.6u
X18 Q a_2682_301# VSS VSUBS nmos_6p0 w=0.795u l=0.6u
X19 VDD a_1356_112# a_1228_476# w_n86_352# pmos_6p0 w=0.76u l=0.5u
X20 VDD a_2682_301# Q w_n86_352# pmos_6p0 w=1.205u l=0.5u
X21 a_2563_527# a_448_472# a_2268_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X22 a_2682_301# a_2268_156# a_3030_156# VSUBS nmos_6p0 w=0.825u l=0.6u
X23 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X24 a_2682_301# RN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X25 Q a_2682_301# VDD w_n86_352# pmos_6p0 w=1.205u l=0.5u
X26 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X27 VSS a_2682_301# Q VSUBS nmos_6p0 w=0.795u l=0.6u
X28 a_2563_527# a_36_124# a_2268_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X29 a_820_476# D VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X30 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X31 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.39u l=0.6u
X32 VSS a_2682_301# Q VSUBS nmos_6p0 w=0.795u l=0.6u
X33 a_820_476# D VDD w_n86_352# pmos_6p0 w=0.76u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 D VDD VSS CLKN SETN RN Q
X0 VDD CLKN a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X1 a_2978_204# a_448_487# a_1356_112# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 a_1476_156# a_1356_112# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X3 a_3202_204# a_36_151# a_2978_204# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X4 a_448_487# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X5 a_1356_112# SETN VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X6 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X7 a_1248_504# RN VDD w_n86_352# pmos_6p0 w=0.805u l=0.5u
X8 Q a_3811_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X9 VSS a_3811_112# a_3763_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 a_1308_156# a_36_151# a_1044_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X11 a_2978_204# a_36_151# a_1356_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VSS CLKN a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X13 a_3811_112# a_2978_204# a_4155_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_3763_156# SETN a_3202_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 VDD a_1044_504# a_1356_112# w_n86_352# pmos_6p0 w=0.805u l=0.5u
X16 a_2544_204# a_1044_504# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1044_504# a_448_487# a_840_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X18 a_3202_204# a_448_487# a_2978_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_4155_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X20 a_840_504# D VDD w_n86_352# pmos_6p0 w=0.41u l=0.5u
X21 a_1356_112# SETN a_2544_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_1044_504# a_36_151# a_840_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X23 VDD a_1356_112# a_1248_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X24 a_3811_112# RN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X25 a_3202_204# SETN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X26 VDD a_2978_204# a_3811_112# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X27 VDD a_3811_112# a_3202_204# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X28 a_448_487# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X29 a_1248_504# a_448_487# a_1044_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X30 Q a_3811_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 a_840_504# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 D Q RN VDD VSS CLKN SETN
X0 VDD CLKN a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X1 a_2978_204# a_448_487# a_1356_112# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 VDD a_3811_112# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_1476_156# a_1356_112# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X4 a_3202_204# a_36_151# a_2978_204# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X5 a_448_487# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X6 a_1356_112# SETN VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X7 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X8 a_1248_504# RN VDD w_n86_352# pmos_6p0 w=0.805u l=0.5u
X9 Q a_3811_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X10 VSS a_3811_112# a_3763_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_1308_156# a_36_151# a_1044_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X12 a_2978_204# a_36_151# a_1356_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 VSS CLKN a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X14 a_3811_112# a_2978_204# a_4155_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_3763_156# SETN a_3202_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 VDD a_1044_504# a_1356_112# w_n86_352# pmos_6p0 w=0.805u l=0.5u
X17 a_2544_204# a_1044_504# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_1044_504# a_448_487# a_840_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 a_3202_204# a_448_487# a_2978_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X20 a_4155_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_840_504# D VDD w_n86_352# pmos_6p0 w=0.41u l=0.5u
X22 a_1356_112# SETN a_2544_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_1044_504# a_36_151# a_840_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X24 VDD a_1356_112# a_1248_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X25 a_3811_112# RN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X26 a_3202_204# SETN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X27 VDD a_2978_204# a_3811_112# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X28 VDD a_3811_112# a_3202_204# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X29 a_448_487# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X30 VSS a_3811_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X31 a_1248_504# a_448_487# a_1044_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X32 Q a_3811_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X33 a_840_504# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 D Q RN SETN VDD VSS CLKN
X0 VDD CLKN a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X1 a_2978_204# a_448_487# a_1356_112# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 VDD a_3811_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 a_1476_156# a_1356_112# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X4 VSS a_3811_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X5 a_3202_204# a_36_151# a_2978_204# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X6 a_448_487# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X7 a_1356_112# SETN VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X8 VSS RN a_1476_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X9 a_1248_504# RN VDD w_n86_352# pmos_6p0 w=0.805u l=0.5u
X10 Q a_3811_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X11 Q a_3811_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 VSS a_3811_112# a_3763_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 a_1308_156# a_36_151# a_1044_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X14 a_2978_204# a_36_151# a_1356_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 VDD a_3811_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X16 VSS CLKN a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X17 a_3811_112# a_2978_204# a_4155_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_3763_156# SETN a_3202_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 VDD a_1044_504# a_1356_112# w_n86_352# pmos_6p0 w=0.805u l=0.5u
X20 a_2544_204# a_1044_504# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_1044_504# a_448_487# a_840_504# VSUBS nmos_6p0 w=0.38u l=0.6u
X22 a_3202_204# a_448_487# a_2978_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_4155_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X24 a_840_504# D VDD w_n86_352# pmos_6p0 w=0.41u l=0.5u
X25 a_1356_112# SETN a_2544_204# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_1044_504# a_36_151# a_840_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X27 VDD a_1356_112# a_1248_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X28 a_3811_112# RN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X29 a_3202_204# SETN VDD w_n86_352# pmos_6p0 w=0.875u l=0.5u
X30 VDD a_2978_204# a_3811_112# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X31 Q a_3811_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X32 VDD a_3811_112# a_3202_204# w_n86_352# pmos_6p0 w=0.875u l=0.5u
X33 a_448_487# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X34 VSS a_3811_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X35 a_1248_504# a_448_487# a_1044_504# w_n86_352# pmos_6p0 w=0.41u l=0.5u
X36 Q a_3811_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X37 a_840_504# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 CLKN Q SETN VDD VSS D
X0 VSS a_1296_336# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X1 a_1708_156# a_1044_472# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X2 Q a_3148_126# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_840_156# D VDD w_n86_352# pmos_6p0 w=0.605u l=0.5u
X4 VDD SETN a_1296_336# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 Q a_3148_126# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 VSS a_3148_126# a_3008_145# VSUBS nmos_6p0 w=0.31u l=0.6u
X7 a_1296_336# a_1044_472# VDD w_n86_352# pmos_6p0 w=0.57u l=0.5u
X8 a_1044_472# a_36_124# a_840_156# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X9 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.54u l=0.6u
X10 a_1308_156# a_36_124# a_1044_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X11 a_2384_156# a_36_124# a_2160_156# w_n86_352# pmos_6p0 w=0.65u l=0.5u
X12 a_2384_156# SETN VDD w_n86_352# pmos_6p0 w=0.705u l=0.5u
X13 a_1248_472# a_448_472# a_1044_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X14 VDD a_3148_126# a_2384_156# w_n86_352# pmos_6p0 w=0.58u l=0.5u
X15 VDD a_1296_336# a_1248_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X16 a_840_156# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X17 a_2384_156# a_448_472# a_2160_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X18 a_1044_472# a_448_472# a_840_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.94u l=0.5u
X20 a_1296_336# SETN a_1708_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X21 a_2160_156# a_448_472# a_1296_336# w_n86_352# pmos_6p0 w=0.535u l=0.5u
X22 a_3148_126# a_2160_156# VSS VSUBS nmos_6p0 w=0.375u l=0.6u
X23 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.94u l=0.5u
X24 a_3148_126# a_2160_156# VDD w_n86_352# pmos_6p0 w=0.655u l=0.5u
X25 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X26 a_3008_145# SETN a_2384_156# VSUBS nmos_6p0 w=0.435u l=0.6u
X27 a_2160_156# a_36_124# a_1296_336# VSUBS nmos_6p0 w=0.38u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 D Q SETN VDD VSS CLKN
X0 VDD a_3148_126# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X1 VSS a_1296_336# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_1708_156# a_1044_472# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X3 Q a_3148_126# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X4 a_840_156# D VDD w_n86_352# pmos_6p0 w=0.605u l=0.5u
X5 VDD SETN a_1296_336# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X6 Q a_3148_126# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 VSS a_3148_126# a_3008_145# VSUBS nmos_6p0 w=0.31u l=0.6u
X8 a_1296_336# a_1044_472# VDD w_n86_352# pmos_6p0 w=0.57u l=0.5u
X9 a_1044_472# a_36_124# a_840_156# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X10 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.54u l=0.6u
X11 a_1308_156# a_36_124# a_1044_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X12 a_2384_156# a_36_124# a_2160_156# w_n86_352# pmos_6p0 w=0.65u l=0.5u
X13 a_2384_156# SETN VDD w_n86_352# pmos_6p0 w=0.705u l=0.5u
X14 a_1248_472# a_448_472# a_1044_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X15 VDD a_3148_126# a_2384_156# w_n86_352# pmos_6p0 w=0.58u l=0.5u
X16 VDD a_1296_336# a_1248_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X17 a_840_156# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X18 a_2384_156# a_448_472# a_2160_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 a_1044_472# a_448_472# a_840_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X20 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.94u l=0.5u
X21 a_1296_336# SETN a_1708_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X22 a_2160_156# a_448_472# a_1296_336# w_n86_352# pmos_6p0 w=0.535u l=0.5u
X23 a_3148_126# a_2160_156# VSS VSUBS nmos_6p0 w=0.375u l=0.6u
X24 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.94u l=0.5u
X25 a_3148_126# a_2160_156# VDD w_n86_352# pmos_6p0 w=0.655u l=0.5u
X26 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X27 a_3008_145# SETN a_2384_156# VSUBS nmos_6p0 w=0.435u l=0.6u
X28 a_2160_156# a_36_124# a_1296_336# VSUBS nmos_6p0 w=0.38u l=0.6u
X29 VSS a_3148_126# Q VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 D Q SETN VDD VSS CLKN
X0 VDD a_3148_126# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X1 VSS a_1296_336# a_1308_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_1708_156# a_1044_472# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X3 Q a_3148_126# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X4 a_840_156# D VDD w_n86_352# pmos_6p0 w=0.605u l=0.5u
X5 VDD SETN a_1296_336# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X6 Q a_3148_126# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 Q a_3148_126# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X8 VSS a_3148_126# a_3008_145# VSUBS nmos_6p0 w=0.31u l=0.6u
X9 a_1296_336# a_1044_472# VDD w_n86_352# pmos_6p0 w=0.57u l=0.5u
X10 VDD a_3148_126# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X11 a_1044_472# a_36_124# a_840_156# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X12 VSS CLKN a_36_124# VSUBS nmos_6p0 w=0.54u l=0.6u
X13 Q a_3148_126# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X14 a_1308_156# a_36_124# a_1044_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X15 a_2384_156# a_36_124# a_2160_156# w_n86_352# pmos_6p0 w=0.65u l=0.5u
X16 a_2384_156# SETN VDD w_n86_352# pmos_6p0 w=0.705u l=0.5u
X17 a_1248_472# a_448_472# a_1044_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X18 VDD a_3148_126# a_2384_156# w_n86_352# pmos_6p0 w=0.58u l=0.5u
X19 VDD a_1296_336# a_1248_472# w_n86_352# pmos_6p0 w=0.605u l=0.5u
X20 a_840_156# D VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X21 a_2384_156# a_448_472# a_2160_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X22 a_1044_472# a_448_472# a_840_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X23 VDD CLKN a_36_124# w_n86_352# pmos_6p0 w=0.94u l=0.5u
X24 a_1296_336# SETN a_1708_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X25 a_2160_156# a_448_472# a_1296_336# w_n86_352# pmos_6p0 w=0.535u l=0.5u
X26 a_3148_126# a_2160_156# VSS VSUBS nmos_6p0 w=0.375u l=0.6u
X27 a_448_472# a_36_124# VDD w_n86_352# pmos_6p0 w=0.94u l=0.5u
X28 a_3148_126# a_2160_156# VDD w_n86_352# pmos_6p0 w=0.655u l=0.5u
X29 a_448_472# a_36_124# VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X30 a_3008_145# SETN a_2384_156# VSUBS nmos_6p0 w=0.435u l=0.6u
X31 a_2160_156# a_36_124# a_1296_336# VSUBS nmos_6p0 w=0.38u l=0.6u
X32 VSS a_3148_126# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X33 VSS a_3148_126# Q VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D
X0 a_880_527# a_448_472# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X1 a_1348_527# a_36_151# a_1004_159# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 a_1328_159# a_448_472# a_1004_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 VDD a_1376_115# a_1348_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_2304_115# a_2296_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 a_2304_115# a_2011_527# VDD w_n86_352# pmos_6p0 w=0.8u l=0.5u
X6 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X7 Q a_2304_115# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_2304_115# a_2011_527# VSS VSUBS nmos_6p0 w=0.4u l=0.6u
X9 a_1004_159# D a_836_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 a_1004_159# D a_880_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 a_2011_527# a_36_151# a_1376_115# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X12 a_2296_527# a_448_472# a_2011_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X13 a_1376_115# a_1004_159# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X15 VSS a_1376_115# a_1328_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2011_527# a_448_472# a_1376_115# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X18 Q a_2304_115# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_1376_115# a_1004_159# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X20 VSS a_2304_115# a_2256_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_836_159# a_36_151# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X23 a_2256_159# a_36_151# a_2011_527# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D VDD VSS CLK Q
X0 a_880_527# a_448_472# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X1 a_1348_527# a_36_151# a_1004_159# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 a_1328_159# a_448_472# a_1004_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 VDD a_1376_115# a_1348_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_2304_115# a_2296_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 a_2304_115# a_2011_527# VDD w_n86_352# pmos_6p0 w=0.8u l=0.5u
X6 VSS a_2304_115# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X8 Q a_2304_115# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_2304_115# a_2011_527# VSS VSUBS nmos_6p0 w=0.4u l=0.6u
X10 a_1004_159# D a_836_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_1004_159# D a_880_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X12 a_2011_527# a_36_151# a_1376_115# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X13 a_2296_527# a_448_472# a_2011_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 a_1376_115# a_1004_159# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X16 VDD a_2304_115# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VSS a_1376_115# a_1328_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_2011_527# a_448_472# a_1376_115# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X20 Q a_2304_115# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_1376_115# a_1004_159# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 VSS a_2304_115# a_2256_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_836_159# a_36_151# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X24 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X25 a_2256_159# a_36_151# a_2011_527# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D Q VDD VSS CLK
X0 a_880_527# a_448_472# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X1 a_1348_527# a_36_151# a_1004_159# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VDD a_2304_115# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_1328_159# a_448_472# a_1004_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD a_1376_115# a_1348_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_2011_527# a_2304_115# VSUBS nmos_6p0 w=0.815u l=0.6u
X6 VDD a_2304_115# a_2296_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 a_2304_115# a_2011_527# VDD w_n86_352# pmos_6p0 w=0.945u l=0.5u
X8 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X9 VDD a_2011_527# a_2304_115# w_n86_352# pmos_6p0 w=0.945u l=0.5u
X10 a_1004_159# D a_836_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VSS a_2304_115# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_2304_115# a_2011_527# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X13 a_1004_159# D a_880_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 a_2011_527# a_36_151# a_1376_115# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_2296_527# a_448_472# a_2011_527# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 Q a_2304_115# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VSS a_2304_115# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X18 a_1376_115# a_1004_159# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X19 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X20 VDD a_2304_115# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 VSS a_1376_115# a_1328_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_2011_527# a_448_472# a_1376_115# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 Q a_2304_115# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X25 Q a_2304_115# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X26 a_1376_115# a_1004_159# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X27 VSS a_2304_115# a_2256_159# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 Q a_2304_115# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X29 a_836_159# a_36_151# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X30 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X31 a_2256_159# a_36_151# a_2011_527# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D Q RN VSS CLK VDD
X0 a_1308_423# a_1000_472# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X1 a_1000_472# a_36_151# a_796_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_796_472# D VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X3 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X4 VSS RN a_1456_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 Q a_2665_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 a_796_472# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X7 VSS a_2665_112# a_2560_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_2665_112# a_2248_156# a_3041_156# VSUBS nmos_6p0 w=0.4u l=0.6u
X9 a_1000_472# a_448_472# a_796_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X10 a_2248_156# a_36_151# a_1308_423# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X11 a_2248_156# a_448_472# a_1308_423# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X13 a_1456_156# a_1308_423# a_1288_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1308_423# a_1000_472# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X15 Q a_2665_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X16 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X17 a_1204_472# a_36_151# a_1000_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X18 a_1204_472# RN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X19 a_2665_112# RN VDD w_n86_352# pmos_6p0 w=1u l=0.5u
X20 a_2560_156# a_36_151# a_2248_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 VDD a_2248_156# a_2665_112# w_n86_352# pmos_6p0 w=1u l=0.5u
X22 a_1288_156# a_448_472# a_1000_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 VDD a_1308_423# a_1204_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X24 a_2560_156# a_448_472# a_2248_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X25 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X26 a_3041_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X27 VDD a_2665_112# a_2560_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D Q RN VDD VSS CLK
X0 a_1308_423# a_1000_472# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X1 a_1000_472# a_36_151# a_796_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_796_472# D VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X3 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X4 Q a_2665_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 VSS RN a_1456_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VDD a_2665_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 a_796_472# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X8 VSS a_2665_112# a_2560_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_1000_472# a_448_472# a_796_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X10 a_2248_156# a_36_151# a_1308_423# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X11 a_2248_156# a_448_472# a_1308_423# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X13 a_1456_156# a_1308_423# a_1288_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1308_423# a_1000_472# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X15 Q a_2665_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X16 a_2665_112# a_2248_156# a_3041_156# VSUBS nmos_6p0 w=0.815u l=0.6u
X17 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X18 a_1204_472# a_36_151# a_1000_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X19 a_1204_472# RN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X20 a_2560_156# a_36_151# a_2248_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_1288_156# a_448_472# a_1000_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_2665_112# RN VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X23 VDD a_1308_423# a_1204_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X24 a_2560_156# a_448_472# a_2248_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X25 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X26 VDD a_2248_156# a_2665_112# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X27 a_3041_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X28 VSS a_2665_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X29 VDD a_2665_112# a_2560_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D Q RN VDD VSS CLK
X0 VSS a_2665_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X1 a_1308_423# a_1000_472# VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X2 a_1000_472# a_36_151# a_796_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_796_472# D VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X4 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X5 Q a_2665_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 VDD a_2665_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 VSS RN a_1456_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 VDD a_2665_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 a_796_472# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X10 VSS a_2665_112# a_2560_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_1000_472# a_448_472# a_796_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X12 a_2248_156# a_36_151# a_1308_423# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X13 a_2248_156# a_448_472# a_1308_423# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X15 Q a_2665_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X16 a_1456_156# a_1308_423# a_1288_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1308_423# a_1000_472# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 Q a_2665_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X19 Q a_2665_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X20 a_2665_112# a_2248_156# a_3041_156# VSUBS nmos_6p0 w=0.815u l=0.6u
X21 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X22 a_1204_472# a_36_151# a_1000_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X23 a_1204_472# RN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X24 a_2560_156# a_36_151# a_2248_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_1288_156# a_448_472# a_1000_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_2665_112# RN VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X27 VDD a_1308_423# a_1204_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X28 a_2560_156# a_448_472# a_2248_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X29 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X30 VDD a_2248_156# a_2665_112# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X31 a_3041_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X32 VSS a_2665_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X33 VDD a_2665_112# a_2560_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 RN D Q CLK VSS VDD SETN
X0 a_1036_517# a_428_472# a_832_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X1 a_832_517# D VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X2 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X3 a_2664_156# a_36_151# a_2440_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X4 a_2664_156# SETN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X5 a_428_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X6 a_1240_517# a_36_151# a_1036_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X7 VDD a_3296_112# a_2664_156# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X8 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X9 a_2036_156# a_1036_517# VSS VSUBS nmos_6p0 w=0.505u l=0.6u
X10 Q a_3296_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X11 VDD a_1344_416# a_1240_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X12 a_3296_112# RN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X13 a_1524_171# a_1344_416# a_1356_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X14 a_1240_517# RN VDD w_n86_352# pmos_6p0 w=0.755u l=0.5u
X15 VDD a_2440_156# a_3296_112# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X16 a_3232_156# SETN a_2664_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X17 a_2440_156# a_428_472# a_1344_416# VSUBS nmos_6p0 w=0.505u l=0.6u
X18 a_1356_171# a_428_472# a_1036_517# VSUBS nmos_6p0 w=0.365u l=0.6u
X19 a_1344_416# SETN a_2036_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X20 a_1344_416# SETN VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X21 Q a_3296_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X22 a_2440_156# a_36_151# a_1344_416# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X23 a_3640_156# RN VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X24 a_2664_156# a_428_472# a_2440_156# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X25 VDD a_1036_517# a_1344_416# w_n86_352# pmos_6p0 w=0.755u l=0.5u
X26 VSS a_3296_112# a_3232_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X27 a_428_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X28 a_832_517# D VDD w_n86_352# pmos_6p0 w=0.365u l=0.5u
X29 VSS RN a_1524_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X30 a_3296_112# a_2440_156# a_3640_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X31 a_1036_517# a_36_151# a_832_517# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 RN D Q CLK VSS VDD SETN
X0 VSS a_3296_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X1 a_1036_517# a_428_472# a_832_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X2 a_832_517# D VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X3 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X4 a_2664_156# a_36_151# a_2440_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X5 a_2664_156# SETN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X6 a_428_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X7 a_1240_517# a_36_151# a_1036_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X8 VDD a_3296_112# a_2664_156# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X9 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X10 a_2036_156# a_1036_517# VSS VSUBS nmos_6p0 w=0.505u l=0.6u
X11 Q a_3296_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 VDD a_1344_416# a_1240_517# w_n86_352# pmos_6p0 w=0.365u l=0.5u
X13 a_3296_112# RN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X14 a_1524_171# a_1344_416# a_1356_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X15 a_1240_517# RN VDD w_n86_352# pmos_6p0 w=0.755u l=0.5u
X16 VDD a_2440_156# a_3296_112# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X17 a_3232_156# SETN a_2664_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X18 a_2440_156# a_428_472# a_1344_416# VSUBS nmos_6p0 w=0.505u l=0.6u
X19 a_1356_171# a_428_472# a_1036_517# VSUBS nmos_6p0 w=0.365u l=0.6u
X20 a_1344_416# SETN a_2036_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X21 a_1344_416# SETN VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X22 Q a_3296_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X23 a_2440_156# a_36_151# a_1344_416# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X24 a_3640_156# RN VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X25 VDD a_3296_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X26 a_2664_156# a_428_472# a_2440_156# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X27 VDD a_1036_517# a_1344_416# w_n86_352# pmos_6p0 w=0.755u l=0.5u
X28 VSS a_3296_112# a_3232_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X29 a_428_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X30 a_832_517# D VDD w_n86_352# pmos_6p0 w=0.365u l=0.5u
X31 VSS RN a_1524_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X32 a_3296_112# a_2440_156# a_3640_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X33 a_1036_517# a_36_151# a_832_517# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 D Q RN SETN VDD VSS CLK
X0 VSS a_3296_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X1 a_832_504# D VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X2 Q a_3296_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X3 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X4 a_2664_156# a_36_151# a_2440_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X5 a_2664_156# SETN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X6 VDD a_3296_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 a_428_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X8 a_832_504# D VDD w_n86_352# pmos_6p0 w=0.475u l=0.5u
X9 VDD a_1036_504# a_1344_416# w_n86_352# pmos_6p0 w=0.69u l=0.5u
X10 VDD a_3296_112# a_2664_156# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X11 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X12 a_2036_156# a_1036_504# VSS VSUBS nmos_6p0 w=0.505u l=0.6u
X13 Q a_3296_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X14 a_1036_504# a_428_472# a_832_504# w_n86_352# pmos_6p0 w=0.475u l=0.5u
X15 a_3296_112# RN VDD w_n86_352# pmos_6p0 w=0.77u l=0.5u
X16 a_1524_171# a_1344_416# a_1356_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X17 VDD a_2440_156# a_3296_112# w_n86_352# pmos_6p0 w=0.77u l=0.5u
X18 a_1240_504# a_36_151# a_1036_504# w_n86_352# pmos_6p0 w=0.475u l=0.5u
X19 a_3232_156# SETN a_2664_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X20 a_2440_156# a_428_472# a_1344_416# VSUBS nmos_6p0 w=0.505u l=0.6u
X21 a_1356_171# a_428_472# a_1036_504# VSUBS nmos_6p0 w=0.365u l=0.6u
X22 a_1344_416# SETN a_2036_156# VSUBS nmos_6p0 w=0.505u l=0.6u
X23 VDD a_1344_416# a_1240_504# w_n86_352# pmos_6p0 w=0.475u l=0.5u
X24 a_1344_416# SETN VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X25 Q a_3296_112# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X26 a_2440_156# a_36_151# a_1344_416# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X27 a_3640_156# RN VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X28 Q a_3296_112# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X29 a_1240_504# RN VDD w_n86_352# pmos_6p0 w=0.69u l=0.5u
X30 VDD a_3296_112# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X31 a_2664_156# a_428_472# a_2440_156# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X32 VSS a_3296_112# a_3232_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X33 a_428_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X34 VSS RN a_1524_171# VSUBS nmos_6p0 w=0.365u l=0.6u
X35 a_3296_112# a_2440_156# a_3640_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X36 VSS a_3296_112# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X37 a_1036_504# a_36_151# a_832_504# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 VSS CLK VDD D Q SETN
X0 a_1353_112# a_1040_527# VDD w_n86_352# pmos_6p0 w=0.585u l=0.5u
X1 a_3129_107# a_2225_156# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X2 VDD SETN a_1353_112# w_n86_352# pmos_6p0 w=0.585u l=0.5u
X3 a_1284_156# a_448_472# a_1040_527# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD a_1353_112# a_1293_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X5 Q a_3129_107# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 a_3129_107# a_2225_156# VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X7 a_1697_156# a_1040_527# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_2449_156# a_36_151# a_2225_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_1293_527# a_36_151# a_1040_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X10 a_3081_151# SETN a_2449_156# VSUBS nmos_6p0 w=0.405u l=0.6u
X11 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X12 a_1353_112# SETN a_1697_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 a_836_156# D VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X14 a_1040_527# a_36_151# a_836_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_1040_527# a_448_472# a_836_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X16 a_2225_156# a_36_151# a_1353_112# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X17 VSS a_1353_112# a_1284_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_2225_156# a_448_472# a_1353_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X20 a_2449_156# a_448_472# a_2225_156# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X21 VDD a_3129_107# a_2449_156# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X22 Q a_3129_107# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X23 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X24 a_2449_156# SETN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X25 VSS a_3129_107# a_3081_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X26 a_836_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X27 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D Q SETN VSS CLK VDD
X0 a_1353_112# a_1040_527# VDD w_n86_352# pmos_6p0 w=0.585u l=0.5u
X1 Q a_3129_107# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X2 VDD SETN a_1353_112# w_n86_352# pmos_6p0 w=0.585u l=0.5u
X3 a_1284_156# a_448_472# a_1040_527# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD a_1353_112# a_1293_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X5 a_1697_156# a_1040_527# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_2449_156# a_36_151# a_2225_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_1293_527# a_36_151# a_1040_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X8 a_3129_107# a_2225_156# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X9 a_3081_151# SETN a_2449_156# VSUBS nmos_6p0 w=0.405u l=0.6u
X10 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X11 a_1353_112# SETN a_1697_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_836_156# D VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X13 a_1040_527# a_36_151# a_836_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1040_527# a_448_472# a_836_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X15 a_2225_156# a_36_151# a_1353_112# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X16 VSS a_1353_112# a_1284_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2225_156# a_448_472# a_1353_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 Q a_3129_107# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X19 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X20 a_2449_156# a_448_472# a_2225_156# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X21 VDD a_3129_107# a_2449_156# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X22 a_3129_107# a_2225_156# VDD w_n86_352# pmos_6p0 w=1.055u l=0.5u
X23 VDD a_3129_107# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X24 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X25 a_2449_156# SETN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X26 VSS a_3129_107# a_3081_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X27 a_836_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X28 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
X29 VSS a_3129_107# Q VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D Q SETN VDD VSS CLK
X0 a_1353_112# a_1040_527# VDD w_n86_352# pmos_6p0 w=0.585u l=0.5u
X1 VDD SETN a_1353_112# w_n86_352# pmos_6p0 w=0.585u l=0.5u
X2 a_1284_156# a_448_472# a_1040_527# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 Q a_3129_107# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 VDD a_1353_112# a_1293_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X5 a_3129_107# a_2225_156# VDD w_n86_352# pmos_6p0 w=1.055u l=0.5u
X6 a_1697_156# a_1040_527# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_2449_156# a_36_151# a_2225_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_1293_527# a_36_151# a_1040_527# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X9 a_3129_107# a_2225_156# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X10 Q a_3129_107# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X11 VDD a_3129_107# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X12 a_3081_151# SETN a_2449_156# VSUBS nmos_6p0 w=0.405u l=0.6u
X13 VDD a_2225_156# a_3129_107# w_n86_352# pmos_6p0 w=1.055u l=0.5u
X14 VSS CLK a_36_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X15 Q a_3129_107# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X16 a_1353_112# SETN a_1697_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_836_156# D VDD w_n86_352# pmos_6p0 w=0.505u l=0.5u
X18 VDD a_3129_107# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X19 VSS a_2225_156# a_3129_107# VSUBS nmos_6p0 w=0.815u l=0.6u
X20 a_1040_527# a_36_151# a_836_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 VSS a_3129_107# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X22 a_1040_527# a_448_472# a_836_156# w_n86_352# pmos_6p0 w=0.505u l=0.5u
X23 a_2225_156# a_36_151# a_1353_112# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X24 VSS a_3129_107# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X25 VSS a_1353_112# a_1284_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_2225_156# a_448_472# a_1353_112# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 Q a_3129_107# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X28 VDD CLK a_36_151# w_n86_352# pmos_6p0 w=0.865u l=0.5u
X29 a_2449_156# a_448_472# a_2225_156# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X30 VDD a_3129_107# a_2449_156# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X31 a_448_472# a_36_151# VDD w_n86_352# pmos_6p0 w=0.865u l=0.5u
X32 a_2449_156# SETN VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X33 VSS a_3129_107# a_3081_151# VSUBS nmos_6p0 w=0.405u l=0.6u
X34 a_836_156# D VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X35 a_448_472# a_36_151# VSS VSUBS nmos_6p0 w=0.405u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dffsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 VSS Z I VDD
X0 Z a_608_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_448_495# a_36_126# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VSS a_448_495# a_608_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 Z a_608_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_448_495# a_36_126# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VDD I a_36_126# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X6 VSS I a_36_126# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 VDD a_448_495# a_608_472# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 VDD I Z VSS
X0 VSS a_608_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_448_495# a_36_126# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VSS a_448_495# a_608_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 Z a_608_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_448_495# a_36_126# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VDD I a_36_126# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X6 VDD a_608_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 Z a_608_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VSS I a_36_126# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 VDD a_448_495# a_608_472# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_4 VSS Z I VDD
X0 VDD a_629_110# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 Z a_629_110# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS a_449_526# a_629_110# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 Z a_629_110# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS a_629_110# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS I a_37_110# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VDD a_449_526# a_629_110# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 a_449_526# a_37_110# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 VDD a_629_110# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VSS a_629_110# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD I a_37_110# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 Z a_629_110# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_449_526# a_37_110# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X13 Z a_629_110# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlya_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 VDD I VSS Z
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X1 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 Z a_895_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X5 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 VDD a_671_644# a_1127_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 Z a_895_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_1147_68# a_671_644# a_895_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X11 a_1127_622# a_671_644# a_895_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_2 VDD I Z VSS
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X1 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X4 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VSS a_895_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X6 Z a_895_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 VDD a_671_644# a_1127_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 VDD a_895_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 Z a_895_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_1147_68# a_671_644# a_895_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X13 a_1127_622# a_671_644# a_895_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_4 VSS Z I VDD
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X1 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X2 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X4 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VSS a_895_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X6 Z a_895_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 VDD a_671_644# a_1127_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 VDD a_895_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 Z a_895_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS a_895_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X12 Z a_895_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 VDD a_895_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 Z a_895_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_1147_68# a_671_644# a_895_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X17 a_1127_622# a_671_644# a_895_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyb_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 Z VSS I VDD
X0 a_518_68# a_42_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X1 a_666_644# a_42_68# a_518_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1142_68# a_666_644# a_870_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_2158_622# a_1702_68# a_1926_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 a_2178_68# a_1702_68# a_1926_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X5 VSS a_666_644# a_1142_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VSS a_1702_68# a_2178_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X7 VDD a_666_644# a_1102_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 a_666_644# a_42_68# a_498_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 VSS I a_42_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 a_1702_68# a_870_562# a_1554_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 Z a_1926_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_498_644# a_42_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X13 a_1554_644# a_870_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 a_1102_644# a_666_644# a_870_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 VDD I a_42_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 a_1534_68# a_870_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1702_68# a_870_562# a_1534_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 Z a_1926_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 VDD a_1702_68# a_2158_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_2 VDD I VSS Z
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 Z a_1931_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_1931_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_671_644# a_1107_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_1707_68# a_875_562# a_1559_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 Z a_1931_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_1559_644# a_875_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X10 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VSS a_1931_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_2183_68# a_1707_68# a_1931_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X13 VSS a_1707_68# a_2183_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X14 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_1107_644# a_671_644# a_875_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 a_1539_68# a_875_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X17 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X18 a_1707_68# a_875_562# a_1539_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 VDD a_1707_68# a_2163_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X20 a_1147_68# a_671_644# a_875_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_2163_622# a_1707_68# a_1931_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_4 Z VSS I VDD
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 Z a_1931_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_1931_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_671_644# a_1107_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 Z a_1931_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 Z a_1931_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_1707_68# a_875_562# a_1559_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 Z a_1931_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_1559_644# a_875_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X12 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 VSS a_1931_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_2183_68# a_1707_68# a_1931_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X15 VSS a_1707_68# a_2183_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X16 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X17 a_1107_644# a_671_644# a_875_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X18 VSS a_1931_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_1539_68# a_875_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X20 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X21 a_1707_68# a_875_562# a_1539_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 VDD a_1931_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VDD a_1707_68# a_2163_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X24 a_1147_68# a_671_644# a_875_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_2163_622# a_1707_68# a_1931_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyc_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 VDD I VSS Z
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 Z a_2987_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_2163_644# a_1707_68# a_1931_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X3 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_671_644# a_1107_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_2615_644# a_1931_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 a_1707_68# a_875_562# a_1559_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 VDD a_2763_68# a_3219_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X10 a_1559_644# a_875_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 Z a_2987_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X14 a_1107_644# a_671_644# a_875_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_2595_68# a_1931_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2763_68# a_1931_562# a_2595_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1539_68# a_875_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X19 a_1707_68# a_875_562# a_1539_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X20 a_2763_68# a_1931_562# a_2615_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X21 a_3219_622# a_2763_68# a_2987_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X22 a_3239_68# a_2763_68# a_2987_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X23 a_2203_68# a_1707_68# a_1931_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X24 VSS a_1707_68# a_2203_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 VDD a_1707_68# a_2163_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X26 VSS a_2763_68# a_3239_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X27 a_1147_68# a_671_644# a_875_562# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_2 VDD I VSS Z
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 Z a_2987_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_2163_644# a_1707_68# a_1931_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X3 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_671_644# a_1107_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 VDD a_2987_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_2615_644# a_1931_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 a_1707_68# a_875_562# a_1559_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X10 VDD a_2763_68# a_3219_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X11 a_1559_644# a_875_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X12 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 Z a_2987_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_1107_644# a_671_644# a_875_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 a_2595_68# a_1931_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2763_68# a_1931_562# a_2595_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 VSS a_2987_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_1539_68# a_875_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X20 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X21 a_1707_68# a_875_562# a_1539_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_2763_68# a_1931_562# a_2615_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X23 a_3219_622# a_2763_68# a_2987_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X24 a_3239_68# a_2763_68# a_2987_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X25 a_2203_68# a_1707_68# a_1931_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 VSS a_1707_68# a_2203_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 VDD a_1707_68# a_2163_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X28 VSS a_2763_68# a_3239_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X29 a_1147_68# a_671_644# a_875_562# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 Z VDD I VSS
X0 VSS a_671_644# a_1147_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 Z a_2987_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_2163_644# a_1707_68# a_1931_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X3 a_671_644# a_47_68# a_503_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_671_644# a_1107_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X5 VDD a_2987_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS I a_47_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_2615_644# a_1931_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X8 a_1707_68# a_875_562# a_1559_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 Z a_2987_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VSS a_2987_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_523_68# a_47_68# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VDD a_2763_68# a_3219_622# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X13 VDD a_2987_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 Z a_2987_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1559_644# a_875_562# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 a_671_644# a_47_68# a_523_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 Z a_2987_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_503_644# a_47_68# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X19 a_1107_644# a_671_644# a_875_562# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X20 a_2595_68# a_1931_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_2763_68# a_1931_562# a_2595_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 VSS a_2987_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_1539_68# a_875_562# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X24 VDD I a_47_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X25 a_1707_68# a_875_562# a_1539_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_2763_68# a_1931_562# a_2615_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X27 a_3219_622# a_2763_68# a_2987_68# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X28 a_3239_68# a_2763_68# a_2987_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X29 a_2203_68# a_1707_68# a_1931_562# VSUBS nmos_6p0 w=0.36u l=0.6u
X30 VSS a_1707_68# a_2203_68# VSUBS nmos_6p0 w=0.36u l=0.6u
X31 VDD a_1707_68# a_2163_644# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X32 VSS a_2763_68# a_3239_68# VSUBS nmos_6p0 w=0.365u l=0.6u
X33 a_1147_68# a_671_644# a_875_562# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__dlyd_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__endcap.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VSS VDD
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__endcap.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_4 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_8 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_16 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_32.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_32 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_32.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_64.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fill_64 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fill_64.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
X0 VDD a_124_375# a_36_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X1 a_124_375# a_36_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
X0 VDD a_124_375# a_36_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X1 VDD a_572_375# a_484_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X3 a_124_375# a_36_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
X0 VDD a_1468_375# a_1380_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X1 VDD a_124_375# a_36_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X2 a_1020_375# a_932_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X3 VDD a_572_375# a_484_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X4 a_572_375# a_484_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X5 a_124_375# a_36_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X7 VDD a_1020_375# a_932_472# w_n86_352# pmos_6p0 w=1.22u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_32.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
X0 VDD a_1468_375# a_1380_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X1 VDD a_124_375# a_36_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X2 a_1020_375# a_932_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X3 VDD a_572_375# a_484_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X4 VDD a_2364_375# a_2276_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X5 a_572_375# a_484_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X6 VDD a_1916_375# a_1828_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X7 a_124_375# a_36_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X8 a_1916_375# a_1828_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X9 a_1468_375# a_1380_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X10 a_2812_375# a_2724_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X11 VDD a_3260_375# a_3172_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X12 a_2364_375# a_2276_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X13 VDD a_2812_375# a_2724_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X14 a_3260_375# a_3172_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X15 VDD a_1020_375# a_932_472# w_n86_352# pmos_6p0 w=1.22u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_32.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_64.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
X0 VDD a_1468_375# a_1380_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X1 VDD a_4156_375# a_4068_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X2 VDD a_5948_375# a_5860_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X3 VDD a_124_375# a_36_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X4 a_3708_375# a_3620_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X5 VDD a_3708_375# a_3620_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X6 a_1020_375# a_932_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X7 a_4604_375# a_4516_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X8 VDD a_572_375# a_484_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X9 VDD a_2364_375# a_2276_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X10 a_4156_375# a_4068_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X11 a_5500_375# a_5412_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X12 VDD a_6844_375# a_6756_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X13 a_572_375# a_484_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X14 VDD a_5052_375# a_4964_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X15 VDD a_1916_375# a_1828_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X16 a_124_375# a_36_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X17 a_5052_375# a_4964_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X18 a_1916_375# a_1828_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X19 VDD a_4604_375# a_4516_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X20 a_1468_375# a_1380_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X21 a_2812_375# a_2724_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X22 VDD a_3260_375# a_3172_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X23 a_2364_375# a_2276_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X24 a_5948_375# a_5860_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X25 VDD a_2812_375# a_2724_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X26 a_3260_375# a_3172_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X27 VDD a_1020_375# a_932_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X28 VDD a_5500_375# a_5412_472# w_n86_352# pmos_6p0 w=1.22u l=1u
X29 a_6844_375# a_6756_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X30 a_6396_375# a_6308_472# VSS VSUBS nmos_6p0 w=0.82u l=1u
X31 VDD a_6396_375# a_6308_472# w_n86_352# pmos_6p0 w=1.22u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__fillcap_64.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__filltie.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__filltie.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__hold.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__hold Z VDD VSS
X0 a_168_69# Z VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VDD a_168_69# Z w_n86_352# pmos_6p0 w=0.32u l=2u
X2 a_168_69# Z VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS a_168_69# Z VSUBS nmos_6p0 w=0.32u l=2u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__hold.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_1 Q TE VDD VSS CLKN E
X0 VDD a_688_515# a_1059_112# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X1 Q a_2739_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_688_515# a_572_109# a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X3 a_2739_93# a_2007_475# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X4 Q a_2739_93# VSS VSUBS nmos_6p0 w=0.625u l=0.6u
X5 VDD CLKN a_588_415# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X6 a_919_153# a_588_415# a_688_515# VSUBS nmos_6p0 w=0.395u l=0.6u
X7 a_2735_472# a_2007_475# VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X8 a_2739_93# CLKN a_2735_472# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X9 VSS CLKN a_2739_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X10 VSS a_1059_112# a_919_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X11 a_987_515# a_572_109# a_688_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X12 a_572_109# a_588_415# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X13 a_36_153# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X14 VSS CLKN a_588_415# VSUBS nmos_6p0 w=0.395u l=0.6u
X15 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X16 a_688_515# a_588_415# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X17 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X18 VDD a_1059_112# a_987_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X19 a_2007_475# a_1059_112# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X20 a_2007_475# a_1059_112# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X21 VSS a_688_515# a_1059_112# VSUBS nmos_6p0 w=0.395u l=0.6u
X22 a_572_109# a_588_415# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X23 VSS TE a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_2 Q TE VDD VSS CLKN E
X0 VDD a_688_515# a_1059_112# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X1 a_688_515# a_572_109# a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 a_2739_93# a_2007_475# VSS VSUBS nmos_6p0 w=0.475u l=0.6u
X3 Q a_2739_93# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X4 VDD CLKN a_588_415# w_n86_352# pmos_6p0 w=1.155u l=0.5u
X5 Q a_2739_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_919_153# a_588_415# a_688_515# VSUBS nmos_6p0 w=0.395u l=0.6u
X7 VDD a_2739_93# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_2735_472# a_2007_475# VDD w_n86_352# pmos_6p0 w=1.155u l=0.5u
X9 a_2739_93# CLKN a_2735_472# w_n86_352# pmos_6p0 w=1.155u l=0.5u
X10 VSS CLKN a_2739_93# VSUBS nmos_6p0 w=0.475u l=0.6u
X11 VSS a_1059_112# a_919_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X12 a_987_515# a_572_109# a_688_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X13 a_572_109# a_588_415# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X14 a_36_153# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X15 VSS CLKN a_588_415# VSUBS nmos_6p0 w=0.475u l=0.6u
X16 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 a_688_515# a_588_415# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X18 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X19 VDD a_1059_112# a_987_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X20 a_2007_475# a_1059_112# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X21 a_2007_475# a_1059_112# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X22 VSS a_688_515# a_1059_112# VSUBS nmos_6p0 w=0.395u l=0.6u
X23 a_572_109# a_588_415# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X24 VSS a_2739_93# Q VSUBS nmos_6p0 w=0.63u l=0.6u
X25 VSS TE a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtn_4 Q TE VDD VSS CLKN E
X0 VDD a_688_515# a_1059_112# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X1 a_688_515# a_572_109# a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 a_2739_93# a_2007_475# VSS VSUBS nmos_6p0 w=0.475u l=0.6u
X3 Q a_2739_93# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X4 VDD CLKN a_588_415# w_n86_352# pmos_6p0 w=1.155u l=0.5u
X5 Q a_2739_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_919_153# a_588_415# a_688_515# VSUBS nmos_6p0 w=0.395u l=0.6u
X7 VDD a_2739_93# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_2735_472# a_2007_475# VDD w_n86_352# pmos_6p0 w=1.155u l=0.5u
X9 a_2739_93# CLKN a_2735_472# w_n86_352# pmos_6p0 w=1.155u l=0.5u
X10 Q a_2739_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS CLKN a_2739_93# VSUBS nmos_6p0 w=0.475u l=0.6u
X12 VSS a_1059_112# a_919_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X13 a_987_515# a_572_109# a_688_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X14 a_572_109# a_588_415# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X15 VDD a_2739_93# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_36_153# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X17 VSS CLKN a_588_415# VSUBS nmos_6p0 w=0.475u l=0.6u
X18 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X19 Q a_2739_93# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X20 a_688_515# a_588_415# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X21 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X22 VDD a_1059_112# a_987_515# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X23 a_2007_475# a_1059_112# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X24 a_2007_475# a_1059_112# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X25 VSS a_688_515# a_1059_112# VSUBS nmos_6p0 w=0.395u l=0.6u
X26 VSS a_2739_93# Q VSUBS nmos_6p0 w=0.63u l=0.6u
X27 a_572_109# a_588_415# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X28 VSS a_2739_93# Q VSUBS nmos_6p0 w=0.63u l=0.6u
X29 VSS TE a_36_153# VSUBS nmos_6p0 w=0.395u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtn_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_1 Q TE VDD VSS CLK E
X0 Q a_2319_91# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X1 a_688_507# a_572_93# a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 a_2319_91# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X3 VDD a_1059_112# a_2319_91# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X4 a_919_137# a_588_407# a_688_507# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 a_572_93# CLK VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X6 VSS a_572_93# a_588_407# VSUBS nmos_6p0 w=0.39u l=0.6u
X7 VSS a_1059_112# a_919_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X8 VSS a_1059_112# a_2527_91# VSUBS nmos_6p0 w=0.39u l=0.6u
X9 VDD a_572_93# a_588_407# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X10 a_572_93# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X11 a_36_137# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X12 a_987_507# a_572_93# a_688_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X13 a_1059_112# a_688_507# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X14 Q a_2319_91# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X16 a_688_507# a_588_407# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X17 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X18 VDD a_1059_112# a_987_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X19 a_1059_112# a_688_507# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X20 VSS TE a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X21 a_2527_91# CLK a_2319_91# VSUBS nmos_6p0 w=0.39u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_2 Q TE VDD VSS CLK E
X0 a_688_507# a_572_93# a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 a_2319_91# CLK VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS a_2319_91# Q VSUBS nmos_6p0 w=0.625u l=0.6u
X3 Q a_2319_91# VSS VSUBS nmos_6p0 w=0.625u l=0.6u
X4 VDD a_1059_112# a_2319_91# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_919_137# a_588_407# a_688_507# VSUBS nmos_6p0 w=0.395u l=0.6u
X6 Q a_2319_91# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_572_93# CLK VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X8 VSS a_572_93# a_588_407# VSUBS nmos_6p0 w=0.39u l=0.6u
X9 VSS a_1059_112# a_919_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X10 VSS a_1059_112# a_2527_91# VSUBS nmos_6p0 w=0.625u l=0.6u
X11 VDD a_572_93# a_588_407# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X12 a_572_93# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X13 a_36_137# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X14 a_987_507# a_572_93# a_688_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X15 a_1059_112# a_688_507# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X16 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 a_688_507# a_588_407# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X18 VDD a_2319_91# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X20 VDD a_1059_112# a_987_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X21 a_1059_112# a_688_507# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X22 VSS TE a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X23 a_2527_91# CLK a_2319_91# VSUBS nmos_6p0 w=0.625u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_4 Q TE VDD VSS CLK E
X0 VSS a_2319_91# Q VSUBS nmos_6p0 w=0.63u l=0.6u
X1 a_688_507# a_572_92# a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 a_2319_91# CLK VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS a_2319_91# Q VSUBS nmos_6p0 w=0.63u l=0.6u
X4 Q a_2319_91# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X5 VDD a_1059_112# a_2319_91# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD a_2319_91# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_919_137# a_588_407# a_688_507# VSUBS nmos_6p0 w=0.395u l=0.6u
X8 Q a_2319_91# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 Q a_2319_91# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD a_2319_91# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 Q a_2319_91# VSS VSUBS nmos_6p0 w=0.63u l=0.6u
X12 a_572_92# CLK VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X13 VSS a_572_92# a_588_407# VSUBS nmos_6p0 w=0.395u l=0.6u
X14 VSS a_1059_112# a_919_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X15 VSS a_1059_112# a_2527_91# VSUBS nmos_6p0 w=0.63u l=0.6u
X16 VDD a_572_92# a_588_407# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X17 a_572_92# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X18 a_36_137# E VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X19 a_987_507# a_572_92# a_688_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X20 a_1059_112# a_688_507# VDD w_n86_352# pmos_6p0 w=0.765u l=0.5u
X21 a_244_475# TE VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X22 a_688_507# a_588_407# a_448_475# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X23 a_448_475# E a_244_475# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X24 VDD a_1059_112# a_987_507# w_n86_352# pmos_6p0 w=0.765u l=0.5u
X25 a_1059_112# a_688_507# VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X26 VSS TE a_36_137# VSUBS nmos_6p0 w=0.395u l=0.6u
X27 a_2527_91# CLK a_2319_91# VSUBS nmos_6p0 w=0.63u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__icgtp_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD
X0 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 VSS ZN I VDD
X0 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_12 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_16 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X20 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X25 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X26 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X28 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X29 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X30 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_20.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_20 VSS ZN I VDD
X0 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X15 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X26 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X29 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X31 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X32 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X33 ZN I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 ZN I VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X35 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X36 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X37 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X38 VDD I ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X39 VSS I ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__inv_20.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 VDD VSS ZN EN I
X0 VSS a_1405_49# a_468_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 VDD a_428_560# ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_1405_49# I VDD w_n86_352# pmos_6p0 w=0.62u l=0.5u
X3 VSS a_468_93# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VDD EN a_36_93# w_n86_352# pmos_6p0 w=0.62u l=0.5u
X5 a_468_93# a_36_93# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_428_560# EN VDD w_n86_352# pmos_6p0 w=0.62u l=0.5u
X7 VDD a_1405_49# a_428_560# w_n86_352# pmos_6p0 w=0.62u l=0.5u
X8 a_468_93# a_36_93# a_428_560# w_n86_352# pmos_6p0 w=0.62u l=0.5u
X9 a_1405_49# I VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X10 a_428_560# EN a_468_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VSS EN a_36_93# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_2 VDD VSS ZN EN I
X0 VDD EN a_38_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 VDD a_986_24# a_479_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X2 a_986_24# I VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X3 ZN a_479_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X4 VSS a_470_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_479_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_470_68# a_38_68# a_479_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 VDD a_479_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X8 a_479_497# EN a_470_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VSS EN a_38_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS a_986_24# a_470_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 ZN a_470_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_470_68# a_38_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_986_24# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_3.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_3 VDD VSS ZN EN I
X0 VSS I a_938_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_479_68# a_47_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS a_938_68# a_479_68# VSUBS nmos_6p0 w=0.54u l=0.6u
X3 VDD I a_938_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 ZN a_488_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X5 ZN a_488_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X6 a_488_497# a_938_68# VDD w_n86_352# pmos_6p0 w=1.005u l=0.5u
X7 ZN a_479_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_488_497# EN a_479_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD a_488_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X10 VDD a_938_68# a_488_497# w_n86_352# pmos_6p0 w=1.005u l=0.5u
X11 VSS EN a_47_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_479_68# a_938_68# VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X13 ZN a_479_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD EN a_47_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 a_488_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_479_68# a_47_68# a_488_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 VSS a_479_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_3.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_4 VDD VSS ZN EN I
X0 VDD a_901_68# a_477_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X1 a_468_68# a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VSS a_468_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS I a_901_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS a_901_68# a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN a_477_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X7 a_477_497# EN a_468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS a_468_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN a_477_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X10 VSS EN a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD a_477_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X12 VDD a_477_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X13 ZN a_468_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_468_68# a_901_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 VDD I a_901_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 VDD EN a_36_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_477_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 a_468_68# a_36_68# a_477_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 a_477_497# a_901_68# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_8.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_8 VDD VSS ZN EN I
X0 VDD a_1221_497# a_494_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X1 ZN a_471_68# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X2 a_471_68# a_1221_497# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X3 VDD a_494_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X4 VSS a_1221_497# a_471_68# VSUBS nmos_6p0 w=0.815u l=0.6u
X5 VDD a_494_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X6 ZN a_471_68# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X7 VSS I a_1221_497# VSUBS nmos_6p0 w=0.815u l=0.6u
X8 ZN a_494_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X9 ZN a_494_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X10 a_494_497# EN a_471_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VSS EN a_39_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_494_497# a_1221_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X13 VDD a_494_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X14 ZN a_471_68# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X15 VDD a_494_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X16 a_471_68# a_39_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X17 ZN a_494_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X18 ZN a_471_68# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X19 VDD EN a_39_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 ZN a_494_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X21 a_494_497# a_1221_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X22 VSS a_471_68# ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X23 a_1221_497# I VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X24 VSS a_1221_497# a_471_68# VSUBS nmos_6p0 w=0.815u l=0.6u
X25 a_494_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X26 VDD a_1221_497# a_494_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X27 VSS a_471_68# ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X28 VDD I a_1221_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X29 a_1221_497# I VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X30 VSS a_471_68# ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X31 a_471_68# a_1221_497# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X32 a_471_68# a_39_68# a_494_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X33 VSS a_471_68# ZN VSUBS nmos_6p0 w=0.815u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_8.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_12.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_12 VDD VSS ZN EN I
X0 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X1 a_918_68# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD I a_918_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X4 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X5 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X6 VSS a_918_68# a_478_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X9 VDD I a_918_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 a_501_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X13 a_478_68# a_46_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD a_918_68# a_501_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X15 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_501_497# a_918_68# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X17 VSS I a_918_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_478_68# a_46_68# a_501_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 VDD a_918_68# a_501_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X21 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X23 a_501_497# EN a_478_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X24 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_501_497# a_918_68# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X26 VSS a_918_68# a_478_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X27 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X28 VSS EN a_46_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X29 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X30 VDD a_918_68# a_501_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X31 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X32 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X33 VSS I a_918_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X34 a_478_68# a_918_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X35 VSS a_918_68# a_478_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X36 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X37 a_501_497# a_918_68# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X38 a_478_68# a_918_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X39 VSS a_478_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X40 VDD a_501_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X41 a_478_68# a_918_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X42 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X43 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X44 VDD EN a_46_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X45 a_918_68# I VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X46 ZN a_501_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X47 ZN a_478_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_12.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_16.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__invz_16 VDD VSS ZN EN I
X0 a_1239_497# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_1239_497# a_512_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X3 a_489_68# a_1239_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD I a_1239_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X8 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD EN a_57_68# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X11 VSS a_1239_497# a_489_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VDD a_1239_497# a_512_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X13 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X15 a_512_497# EN VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 VDD a_1239_497# a_512_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X17 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD I a_1239_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X20 a_489_68# a_1239_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_489_68# a_57_68# a_512_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X22 a_1239_497# I VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X24 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X25 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X26 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X27 a_512_497# a_1239_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X28 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X29 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X30 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X31 a_512_497# a_1239_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X32 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X33 a_489_68# a_57_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 VSS a_1239_497# a_489_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X35 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X36 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X37 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X38 VDD a_1239_497# a_512_497# w_n86_352# pmos_6p0 w=1.18u l=0.5u
X39 VSS I a_1239_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X40 VSS I a_1239_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X41 a_512_497# EN a_489_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X42 VSS a_1239_497# a_489_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X43 a_512_497# a_1239_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X44 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X45 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X46 VSS EN a_57_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X47 a_1239_497# I VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X48 VSS a_1239_497# a_489_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X49 a_512_497# a_1239_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X50 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X51 a_489_68# a_1239_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X52 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X53 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X54 VSS a_489_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X55 VDD a_512_497# ZN w_n86_352# pmos_6p0 w=1.18u l=0.5u
X56 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X57 ZN a_489_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X58 a_1239_497# I VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X59 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
X60 a_489_68# a_1239_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X61 ZN a_512_497# VDD w_n86_352# pmos_6p0 w=1.18u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__invz_16.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 Q VDD VSS D E
X0 a_1404_42# a_1020_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X1 VDD E a_36_87# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X2 a_484_591# a_36_87# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X3 a_1404_42# a_1020_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 a_872_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_872_86# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X6 a_1020_590# a_484_591# a_872_86# VSUBS nmos_6p0 w=0.395u l=0.6u
X7 VSS a_1404_42# a_1264_86# VSUBS nmos_6p0 w=0.465u l=0.6u
X8 VDD a_1020_590# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_1020_590# a_36_87# a_872_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 VDD a_1404_42# a_1224_590# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X11 VSS E a_36_87# VSUBS nmos_6p0 w=0.46u l=0.6u
X12 a_1224_590# a_484_591# a_1020_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 a_484_591# a_36_87# VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X14 a_1264_86# a_36_87# a_1020_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X15 VSS a_1020_590# Q VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latq_2 Q VDD VSS D E
X0 VDD E a_36_87# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X1 a_484_591# a_36_87# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X2 a_1364_316# a_1020_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_872_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X4 VDD a_1364_316# a_1224_590# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X5 a_872_86# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X6 a_1020_590# a_484_591# a_872_86# VSUBS nmos_6p0 w=0.395u l=0.6u
X7 a_1364_316# a_1020_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X8 VSS a_1364_316# a_1264_86# VSUBS nmos_6p0 w=0.465u l=0.6u
X9 VSS a_1020_590# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_1020_590# a_36_87# a_872_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X11 VSS E a_36_87# VSUBS nmos_6p0 w=0.46u l=0.6u
X12 a_1224_590# a_484_591# a_1020_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 a_484_591# a_36_87# VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X14 a_1264_86# a_36_87# a_1020_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X15 Q a_1020_590# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 Q a_1020_590# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VDD a_1020_590# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latq_4 Q VDD VSS D E
X0 a_1404_42# a_1020_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X1 a_484_591# a_36_87# VSS VSUBS nmos_6p0 w=0.39u l=0.6u
X2 Q a_1020_590# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_1404_42# a_1020_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 a_872_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 VDD a_1020_590# a_1404_42# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X6 a_872_86# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X7 Q a_1020_590# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_1020_590# a_484_591# a_872_86# VSUBS nmos_6p0 w=0.395u l=0.6u
X9 VSS a_1020_590# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS a_1020_590# a_1404_42# VSUBS nmos_6p0 w=0.465u l=0.6u
X11 VSS a_1020_590# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VSS a_1404_42# a_1264_86# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VDD a_1020_590# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_1020_590# a_36_87# a_872_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X15 VSS E a_36_87# VSUBS nmos_6p0 w=0.46u l=0.6u
X16 Q a_1020_590# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VDD E a_36_87# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X18 VDD a_1020_590# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_1224_590# a_484_591# a_1020_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 Q a_1020_590# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_484_591# a_36_87# VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X22 a_1264_86# a_36_87# a_1020_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X23 VDD a_1404_42# a_1224_590# w_n86_352# pmos_6p0 w=0.925u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 Q RN VSS E VDD D
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 Q a_1820_139# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X3 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X4 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 Q a_1820_139# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X7 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X8 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X9 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X10 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X11 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X12 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VSS a_1112_24# a_1820_139# VSUBS nmos_6p0 w=0.465u l=0.6u
X14 VDD a_1112_24# a_1820_139# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X15 a_1112_24# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_2 RN Q D VDD E VSS
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 Q a_1820_139# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X3 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X4 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 Q a_1820_139# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD a_1820_139# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X8 VSS a_1820_139# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X10 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X11 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X12 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X13 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X14 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X15 VSS a_1112_24# a_1820_139# VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VDD a_1112_24# a_1820_139# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 a_1112_24# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X18 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X19 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_4 Q RN VDD VSS D E
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 a_2108_93# a_1112_24# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X2 a_2108_93# a_1112_24# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X3 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X4 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X6 VDD a_1112_24# a_2108_93# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X7 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X8 VSS a_388_590# a_1112_24# VSUBS nmos_6p0 w=0.465u l=0.6u
X9 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X10 VSS a_2108_93# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X12 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X13 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X14 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X15 VSS a_1112_24# a_2108_93# VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VSS a_2108_93# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X17 Q a_2108_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_1112_24# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X19 Q a_2108_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X20 Q a_2108_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X22 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 VDD a_2108_93# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X25 VDD a_2108_93# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X26 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X27 Q a_2108_93# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 VDD a_388_590# a_1112_24# w_n86_352# pmos_6p0 w=0.925u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 SETN Q RN VSS E VDD D
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X3 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X4 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X6 Q a_2044_139# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X8 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X9 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X10 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X11 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X12 a_1112_24# SETN a_1660_93# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 a_1660_93# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X14 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X15 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X16 VDD SETN a_1112_24# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 VSS a_1112_24# a_2044_139# VSUBS nmos_6p0 w=0.465u l=0.6u
X19 VDD a_1112_24# a_2044_139# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X20 Q a_2044_139# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 RN SETN Q D VSS VDD E
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 VSS a_2016_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X3 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X4 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 VSS a_1112_24# a_2016_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X7 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X8 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X9 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X10 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X11 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X12 Q a_2016_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_1660_93# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X14 VDD a_2016_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X16 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X17 a_1112_24# SETN a_1660_93# VSUBS nmos_6p0 w=0.465u l=0.6u
X18 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X19 VDD SETN a_1112_24# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X20 Q a_2016_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X22 VDD a_1112_24# a_2016_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 RN SETN Q D VSS VDD E
X0 a_1232_93# a_1112_24# a_1064_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X1 Q a_2224_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD a_1112_24# a_2224_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_388_590# a_36_79# a_780_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X4 a_1064_93# a_36_79# a_388_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 VSS RN a_1232_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X6 a_2224_68# a_1112_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 Q a_2224_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_1132_590# E a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 a_504_93# RN VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X10 a_672_93# D a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X11 a_388_590# E a_672_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X12 VDD a_1112_24# a_1132_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X14 Q a_2224_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_1660_93# a_388_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X17 VDD RN a_388_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 VDD a_2224_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_1112_24# SETN a_1660_93# VSUBS nmos_6p0 w=0.465u l=0.6u
X20 VSS a_2224_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_780_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X22 VDD SETN a_1112_24# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X23 Q a_2224_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 VSS a_1112_24# a_2224_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_1112_24# a_388_590# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X26 VSS a_2224_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X27 VDD a_2224_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X28 a_2224_68# a_1112_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latrsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_1 Q VSS SETN VDD D E
X0 a_944_35# a_632_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X1 a_896_93# a_36_79# a_632_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 VDD SETN a_944_35# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X3 VSS a_944_35# a_896_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X4 a_1324_79# a_632_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X5 Q a_1708_139# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_944_35# SETN a_1324_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X7 Q a_1708_139# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_484_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 a_504_93# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X10 a_632_590# E a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X11 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X12 VSS a_944_35# a_1708_139# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VDD a_944_35# a_1708_139# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X14 VDD a_944_35# a_836_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X15 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X16 a_632_590# a_36_79# a_484_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X17 a_836_590# E a_632_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_2 Q VSS SETN VDD D E
X0 a_944_35# a_632_590# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X1 Q a_1668_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_896_93# a_36_79# a_632_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X3 VDD SETN a_944_35# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X4 VSS a_944_35# a_896_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X5 VDD E a_36_79# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X6 VDD a_1668_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_1324_79# a_632_590# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X8 a_944_35# SETN a_1324_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X9 a_484_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 a_504_93# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X11 a_632_590# E a_504_93# VSUBS nmos_6p0 w=0.395u l=0.6u
X12 VSS E a_36_79# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VDD a_944_35# a_1668_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD a_944_35# a_836_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X15 VSS a_944_35# a_1668_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_632_590# a_36_79# a_484_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X17 a_836_590# E a_632_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 VSS a_1668_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X19 Q a_1668_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__latsnq_4 Q D VDD SETN VSS E
X0 VSS a_944_35# a_1888_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VSS a_944_35# a_896_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X2 a_1324_68# a_632_590# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VDD E a_36_139# w_n86_352# pmos_6p0 w=0.925u l=0.5u
X4 a_944_35# SETN a_1324_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS a_1888_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X6 Q a_1888_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 a_896_153# a_36_139# a_632_590# VSUBS nmos_6p0 w=0.395u l=0.6u
X8 VDD a_1888_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_484_590# D VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 a_944_35# a_632_590# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 Q a_1888_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 VDD SETN a_944_35# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VDD a_1888_68# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_1888_68# a_944_35# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VDD a_944_35# a_836_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X16 VSS E a_36_139# VSUBS nmos_6p0 w=0.465u l=0.6u
X17 VSS a_1888_68# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD a_944_35# a_1888_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_632_590# E a_504_153# VSUBS nmos_6p0 w=0.395u l=0.6u
X20 a_632_590# a_36_139# a_484_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X21 a_836_590# E a_632_590# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X22 a_1888_68# a_944_35# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_504_153# D VSS VSUBS nmos_6p0 w=0.395u l=0.6u
X24 Q a_1888_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 Q a_1888_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__latsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_1 S VDD VSS Z I0 I1
X0 a_896_104# a_592_407# a_124_24# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 a_124_24# a_592_407# a_537_593# w_n86_352# pmos_6p0 w=0.615u l=0.5u
X2 a_896_593# S a_124_24# w_n86_352# pmos_6p0 w=0.615u l=0.5u
X3 VSS a_124_24# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_124_24# S a_504_104# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VDD a_124_24# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD I0 a_896_593# w_n86_352# pmos_6p0 w=0.615u l=0.5u
X7 a_592_407# S VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_504_104# I1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_592_407# S VDD w_n86_352# pmos_6p0 w=0.615u l=0.5u
X10 a_537_593# I1 VDD w_n86_352# pmos_6p0 w=0.615u l=0.5u
X11 VSS I0 a_896_104# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1
X0 VSS I0 a_1084_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_1084_68# a_848_380# a_124_24# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS a_124_24# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_124_24# a_848_380# a_692_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_1152_472# S a_124_24# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_692_68# I1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_124_24# S a_692_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 Z a_124_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_848_380# S VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD a_124_24# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VDD I0 a_1152_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_692_472# I1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_848_380# S VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 Z a_124_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 S VDD VSS Z I0 I1
X0 a_1543_68# a_1307_380# a_135_24# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VDD a_135_24# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS a_135_24# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_1151_472# I1 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS a_135_24# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_1151_68# I1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD a_135_24# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 Z a_135_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS I0 a_1543_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 Z a_135_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_135_24# a_1307_380# a_1151_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 a_1307_380# S VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_1611_472# S a_135_24# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 Z a_135_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD I0 a_1611_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_135_24# S a_1151_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_1307_380# S VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 Z a_135_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 VSS VDD I2 I1 S0 I3 S1 Z
X0 a_224_515# I2 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X1 a_348_112# S0 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X2 a_2521_156# I1 VDD w_n86_352# pmos_6p0 w=0.565u l=0.5u
X3 VSS S1 a_1525_369# VSUBS nmos_6p0 w=0.365u l=0.6u
X4 VDD I0 a_2929_515# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X5 a_2929_515# a_348_112# a_1901_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X6 a_1081_112# S1 a_468_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X7 a_1901_156# a_348_112# a_2521_156# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X8 a_1901_156# a_1525_369# a_1081_112# VSUBS nmos_6p0 w=0.365u l=0.6u
X9 VDD S1 a_1525_369# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X10 a_2929_515# S0 a_1901_156# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X11 Z a_1081_112# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X12 VSS I3 a_712_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X13 Z a_1081_112# VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X14 VSS I0 a_2929_515# VSUBS nmos_6p0 w=0.365u l=0.6u
X15 VDD I3 a_712_156# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X16 a_1901_156# S0 a_2521_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X17 a_468_156# a_348_112# a_224_515# VSUBS nmos_6p0 w=0.365u l=0.6u
X18 a_468_156# S0 a_224_515# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X19 a_224_515# I2 VDD w_n86_352# pmos_6p0 w=0.565u l=0.5u
X20 a_1901_156# S1 a_1081_112# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X21 a_712_156# S0 a_468_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X22 a_348_112# S0 VDD w_n86_352# pmos_6p0 w=0.565u l=0.5u
X23 a_1081_112# a_1525_369# a_468_156# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X24 a_712_156# a_348_112# a_468_156# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X25 a_2521_156# I1 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 VSS VDD I2 I1 S0 I3 S1 Z
X0 a_1108_112# a_1772_369# a_468_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X1 a_224_472# I2 VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_2147_156# S0 a_2768_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X3 a_224_472# I2 VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X4 a_468_156# S0 a_224_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X5 a_348_112# S0 VDD w_n86_352# pmos_6p0 w=0.595u l=0.5u
X6 VSS I0 a_3176_509# VSUBS nmos_6p0 w=0.365u l=0.6u
X7 a_3176_509# S0 a_2147_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X8 Z a_1108_112# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X9 a_728_472# a_348_112# a_468_156# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X10 VSS I3 a_728_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X11 a_2768_156# I1 VDD w_n86_352# pmos_6p0 w=0.595u l=0.5u
X12 Z a_1108_112# VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X13 a_2147_156# a_348_112# a_2768_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X14 a_3176_509# a_348_112# a_2147_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X15 VDD I3 a_728_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X16 VDD a_1108_112# Z w_n86_352# pmos_6p0 w=0.78u l=0.5u
X17 a_2768_156# I1 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X18 a_468_156# a_348_112# a_224_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X19 VDD I0 a_3176_509# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X20 a_2147_156# S1 a_1108_112# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X21 a_2147_156# a_1772_369# a_1108_112# VSUBS nmos_6p0 w=0.365u l=0.6u
X22 a_728_472# S0 a_468_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X23 a_1108_112# S1 a_468_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X24 VDD S1 a_1772_369# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X25 VSS a_1108_112# Z VSUBS nmos_6p0 w=0.38u l=0.6u
X26 a_348_112# S0 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X27 VSS S1 a_1772_369# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 VSS VDD I2 I1 S0 I3 S1 Z
X0 a_224_472# I2 VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X1 VSS a_1108_112# Z VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_348_112# S0 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X3 VSS S1 a_2220_369# VSUBS nmos_6p0 w=0.365u l=0.6u
X4 a_224_472# I2 VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X5 a_1108_112# a_2220_369# a_468_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X6 a_468_156# S0 a_224_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X7 a_2595_156# S0 a_3216_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X8 Z a_1108_112# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X9 a_728_472# a_348_112# a_468_156# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X10 VSS I3 a_728_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X11 Z a_1108_112# VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X12 a_348_112# S0 VDD w_n86_352# pmos_6p0 w=0.595u l=0.5u
X13 Z a_1108_112# VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X14 a_3216_156# I1 VSS VSUBS nmos_6p0 w=0.365u l=0.6u
X15 VDD I3 a_728_472# w_n86_352# pmos_6p0 w=0.78u l=0.5u
X16 VDD a_1108_112# Z w_n86_352# pmos_6p0 w=0.78u l=0.5u
X17 VSS I0 a_3624_509# VSUBS nmos_6p0 w=0.365u l=0.6u
X18 a_3216_156# I1 VDD w_n86_352# pmos_6p0 w=0.595u l=0.5u
X19 Z a_1108_112# VDD w_n86_352# pmos_6p0 w=0.78u l=0.5u
X20 a_468_156# a_348_112# a_224_472# VSUBS nmos_6p0 w=0.38u l=0.6u
X21 a_2595_156# a_348_112# a_3216_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X22 VDD a_1108_112# Z w_n86_352# pmos_6p0 w=0.78u l=0.5u
X23 a_3624_509# S0 a_2595_156# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X24 a_728_472# S0 a_468_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X25 a_2595_156# S1 a_1108_112# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X26 VDD I0 a_3624_509# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X27 a_2595_156# a_2220_369# a_1108_112# VSUBS nmos_6p0 w=0.365u l=0.6u
X28 VSS a_1108_112# Z VSUBS nmos_6p0 w=0.38u l=0.6u
X29 a_3624_509# a_348_112# a_2595_156# VSUBS nmos_6p0 w=0.365u l=0.6u
X30 VDD S1 a_2220_369# w_n86_352# pmos_6p0 w=0.595u l=0.5u
X31 a_1108_112# S1 a_468_156# VSUBS nmos_6p0 w=0.365u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__mux4_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2
X0 ZN A2 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X1 ZN A1 a_245_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD A1 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X3 a_245_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2
X0 ZN A1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_244_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A2 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X3 VDD A1 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X4 a_652_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS A2 a_652_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN A1 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X7 VDD A2 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 VDD VSS ZN A1 A2
X0 VSS A2 a_1468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN A2 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X2 VDD A1 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X3 ZN A1 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X4 VSS A2 a_661_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN A1 a_260_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD A2 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X7 a_1468_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X8 ZN A2 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X9 VDD A1 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X10 ZN A1 a_1060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 ZN A1 VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
X12 VDD A2 ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X13 a_661_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_1060_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_260_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2
X0 a_271_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_455_68# A2 a_271_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A1 a_455_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A3 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X4 VDD A2 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X5 ZN A1 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2
X0 ZN A3 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X1 VDD A2 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X2 a_452_68# A2 a_276_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A1 a_452_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN A1 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X5 VDD A1 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X6 a_1044_68# A2 a_860_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_860_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X8 ZN A2 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X9 VDD A3 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X10 VSS A3 a_1044_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_276_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2
X0 ZN A2 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X1 a_672_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD A3 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X3 ZN A1 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X4 VDD A1 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X5 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN A2 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X7 a_36_68# A2 a_672_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_1732_68# A2 a_1528_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN A3 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X10 a_244_68# A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_1528_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VDD A2 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X13 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A3 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X15 VDD A1 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X16 a_1100_68# A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 ZN A1 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X18 ZN A3 VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X19 ZN A1 a_1732_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VSS A3 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X21 VDD A2 ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X22 VSS A3 a_1100_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand3_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A3 A4 VDD VSS ZN A1 A2
X0 a_469_68# A3 a_275_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN A1 a_673_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A4 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X3 VDD A3 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X4 ZN A2 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X5 VDD A1 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X6 a_275_68# A4 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_673_68# A2 a_469_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2
X0 ZN A2 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X1 VSS A4 a_1458_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD A3 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X3 ZN A4 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X4 a_1458_68# A3 a_1254_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_632_68# A2 a_438_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD A4 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X7 a_244_68# A4 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 ZN A3 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X9 a_438_68# A3 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD A2 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X11 ZN A1 a_632_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN A1 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X13 VDD A1 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X14 a_1060_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1254_68# A2 a_1060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A3 A4 VDD VSS ZN A1 A2
X0 VDD A4 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X1 ZN A2 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X2 ZN A1 a_2780_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_2780_68# A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN A4 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X5 VDD A1 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X6 a_36_68# A2 a_3276_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD A3 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X8 a_1662_68# A3 a_1468_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN A1 a_1866_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 ZN A2 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X11 VDD A1 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X12 VSS A4 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X13 ZN A3 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X14 a_244_68# A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1468_68# A4 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD A4 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X17 a_1866_68# A2 a_1662_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 ZN A4 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X19 ZN A1 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X20 a_3276_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_652_68# A4 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_36_68# A3 a_652_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 VDD A2 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X24 VDD A3 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
X25 VSS A4 a_1060_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X26 ZN A3 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X27 a_2372_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X28 a_36_68# A2 a_2372_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X29 ZN A1 VDD w_n86_352# pmos_6p0 w=0.845u l=0.5u
X30 a_1060_68# A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X31 VDD A2 ZN w_n86_352# pmos_6p0 w=0.845u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nand4_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2
X0 a_224_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 ZN A2 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X2 ZN A1 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS A1 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2
X0 ZN A2 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X1 a_672_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X3 ZN A1 a_234_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS A1 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
X5 a_234_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD A2 a_672_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VSS A2 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 VDD VSS ZN A1 A2
X0 VSS A2 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
X1 VSS A1 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
X2 ZN A2 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X3 a_1140_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN A1 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X5 ZN A1 a_1140_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 ZN A2 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X7 a_1588_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VDD A2 a_1588_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 ZN A1 VSS VSUBS nmos_6p0 w=0.565u l=0.6u
X10 a_244_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN A1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_692_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS A2 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
X14 VDD A2 a_692_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VSS A1 ZN VSUBS nmos_6p0 w=0.565u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2
X0 ZN A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X1 ZN A1 a_448_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 ZN A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_244_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_448_472# A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS A2 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2
X0 ZN A1 a_468_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X2 VSS A3 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_468_472# A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD A3 a_1130_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_1130_472# A2 a_906_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 ZN A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X7 a_244_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X9 ZN A2 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X10 VSS A2 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X11 a_906_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2
X0 a_1568_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 ZN A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X2 VSS A1 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X3 ZN A2 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 a_224_472# A2 a_36_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X6 ZN A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X7 a_672_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 ZN A1 a_36_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 ZN A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X10 VDD A3 a_1120_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 ZN A1 a_1792_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 VSS A2 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VSS A3 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X14 a_1792_472# A2 a_1568_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VSS A1 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VDD A3 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VSS A2 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X18 a_36_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 VSS A3 ZN VSUBS nmos_6p0 w=0.465u l=0.6u
X20 a_1120_472# A2 a_36_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 ZN A2 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X22 a_36_472# A2 a_672_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 a_36_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor3_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A3 A4 VDD VSS ZN A1 A2
X0 a_672_472# A2 a_448_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS A1 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X2 VSS A3 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_244_472# A4 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 a_448_472# A3 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X6 ZN A4 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X7 ZN A1 a_672_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A3 A4 VDD VSS ZN A1 A2
X0 ZN A1 a_1213_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_683_472# A4 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS A3 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_1213_472# A2 a_943_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS A2 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X5 a_943_472# A3 a_683_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS A1 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_1661_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VSS A4 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_57_472# A2 a_1661_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 ZN A1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VDD A4 a_245_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X13 ZN A4 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_245_472# A3 a_57_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 ZN A3 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2
X0 ZN A3 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X1 VDD A4 a_1212_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X2 VSS A1 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_692_473# A4 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 ZN A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VSS A2 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X6 ZN A1 a_3220_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 ZN A1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_66_473# A3 a_692_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 VSS A3 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X10 a_2180_473# A2 a_1920_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X11 a_3220_473# A2 a_66_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X12 a_3740_473# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X13 a_1212_473# A3 a_66_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X14 VSS A3 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X15 ZN A1 a_2180_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X16 a_66_473# A2 a_2700_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X17 a_66_473# A2 a_3740_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X18 ZN A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X19 VDD A4 a_254_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X20 VSS A4 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X21 ZN A1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_1660_473# A4 VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X23 a_2700_473# A1 ZN w_n86_352# pmos_6p0 w=1.215u l=0.5u
X24 VSS A1 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_254_473# A3 a_66_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X26 VSS A4 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X27 a_1920_473# A3 a_1660_473# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X28 VSS A2 ZN VSUBS nmos_6p0 w=0.36u l=0.6u
X29 ZN A4 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X30 ZN A3 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X31 ZN A4 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__nor4_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS
X0 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VDD B ZN w_n86_352# pmos_6p0 w=1.13u l=0.5u
X4 a_244_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN A1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A2 ZN A1 VSS B VDD
X0 VDD A2 a_1164_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A1 a_692_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_1164_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 ZN B VDD w_n86_352# pmos_6p0 w=0.955u l=0.5u
X10 a_692_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 VDD B ZN w_n86_352# pmos_6p0 w=0.955u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 B VDD VSS A1 ZN A2
X0 a_1612_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN B VDD w_n86_352# pmos_6p0 w=0.955u l=0.5u
X2 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VDD B ZN w_n86_352# pmos_6p0 w=0.955u l=0.5u
X6 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_224_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 ZN B VDD w_n86_352# pmos_6p0 w=0.955u l=0.5u
X9 ZN A1 a_224_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_716_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 VDD B ZN w_n86_352# pmos_6p0 w=0.955u l=0.5u
X13 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A2 a_716_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_1164_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 VDD A2 a_1612_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X23 ZN A1 a_1164_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai21_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1
X0 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN B1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_244_472# B2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_692_472# A1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD A2 a_692_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 B2 VDD VSS ZN A1 A2 B1
X0 a_1612_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VDD A2 a_1612_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 ZN B1 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_672_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 a_1140_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_244_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 ZN A1 a_1140_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 VDD B2 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 B1 VDD VSS ZN A1 A2 B2
X0 a_2036_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_1568_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 ZN A1 a_2036_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 ZN B1 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 a_672_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 a_2508_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VDD A2 a_2508_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X15 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_2956_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 ZN A1 a_2956_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD B2 a_1568_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X21 a_244_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X22 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 VDD B2 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X24 a_3404_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X25 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X26 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X27 a_1120_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X28 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X29 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X30 ZN B1 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X31 VDD A2 a_3404_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai22_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 VDD ZN B A1 A2 VSS A3
X0 ZN A3 a_244_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X1 a_468_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_244_69# A2 ZN VSUBS nmos_6p0 w=0.815u l=0.6u
X3 a_780_497# A2 a_468_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 ZN A1 a_244_69# VSUBS nmos_6p0 w=0.815u l=0.6u
X5 VDD A3 a_780_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_244_69# B VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X7 ZN B VDD w_n86_352# pmos_6p0 w=1.13u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1
X0 a_1612_497# A2 a_1388_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A1 a_960_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_1388_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 VDD A3 a_1612_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_960_497# A2 a_692_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN B VDD w_n86_352# pmos_6p0 w=1.08u l=0.5u
X13 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_692_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 VDD B ZN w_n86_352# pmos_6p0 w=1.08u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A3 B VDD VSS ZN A1 A2
X0 a_1612_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_1184_497# A2 a_940_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_56_497# A2 a_1612_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_2060_497# A2 a_56_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 ZN A1 a_2060_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 a_36_68# B VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD B ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_2508_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 ZN B VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_56_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 ZN B VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X20 VDD A3 a_56_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X21 VDD B ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X22 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X23 VDD A3 a_56_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X24 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X26 a_940_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X27 VSS B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X28 ZN A1 a_1184_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X29 a_56_497# A2 a_2508_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X30 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X31 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai31_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2
X0 ZN B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_224_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS A2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_244_68# B2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_468_472# A2 a_224_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 ZN A1 a_468_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_244_68# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_244_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_916_472# B1 ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VDD B2 a_916_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A3 B1 B2 VDD VSS ZN A1 A2
X0 a_36_68# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_36_68# B2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN B1 a_1588_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_36_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_2060_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 VSS A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_468_497# A2 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 VSS A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD B2 a_2060_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 VDD A3 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 a_1588_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 ZN B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_244_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 a_36_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X15 ZN A1 a_468_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_1120_497# A2 a_896_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_36_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_896_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 ZN B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A3 B1 B2 VDD VSS ZN A1 A2
X0 VSS A3 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_77_68# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_1161_497# A2 a_87_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_77_68# B2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS A2 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN A1 a_1853_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 VSS A1 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VSS A3 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD B2 a_4401_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 ZN B2 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS A1 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_77_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN A1 a_87_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 ZN B2 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A3 a_1161_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 a_77_68# B2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X16 ZN B1 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_87_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 a_77_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_1609_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 ZN B1 a_3077_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X21 ZN B1 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_1853_497# A2 a_1609_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 a_77_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X24 a_3505_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X25 ZN B1 a_3953_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X26 a_77_68# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X27 VDD B2 a_3505_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X28 VDD A3 a_285_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X29 a_77_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X30 a_77_68# B1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X31 a_713_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X32 a_3953_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X33 a_77_68# A3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 a_285_497# A2 a_87_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X35 VSS A2 a_77_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X36 a_87_497# A2 a_713_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X37 a_3077_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X38 a_4401_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X39 a_87_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai32_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A3 B1 B2 B3 VDD VSS ZN A1 A2
X0 a_1228_497# A2 a_896_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN A1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD A3 a_1228_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VSS B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_224_497# B3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_244_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN B1 a_448_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_244_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_244_68# B3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN A3 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_448_497# B2 a_224_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 a_896_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_2 A3 B1 B2 B3 VDD VSS ZN A1 A2
X0 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_1856_497# A2 a_1588_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_468_497# B2 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_2508_497# A2 a_2284_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VSS B3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD B3 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 a_2284_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 a_1588_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X13 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A3 a_2508_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 ZN A1 a_1856_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_244_497# B3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X18 ZN B1 a_468_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 a_1120_497# B2 a_896_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X20 a_36_68# B3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_896_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A3 B1 B2 B3 VDD VSS ZN A1 A2
X0 ZN B1 a_1792_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 a_4808_497# A2 a_2848_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_46_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VDD A3 a_4808_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_1568_497# B3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_3932_497# A2 a_3688_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 a_36_68# B3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD B3 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 a_672_497# B3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 VSS B3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_2848_497# A2 a_5256_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD A3 a_3932_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X20 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_4360_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 VSS B3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X24 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X26 a_2848_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X27 a_36_68# A3 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X28 a_1792_497# B2 a_1568_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X29 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X30 a_244_497# B2 a_46_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X31 ZN A1 a_2848_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X32 VSS B1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X33 a_46_497# B2 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X34 ZN A1 a_2848_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X35 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X36 a_3688_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X37 a_46_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X38 a_36_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X39 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X40 ZN A3 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X41 a_1120_497# B2 a_46_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X42 a_2848_497# A2 a_4360_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X43 a_36_68# B3 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X44 ZN B1 a_46_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X45 a_5256_497# A3 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X46 VDD B3 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X47 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai33_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2
X0 VSS C a_692_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_692_68# B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_244_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VDD B ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X6 ZN A1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 ZN C VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS
X0 ZN B VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X1 VDD C ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X2 VSS C a_1229_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN A1 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 ZN C VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X5 a_1229_68# B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD B ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X7 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_716_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 a_36_68# B a_1657_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD A2 a_716_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_244_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_1657_68# C VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2
X0 a_1612_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_3368_68# C VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 ZN B VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X5 a_2960_68# B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN A1 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 VDD A2 a_1612_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 VDD C ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X9 ZN A1 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_716_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 VDD A2 a_716_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X12 ZN C VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X13 a_2124_68# B a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD C ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X15 ZN A2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VSS C a_2960_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VDD B ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X19 ZN C VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X20 a_36_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_1164_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X22 ZN B VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X23 VDD B ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X24 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_36_68# B a_3368_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X26 a_244_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X27 VSS C a_2124_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X28 a_36_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X29 ZN A1 a_1164_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X30 a_36_68# B a_2552_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X31 a_2552_68# C VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai211_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 B1 C VDD VSS ZN A1 A2 B2
X0 a_36_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_692_68# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_692_68# C a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_932_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS B2 a_36_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 ZN A2 a_692_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_244_472# B2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 ZN A1 a_932_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 VDD C ZN w_n86_352# pmos_6p0 w=0.945u l=0.5u
X9 ZN B1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A2 A1 B1 C B2 ZN VSS VDD
X0 VSS B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VSS B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN A1 a_2160_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 a_224_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_1732_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 ZN B1 a_224_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_672_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_244_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_244_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_1076_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_1076_93# C a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD C ZN w_n86_352# pmos_6p0 w=0.985u l=0.5u
X12 a_2160_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 ZN C VDD w_n86_352# pmos_6p0 w=0.985u l=0.5u
X14 VDD B2 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 VDD A2 a_1732_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 ZN A1 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 a_1076_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X18 a_244_68# C a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 ZN A2 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 B1 B2 C VDD VSS ZN A2
X0 ZN A1 a_4400_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 VSS B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_1568_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VDD C ZN w_n86_352# pmos_6p0 w=0.935u l=0.5u
X4 VSS B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_1972_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN C VDD w_n86_352# pmos_6p0 w=0.935u l=0.5u
X7 a_244_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 VDD B2 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 ZN A1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD A2 a_3076_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 a_244_68# C a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_1972_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_672_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 a_244_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X15 ZN A1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 ZN B1 a_1568_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_3504_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 VDD A2 a_3952_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 a_244_68# B1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X20 ZN A2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_1972_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 ZN A1 a_3504_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 ZN A2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X24 a_244_68# B2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X25 a_1972_93# C a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X26 a_3952_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X27 VDD C ZN w_n86_352# pmos_6p0 w=0.935u l=0.5u
X28 a_1972_93# C a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X29 a_244_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X30 ZN B1 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X31 ZN C VDD w_n86_352# pmos_6p0 w=0.935u l=0.5u
X32 a_3076_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X33 a_4400_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X34 a_1972_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X35 VSS B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X36 a_1120_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X37 VSS B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X38 VDD B2 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X39 a_244_68# C a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai221_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 B1 B2 C1 C2 VDD VSS ZN A1 A2
X0 a_816_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 a_244_68# B1 a_628_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS C1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_628_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_628_93# B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_244_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VDD B2 a_816_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 a_244_497# C2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 a_1284_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 ZN A1 a_1284_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 ZN C1 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 ZN A2 a_628_93# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 B1 B2 C1 C2 VDD VSS ZN A1 A2
X0 VSS C1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_2180_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_2608_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 VSS C2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VDD C2 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 ZN B1 a_1712_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 ZN A1 a_2608_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 ZN A2 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_672_497# C2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X9 a_244_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 a_244_68# C1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_1076_93# B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_1076_93# B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD B2 a_1284_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 a_1076_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X15 a_244_497# C1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_1712_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 ZN C1 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 a_1284_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X19 a_1076_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X20 a_244_68# B2 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X21 a_244_68# B1 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X22 VDD A2 a_2180_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X23 ZN A1 a_1076_93# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 B1 B2 C1 C2 VDD VSS ZN A1 A2
X0 ZN B1 a_3504_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 VDD A2 a_4848_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 VSS C1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_1568_497# C2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_2180_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_2608_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X6 a_3972_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X7 ZN B1 a_2608_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 VSS C2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_1972_93# B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X10 ZN A2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_244_68# C1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 a_1972_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_1972_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_3056_497# B1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X15 VDD C2 a_244_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X16 a_244_68# B1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X17 VDD B2 a_3056_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X18 a_244_68# B2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 a_1972_93# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X20 a_672_497# C2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X21 a_244_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 ZN A1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 ZN C1 a_1568_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X24 ZN A1 a_5296_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X25 a_3504_497# B2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X26 VDD A2 a_3972_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X27 a_244_68# C1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X28 a_244_68# B2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X29 ZN A2 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X30 a_1972_93# A1 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X31 a_244_68# C2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X32 a_1972_93# B1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X33 a_1972_93# B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X34 a_244_497# C1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X35 ZN C1 a_672_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X36 a_4400_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X37 a_1972_93# B2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X38 VSS C1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X39 ZN A1 a_4400_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X40 a_1120_497# C1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X41 a_5296_497# A2 VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X42 VSS C2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X43 ZN A1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
X44 VDD C2 a_1120_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X45 VDD B2 a_2180_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X46 a_4848_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X47 a_244_68# B1 a_1972_93# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__oai222_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2
X0 a_255_603# A1 a_67_603# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X1 Z a_67_603# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VDD A2 a_255_603# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X3 VSS A2 a_67_603# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 Z a_67_603# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_67_603# A1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 VDD VSS Z A1 A2
X0 Z a_56_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_56_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS A2 a_56_472# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 Z a_56_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_56_472# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_244_472# A1 a_56_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD a_56_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 VDD VSS Z A1 A2
X0 a_682_472# A1 a_244_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS A2 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X2 VSS A1 a_244_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X3 Z a_244_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 Z a_244_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_244_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_244_68# A1 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VSS a_244_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_244_68# A2 VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_244_68# A1 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VSS a_244_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_244_472# A2 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 VDD a_244_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VDD a_244_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD A2 a_682_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 Z a_244_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A3 VDD VSS Z A1 A2
X0 VSS A3 a_36_88# VSUBS nmos_6p0 w=0.4u l=0.6u
X1 VDD A3 a_448_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 Z a_36_88# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_224_604# A1 a_36_88# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X4 a_36_88# A2 VSS VSUBS nmos_6p0 w=0.4u l=0.6u
X5 Z a_36_88# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS A1 a_36_88# VSUBS nmos_6p0 w=0.4u l=0.6u
X7 a_448_604# A2 a_224_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A3 VDD VSS Z A1 A2
X0 VDD a_36_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_36_68# A2 VSS VSUBS nmos_6p0 w=0.665u l=0.6u
X2 VDD A3 a_448_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS A3 a_36_68# VSUBS nmos_6p0 w=0.665u l=0.6u
X4 Z a_36_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VSS A1 a_36_68# VSUBS nmos_6p0 w=0.665u l=0.6u
X6 VSS a_36_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_244_472# A1 a_36_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_448_472# A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 Z a_36_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A3 VDD VSS Z A1 A2
X0 Z a_244_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_244_68# A1 a_458_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VDD a_244_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS A1 a_244_68# VSUBS nmos_6p0 w=0.665u l=0.6u
X4 VSS a_244_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS A2 a_244_68# VSUBS nmos_6p0 w=0.665u l=0.6u
X6 a_244_68# A2 VSS VSUBS nmos_6p0 w=0.665u l=0.6u
X7 VSS a_244_68# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X8 Z a_244_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_244_68# A1 VSS VSUBS nmos_6p0 w=0.665u l=0.6u
X10 VDD A3 a_1120_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 Z a_244_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 Z a_244_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_244_68# A3 VSS VSUBS nmos_6p0 w=0.665u l=0.6u
X14 a_458_472# A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_244_472# A3 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_1120_472# A2 a_906_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X17 VDD a_244_68# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VSS A3 a_244_68# VSUBS nmos_6p0 w=0.665u l=0.6u
X19 a_906_472# A1 a_244_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or3_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A3 A4 VDD VSS Z A1 A2
X0 a_56_604# A3 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X1 a_708_604# A3 a_484_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 a_484_604# A2 a_244_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X3 VSS A4 a_56_604# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 Z a_56_604# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 Z a_56_604# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VSS A2 a_56_604# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 VDD A4 a_708_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X8 a_244_604# A1 a_56_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X9 a_56_604# A1 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A3 A4 VDD VSS Z A2
X0 a_56_472# A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X1 a_56_472# A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X2 a_468_472# A2 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 Z a_56_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_244_472# A1 a_56_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VDD A4 a_692_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD a_56_472# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VSS A4 a_56_472# VSUBS nmos_6p0 w=0.465u l=0.6u
X8 VSS a_56_472# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_692_472# A3 a_468_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VSS A2 a_56_472# VSUBS nmos_6p0 w=0.465u l=0.6u
X11 Z a_56_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A3 A4 VDD VSS Z A1 A2
X0 a_682_472# A2 a_458_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_244_72# A2 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X2 a_244_72# A4 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 Z a_244_72# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VSS a_244_72# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_244_72# A3 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X6 VSS a_244_72# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X7 Z a_244_72# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_458_472# A3 a_244_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 VDD a_244_72# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VSS A4 a_244_72# VSUBS nmos_6p0 w=0.465u l=0.6u
X11 Z a_244_72# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 VSS A2 a_244_72# VSUBS nmos_6p0 w=0.465u l=0.6u
X13 VDD A4 a_1578_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_244_472# A4 VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_244_72# A1 a_682_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 VSS A1 a_244_72# VSUBS nmos_6p0 w=0.465u l=0.6u
X17 a_1578_472# A3 a_1364_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VDD a_244_72# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 VSS A3 a_244_72# VSUBS nmos_6p0 w=0.465u l=0.6u
X20 a_1120_472# A1 a_244_72# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_244_72# A1 VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X22 a_1364_472# A2 a_1120_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 Z a_244_72# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__or4_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 Q SE SI VDD VSS CLK D
X0 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 VDD D a_800_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 a_1288_135# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 VSS a_3312_458# a_3284_158# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 a_2132_502# a_1288_135# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 Q a_3312_458# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X6 a_1288_135# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X7 a_3284_158# a_1288_135# a_3050_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_2346_502# a_1288_135# a_2132_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 a_2424_386# a_2132_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X10 Q a_3312_458# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X11 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_1751_139# a_1288_135# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X13 a_1751_139# a_1288_135# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X14 a_2132_502# a_1751_139# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X15 a_3264_502# a_1751_139# a_3050_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X16 VSS a_2424_386# a_2387_158# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_2424_386# a_2132_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.51u
X21 a_2387_158# a_1751_139# a_2132_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 VSS D a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 VDD a_3312_458# a_3264_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X24 a_3312_458# a_3050_502# VSS VSUBS nmos_6p0 w=0.435u l=0.6u
X25 VDD a_2424_386# a_2346_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X26 a_3312_458# a_3050_502# VDD w_n86_352# pmos_6p0 w=0.705u l=0.5u
X27 a_3050_502# a_1751_139# a_2424_386# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 a_3050_502# a_1288_135# a_2424_386# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X29 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X30 a_800_502# SE a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X31 a_860_156# a_36_156# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_2 Q SE SI VDD VSS CLK D
X0 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 VDD D a_800_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 a_1288_135# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 VDD a_3404_428# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X4 VSS a_3404_428# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X5 a_2132_502# a_1288_135# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 Q a_3404_428# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X7 a_1288_135# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X8 a_3050_502# a_1751_139# a_2424_386# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2346_502# a_1288_135# a_2132_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 VDD a_3404_428# a_3264_502# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X11 Q a_3404_428# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 a_1751_139# a_1288_135# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X14 a_1751_139# a_1288_135# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X15 a_2132_502# a_1751_139# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X16 a_3264_502# a_1751_139# a_3050_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X17 VSS a_2424_386# a_2387_158# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_3280_158# a_1288_135# a_3050_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_3404_428# a_3050_502# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X22 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 a_2424_386# a_2132_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.51u
X24 a_3404_428# a_3050_502# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X25 a_2387_158# a_1751_139# a_2132_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 VSS D a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 VSS a_3404_428# a_3280_158# VSUBS nmos_6p0 w=0.815u l=0.6u
X28 VDD a_2424_386# a_2346_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X29 a_3050_502# a_1288_135# a_2424_386# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X30 a_2424_386# a_2132_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X31 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X32 a_800_502# SE a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X33 a_860_156# a_36_156# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_4 Q SE SI VDD CLK D VSS
X0 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X1 VSS a_3404_428# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X2 VDD D a_800_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X3 a_1288_135# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 VDD a_3404_428# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X5 VSS a_3404_428# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X6 a_2132_502# a_1288_135# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 Q a_3404_428# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X8 VDD a_3404_428# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X9 a_1288_135# CLK VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X10 a_3050_502# a_1751_139# a_2424_386# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 Q a_3404_428# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 a_2346_502# a_1288_135# a_2132_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 VDD a_3404_428# a_3264_502# w_n86_352# pmos_6p0 w=1.215u l=0.5u
X14 Q a_3404_428# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X15 Q a_3404_428# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X16 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1751_139# a_1288_135# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X18 a_1751_139# a_1288_135# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X19 a_2132_502# a_1751_139# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_3264_502# a_1751_139# a_3050_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X21 VSS a_2424_386# a_2387_158# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_3280_158# a_1288_135# a_3050_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X24 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_3404_428# a_3050_502# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X26 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X27 a_2424_386# a_2132_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.51u
X28 a_3404_428# a_3050_502# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X29 a_2387_158# a_1751_139# a_2132_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X30 VSS D a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X31 VSS a_3404_428# a_3280_158# VSUBS nmos_6p0 w=0.815u l=0.6u
X32 VDD a_2424_386# a_2346_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X33 a_3050_502# a_1288_135# a_2424_386# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 a_2424_386# a_2132_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X35 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X36 a_800_502# SE a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X37 a_860_156# a_36_156# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 Q RN SE SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 a_3572_185# a_1748_497# a_3348_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_2572_124# a_2452_80# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VDD a_3690_141# a_3572_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X7 Q a_3690_141# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X8 a_2452_80# a_2154_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2358_502# RN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 a_2404_124# a_1748_497# a_2154_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_3572_185# a_1285_502# a_3348_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_2154_502# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 VSS a_3690_141# a_3572_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X16 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2358_502# a_1285_502# a_2154_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 a_4122_160# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X19 VDD a_2452_80# a_2358_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X21 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 a_2154_502# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X24 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X25 a_2452_80# a_2154_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X26 a_3348_185# a_1748_497# a_2452_80# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 a_3690_141# RN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X28 Q a_3690_141# VSS VSUBS nmos_6p0 w=0.81u l=0.6u
X29 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X30 a_3348_185# a_1285_502# a_2452_80# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X31 a_3690_141# a_3348_185# a_4122_160# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 VDD a_3348_185# a_3690_141# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X33 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X35 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 Q RN SE SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 a_3572_185# a_1748_497# a_3348_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_2572_124# a_2452_80# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_4122_124# RN VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X7 VSS a_3690_141# Q VSUBS nmos_6p0 w=0.81u l=0.6u
X8 VDD a_3690_141# a_3572_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 VDD a_3690_141# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X10 a_2452_80# a_2154_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_2358_502# RN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X12 Q a_3690_141# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X13 a_2404_124# a_1748_497# a_2154_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_3572_185# a_1285_502# a_3348_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_2154_502# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X16 VSS a_3690_141# a_3572_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 Q a_3690_141# VSS VSUBS nmos_6p0 w=0.81u l=0.6u
X18 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X20 a_3690_141# a_3348_185# a_4122_124# VSUBS nmos_6p0 w=0.54u l=0.6u
X21 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_2358_502# a_1285_502# a_2154_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 VDD a_2452_80# a_2358_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X24 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X25 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X27 a_2154_502# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X29 a_2452_80# a_2154_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X30 a_3348_185# a_1748_497# a_2452_80# VSUBS nmos_6p0 w=0.36u l=0.6u
X31 a_3690_141# RN VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X32 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X33 a_3348_185# a_1285_502# a_2452_80# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 VDD a_3348_185# a_3690_141# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X35 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X36 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X37 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 Q RN SE SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 a_3572_185# a_1748_497# a_3348_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X2 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_2572_124# a_2452_80# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_4122_124# RN VSS VSUBS nmos_6p0 w=0.54u l=0.6u
X7 VSS a_3690_141# Q VSUBS nmos_6p0 w=0.81u l=0.6u
X8 VDD a_3690_141# a_3572_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 VDD a_3690_141# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X10 a_2452_80# a_2154_502# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VSS a_3690_141# Q VSUBS nmos_6p0 w=0.81u l=0.6u
X12 a_2358_502# RN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X13 Q a_3690_141# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X14 a_2404_124# a_1748_497# a_2154_502# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 VDD a_3690_141# Q w_n86_352# pmos_6p0 w=1.215u l=0.5u
X16 a_3572_185# a_1285_502# a_3348_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2154_502# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X18 VSS a_3690_141# a_3572_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X19 Q a_3690_141# VSS VSUBS nmos_6p0 w=0.81u l=0.6u
X20 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X22 a_3690_141# a_3348_185# a_4122_124# VSUBS nmos_6p0 w=0.54u l=0.6u
X23 Q a_3690_141# VDD w_n86_352# pmos_6p0 w=1.215u l=0.5u
X24 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_2358_502# a_1285_502# a_2154_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X26 VDD a_2452_80# a_2358_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X27 Q a_3690_141# VSS VSUBS nmos_6p0 w=0.81u l=0.6u
X28 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X29 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X30 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X31 a_2154_502# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X33 a_2452_80# a_2154_502# VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 a_3348_185# a_1748_497# a_2452_80# VSUBS nmos_6p0 w=0.36u l=0.6u
X35 a_3690_141# RN VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X36 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X37 a_3348_185# a_1285_502# a_2452_80# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X38 VDD a_3348_185# a_3690_141# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X39 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X40 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X41 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 Q RN SE SETN SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_4186_156# SETN a_3696_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_2572_124# a_2440_430# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_3696_185# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X7 VDD a_4234_112# a_3696_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X8 a_3696_185# a_1285_502# a_3471_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2404_124# a_1748_497# a_2096_497# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 VDD a_3471_185# a_4234_112# w_n86_352# pmos_6p0 w=0.92u l=0.5u
X11 a_3079_185# a_2096_497# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X12 Q a_4234_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X15 a_4578_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2336_474# a_1285_502# a_2096_497# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X17 a_3471_185# a_1748_497# a_2440_430# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_2096_497# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X19 VDD a_2440_430# a_2336_474# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X20 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X21 a_2440_430# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X22 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X23 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X24 a_2336_474# RN VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X25 a_2096_497# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X27 a_3471_185# a_1285_502# a_2440_430# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X28 a_3696_185# a_1748_497# a_3471_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X29 a_4234_112# RN VDD w_n86_352# pmos_6p0 w=0.92u l=0.5u
X30 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X31 VSS a_4234_112# a_4186_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 a_4234_112# a_3471_185# a_4578_156# VSUBS nmos_6p0 w=0.465u l=0.6u
X33 Q a_4234_112# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 VDD a_2096_497# a_2440_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X35 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X36 a_2440_430# SETN a_3079_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X37 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X38 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X39 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 Q RN SE SETN SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_4186_156# SETN a_3696_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_4234_112# a_3471_185# a_4578_156# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VSS a_4234_112# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD a_4234_112# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X8 a_2572_124# a_2440_430# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_3696_185# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 VDD a_4234_112# a_3696_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X11 a_3696_185# a_1285_502# a_3471_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_2404_124# a_1748_497# a_2096_497# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 a_3079_185# a_2096_497# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VDD a_3471_185# a_4234_112# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X17 a_4578_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_2336_474# a_1285_502# a_2096_497# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X19 a_3471_185# a_1748_497# a_2440_430# VSUBS nmos_6p0 w=0.36u l=0.6u
X20 a_2096_497# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X21 VDD a_2440_430# a_2336_474# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X22 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 a_2440_430# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X24 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X26 a_2336_474# RN VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X27 a_2096_497# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X29 a_3471_185# a_1285_502# a_2440_430# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X30 a_3696_185# a_1748_497# a_3471_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X31 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 VSS a_4234_112# a_4186_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X33 Q a_4234_112# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X34 VDD a_2096_497# a_2440_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X35 a_4234_112# RN VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X36 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X37 a_2440_430# SETN a_3079_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X38 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X39 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X40 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X41 Q a_4234_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 Q RN SE SETN SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 a_4186_156# SETN a_3696_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X5 a_4234_112# a_3471_185# a_4578_156# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 VSS a_4234_112# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_2572_124# a_2440_430# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_3696_185# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X9 VDD a_4234_112# a_3696_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X10 a_3696_185# a_1285_502# a_3471_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 Q a_4234_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_2404_124# a_1748_497# a_2096_497# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 VDD a_4234_112# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 a_3079_185# a_2096_497# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X15 VDD a_3471_185# a_4234_112# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X18 a_4578_156# RN VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_2336_474# a_1285_502# a_2096_497# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X20 Q a_4234_112# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_3471_185# a_1748_497# a_2440_430# VSUBS nmos_6p0 w=0.36u l=0.6u
X22 VSS a_4234_112# Q VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_2096_497# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X24 VDD a_2440_430# a_2336_474# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X25 VDD a_4234_112# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X26 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X27 a_2440_430# SETN VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X28 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X29 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X30 a_2336_474# RN VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X31 a_2096_497# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X33 a_3471_185# a_1285_502# a_2440_430# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 Q a_4234_112# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X35 a_3696_185# a_1748_497# a_3471_185# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X36 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X37 VSS a_4234_112# a_4186_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X38 Q a_4234_112# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X39 VDD a_2096_497# a_2440_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X40 a_4234_112# RN VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X41 VSS RN a_2572_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X42 a_2440_430# SETN a_3079_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X43 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X44 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X45 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 Q SE SETN SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X4 VDD a_2476_430# a_2336_474# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X5 a_3300_185# a_1748_497# a_2476_430# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 Q a_4110_62# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X7 VDD a_4110_62# a_3524_185# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X8 a_2404_124# a_1748_497# a_2096_497# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_4110_62# a_3300_185# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X10 a_3524_185# SETN VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X11 VSS a_2476_430# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 Q a_4110_62# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X15 a_2336_474# a_1285_502# a_2096_497# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X16 VSS a_4110_62# a_4005_106# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2096_497# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X18 VDD SETN a_2476_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X19 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X20 a_3300_185# a_1285_502# a_2476_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X21 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 a_3524_185# a_1748_497# a_3300_185# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X24 a_2096_497# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X25 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X26 a_4005_106# SETN a_3524_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X27 a_2476_430# a_2096_497# VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X28 a_2476_430# SETN a_2908_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X29 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X30 a_4110_62# a_3300_185# VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X31 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X32 a_3524_185# a_1285_502# a_3300_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X33 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X34 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X35 a_2908_185# a_2096_497# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 Q SE SETN SI VDD VSS CLK D
X0 a_1748_497# a_1285_502# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1285_502# CLK VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X3 VDD SE a_840_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X4 VDD a_2476_430# a_2336_474# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X5 VDD a_4110_62# a_3524_185# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X6 a_3300_185# a_1748_497# a_2476_430# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_3524_185# SETN VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X8 a_2404_124# a_1748_497# a_2096_497# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 VSS a_2476_430# a_2404_124# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 Q a_4110_62# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_1748_497# a_1285_502# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X13 a_4110_62# a_3300_185# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X14 a_2336_474# a_1285_502# a_2096_497# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X15 VSS a_4110_62# a_4005_106# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_2096_497# a_1748_497# a_596_502# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X17 VDD SETN a_2476_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X18 a_448_502# SI VDD w_n86_352# pmos_6p0 w=0.63u l=0.5u
X19 a_3300_185# a_1285_502# a_2476_430# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X20 a_468_156# SI VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 VDD a_4110_62# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 a_596_502# a_36_156# a_448_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X23 a_3524_185# a_1748_497# a_3300_185# w_n86_352# pmos_6p0 w=0.625u l=0.5u
X24 VSS a_4110_62# Q VSUBS nmos_6p0 w=0.82u l=0.64u
X25 a_2096_497# a_1285_502# a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X26 a_1285_502# CLK VDD w_n86_352# pmos_6p0 w=0.925u l=0.5u
X27 a_4005_106# SETN a_3524_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 a_2476_430# a_2096_497# VDD w_n86_352# pmos_6p0 w=0.625u l=0.5u
X29 a_4110_62# a_3300_185# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X30 a_2476_430# SETN a_2908_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X31 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X32 a_840_502# D a_596_502# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X33 a_3524_185# a_1285_502# a_3300_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X34 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.63u l=0.5u
X35 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.36u l=0.6u
X36 Q a_4110_62# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X37 a_2908_185# a_2096_497# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 D Q SE SETN SI VDD VSS CLK
X0 a_3636_185# a_1850_497# a_3412_185# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X1 VSS SE a_36_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X2 a_2288_518# a_1300_144# a_636_156# VSUBS nmos_6p0 w=0.475u l=0.6u
X3 VSS a_4197_114# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X4 a_1850_497# a_1300_144# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X5 Q a_4197_114# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X6 VDD a_2540_426# a_2492_518# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 a_4197_114# a_3412_185# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X8 VSS CLK a_1300_144# VSUBS nmos_6p0 w=0.465u l=0.6u
X9 a_3636_185# SETN VDD w_n86_352# pmos_6p0 w=0.47u l=0.5u
X10 a_4149_158# SETN a_3636_185# VSUBS nmos_6p0 w=0.37u l=0.6u
X11 Q a_4197_114# VSS VSUBS nmos_6p0 w=0.815u l=0.6u
X12 VDD a_4197_114# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_2540_426# SETN a_3020_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VDD a_4197_114# a_3636_185# w_n86_352# pmos_6p0 w=0.47u l=0.5u
X15 a_448_556# SI VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X16 VSS a_2540_426# a_2552_124# VSUBS nmos_6p0 w=0.475u l=0.6u
X17 a_636_156# SE a_468_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X18 a_596_556# a_36_156# a_448_556# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X19 a_1850_497# a_1300_144# VSS VSUBS nmos_6p0 w=0.465u l=0.6u
X20 a_2552_124# a_1850_497# a_2288_518# VSUBS nmos_6p0 w=0.475u l=0.6u
X21 a_468_156# SI VSS VSUBS nmos_6p0 w=0.38u l=0.6u
X22 a_4197_114# a_3412_185# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 Q a_4197_114# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X24 VDD a_4197_114# Q w_n86_352# pmos_6p0 w=1.22u l=0.5u
X25 a_2288_518# a_1850_497# a_596_556# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X26 a_840_556# D a_596_556# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X27 a_3636_185# a_1300_144# a_3412_185# VSUBS nmos_6p0 w=0.36u l=0.6u
X28 VDD SE a_36_156# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X29 VDD CLK a_1300_144# w_n86_352# pmos_6p0 w=0.815u l=0.5u
X30 a_2492_518# a_1300_144# a_2288_518# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X31 VDD a_3412_185# a_4197_114# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X32 VSS a_4197_114# a_4149_158# VSUBS nmos_6p0 w=0.37u l=0.6u
X33 VDD SETN a_2540_426# w_n86_352# pmos_6p0 w=0.815u l=0.5u
X34 VSS a_36_156# a_860_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X35 VSS a_3412_185# a_4197_114# VSUBS nmos_6p0 w=0.815u l=0.6u
X36 VDD SE a_840_556# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X37 a_3412_185# a_1850_497# a_2540_426# VSUBS nmos_6p0 w=0.36u l=0.6u
X38 Q a_4197_114# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X39 a_3412_185# a_1300_144# a_2540_426# w_n86_352# pmos_6p0 w=0.415u l=0.5u
X40 a_2540_426# a_2288_518# VDD w_n86_352# pmos_6p0 w=0.815u l=0.5u
X41 VSS a_4197_114# Q VSUBS nmos_6p0 w=0.815u l=0.6u
X42 a_860_156# D a_636_156# VSUBS nmos_6p0 w=0.38u l=0.6u
X43 a_3020_185# a_2288_518# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__tieh.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
X0 Z a_125_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_125_24# a_125_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__tieh.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__tiel.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
X0 ZN a_124_24# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X1 a_124_24# a_124_24# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__tiel.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 VDD VSS ZN A1 A2
X0 a_716_68# A2 ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VDD A1 a_64_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X2 a_930_497# A1 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 ZN a_64_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X4 a_272_93# A2 a_64_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VSS A1 a_272_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_716_68# a_64_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 VDD A2 a_930_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 ZN A1 a_716_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 a_64_93# A2 VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 VDD VSS ZN A1 A2
X0 VSS a_728_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 ZN a_728_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 a_728_472# a_56_565# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 ZN a_728_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_728_68# A1 a_728_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 VDD A1 a_244_565# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X6 VSS A1 a_56_565# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_244_565# A2 a_56_565# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X8 a_728_472# A2 a_728_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_728_68# a_56_565# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VSS A2 a_952_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_56_565# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X12 a_952_68# A1 a_728_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X13 VDD a_728_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 VDD VSS ZN A1 A2
X0 VSS a_728_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VSS a_728_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X2 ZN a_728_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 ZN a_728_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 ZN a_728_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_728_68# A1 a_708_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 VDD A1 a_234_472# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 VSS A1 a_46_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_708_472# A2 a_728_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_728_68# a_46_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X10 VDD a_728_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X11 VSS A2 a_952_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN a_728_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 a_46_472# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_708_472# a_46_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X15 VDD a_728_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_234_472# A2 a_46_472# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X17 a_952_68# A1 a_728_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A3 VDD VSS ZN A1 A2
X0 a_1296_93# a_728_93# VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X1 a_728_93# a_56_567# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X2 VDD A3 a_1296_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X3 VDD A1 a_244_567# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X4 VSS A2 a_952_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 a_952_93# A1 a_728_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_244_567# A2 a_56_567# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X7 a_728_93# A1 a_718_527# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X8 ZN A3 a_1948_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X9 ZN a_1296_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 VDD a_728_93# a_2172_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 a_718_527# a_56_567# VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X12 a_718_527# A2 a_728_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X13 VSS A1 a_56_567# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VSS A3 a_1504_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X15 a_1948_68# a_728_93# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X16 a_2172_497# A3 ZN w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_1504_93# a_728_93# a_1296_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X18 a_56_567# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X19 a_1948_68# a_1296_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A3 VDD VSS ZN A1 A2
X0 a_728_93# A1 a_728_526# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X1 ZN a_2004_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_728_93# a_56_561# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_2004_68# a_1347_526# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS A2 a_952_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 a_1347_526# a_728_93# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X6 a_728_526# A2 a_728_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X7 a_244_561# A2 a_56_561# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X8 a_952_93# A1 a_728_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X9 a_2004_472# a_1347_526# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X10 VSS A1 a_56_561# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 VSS a_728_93# a_2228_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X12 ZN a_2004_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS a_2004_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A3 a_1535_526# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X15 a_2004_68# A3 a_2004_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_1535_526# a_728_93# a_1347_526# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X17 a_56_561# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 VDD A1 a_244_561# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X19 VSS A3 a_1347_526# VSUBS nmos_6p0 w=0.36u l=0.6u
X20 a_728_526# a_56_561# VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X21 a_2004_472# a_728_93# a_2004_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X22 VDD a_2004_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X23 a_2228_68# A3 a_2004_68# VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_4 A3 VDD VSS ZN A1 A2
X0 ZN a_1979_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_692_527# A2 a_692_93# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X2 VDD a_1979_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 a_1379_527# a_692_93# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X4 ZN a_1979_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 a_1979_68# a_1379_527# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X6 ZN a_1979_68# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_916_93# A1 a_692_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_244_532# A2 a_56_532# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 VSS A1 a_56_532# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 VSS A3 a_1379_527# VSUBS nmos_6p0 w=0.36u l=0.6u
X11 a_1979_68# A3 a_1979_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 ZN a_1979_68# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS a_1979_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X14 VDD A1 a_244_532# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_1979_472# a_692_93# a_1979_68# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X16 a_692_527# a_56_532# VDD w_n86_352# pmos_6p0 w=0.385u l=0.5u
X17 VDD a_1979_68# ZN w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 a_1979_472# a_1379_527# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_1567_527# a_692_93# a_1379_527# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X20 a_692_93# a_56_532# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X21 VSS a_1979_68# ZN VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_692_93# A1 a_692_527# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X23 a_56_532# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X24 VSS a_692_93# a_2203_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X25 VDD A3 a_1567_527# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X26 a_2203_68# A3 a_1979_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X27 VSS A2 a_916_93# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xnor3_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 VDD VSS Z A1 A2
X0 a_728_472# a_56_604# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 Z A1 a_728_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X2 VSS A1 a_56_604# VSUBS nmos_6p0 w=0.36u l=0.6u
X3 a_728_472# A2 Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 Z a_56_604# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X5 VSS A2 a_952_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_244_604# A2 a_56_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X7 a_56_604# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X8 a_952_68# A1 Z VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD A1 a_244_604# w_n86_352# pmos_6p0 w=0.56u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 VDD VSS Z A1 A2
X0 a_730_68# A2 a_730_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X1 VDD A2 a_954_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_730_68# a_78_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X3 VSS a_730_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X4 a_954_497# A1 a_730_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_286_93# A2 a_78_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 Z a_730_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X7 a_730_497# a_78_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X8 Z a_730_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_78_93# A2 VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X10 a_730_497# A1 a_730_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 VDD A1 a_78_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X12 VDD a_730_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X13 VSS A1 a_286_93# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 VDD VSS Z A1 A2
X0 VDD a_721_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 VSS a_721_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X2 a_721_497# a_69_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X3 Z a_721_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X4 VDD a_721_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X5 a_277_93# A2 a_69_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VSS a_721_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X7 Z a_721_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X8 Z a_721_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X9 VDD A2 a_945_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X10 a_721_497# A1 a_721_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X11 Z a_721_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X12 a_945_497# A1 a_721_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X13 VSS A1 a_277_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X14 a_69_93# A2 VDD w_n86_352# pmos_6p0 w=0.385u l=0.5u
X15 a_721_68# A2 a_721_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X16 VDD A1 a_69_93# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X17 a_721_68# a_69_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor2_4.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_1.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2
X0 Z A3 a_1936_472# w_n86_352# pmos_6p0 w=1.22u l=0.5u
X1 a_728_93# a_56_524# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X2 a_1936_472# a_728_93# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X3 VSS A2 a_952_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X4 VDD A3 a_1524_472# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X5 a_1936_472# a_1336_472# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X6 a_952_93# A1 a_728_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_728_93# A1 a_718_524# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X8 a_1524_472# a_728_93# a_1336_472# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X9 a_244_524# A2 a_56_524# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X10 a_718_524# a_56_524# VDD w_n86_352# pmos_6p0 w=0.565u l=0.5u
X11 a_718_524# A2 a_728_93# w_n86_352# pmos_6p0 w=0.565u l=0.5u
X12 VSS A1 a_56_524# VSUBS nmos_6p0 w=0.36u l=0.6u
X13 a_1336_472# a_728_93# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X14 VDD A1 a_244_524# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_56_524# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X16 VSS A3 a_1336_472# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 a_2215_68# A3 Z VSUBS nmos_6p0 w=0.82u l=0.6u
X18 VSS a_728_93# a_2215_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X19 Z a_1336_472# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_1.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_2.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A3 VDD VSS Z A1 A2
X0 a_725_93# A1 a_731_494# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X1 a_725_93# a_89_534# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X2 VSS a_1943_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X3 a_731_494# A2 a_725_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X4 VDD a_725_93# a_2153_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X5 a_89_534# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X6 VSS A2 a_949_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_1943_497# A3 a_1949_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 Z a_1943_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X9 a_1297_93# a_725_93# VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X10 a_2153_497# A3 a_1943_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X11 VSS A1 a_89_534# VSUBS nmos_6p0 w=0.36u l=0.6u
X12 VDD A3 a_1297_93# w_n86_352# pmos_6p0 w=0.56u l=0.5u
X13 a_1943_497# a_1297_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X14 a_1949_68# a_725_93# a_1943_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X15 VSS A3 a_1505_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X16 a_1505_93# a_725_93# a_1297_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X17 VDD a_1943_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X18 VDD A1 a_277_534# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X19 a_1949_68# a_1297_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X20 a_949_93# A1 a_725_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X21 Z a_1943_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X22 a_731_494# a_89_534# VDD w_n86_352# pmos_6p0 w=0.56u l=0.5u
X23 a_277_534# A2 a_89_534# w_n86_352# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_2.ext - technology: gf180mcuB



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_4.ext - technology: gf180mcuB

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_4 A3 VDD VSS Z A1 A2
X0 a_1912_497# a_1260_93# VDD w_n86_352# pmos_6p0 w=1.095u l=0.5u
X1 VDD a_692_93# a_2126_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X2 a_692_519# A2 a_692_93# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X3 Z a_1912_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X4 VSS A3 a_1468_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X5 VSS a_1912_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X6 a_916_93# A1 a_692_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X7 a_1912_497# A3 a_1912_68# VSUBS nmos_6p0 w=0.82u l=0.6u
X8 a_244_524# A2 a_56_524# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X9 VSS A1 a_56_524# VSUBS nmos_6p0 w=0.36u l=0.6u
X10 VSS a_1912_497# Z VSUBS nmos_6p0 w=0.82u l=0.6u
X11 a_1912_68# a_1260_93# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X12 Z a_1912_497# VSS VSUBS nmos_6p0 w=0.82u l=0.6u
X13 Z a_1912_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X14 VDD A1 a_244_524# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X15 a_692_519# a_56_524# VDD w_n86_352# pmos_6p0 w=0.385u l=0.5u
X16 a_2126_497# A3 a_1912_497# w_n86_352# pmos_6p0 w=1.095u l=0.5u
X17 a_692_93# a_56_524# VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X18 VDD a_1912_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X19 a_692_93# A1 a_692_519# w_n86_352# pmos_6p0 w=0.385u l=0.5u
X20 Z a_1912_497# VDD w_n86_352# pmos_6p0 w=1.22u l=0.5u
X21 a_56_524# A2 VSS VSUBS nmos_6p0 w=0.36u l=0.6u
X22 a_1912_68# a_692_93# a_1912_497# VSUBS nmos_6p0 w=0.82u l=0.6u
X23 a_1468_93# a_692_93# a_1260_93# VSUBS nmos_6p0 w=0.36u l=0.6u
X24 a_1260_93# a_692_93# VDD w_n86_352# pmos_6p0 w=0.36u l=0.5u
X25 VDD A3 a_1260_93# w_n86_352# pmos_6p0 w=0.36u l=0.5u
X26 VDD a_1912_497# Z w_n86_352# pmos_6p0 w=1.22u l=0.5u
X27 VSS A2 a_916_93# VSUBS nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu7t5v0__xor3_4.ext - technology: gf180mcuB



******* EOF

