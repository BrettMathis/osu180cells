magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 552 1254
<< mvpmos >>
rect 0 0 120 1134
rect 224 0 344 1134
<< mvpdiff >>
rect -88 1121 0 1134
rect -88 1075 -75 1121
rect -29 1075 0 1121
rect -88 1015 0 1075
rect -88 969 -75 1015
rect -29 969 0 1015
rect -88 909 0 969
rect -88 863 -75 909
rect -29 863 0 909
rect -88 803 0 863
rect -88 757 -75 803
rect -29 757 0 803
rect -88 697 0 757
rect -88 651 -75 697
rect -29 651 0 697
rect -88 591 0 651
rect -88 545 -75 591
rect -29 545 0 591
rect -88 485 0 545
rect -88 439 -75 485
rect -29 439 0 485
rect -88 379 0 439
rect -88 333 -75 379
rect -29 333 0 379
rect -88 273 0 333
rect -88 227 -75 273
rect -29 227 0 273
rect -88 166 0 227
rect -88 120 -75 166
rect -29 120 0 166
rect -88 59 0 120
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1121 224 1134
rect 120 1075 149 1121
rect 195 1075 224 1121
rect 120 1015 224 1075
rect 120 969 149 1015
rect 195 969 224 1015
rect 120 909 224 969
rect 120 863 149 909
rect 195 863 224 909
rect 120 803 224 863
rect 120 757 149 803
rect 195 757 224 803
rect 120 697 224 757
rect 120 651 149 697
rect 195 651 224 697
rect 120 591 224 651
rect 120 545 149 591
rect 195 545 224 591
rect 120 485 224 545
rect 120 439 149 485
rect 195 439 224 485
rect 120 379 224 439
rect 120 333 149 379
rect 195 333 224 379
rect 120 273 224 333
rect 120 227 149 273
rect 195 227 224 273
rect 120 166 224 227
rect 120 120 149 166
rect 195 120 224 166
rect 120 59 224 120
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 1121 432 1134
rect 344 1075 373 1121
rect 419 1075 432 1121
rect 344 1015 432 1075
rect 344 969 373 1015
rect 419 969 432 1015
rect 344 909 432 969
rect 344 863 373 909
rect 419 863 432 909
rect 344 803 432 863
rect 344 757 373 803
rect 419 757 432 803
rect 344 697 432 757
rect 344 651 373 697
rect 419 651 432 697
rect 344 591 432 651
rect 344 545 373 591
rect 419 545 432 591
rect 344 485 432 545
rect 344 439 373 485
rect 419 439 432 485
rect 344 379 432 439
rect 344 333 373 379
rect 419 333 432 379
rect 344 273 432 333
rect 344 227 373 273
rect 419 227 432 273
rect 344 166 432 227
rect 344 120 373 166
rect 419 120 432 166
rect 344 59 432 120
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 1075 -29 1121
rect -75 969 -29 1015
rect -75 863 -29 909
rect -75 757 -29 803
rect -75 651 -29 697
rect -75 545 -29 591
rect -75 439 -29 485
rect -75 333 -29 379
rect -75 227 -29 273
rect -75 120 -29 166
rect -75 13 -29 59
rect 149 1075 195 1121
rect 149 969 195 1015
rect 149 863 195 909
rect 149 757 195 803
rect 149 651 195 697
rect 149 545 195 591
rect 149 439 195 485
rect 149 333 195 379
rect 149 227 195 273
rect 149 120 195 166
rect 149 13 195 59
rect 373 1075 419 1121
rect 373 969 419 1015
rect 373 863 419 909
rect 373 757 419 803
rect 373 651 419 697
rect 373 545 419 591
rect 373 439 419 485
rect 373 333 419 379
rect 373 227 419 273
rect 373 120 419 166
rect 373 13 419 59
<< polysilicon >>
rect 0 1134 120 1178
rect 224 1134 344 1178
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 1121 -29 1134
rect -75 1015 -29 1075
rect -75 909 -29 969
rect -75 803 -29 863
rect -75 697 -29 757
rect -75 591 -29 651
rect -75 485 -29 545
rect -75 379 -29 439
rect -75 273 -29 333
rect -75 166 -29 227
rect -75 59 -29 120
rect -75 0 -29 13
rect 149 1121 195 1134
rect 149 1015 195 1075
rect 149 909 195 969
rect 149 803 195 863
rect 149 697 195 757
rect 149 591 195 651
rect 149 485 195 545
rect 149 379 195 439
rect 149 273 195 333
rect 149 166 195 227
rect 149 59 195 120
rect 149 0 195 13
rect 373 1121 419 1134
rect 373 1015 419 1075
rect 373 909 419 969
rect 373 803 419 863
rect 373 697 419 757
rect 373 591 419 651
rect 373 485 419 545
rect 373 379 419 439
rect 373 273 419 333
rect 373 166 419 227
rect 373 59 419 120
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 567 -52 567 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 567 396 567 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 567 172 567 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 296444
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 292990
<< end >>
