magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 682
<< mvndiff >>
rect -88 669 0 682
rect -88 13 -75 669
rect -29 13 0 669
rect -88 0 0 13
rect 120 669 208 682
rect 120 13 149 669
rect 195 13 208 669
rect 120 0 208 13
<< mvndiffc >>
rect -75 13 -29 669
rect 149 13 195 669
<< polysilicon >>
rect 0 682 120 726
rect 0 -44 120 0
<< metal1 >>
rect -75 669 -29 682
rect -75 0 -29 13
rect 149 669 195 682
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 341 -52 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 341 172 341 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 140028
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 138236
<< end >>
