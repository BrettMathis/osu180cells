magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 3000 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
rect 1550 190 1610 360
rect 1720 190 1780 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2230 190 2290 360
rect 2400 190 2460 360
rect 2570 190 2630 360
rect 2740 190 2800 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
rect 870 1090 930 1430
rect 1040 1090 1100 1430
rect 1210 1090 1270 1430
rect 1380 1090 1440 1430
rect 1550 1090 1610 1430
rect 1720 1090 1780 1430
rect 1890 1090 1950 1430
rect 2060 1090 2120 1430
rect 2230 1090 2290 1430
rect 2400 1090 2460 1430
rect 2570 1090 2630 1430
rect 2740 1090 2800 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 870 360
rect 760 252 792 298
rect 838 252 870 298
rect 760 190 870 252
rect 930 298 1040 360
rect 930 252 962 298
rect 1008 252 1040 298
rect 930 190 1040 252
rect 1100 298 1210 360
rect 1100 252 1132 298
rect 1178 252 1210 298
rect 1100 190 1210 252
rect 1270 298 1380 360
rect 1270 252 1302 298
rect 1348 252 1380 298
rect 1270 190 1380 252
rect 1440 298 1550 360
rect 1440 252 1472 298
rect 1518 252 1550 298
rect 1440 190 1550 252
rect 1610 298 1720 360
rect 1610 252 1642 298
rect 1688 252 1720 298
rect 1610 190 1720 252
rect 1780 298 1890 360
rect 1780 252 1812 298
rect 1858 252 1890 298
rect 1780 190 1890 252
rect 1950 298 2060 360
rect 1950 252 1982 298
rect 2028 252 2060 298
rect 1950 190 2060 252
rect 2120 298 2230 360
rect 2120 252 2152 298
rect 2198 252 2230 298
rect 2120 190 2230 252
rect 2290 298 2400 360
rect 2290 252 2322 298
rect 2368 252 2400 298
rect 2290 190 2400 252
rect 2460 298 2570 360
rect 2460 252 2492 298
rect 2538 252 2570 298
rect 2460 190 2570 252
rect 2630 298 2740 360
rect 2630 252 2662 298
rect 2708 252 2740 298
rect 2630 190 2740 252
rect 2800 298 2900 360
rect 2800 252 2832 298
rect 2878 252 2900 298
rect 2800 190 2900 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 870 1430
rect 760 1143 792 1377
rect 838 1143 870 1377
rect 760 1090 870 1143
rect 930 1377 1040 1430
rect 930 1143 962 1377
rect 1008 1143 1040 1377
rect 930 1090 1040 1143
rect 1100 1377 1210 1430
rect 1100 1143 1132 1377
rect 1178 1143 1210 1377
rect 1100 1090 1210 1143
rect 1270 1377 1380 1430
rect 1270 1143 1302 1377
rect 1348 1143 1380 1377
rect 1270 1090 1380 1143
rect 1440 1377 1550 1430
rect 1440 1143 1472 1377
rect 1518 1143 1550 1377
rect 1440 1090 1550 1143
rect 1610 1377 1720 1430
rect 1610 1143 1642 1377
rect 1688 1143 1720 1377
rect 1610 1090 1720 1143
rect 1780 1377 1890 1430
rect 1780 1143 1812 1377
rect 1858 1143 1890 1377
rect 1780 1090 1890 1143
rect 1950 1377 2060 1430
rect 1950 1143 1982 1377
rect 2028 1143 2060 1377
rect 1950 1090 2060 1143
rect 2120 1377 2230 1430
rect 2120 1143 2152 1377
rect 2198 1143 2230 1377
rect 2120 1090 2230 1143
rect 2290 1377 2400 1430
rect 2290 1143 2322 1377
rect 2368 1143 2400 1377
rect 2290 1090 2400 1143
rect 2460 1377 2570 1430
rect 2460 1143 2492 1377
rect 2538 1143 2570 1377
rect 2460 1090 2570 1143
rect 2630 1377 2740 1430
rect 2630 1143 2662 1377
rect 2708 1143 2740 1377
rect 2630 1090 2740 1143
rect 2800 1377 2900 1430
rect 2800 1143 2832 1377
rect 2878 1143 2900 1377
rect 2800 1090 2900 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
rect 962 252 1008 298
rect 1132 252 1178 298
rect 1302 252 1348 298
rect 1472 252 1518 298
rect 1642 252 1688 298
rect 1812 252 1858 298
rect 1982 252 2028 298
rect 2152 252 2198 298
rect 2322 252 2368 298
rect 2492 252 2538 298
rect 2662 252 2708 298
rect 2832 252 2878 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
rect 962 1143 1008 1377
rect 1132 1143 1178 1377
rect 1302 1143 1348 1377
rect 1472 1143 1518 1377
rect 1642 1143 1688 1377
rect 1812 1143 1858 1377
rect 1982 1143 2028 1377
rect 2152 1143 2198 1377
rect 2322 1143 2368 1377
rect 2492 1143 2538 1377
rect 2662 1143 2708 1377
rect 2832 1143 2878 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
rect 2730 98 2820 120
rect 2730 52 2752 98
rect 2798 52 2820 98
rect 2730 30 2820 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
rect 1290 1568 1380 1590
rect 1290 1522 1312 1568
rect 1358 1522 1380 1568
rect 1290 1500 1380 1522
rect 1530 1568 1620 1590
rect 1530 1522 1552 1568
rect 1598 1522 1620 1568
rect 1530 1500 1620 1522
rect 1770 1568 1860 1590
rect 1770 1522 1792 1568
rect 1838 1522 1860 1568
rect 1770 1500 1860 1522
rect 2010 1568 2100 1590
rect 2010 1522 2032 1568
rect 2078 1522 2100 1568
rect 2010 1500 2100 1522
rect 2250 1568 2340 1590
rect 2250 1522 2272 1568
rect 2318 1522 2340 1568
rect 2250 1500 2340 1522
rect 2490 1568 2580 1590
rect 2490 1522 2512 1568
rect 2558 1522 2580 1568
rect 2490 1500 2580 1522
rect 2730 1568 2820 1590
rect 2730 1522 2752 1568
rect 2798 1522 2820 1568
rect 2730 1500 2820 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
rect 2752 52 2798 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
rect 1552 1522 1598 1568
rect 1792 1522 1838 1568
rect 2032 1522 2078 1568
rect 2272 1522 2318 1568
rect 2512 1522 2558 1568
rect 2752 1522 2798 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 870 1430 930 1480
rect 1040 1430 1100 1480
rect 1210 1430 1270 1480
rect 1380 1430 1440 1480
rect 1550 1430 1610 1480
rect 1720 1430 1780 1480
rect 1890 1430 1950 1480
rect 2060 1430 2120 1480
rect 2230 1430 2290 1480
rect 2400 1430 2460 1480
rect 2570 1430 2630 1480
rect 2740 1430 2800 1480
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 870 1040 930 1090
rect 1040 1040 1100 1090
rect 1210 1040 1270 1090
rect 1380 1040 1440 1090
rect 1550 1040 1610 1090
rect 1720 1040 1780 1090
rect 1890 1040 1950 1090
rect 2060 1040 2120 1090
rect 2230 1040 2290 1090
rect 2400 1040 2460 1090
rect 2570 1040 2630 1090
rect 2740 1040 2800 1090
rect 190 990 2800 1040
rect 190 800 250 990
rect 160 780 250 800
rect 90 758 250 780
rect 90 712 112 758
rect 158 712 250 758
rect 90 690 250 712
rect 160 680 250 690
rect 190 450 250 680
rect 190 400 2800 450
rect 190 360 250 400
rect 360 360 420 400
rect 530 360 590 400
rect 700 360 760 400
rect 870 360 930 400
rect 1040 360 1100 400
rect 1210 360 1270 400
rect 1380 360 1440 400
rect 1550 360 1610 400
rect 1720 360 1780 400
rect 1890 360 1950 400
rect 2060 360 2120 400
rect 2230 360 2290 400
rect 2400 360 2460 400
rect 2570 360 2630 400
rect 2740 360 2800 400
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
rect 1550 140 1610 190
rect 1720 140 1780 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2230 140 2290 190
rect 2400 140 2460 190
rect 2570 140 2630 190
rect 2740 140 2800 190
<< polycontact >>
rect 112 712 158 758
<< metal1 >>
rect 0 1568 3000 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1552 1568
rect 1598 1566 1792 1568
rect 1838 1566 2032 1568
rect 2078 1566 2272 1568
rect 2318 1566 2512 1568
rect 2558 1566 2752 1568
rect 2798 1566 3000 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 1366 1522 1552 1566
rect 1606 1522 1792 1566
rect 1846 1522 2032 1566
rect 2086 1522 2272 1566
rect 2326 1522 2512 1566
rect 2566 1522 2752 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1554 1522
rect 1606 1514 1794 1522
rect 1846 1514 2034 1522
rect 2086 1514 2274 1522
rect 2326 1514 2514 1522
rect 2566 1514 2754 1522
rect 2806 1514 3000 1566
rect 0 1470 3000 1514
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1060 160 1143
rect 280 1377 330 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 940 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1060 500 1143
rect 620 1377 670 1430
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 940 670 1143
rect 790 1377 840 1470
rect 790 1143 792 1377
rect 838 1143 840 1377
rect 790 1060 840 1143
rect 960 1377 1010 1430
rect 960 1143 962 1377
rect 1008 1143 1010 1377
rect 960 940 1010 1143
rect 1130 1377 1180 1470
rect 1130 1143 1132 1377
rect 1178 1143 1180 1377
rect 1130 1060 1180 1143
rect 1300 1377 1350 1430
rect 1300 1143 1302 1377
rect 1348 1143 1350 1377
rect 1300 940 1350 1143
rect 1470 1377 1520 1470
rect 1470 1143 1472 1377
rect 1518 1143 1520 1377
rect 1470 1060 1520 1143
rect 1640 1377 1690 1430
rect 1640 1143 1642 1377
rect 1688 1143 1690 1377
rect 1640 940 1690 1143
rect 1810 1377 1860 1470
rect 1810 1143 1812 1377
rect 1858 1143 1860 1377
rect 1810 1060 1860 1143
rect 1980 1377 2030 1430
rect 1980 1143 1982 1377
rect 2028 1143 2030 1377
rect 1980 940 2030 1143
rect 2150 1377 2200 1470
rect 2150 1143 2152 1377
rect 2198 1143 2200 1377
rect 2150 1060 2200 1143
rect 2320 1377 2370 1430
rect 2320 1143 2322 1377
rect 2368 1143 2370 1377
rect 2320 940 2370 1143
rect 2490 1377 2540 1470
rect 2490 1143 2492 1377
rect 2538 1143 2540 1377
rect 2490 1060 2540 1143
rect 2660 1377 2710 1430
rect 2660 1143 2662 1377
rect 2708 1143 2710 1377
rect 2660 940 2710 1143
rect 2830 1377 2880 1470
rect 2830 1143 2832 1377
rect 2878 1143 2880 1377
rect 2830 1060 2880 1143
rect 280 936 2710 940
rect 280 884 2654 936
rect 2706 884 2710 936
rect 280 860 2710 884
rect 80 758 180 760
rect 80 756 112 758
rect 80 704 104 756
rect 158 712 180 758
rect 156 704 180 712
rect 80 670 180 704
rect 280 460 330 860
rect 620 460 670 860
rect 960 460 1010 860
rect 1300 460 1350 860
rect 1640 460 1690 860
rect 1980 460 2030 860
rect 2320 460 2370 860
rect 2630 840 2710 860
rect 2660 460 2710 840
rect 280 380 2710 460
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 380
rect 280 252 282 298
rect 328 252 330 298
rect 280 160 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 380
rect 620 252 622 298
rect 668 252 670 298
rect 620 160 670 252
rect 790 298 840 360
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 960 298 1010 380
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 160 1010 252
rect 1130 298 1180 360
rect 1130 252 1132 298
rect 1178 252 1180 298
rect 1130 120 1180 252
rect 1300 298 1350 380
rect 1300 252 1302 298
rect 1348 252 1350 298
rect 1300 160 1350 252
rect 1470 298 1520 360
rect 1470 252 1472 298
rect 1518 252 1520 298
rect 1470 120 1520 252
rect 1640 298 1690 380
rect 1640 252 1642 298
rect 1688 252 1690 298
rect 1640 160 1690 252
rect 1810 298 1860 360
rect 1810 252 1812 298
rect 1858 252 1860 298
rect 1810 120 1860 252
rect 1980 298 2030 380
rect 1980 252 1982 298
rect 2028 252 2030 298
rect 1980 160 2030 252
rect 2150 298 2200 360
rect 2150 252 2152 298
rect 2198 252 2200 298
rect 2150 120 2200 252
rect 2320 298 2370 380
rect 2320 252 2322 298
rect 2368 252 2370 298
rect 2320 160 2370 252
rect 2490 298 2540 360
rect 2490 252 2492 298
rect 2538 252 2540 298
rect 2490 120 2540 252
rect 2660 298 2710 380
rect 2660 252 2662 298
rect 2708 252 2710 298
rect 2660 160 2710 252
rect 2830 298 2880 360
rect 2830 252 2832 298
rect 2878 252 2880 298
rect 2830 120 2880 252
rect 0 106 3000 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 2566 98 2754 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2752 98
rect 2806 54 3000 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2752 54
rect 2798 52 3000 54
rect 0 -30 3000 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 1554 1522 1598 1566
rect 1598 1522 1606 1566
rect 1794 1522 1838 1566
rect 1838 1522 1846 1566
rect 2034 1522 2078 1566
rect 2078 1522 2086 1566
rect 2274 1522 2318 1566
rect 2318 1522 2326 1566
rect 2514 1522 2558 1566
rect 2558 1522 2566 1566
rect 2754 1522 2798 1566
rect 2798 1522 2806 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1554 1514 1606 1522
rect 1794 1514 1846 1522
rect 2034 1514 2086 1522
rect 2274 1514 2326 1522
rect 2514 1514 2566 1522
rect 2754 1514 2806 1522
rect 2654 884 2706 936
rect 104 712 112 756
rect 112 712 156 756
rect 104 704 156 712
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 2754 98 2806 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
rect 2754 54 2798 98
rect 2798 54 2806 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 1540 1570 1620 1580
rect 1780 1570 1860 1580
rect 2020 1570 2100 1580
rect 2260 1570 2340 1580
rect 2500 1570 2580 1580
rect 2740 1570 2820 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1480 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1480 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1480 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1480 1390 1514
rect 1530 1566 1630 1570
rect 1530 1514 1554 1566
rect 1606 1514 1630 1566
rect 1530 1480 1630 1514
rect 1770 1566 1870 1570
rect 1770 1514 1794 1566
rect 1846 1514 1870 1566
rect 1770 1480 1870 1514
rect 2010 1566 2110 1570
rect 2010 1514 2034 1566
rect 2086 1514 2110 1566
rect 2010 1480 2110 1514
rect 2250 1566 2350 1570
rect 2250 1514 2274 1566
rect 2326 1514 2350 1566
rect 2250 1480 2350 1514
rect 2490 1566 2590 1570
rect 2490 1514 2514 1566
rect 2566 1514 2590 1566
rect 2490 1480 2590 1514
rect 2730 1566 2830 1570
rect 2730 1514 2754 1566
rect 2806 1514 2830 1566
rect 2730 1480 2830 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 580 1470 660 1480
rect 820 1470 900 1480
rect 1060 1470 1140 1480
rect 1300 1470 1380 1480
rect 1540 1470 1620 1480
rect 1780 1470 1860 1480
rect 2020 1470 2100 1480
rect 2260 1470 2340 1480
rect 2500 1470 2580 1480
rect 2740 1470 2820 1480
rect 2630 936 2730 950
rect 2630 884 2654 936
rect 2706 884 2730 936
rect 2630 840 2730 884
rect 80 756 180 770
rect 80 704 104 756
rect 156 704 180 756
rect 80 660 180 704
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 2740 110 2820 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 20 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 20 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 20 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 20 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 20 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 20 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 20 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 20 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 20 2590 54
rect 2730 106 2830 110
rect 2730 54 2754 106
rect 2806 54 2830 106
rect 2730 20 2830 54
rect 100 10 180 20
rect 340 10 420 20
rect 580 10 660 20
rect 820 10 900 20
rect 1060 10 1140 20
rect 1300 10 1380 20
rect 1540 10 1620 20
rect 1780 10 1860 20
rect 2020 10 2100 20
rect 2260 10 2340 20
rect 2500 10 2580 20
rect 2740 10 2820 20
<< labels >>
rlabel metal2 s 100 1470 180 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 100 10 180 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 80 660 180 740 4 A
port 1 nsew signal input
rlabel metal2 s 2630 840 2730 920 4 Y
port 2 nsew signal output
rlabel metal1 s 80 670 180 730 1 A
port 1 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 580 1470 660 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 570 1480 670 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 820 1470 900 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 810 1480 910 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1060 1470 1140 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1050 1480 1150 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1300 1470 1380 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1290 1480 1390 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1540 1470 1620 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1530 1480 1630 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1780 1470 1860 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1770 1480 1870 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2020 1470 2100 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2010 1480 2110 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2260 1470 2340 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2250 1480 2350 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2500 1470 2580 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2490 1480 2590 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2740 1470 2820 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2730 1480 2830 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 1060 840 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1130 1060 1180 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1470 1060 1520 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1810 1060 1860 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 1060 2200 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2490 1060 2540 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2830 1060 2880 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1470 3000 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 580 10 660 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 570 20 670 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 820 10 900 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 810 20 910 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1060 10 1140 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1050 20 1150 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1300 10 1380 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1290 20 1390 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1540 10 1620 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1530 20 1630 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1780 10 1860 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1770 20 1870 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2020 10 2100 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2010 20 2110 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2260 10 2340 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2250 20 2350 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2500 10 2580 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2490 20 2590 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2740 10 2820 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2730 20 2830 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 -30 840 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1130 -30 1180 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1470 -30 1520 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1810 -30 1860 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2150 -30 2200 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2490 -30 2540 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2830 -30 2880 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 -30 3000 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 620 160 670 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 960 160 1010 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 160 1350 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1640 160 1690 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 1980 160 2030 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 2320 160 2370 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 380 2710 430 1 Y
port 2 nsew signal output
rlabel metal1 s 2630 840 2710 910 1 Y
port 2 nsew signal output
rlabel metal1 s 280 860 2710 910 1 Y
port 2 nsew signal output
rlabel metal1 s 2660 160 2710 1400 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 3000 1590
string GDS_END 216518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 194022
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
