magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 111 78 123
rect 28 85 33 111
rect 62 76 67 104
rect 60 70 70 76
rect 32 57 42 63
rect 12 44 22 50
rect 47 44 57 50
rect 62 38 67 70
rect 14 12 19 36
rect 42 33 67 38
rect 42 19 47 33
rect 59 12 64 28
rect 0 0 78 12
<< obsm1 >>
rect 11 80 16 104
rect 45 80 50 104
rect 11 75 50 80
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 60 69 70 77
rect 32 56 42 64
rect 12 43 22 51
rect 47 43 57 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 s 12 43 22 51 6 A0
port 2 nsew signal input
rlabel metal1 s 12 44 22 50 6 A0
port 2 nsew signal input
rlabel metal2 s 32 56 42 64 6 A1
port 3 nsew signal input
rlabel metal1 s 32 57 42 63 6 A1
port 3 nsew signal input
rlabel metal2 s 47 43 57 51 6 B
port 4 nsew signal input
rlabel metal1 s 47 44 57 50 6 B
port 4 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal1 s 28 85 33 123 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 111 78 123 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal1 s 14 0 19 36 6 VSS
port 10 nsew ground bidirectional
rlabel metal1 s 59 0 64 28 6 VSS
port 10 nsew ground bidirectional
rlabel metal1 s 0 0 78 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 60 69 70 77 6 Y
port 1 nsew signal output
rlabel metal1 s 42 19 47 38 6 Y
port 1 nsew signal output
rlabel metal1 s 42 33 67 38 6 Y
port 1 nsew signal output
rlabel metal1 s 62 33 67 104 6 Y
port 1 nsew signal output
rlabel metal1 s 60 70 70 76 6 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 78 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 55012
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 48056
<< end >>
