magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3894 1094
<< pwell >>
rect -86 -86 3894 453
<< mvnmos >>
rect 124 170 244 328
rect 348 170 468 328
rect 716 169 836 309
rect 940 169 1060 309
rect 1164 169 1284 309
rect 1332 169 1452 309
rect 1536 169 1656 309
rect 1804 169 1924 309
rect 2030 169 2150 309
rect 2254 169 2374 309
rect 2478 169 2598 309
rect 2702 169 2822 309
rect 2962 73 3082 309
rect 3340 83 3460 333
rect 3564 83 3684 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 720 593 820 793
rect 924 593 1024 793
rect 1128 593 1228 793
rect 1332 593 1432 793
rect 1536 593 1636 793
rect 1884 628 1984 828
rect 2088 628 2188 828
rect 2292 628 2392 828
rect 2496 628 2596 828
rect 2744 573 2844 939
rect 2948 573 3048 939
rect 3360 573 3460 939
rect 3564 573 3664 939
<< mvndiff >>
rect 36 315 124 328
rect 36 269 49 315
rect 95 269 124 315
rect 36 170 124 269
rect 244 229 348 328
rect 244 183 273 229
rect 319 183 348 229
rect 244 170 348 183
rect 468 315 556 328
rect 468 269 497 315
rect 543 269 556 315
rect 468 170 556 269
rect 628 228 716 309
rect 628 182 641 228
rect 687 182 716 228
rect 628 169 716 182
rect 836 296 940 309
rect 836 250 865 296
rect 911 250 940 296
rect 836 169 940 250
rect 1060 294 1164 309
rect 1060 248 1089 294
rect 1135 248 1164 294
rect 1060 169 1164 248
rect 1284 169 1332 309
rect 1452 169 1536 309
rect 1656 228 1804 309
rect 1656 182 1685 228
rect 1731 182 1804 228
rect 1656 169 1804 182
rect 1924 296 2030 309
rect 1924 250 1953 296
rect 1999 250 2030 296
rect 1924 169 2030 250
rect 2150 296 2254 309
rect 2150 250 2179 296
rect 2225 250 2254 296
rect 2150 169 2254 250
rect 2374 296 2478 309
rect 2374 250 2403 296
rect 2449 250 2478 296
rect 2374 169 2478 250
rect 2598 228 2702 309
rect 2598 182 2627 228
rect 2673 182 2702 228
rect 2598 169 2702 182
rect 2822 169 2962 309
rect 2882 73 2962 169
rect 3082 296 3170 309
rect 3082 156 3111 296
rect 3157 156 3170 296
rect 3082 73 3170 156
rect 3252 236 3340 333
rect 3252 96 3265 236
rect 3311 96 3340 236
rect 3252 83 3340 96
rect 3460 320 3564 333
rect 3460 180 3489 320
rect 3535 180 3564 320
rect 3460 83 3564 180
rect 3684 236 3772 333
rect 3684 96 3713 236
rect 3759 96 3772 236
rect 3684 83 3772 96
<< mvpdiff >>
rect 56 736 144 849
rect 56 596 69 736
rect 115 596 144 736
rect 56 573 144 596
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 2656 926 2744 939
rect 2656 880 2669 926
rect 2715 880 2744 926
rect 2656 828 2744 880
rect 1796 815 1884 828
rect 448 586 477 726
rect 523 586 536 726
rect 632 780 720 793
rect 632 734 645 780
rect 691 734 720 780
rect 632 593 720 734
rect 820 746 924 793
rect 820 606 849 746
rect 895 606 924 746
rect 820 593 924 606
rect 1024 746 1128 793
rect 1024 606 1053 746
rect 1099 606 1128 746
rect 1024 593 1128 606
rect 1228 780 1332 793
rect 1228 640 1257 780
rect 1303 640 1332 780
rect 1228 593 1332 640
rect 1432 780 1536 793
rect 1432 734 1461 780
rect 1507 734 1536 780
rect 1432 593 1536 734
rect 1636 780 1724 793
rect 1636 640 1665 780
rect 1711 640 1724 780
rect 1636 593 1724 640
rect 1796 675 1809 815
rect 1855 675 1884 815
rect 1796 628 1884 675
rect 1984 781 2088 828
rect 1984 641 2013 781
rect 2059 641 2088 781
rect 1984 628 2088 641
rect 2188 781 2292 828
rect 2188 641 2217 781
rect 2263 641 2292 781
rect 2188 628 2292 641
rect 2392 687 2496 828
rect 2392 641 2421 687
rect 2467 641 2496 687
rect 2392 628 2496 641
rect 2596 628 2744 828
rect 448 573 536 586
rect 2664 573 2744 628
rect 2844 634 2948 939
rect 2844 588 2873 634
rect 2919 588 2948 634
rect 2844 573 2948 588
rect 3048 926 3136 939
rect 3048 786 3077 926
rect 3123 786 3136 926
rect 3048 573 3136 786
rect 3272 926 3360 939
rect 3272 786 3285 926
rect 3331 786 3360 926
rect 3272 573 3360 786
rect 3460 726 3564 939
rect 3460 586 3489 726
rect 3535 586 3564 726
rect 3460 573 3564 586
rect 3664 926 3752 939
rect 3664 786 3693 926
rect 3739 786 3752 926
rect 3664 573 3752 786
<< mvndiffc >>
rect 49 269 95 315
rect 273 183 319 229
rect 497 269 543 315
rect 641 182 687 228
rect 865 250 911 296
rect 1089 248 1135 294
rect 1685 182 1731 228
rect 1953 250 1999 296
rect 2179 250 2225 296
rect 2403 250 2449 296
rect 2627 182 2673 228
rect 3111 156 3157 296
rect 3265 96 3311 236
rect 3489 180 3535 320
rect 3713 96 3759 236
<< mvpdiffc >>
rect 69 596 115 736
rect 273 696 319 836
rect 2669 880 2715 926
rect 477 586 523 726
rect 645 734 691 780
rect 849 606 895 746
rect 1053 606 1099 746
rect 1257 640 1303 780
rect 1461 734 1507 780
rect 1665 640 1711 780
rect 1809 675 1855 815
rect 2013 641 2059 781
rect 2217 641 2263 781
rect 2421 641 2467 687
rect 2873 588 2919 634
rect 3077 786 3123 926
rect 3285 786 3331 926
rect 3489 586 3535 726
rect 3693 786 3739 926
<< polysilicon >>
rect 348 933 2188 973
rect 2744 939 2844 983
rect 2948 939 3048 983
rect 3360 939 3460 983
rect 3564 939 3664 983
rect 144 849 244 893
rect 348 849 448 933
rect 924 872 1024 885
rect 720 793 820 837
rect 924 826 937 872
rect 983 826 1024 872
rect 924 793 1024 826
rect 1128 793 1228 933
rect 1332 793 1432 837
rect 1536 793 1636 837
rect 1884 828 1984 872
rect 2088 828 2188 933
rect 2292 828 2392 872
rect 2496 828 2596 872
rect 144 499 244 573
rect 144 453 157 499
rect 203 453 244 499
rect 144 372 244 453
rect 124 328 244 372
rect 348 407 448 573
rect 348 361 361 407
rect 407 372 448 407
rect 720 523 820 593
rect 720 477 733 523
rect 779 477 820 523
rect 407 361 468 372
rect 348 328 468 361
rect 720 353 820 477
rect 924 501 1024 593
rect 1128 549 1228 593
rect 924 461 1284 501
rect 1164 388 1284 461
rect 716 309 836 353
rect 940 309 1060 353
rect 1164 342 1182 388
rect 1228 342 1284 388
rect 1164 309 1284 342
rect 1332 491 1432 593
rect 1332 445 1373 491
rect 1419 445 1432 491
rect 1332 353 1432 445
rect 1536 353 1636 593
rect 1884 583 1984 628
rect 1884 537 1897 583
rect 1943 537 1984 583
rect 1884 369 1984 537
rect 2088 489 2188 628
rect 2292 595 2392 628
rect 2292 549 2317 595
rect 2363 549 2392 595
rect 2292 536 2392 549
rect 2496 595 2596 628
rect 2496 549 2537 595
rect 2583 549 2596 595
rect 2088 486 2274 489
rect 2088 449 2374 486
rect 2032 388 2150 401
rect 1332 309 1452 353
rect 1536 309 1656 353
rect 1804 309 1924 369
rect 2032 353 2045 388
rect 2030 342 2045 353
rect 2091 342 2150 388
rect 2030 309 2150 342
rect 2254 309 2374 449
rect 2496 353 2596 549
rect 2744 523 2844 573
rect 2948 540 3048 573
rect 2948 529 2985 540
rect 2744 477 2757 523
rect 2803 477 2844 523
rect 2744 369 2844 477
rect 2962 494 2985 529
rect 3031 494 3048 540
rect 2478 309 2598 353
rect 2702 309 2822 369
rect 2962 353 3048 494
rect 3360 464 3460 573
rect 3564 464 3664 573
rect 3360 425 3664 464
rect 3340 412 3664 425
rect 3340 366 3353 412
rect 3399 393 3664 412
rect 3399 366 3460 393
rect 2962 309 3082 353
rect 3340 333 3460 366
rect 3564 377 3664 393
rect 3564 333 3684 377
rect 124 126 244 170
rect 348 77 468 170
rect 716 125 836 169
rect 940 77 1060 169
rect 1164 125 1284 169
rect 1332 125 1452 169
rect 348 37 1060 77
rect 1536 77 1656 169
rect 1804 125 1924 169
rect 2030 125 2150 169
rect 2254 125 2374 169
rect 2478 125 2598 169
rect 2702 77 2822 169
rect 1536 37 2822 77
rect 2962 29 3082 73
rect 3340 39 3460 83
rect 3564 39 3684 83
<< polycontact >>
rect 937 826 983 872
rect 157 453 203 499
rect 361 361 407 407
rect 733 477 779 523
rect 1182 342 1228 388
rect 1373 445 1419 491
rect 1897 537 1943 583
rect 2317 549 2363 595
rect 2537 549 2583 595
rect 2045 342 2091 388
rect 2757 477 2803 523
rect 2985 494 3031 540
rect 3353 366 3399 412
<< metal1 >>
rect 0 926 3808 1098
rect 0 918 2669 926
rect 273 836 319 918
rect 69 736 115 747
rect 645 780 691 918
rect 273 685 319 696
rect 477 726 523 737
rect 115 596 418 639
rect 69 593 418 596
rect 69 585 115 593
rect 142 499 318 542
rect 142 453 157 499
rect 203 453 318 499
rect 372 407 418 593
rect 49 361 361 407
rect 407 361 418 407
rect 645 723 691 734
rect 737 826 937 872
rect 983 826 994 872
rect 737 677 783 826
rect 1257 780 1303 791
rect 523 631 783 677
rect 849 746 911 757
rect 523 586 543 631
rect 49 315 95 361
rect 49 258 95 269
rect 477 315 543 586
rect 895 606 911 746
rect 592 523 779 542
rect 592 477 733 523
rect 592 466 779 477
rect 477 269 497 315
rect 477 258 543 269
rect 849 296 911 606
rect 849 250 865 296
rect 273 229 319 240
rect 849 239 911 250
rect 1053 746 1099 757
rect 1461 780 1507 918
rect 1809 815 1855 918
rect 2715 918 3077 926
rect 2669 869 2715 880
rect 1461 723 1507 734
rect 1665 780 1711 791
rect 1303 640 1665 675
rect 1809 664 1855 675
rect 2013 781 2059 792
rect 1257 629 1711 640
rect 1053 583 1099 606
rect 1053 537 1897 583
rect 1943 537 1954 583
rect 1053 305 1099 537
rect 2013 491 2059 641
rect 1362 445 1373 491
rect 1419 445 2059 491
rect 2179 781 3031 792
rect 2179 641 2217 781
rect 2263 746 3031 781
rect 3123 918 3285 926
rect 3077 775 3123 786
rect 3331 918 3693 926
rect 3285 775 3331 786
rect 3739 918 3808 926
rect 3693 775 3739 786
rect 1171 342 1182 388
rect 1228 342 1907 388
rect 1053 294 1135 305
rect 1053 248 1089 294
rect 273 90 319 183
rect 641 228 687 239
rect 1053 237 1135 248
rect 641 90 687 182
rect 1685 228 1731 239
rect 1685 90 1731 182
rect 1861 193 1907 342
rect 1953 296 1999 445
rect 1953 239 1999 250
rect 2045 388 2091 399
rect 2045 193 2091 342
rect 2179 296 2263 641
rect 2421 687 2467 698
rect 2225 250 2263 296
rect 2179 239 2263 250
rect 2311 595 2363 606
rect 2311 549 2317 595
rect 2311 538 2363 549
rect 2311 193 2357 538
rect 2421 307 2467 641
rect 2526 595 2873 634
rect 2526 549 2537 595
rect 2583 588 2873 595
rect 2919 588 2939 634
rect 2583 549 2594 588
rect 2718 523 2803 542
rect 2718 477 2757 523
rect 2718 466 2803 477
rect 2893 437 2939 588
rect 2985 540 3031 746
rect 2985 483 3031 494
rect 3489 726 3554 737
rect 3535 586 3554 726
rect 2893 412 3410 437
rect 2893 391 3353 412
rect 2403 296 2467 307
rect 2449 250 2467 296
rect 2403 239 2467 250
rect 3111 366 3353 391
rect 3399 366 3410 412
rect 3111 296 3157 366
rect 1861 147 2357 193
rect 2627 228 2673 239
rect 2627 90 2673 182
rect 3489 320 3554 586
rect 3111 145 3157 156
rect 3265 236 3311 247
rect 3535 180 3554 320
rect 3489 169 3554 180
rect 3713 236 3759 247
rect 3265 90 3311 96
rect 3713 90 3759 96
rect 0 -90 3808 90
<< labels >>
flabel metal1 s 142 453 318 542 0 FreeSans 200 0 0 0 CLK
port 3 nsew clock input
flabel metal1 s 592 466 779 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3489 169 3554 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2718 466 2803 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 0 918 3808 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3713 240 3759 247 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3693 869 3739 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3285 869 3331 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3077 869 3123 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2669 869 2715 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 869 1855 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 869 1507 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 869 691 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 869 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3693 775 3739 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3285 775 3331 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3077 775 3123 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 775 1855 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 775 1507 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 775 691 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 869 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 723 1855 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1461 723 1507 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 723 691 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 723 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 685 1855 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1809 664 1855 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3265 240 3311 247 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3713 239 3759 240 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3265 239 3311 240 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 239 319 240 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3713 90 3759 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3265 90 3311 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2627 90 2673 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1685 90 1731 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 239 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3808 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 1008
string GDS_END 611138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 602046
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
