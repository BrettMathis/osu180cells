****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__addf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__addf_1 A B CI S CO VDD VSS
X0 a_9_70# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_110_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 S a_161_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 S a_161_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_195_19# B a_178_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_178_19# A a_161_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_195_70# B a_178_70# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_110_19# CI VSS VSS nmos_3p3 w=0.85u l=0.3u
X8 a_178_70# A a_161_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_59_19# CI a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS B a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_110_70# CI VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_59_19# CI a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD B a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X15 CO a_59_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VDD A a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS CI a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 CO a_59_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 VDD CI a_195_70# VDD pmos_3p3 w=1.7u l=0.3u
X20 VSS A a_76_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_161_19# a_59_19# a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X22 a_76_19# B a_59_19# VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD A a_76_70# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_161_19# a_59_19# a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X25 a_9_19# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X26 a_110_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X27 a_76_70# B a_59_19# VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__addf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__addh_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__addh_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__addh_1 A B S CO VDD VSS
X0 a_19_14# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_91_19# B a_91_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS a_19_14# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_19_14# a_91_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_19_14# B a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS a_19_14# CO VSS nmos_3p3 w=0.85u l=0.3u
X6 VDD B a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD a_19_14# CO VDD pmos_3p3 w=1.7u l=0.3u
X8 S a_91_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 a_91_19# A a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 S a_91_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X11 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 a_91_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 a_75_19# B a_91_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__addh_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__and2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__and2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__and2_1 A B Y VDD VSS
X0 VDD B a_12_19# VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_12_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y a_12_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_12_19# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_28_19# A a_12_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS B a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__and2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__aoi21_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__aoi21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__aoi21_1 Y A0 A1 B VDD VSS
X0 a_9_70# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS B Y VSS nmos_3p3 w=0.85u l=0.3u
X2 Y B a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD A0 a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_28_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 Y A1 a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__aoi21_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__aoi22_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__aoi22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__aoi22_1 A0 A1 B0 B1 Y VDD VSS
X0 a_9_70# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_56_19# B0 Y VSS nmos_3p3 w=0.85u l=0.3u
X2 Y B0 a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD A0 a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS B1 a_56_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_28_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_9_70# B1 Y VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A1 a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__aoi22_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__buf_1 A Y VDD VSS
X0 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__buf_16 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X13 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X16 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X17 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X18 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X19 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X20 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X21 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X22 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X25 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X26 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X27 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X29 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X30 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X31 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X32 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X33 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__buf_2 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__buf_4 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__buf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__buf_8 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X15 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__buf_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkbuf_1 A Y VDD VSS
X0 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X1 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkbuf_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkbuf_16 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X13 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X16 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X17 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X18 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X19 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X20 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X21 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X22 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X25 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X26 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X27 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X29 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X30 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X31 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X32 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X33 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkbuf_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkbuf_2 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkbuf_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkbuf_4 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkbuf_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkbuf_8 A Y VDD VSS
X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X15 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 Y a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkbuf_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_1 A Y VDD VSS
X0 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_16 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X13 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X18 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X20 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X22 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X23 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X24 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X26 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X27 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X28 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X29 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X30 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X31 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
C0 Y VDD 2.058360fF
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_2 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_4 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_8 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X3 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X6 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X14 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X15 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__clkinv_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__dff_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dff_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dff_1 D Q QN CLK VDD VSS
X0 a_42_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_125_19# a_53_38# a_114_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_86_70# a_53_38# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD a_161_42# a_148_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS a_9_19# a_86_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_19_14# a_53_38# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS a_161_42# QN VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# a_86_70# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_19_14# CLK a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD a_161_42# QN VDD pmos_3p3 w=1.7u l=0.3u
X10 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_53_38# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X13 a_53_38# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 a_148_19# a_53_38# a_125_19# VSS nmos_3p3 w=0.85u l=0.3u
X15 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 a_114_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X17 a_161_42# a_125_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X18 a_148_70# CLK a_125_19# VDD pmos_3p3 w=1.7u l=0.3u
X19 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X20 a_114_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X21 a_161_42# a_125_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 a_125_19# CLK a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X24 a_86_19# CLK a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS a_161_42# a_148_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__dff_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__dffn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dffn_1 D Q QN CLK VDD VSS
X0 a_42_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_125_19# a_53_38# a_114_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 a_161_42# a_125_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 a_86_70# a_53_38# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X5 VDD a_161_42# a_148_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS a_9_19# a_86_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_19_14# a_53_38# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X9 a_161_42# a_125_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_9_19# a_86_70# VDD pmos_3p3 w=1.7u l=0.3u
X11 a_19_14# a_50_59# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_53_38# a_50_59# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS a_161_42# QN VSS nmos_3p3 w=0.85u l=0.3u
X16 a_53_38# a_50_59# VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS CLK a_50_59# VSS nmos_3p3 w=0.85u l=0.3u
X18 VDD a_161_42# QN VDD pmos_3p3 w=1.7u l=0.3u
X19 a_148_19# a_53_38# a_125_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_114_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD CLK a_50_59# VDD pmos_3p3 w=1.7u l=0.3u
X22 a_148_70# a_50_59# a_125_19# VDD pmos_3p3 w=1.7u l=0.3u
X23 a_114_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 a_125_19# a_50_59# a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X26 a_86_19# a_50_59# a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X27 VSS a_161_42# a_148_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__dffn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__dffsr_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dffsr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dffsr_1 D Q QN SN RN CLK VDD VSS
X0 a_172_70# a_139_41# a_82_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_247_47# a_25_19# a_291_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS a_41_70# a_172_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_41_70# a_172_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS a_247_47# a_234_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD a_247_47# a_234_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_41_70# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_128_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X8 VSS a_247_47# QN VSS nmos_3p3 w=0.85u l=0.3u
X9 a_310_19# a_211_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 a_128_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 VDD a_247_47# QN VDD pmos_3p3 w=1.7u l=0.3u
X13 VDD SN a_57_70# VDD pmos_3p3 w=1.7u l=0.3u
X14 a_200_19# a_41_70# VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 a_247_47# SN a_310_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 a_57_70# a_25_19# a_41_70# VDD pmos_3p3 w=1.7u l=0.3u
X18 a_291_70# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 a_211_19# CLK a_200_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_200_70# a_41_70# VDD VDD pmos_3p3 w=1.7u l=0.3u
X21 VDD a_211_19# a_291_70# VDD pmos_3p3 w=1.7u l=0.3u
X22 a_82_14# a_139_41# a_128_19# VSS nmos_3p3 w=0.85u l=0.3u
X23 a_139_41# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X24 a_211_19# a_139_41# a_200_70# VDD pmos_3p3 w=1.7u l=0.3u
X25 a_82_14# CLK a_128_70# VDD pmos_3p3 w=1.7u l=0.3u
X26 a_139_41# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X27 a_77_19# SN a_41_70# VSS nmos_3p3 w=0.85u l=0.3u
X28 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X29 a_234_19# a_139_41# a_211_19# VSS nmos_3p3 w=0.85u l=0.3u
X30 a_172_19# CLK a_82_14# VSS nmos_3p3 w=0.85u l=0.3u
X31 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X32 VSS a_82_14# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X33 a_57_70# a_82_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X34 a_234_70# CLK a_211_19# VDD pmos_3p3 w=1.7u l=0.3u
X35 VSS a_25_19# a_247_47# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__dffsr_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__dlat_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dlat_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dlat_1 D Q CLK VDD VSS
X0 VDD a_10_19# a_77_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_52_58# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 VDD a_20_14# a_10_19# VDD pmos_3p3 w=1.7u l=0.3u
X3 Q a_137_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_52_58# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 a_46_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_20_14# CLK a_46_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 a_20_14# a_52_58# a_43_70# VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS a_10_19# a_137_19# VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD a_10_19# a_137_19# VDD pmos_3p3 w=1.7u l=0.3u
X10 a_77_19# a_52_58# a_20_14# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_77_70# CLK a_20_14# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_20_14# a_10_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 Q a_137_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 a_43_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS a_10_19# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__dlat_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__dlatn_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dlatn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dlatn_1 D Q CLK VDD VSS
X0 VDD a_10_19# a_77_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD CLK a_54_14# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_52_58# a_54_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD a_20_14# a_10_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_52_58# a_54_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 a_46_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_20_14# a_54_14# a_46_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 VSS a_10_19# a_173_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_20_14# a_52_58# a_43_70# VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD a_10_19# a_173_19# VDD pmos_3p3 w=1.7u l=0.3u
X10 a_77_19# a_52_58# a_20_14# VSS nmos_3p3 w=0.85u l=0.3u
X11 Q a_173_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 a_77_70# a_54_14# a_20_14# VDD pmos_3p3 w=1.7u l=0.3u
X13 Q a_173_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 VSS CLK a_54_14# VSS nmos_3p3 w=0.85u l=0.3u
X15 VSS a_20_14# a_10_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 a_43_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS a_10_19# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__dlatn_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__fill_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__fill_1 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__fill_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__fill_16 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__fill_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__fill_2 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__fill_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__fill_4 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__fill_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__fill_8 VDD VSS
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__fill_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__inv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__inv_1 A Y VDD VSS
X0 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_16.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__inv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__inv_16 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X3 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X13 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X18 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X20 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X22 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X23 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X24 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X26 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X27 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X28 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X29 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X30 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X31 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
C0 Y VDD 2.058360fF
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_16.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_2.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__inv_2.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__inv_2 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_2.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_4.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__inv_4.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__inv_4 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X7 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_4.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_8.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__inv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__inv_8 A Y VDD VSS
X0 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X3 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
X6 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X12 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X14 VSS A Y VSS nmos_3p3 w=0.85u l=0.3u
X15 VDD A Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__inv_8.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__lshifdown.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__lshifdown.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__lshifdown A Y VDDH VDD VSS
X0 a_26_19# A VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X1 Y a_26_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y a_26_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_26_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__lshifdown.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__lshifup.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__lshifup.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__lshifup A Y VDDH VDD VSS
X0 a_77_55# a_26_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 a_26_19# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_77_55# a_67_19# VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X3 Y a_67_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 Y a_67_19# VDDH VDDH pmos_3p3 w=1.7u l=0.3u
X5 VSS A a_67_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 VDDH a_77_55# a_67_19# VDDH pmos_3p3 w=1.7u l=0.3u
X7 a_26_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__lshifup.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__mux2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__mux2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__mux2_1 A B Sel Y VDD VSS
X0 Y a_25_19# A VSS nmos_3p3 w=0.85u l=0.3u
X1 a_25_19# Sel VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y Sel A VDD pmos_3p3 w=1.7u l=0.3u
X3 a_25_19# Sel VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 B Sel Y VSS nmos_3p3 w=0.85u l=0.3u
X5 B a_25_19# Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__mux2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__nand2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nand2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__nand2_1 A B Y VDD VSS
X0 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_28_19# A Y VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS B a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__nand2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__nor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__nor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__nor2_1 A B Y VDD VSS
X0 Y B a_25_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_25_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS B Y VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__nor2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__oai21_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__oai21_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__oai21_1 A0 A1 B Y VDD VSS
X0 a_27_70# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A1 a_27_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y B a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS A0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X5 a_8_19# A1 VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__oai21_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__oai22_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__oai22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__oai22_1 A1 A0 B1 B0 Y VDD VSS
X0 a_27_70# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y A1 a_27_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y B0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VSS A0 a_8_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 a_58_70# B0 Y VDD pmos_3p3 w=1.7u l=0.3u
X5 VDD B1 a_58_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_8_19# B1 Y VSS nmos_3p3 w=0.85u l=0.3u
X7 a_8_19# A1 VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__oai22_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__oai31_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__oai31_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__oai31_1 A0 A1 A2 B Y VDD VSS
X0 a_25_19# A1 VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 a_25_19# A2 VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 Y A1 a_45_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 Y B a_25_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 a_34_70# A2 VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS A0 a_25_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_45_70# A0 a_34_70# VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__oai31_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__or2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__or2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__or2_1 A B Y VDD VSS
X0 VDD B a_25_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_9_70# VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 a_9_70# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 a_25_70# A a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 Y a_9_70# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 VSS B a_9_70# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__or2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__tbuf_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__tbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__tbuf_1 A Y EN VDD VSS
X0 Y a_49_56# a_44_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_49_56# EN VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_44_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 a_44_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 Y EN a_44_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 a_49_56# EN VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__tbuf_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__tieh.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__tieh.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__tieh Y VDD VSS
X0 a_19_14# a_19_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 Y a_19_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__tieh.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__tiel.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__tiel.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__tiel Y VDD VSS
X0 Y a_19_14# VSS VSS nmos_3p3 w=0.85u l=0.3u
X1 a_19_14# a_19_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__tiel.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__tinv_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__tinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__tinv_1 A Y EN VDD VSS
X0 Y a_9_19# a_44_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X3 a_44_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 a_44_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 Y EN a_44_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__tinv_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__xnor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__xnor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__xnor2_1 A B Y VDD VSS
X0 a_42_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_49_14# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_49_14# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_78_19# a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X6 VSS B a_78_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 a_78_70# A Y VDD pmos_3p3 w=1.7u l=0.3u
X8 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD B a_78_70# VDD pmos_3p3 w=1.7u l=0.3u
X10 Y a_49_14# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_49_14# B VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__xnor2_1.spice
****BEGIN OF FILE - gf180mcu_osu_sc_gp9t3v3__xor2_1.spice

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__xor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__xor2_1 A B Y VDD VSS
X0 a_42_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_52_59# a_81_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 VDD B a_81_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 Y B a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 Y a_52_59# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_81_19# a_9_19# Y VSS nmos_3p3 w=0.85u l=0.3u
X8 a_52_59# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 a_81_70# a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X10 a_52_59# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X11 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
.ends


****END OF FILE - gf180mcu_osu_sc_gp9t3v3__xor2_1.spice
