magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1120 844
rect 59 584 105 724
rect 710 657 778 724
rect 486 540 554 586
rect 248 519 554 540
rect 916 519 984 586
rect 248 473 984 519
rect 141 110 200 446
rect 248 110 319 473
rect 365 110 424 427
rect 472 360 674 424
rect 730 360 994 424
rect 472 232 532 360
rect 730 312 788 360
rect 578 248 788 312
rect 945 60 991 178
rect 0 -60 1120 60
<< obsm1 >>
rect 151 632 658 678
rect 151 538 197 632
rect 612 611 658 632
rect 824 632 1090 678
rect 824 611 870 632
rect 612 565 870 611
rect 49 492 197 538
rect 49 110 95 492
rect 1044 274 1090 632
rect 848 228 1090 274
rect 848 167 894 228
rect 486 121 894 167
rect 848 120 894 121
<< labels >>
rlabel metal1 s 365 110 424 427 6 A1
port 1 nsew default input
rlabel metal1 s 141 110 200 446 6 A2
port 2 nsew default input
rlabel metal1 s 472 360 674 424 6 B
port 3 nsew default input
rlabel metal1 s 472 232 532 360 6 B
port 3 nsew default input
rlabel metal1 s 730 360 994 424 6 C
port 4 nsew default input
rlabel metal1 s 730 312 788 360 6 C
port 4 nsew default input
rlabel metal1 s 578 248 788 312 6 C
port 4 nsew default input
rlabel metal1 s 916 540 984 586 6 ZN
port 5 nsew default output
rlabel metal1 s 486 540 554 586 6 ZN
port 5 nsew default output
rlabel metal1 s 916 519 984 540 6 ZN
port 5 nsew default output
rlabel metal1 s 248 519 554 540 6 ZN
port 5 nsew default output
rlabel metal1 s 248 473 984 519 6 ZN
port 5 nsew default output
rlabel metal1 s 248 110 319 473 6 ZN
port 5 nsew default output
rlabel metal1 s 0 724 1120 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 710 657 778 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 657 105 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 584 105 657 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 945 60 991 178 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1120 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 90518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 87160
<< end >>
