magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 2344 2616
<< mvpmos >>
rect 0 0 120 2496
rect 224 0 344 2496
rect 448 0 568 2496
rect 672 0 792 2496
rect 896 0 1016 2496
rect 1120 0 1240 2496
rect 1344 0 1464 2496
rect 1568 0 1688 2496
rect 1792 0 1912 2496
rect 2016 0 2136 2496
<< mvpdiff >>
rect -88 2483 0 2496
rect -88 13 -75 2483
rect -29 13 0 2483
rect -88 0 0 13
rect 120 2483 224 2496
rect 120 13 149 2483
rect 195 13 224 2483
rect 120 0 224 13
rect 344 2483 448 2496
rect 344 13 373 2483
rect 419 13 448 2483
rect 344 0 448 13
rect 568 2483 672 2496
rect 568 13 597 2483
rect 643 13 672 2483
rect 568 0 672 13
rect 792 2483 896 2496
rect 792 13 821 2483
rect 867 13 896 2483
rect 792 0 896 13
rect 1016 2483 1120 2496
rect 1016 13 1045 2483
rect 1091 13 1120 2483
rect 1016 0 1120 13
rect 1240 2483 1344 2496
rect 1240 13 1269 2483
rect 1315 13 1344 2483
rect 1240 0 1344 13
rect 1464 2483 1568 2496
rect 1464 13 1493 2483
rect 1539 13 1568 2483
rect 1464 0 1568 13
rect 1688 2483 1792 2496
rect 1688 13 1717 2483
rect 1763 13 1792 2483
rect 1688 0 1792 13
rect 1912 2483 2016 2496
rect 1912 13 1941 2483
rect 1987 13 2016 2483
rect 1912 0 2016 13
rect 2136 2483 2224 2496
rect 2136 13 2165 2483
rect 2211 13 2224 2483
rect 2136 0 2224 13
<< mvpdiffc >>
rect -75 13 -29 2483
rect 149 13 195 2483
rect 373 13 419 2483
rect 597 13 643 2483
rect 821 13 867 2483
rect 1045 13 1091 2483
rect 1269 13 1315 2483
rect 1493 13 1539 2483
rect 1717 13 1763 2483
rect 1941 13 1987 2483
rect 2165 13 2211 2483
<< polysilicon >>
rect 0 2496 120 2540
rect 224 2496 344 2540
rect 448 2496 568 2540
rect 672 2496 792 2540
rect 896 2496 1016 2540
rect 1120 2496 1240 2540
rect 1344 2496 1464 2540
rect 1568 2496 1688 2540
rect 1792 2496 1912 2540
rect 2016 2496 2136 2540
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
<< metal1 >>
rect -75 2483 -29 2496
rect -75 0 -29 13
rect 149 2483 195 2496
rect 149 0 195 13
rect 373 2483 419 2496
rect 373 0 419 13
rect 597 2483 643 2496
rect 597 0 643 13
rect 821 2483 867 2496
rect 821 0 867 13
rect 1045 2483 1091 2496
rect 1045 0 1091 13
rect 1269 2483 1315 2496
rect 1269 0 1315 13
rect 1493 2483 1539 2496
rect 1493 0 1539 13
rect 1717 2483 1763 2496
rect 1717 0 1763 13
rect 1941 2483 1987 2496
rect 1941 0 1987 13
rect 2165 2483 2211 2496
rect 2165 0 2211 13
<< labels >>
flabel metal1 s -52 1248 -52 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 2188 1248 2188 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1248 172 1248 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 1248 396 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 1248 620 1248 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 1248 844 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 1248 1068 1248 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 1248 1292 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 1248 1516 1248 0 FreeSans 400 0 0 0 D
flabel metal1 s 1740 1248 1740 1248 0 FreeSans 400 0 0 0 S
flabel metal1 s 1964 1248 1964 1248 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 769260
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 747902
<< end >>
