magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect 751 7142 870 7183
rect 1265 7142 1384 7183
rect 465 7096 870 7142
rect 465 7050 539 7096
rect 585 7050 697 7096
rect 743 7050 870 7096
rect 465 7004 870 7050
rect 975 7096 1384 7142
rect 975 7050 1049 7096
rect 1095 7050 1207 7096
rect 1253 7050 1384 7096
rect 975 7004 1384 7050
rect 751 6963 870 7004
rect 1265 6963 1384 7004
<< polycontact >>
rect 539 7050 585 7096
rect 697 7050 743 7096
rect 1049 7050 1095 7096
rect 1207 7050 1253 7096
<< metal1 >>
rect 325 8322 756 8520
rect 325 8270 459 8322
rect 511 8270 666 8322
rect 718 8270 756 8322
rect 325 8104 756 8270
rect 325 8052 459 8104
rect 511 8052 666 8104
rect 718 8052 756 8104
rect 325 7886 756 8052
rect 325 7834 459 7886
rect 511 7834 666 7886
rect 718 7834 756 7886
rect 325 7668 756 7834
rect 325 7616 459 7668
rect 511 7616 666 7668
rect 718 7616 756 7668
rect 325 7222 756 7616
rect 1148 8322 1276 8362
rect 1148 8270 1186 8322
rect 1238 8270 1276 8322
rect 1148 8104 1276 8270
rect 1148 8052 1186 8104
rect 1238 8052 1276 8104
rect 1148 7886 1276 8052
rect 1148 7834 1186 7886
rect 1238 7834 1276 7886
rect 1148 7668 1276 7834
rect 1148 7616 1186 7668
rect 1238 7616 1276 7668
rect 1148 7576 1276 7616
rect 421 7133 761 7140
rect 865 7133 980 7283
rect 421 7099 778 7133
rect 421 7047 459 7099
rect 511 7096 671 7099
rect 723 7096 778 7099
rect 511 7050 539 7096
rect 585 7050 671 7096
rect 743 7050 778 7096
rect 511 7047 671 7050
rect 723 7047 778 7050
rect 421 7013 778 7047
rect 865 7096 1288 7133
rect 865 7050 1049 7096
rect 1095 7050 1207 7096
rect 1253 7050 1288 7096
rect 865 7013 1288 7050
rect 421 7007 761 7013
rect 351 6825 756 6924
rect 865 6859 980 7013
rect 1379 6859 1494 7283
rect 351 6784 769 6825
rect 351 6732 679 6784
rect 731 6732 769 6784
rect 351 6589 769 6732
rect 350 6567 769 6589
rect 350 6515 679 6567
rect 731 6515 769 6567
rect 350 6349 769 6515
rect 350 6297 679 6349
rect 731 6297 769 6349
rect 350 6131 769 6297
rect 350 6079 679 6131
rect 731 6079 769 6131
rect 350 5913 769 6079
rect 350 5861 679 5913
rect 731 5861 769 5913
rect 350 5696 769 5861
rect 350 5644 679 5696
rect 731 5644 769 5696
rect 350 5604 769 5644
rect 1155 6784 1283 6825
rect 1155 6732 1193 6784
rect 1245 6732 1283 6784
rect 1155 6567 1283 6732
rect 1155 6515 1193 6567
rect 1245 6515 1283 6567
rect 1155 6349 1283 6515
rect 1155 6297 1193 6349
rect 1245 6297 1283 6349
rect 1155 6131 1283 6297
rect 1155 6079 1193 6131
rect 1245 6079 1283 6131
rect 1155 5913 1283 6079
rect 1155 5861 1193 5913
rect 1245 5861 1283 5913
rect 1155 5696 1283 5861
rect 1155 5644 1193 5696
rect 1245 5644 1283 5696
rect 1155 5604 1283 5644
rect 350 5603 763 5604
rect 1161 5603 1277 5604
rect 350 3694 756 5603
rect 351 3676 756 3694
rect 860 3987 984 4027
rect 860 3935 896 3987
rect 948 3935 984 3987
rect 860 3769 984 3935
rect 860 3717 896 3769
rect 948 3717 984 3769
rect 860 3677 984 3717
rect 1374 3987 1498 4027
rect 1374 3935 1410 3987
rect 1462 3935 1498 3987
rect 1374 3769 1498 3935
rect 1374 3717 1410 3769
rect 1462 3717 1498 3769
rect 1374 3677 1498 3717
rect -106 3481 1824 3574
rect -106 3279 1824 3372
rect -106 3078 1824 3170
rect -106 2876 1824 2969
rect -106 2674 1824 2767
rect -106 2472 1824 2565
rect 423 1624 547 1664
rect 423 1572 459 1624
rect 511 1572 547 1624
rect 423 1406 547 1572
rect 423 1354 459 1406
rect 511 1354 547 1406
rect 423 1314 547 1354
<< via1 >>
rect 459 8270 511 8322
rect 666 8270 718 8322
rect 459 8052 511 8104
rect 666 8052 718 8104
rect 459 7834 511 7886
rect 666 7834 718 7886
rect 459 7616 511 7668
rect 666 7616 718 7668
rect 1186 8270 1238 8322
rect 1186 8052 1238 8104
rect 1186 7834 1238 7886
rect 1186 7616 1238 7668
rect 459 7047 511 7099
rect 671 7096 723 7099
rect 671 7050 697 7096
rect 697 7050 723 7096
rect 671 7047 723 7050
rect 679 6732 731 6784
rect 679 6515 731 6567
rect 679 6297 731 6349
rect 679 6079 731 6131
rect 679 5861 731 5913
rect 679 5644 731 5696
rect 1193 6732 1245 6784
rect 1193 6515 1245 6567
rect 1193 6297 1245 6349
rect 1193 6079 1245 6131
rect 1193 5861 1245 5913
rect 1193 5644 1245 5696
rect 896 3935 948 3987
rect 896 3717 948 3769
rect 1410 3935 1462 3987
rect 1410 3717 1462 3769
rect 459 1572 511 1624
rect 459 1354 511 1406
<< metal2 >>
rect 421 8324 756 8362
rect 421 8268 457 8324
rect 513 8268 664 8324
rect 720 8268 756 8324
rect 421 8106 756 8268
rect 421 8050 457 8106
rect 513 8050 664 8106
rect 720 8050 756 8106
rect 421 7888 756 8050
rect 421 7832 457 7888
rect 513 7832 664 7888
rect 720 7832 756 7888
rect 421 7670 756 7832
rect 421 7614 457 7670
rect 513 7614 664 7670
rect 720 7614 756 7670
rect 421 7575 756 7614
rect 1148 8324 1276 8361
rect 1148 8268 1184 8324
rect 1240 8268 1276 8324
rect 1148 8106 1276 8268
rect 1148 8050 1184 8106
rect 1240 8050 1276 8106
rect 1148 7888 1276 8050
rect 1148 7832 1184 7888
rect 1240 7832 1276 7888
rect 1148 7670 1276 7832
rect 1148 7614 1184 7670
rect 1240 7614 1276 7670
rect 1148 7576 1276 7614
rect 421 7099 761 7140
rect 421 7047 459 7099
rect 511 7047 671 7099
rect 723 7047 761 7099
rect 421 7007 761 7047
rect 421 1624 550 7007
rect 641 6786 769 6825
rect 641 6730 677 6786
rect 733 6730 769 6786
rect 641 6569 769 6730
rect 641 6513 677 6569
rect 733 6513 769 6569
rect 641 6351 769 6513
rect 641 6295 677 6351
rect 733 6295 769 6351
rect 641 6133 769 6295
rect 641 6077 677 6133
rect 733 6077 769 6133
rect 641 5915 769 6077
rect 641 5859 677 5915
rect 733 5859 769 5915
rect 641 5698 769 5859
rect 641 5642 677 5698
rect 733 5642 769 5698
rect 641 5603 769 5642
rect 1155 6786 1283 6825
rect 1155 6730 1191 6786
rect 1247 6730 1283 6786
rect 1155 6569 1283 6730
rect 1155 6513 1191 6569
rect 1247 6513 1283 6569
rect 1155 6351 1283 6513
rect 1155 6295 1191 6351
rect 1247 6295 1283 6351
rect 1155 6133 1283 6295
rect 1155 6077 1191 6133
rect 1247 6077 1283 6133
rect 1155 5915 1283 6077
rect 1155 5859 1191 5915
rect 1247 5859 1283 5915
rect 1155 5698 1283 5859
rect 1155 5642 1191 5698
rect 1247 5642 1283 5698
rect 1155 5603 1283 5642
rect 1635 4233 1760 4272
rect 1635 4177 1670 4233
rect 1726 4177 1760 4233
rect 1635 4057 1760 4177
rect 860 3987 984 4027
rect 860 3935 896 3987
rect 948 3935 984 3987
rect 860 3769 984 3935
rect 1374 3987 1498 4027
rect 1374 3935 1410 3987
rect 1462 3935 1498 3987
rect 860 3717 896 3769
rect 948 3717 984 3769
rect 860 3677 984 3717
rect 1144 3757 1272 3796
rect 1144 3701 1180 3757
rect 1236 3701 1272 3757
rect 421 1572 459 1624
rect 511 1572 550 1624
rect 421 1406 550 1572
rect 421 1359 459 1406
rect 423 1354 459 1359
rect 511 1359 550 1406
rect 1144 3539 1272 3701
rect 1374 3769 1498 3935
rect 1374 3717 1410 3769
rect 1462 3717 1498 3769
rect 1374 3677 1498 3717
rect 1634 4015 1762 4057
rect 1634 3959 1670 4015
rect 1726 3959 1762 4015
rect 1144 3483 1180 3539
rect 1236 3483 1272 3539
rect 1144 1413 1272 3483
rect 1634 1615 1762 3959
rect 511 1354 547 1359
rect 423 1314 547 1354
rect 1144 1280 1762 1413
<< via2 >>
rect 457 8322 513 8324
rect 457 8270 459 8322
rect 459 8270 511 8322
rect 511 8270 513 8322
rect 457 8268 513 8270
rect 664 8322 720 8324
rect 664 8270 666 8322
rect 666 8270 718 8322
rect 718 8270 720 8322
rect 664 8268 720 8270
rect 457 8104 513 8106
rect 457 8052 459 8104
rect 459 8052 511 8104
rect 511 8052 513 8104
rect 457 8050 513 8052
rect 664 8104 720 8106
rect 664 8052 666 8104
rect 666 8052 718 8104
rect 718 8052 720 8104
rect 664 8050 720 8052
rect 457 7886 513 7888
rect 457 7834 459 7886
rect 459 7834 511 7886
rect 511 7834 513 7886
rect 457 7832 513 7834
rect 664 7886 720 7888
rect 664 7834 666 7886
rect 666 7834 718 7886
rect 718 7834 720 7886
rect 664 7832 720 7834
rect 457 7668 513 7670
rect 457 7616 459 7668
rect 459 7616 511 7668
rect 511 7616 513 7668
rect 457 7614 513 7616
rect 664 7668 720 7670
rect 664 7616 666 7668
rect 666 7616 718 7668
rect 718 7616 720 7668
rect 664 7614 720 7616
rect 1184 8322 1240 8324
rect 1184 8270 1186 8322
rect 1186 8270 1238 8322
rect 1238 8270 1240 8322
rect 1184 8268 1240 8270
rect 1184 8104 1240 8106
rect 1184 8052 1186 8104
rect 1186 8052 1238 8104
rect 1238 8052 1240 8104
rect 1184 8050 1240 8052
rect 1184 7886 1240 7888
rect 1184 7834 1186 7886
rect 1186 7834 1238 7886
rect 1238 7834 1240 7886
rect 1184 7832 1240 7834
rect 1184 7668 1240 7670
rect 1184 7616 1186 7668
rect 1186 7616 1238 7668
rect 1238 7616 1240 7668
rect 1184 7614 1240 7616
rect 677 6784 733 6786
rect 677 6732 679 6784
rect 679 6732 731 6784
rect 731 6732 733 6784
rect 677 6730 733 6732
rect 677 6567 733 6569
rect 677 6515 679 6567
rect 679 6515 731 6567
rect 731 6515 733 6567
rect 677 6513 733 6515
rect 677 6349 733 6351
rect 677 6297 679 6349
rect 679 6297 731 6349
rect 731 6297 733 6349
rect 677 6295 733 6297
rect 677 6131 733 6133
rect 677 6079 679 6131
rect 679 6079 731 6131
rect 731 6079 733 6131
rect 677 6077 733 6079
rect 677 5913 733 5915
rect 677 5861 679 5913
rect 679 5861 731 5913
rect 731 5861 733 5913
rect 677 5859 733 5861
rect 677 5696 733 5698
rect 677 5644 679 5696
rect 679 5644 731 5696
rect 731 5644 733 5696
rect 677 5642 733 5644
rect 1191 6784 1247 6786
rect 1191 6732 1193 6784
rect 1193 6732 1245 6784
rect 1245 6732 1247 6784
rect 1191 6730 1247 6732
rect 1191 6567 1247 6569
rect 1191 6515 1193 6567
rect 1193 6515 1245 6567
rect 1245 6515 1247 6567
rect 1191 6513 1247 6515
rect 1191 6349 1247 6351
rect 1191 6297 1193 6349
rect 1193 6297 1245 6349
rect 1245 6297 1247 6349
rect 1191 6295 1247 6297
rect 1191 6131 1247 6133
rect 1191 6079 1193 6131
rect 1193 6079 1245 6131
rect 1245 6079 1247 6131
rect 1191 6077 1247 6079
rect 1191 5913 1247 5915
rect 1191 5861 1193 5913
rect 1193 5861 1245 5913
rect 1245 5861 1247 5913
rect 1191 5859 1247 5861
rect 1191 5696 1247 5698
rect 1191 5644 1193 5696
rect 1193 5644 1245 5696
rect 1245 5644 1247 5696
rect 1191 5642 1247 5644
rect 1670 4177 1726 4233
rect 1180 3701 1236 3757
rect 1670 3959 1726 4015
rect 1180 3483 1236 3539
<< metal3 >>
rect -1 8324 1824 8427
rect -1 8268 457 8324
rect 513 8268 664 8324
rect 720 8268 1184 8324
rect 1240 8268 1824 8324
rect -1 8106 1824 8268
rect -1 8050 457 8106
rect 513 8050 664 8106
rect 720 8050 1184 8106
rect 1240 8050 1824 8106
rect -1 7888 1824 8050
rect -1 7832 457 7888
rect 513 7832 664 7888
rect 720 7832 1184 7888
rect 1240 7832 1824 7888
rect -1 7670 1824 7832
rect -1 7614 457 7670
rect 513 7614 664 7670
rect 720 7614 1184 7670
rect 1240 7614 1824 7670
rect -1 7519 1824 7614
rect -1 6786 1685 7181
rect -1 6730 677 6786
rect 733 6730 1191 6786
rect 1247 6730 1685 6786
rect -1 6569 1685 6730
rect -1 6513 677 6569
rect 733 6513 1191 6569
rect 1247 6513 1685 6569
rect -1 6351 1685 6513
rect -1 6295 677 6351
rect 733 6295 1191 6351
rect 1247 6295 1685 6351
rect -1 6133 1685 6295
rect -1 6077 677 6133
rect 733 6077 1191 6133
rect 1247 6077 1685 6133
rect -1 5915 1685 6077
rect -1 5859 677 5915
rect 733 5859 1191 5915
rect 1247 5859 1685 5915
rect -1 5698 1685 5859
rect -1 5642 677 5698
rect 733 5642 1191 5698
rect 1247 5642 1685 5698
rect -1 4458 1685 5642
rect 1635 4233 1761 4272
rect 1635 4177 1670 4233
rect 1726 4177 1761 4233
rect 1635 4163 1761 4177
rect 6 4030 1762 4163
rect 1635 4015 1761 4030
rect 1635 3959 1670 4015
rect 1726 3959 1761 4015
rect 1635 3920 1761 3959
rect 14 3757 1815 3796
rect 14 3701 1180 3757
rect 1236 3701 1815 3757
rect 14 3663 1815 3701
rect 1144 3662 1272 3663
rect 1145 3539 1271 3662
rect 1145 3483 1180 3539
rect 1236 3483 1271 3539
rect 1145 3444 1271 3483
use M1_NWELL10_512x8m81  M1_NWELL10_512x8m81_0
timestamp 1669390400
transform 1 0 334 0 1 5142
box -221 -1615 221 1615
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_0
timestamp 1669390400
transform 1 0 1151 0 1 7073
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_1
timestamp 1669390400
transform 1 0 641 0 1 7073
box 0 0 1 1
use M1_PSUB$$47335468_512x8m81  M1_PSUB$$47335468_512x8m81_0
timestamp 1669390400
transform 1 0 395 0 1 7910
box -79 -572 80 572
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1669390400
transform 1 0 591 0 1 7073
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 1489
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1669390400
transform 1 0 922 0 1 3852
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1669390400
transform 1 0 1436 0 1 3852
box 0 0 1 1
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 6214
box 0 0 1 1
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_1
timestamp 1669390400
transform 1 0 705 0 1 6214
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7969
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7969
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7969
box 0 0 1 1
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1669390400
transform 1 0 1698 0 1 4096
box 0 0 1 1
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1669390400
transform 1 0 1208 0 1 3620
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7969
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7969
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7969
box 0 0 1 1
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 6214
box 0 0 1 1
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_1
timestamp 1669390400
transform 1 0 705 0 1 6214
box 0 0 1 1
use alatch_512x8m81  alatch_512x8m81_0
timestamp 1669390400
transform 1 0 70 0 1 -632
box -90 -1 1692 2968
use nmos_1p2$$47336492_512x8m81  nmos_1p2$$47336492_512x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 7214
box -119 -74 177 1388
use nmos_1p2$$47336492_512x8m81  nmos_1p2$$47336492_512x8m81_1
timestamp 1669390400
transform 1 0 782 0 1 7214
box -119 -74 177 1388
use pmos_1p2$$47337516_512x8m81  pmos_1p2$$47337516_512x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 3668
box -286 -141 344 3406
use pmos_1p2$$47337516_512x8m81  pmos_1p2$$47337516_512x8m81_1
timestamp 1669390400
transform 1 0 782 0 1 3668
box -286 -141 344 3406
<< properties >>
string GDS_END 523012
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 520338
<< end >>
