magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 1316 88 1388
rect -31 -74 88 -1
use nmos_5p04310590548775_128x8m81  nmos_5p04310590548775_128x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 1360
<< properties >>
string GDS_END 269514
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 269264
<< end >>
