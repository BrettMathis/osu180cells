magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -2884 1125 2884 1144
rect -2884 1079 -2865 1125
rect -2819 1079 -2749 1125
rect -2703 1079 -2633 1125
rect -2587 1079 -2517 1125
rect -2471 1079 -2401 1125
rect -2355 1079 -2285 1125
rect -2239 1079 -2169 1125
rect -2123 1079 -2053 1125
rect -2007 1079 -1937 1125
rect -1891 1079 -1821 1125
rect -1775 1079 -1705 1125
rect -1659 1079 -1589 1125
rect -1543 1079 -1473 1125
rect -1427 1079 -1357 1125
rect -1311 1079 -1241 1125
rect -1195 1079 -1125 1125
rect -1079 1079 -1009 1125
rect -963 1079 -893 1125
rect -847 1079 -777 1125
rect -731 1079 -661 1125
rect -615 1079 -545 1125
rect -499 1079 -429 1125
rect -383 1079 -313 1125
rect -267 1079 -197 1125
rect -151 1079 -81 1125
rect -35 1079 35 1125
rect 81 1079 151 1125
rect 197 1079 267 1125
rect 313 1079 383 1125
rect 429 1079 499 1125
rect 545 1079 615 1125
rect 661 1079 731 1125
rect 777 1079 847 1125
rect 893 1079 963 1125
rect 1009 1079 1079 1125
rect 1125 1079 1195 1125
rect 1241 1079 1311 1125
rect 1357 1079 1427 1125
rect 1473 1079 1543 1125
rect 1589 1079 1659 1125
rect 1705 1079 1775 1125
rect 1821 1079 1891 1125
rect 1937 1079 2007 1125
rect 2053 1079 2123 1125
rect 2169 1079 2239 1125
rect 2285 1079 2355 1125
rect 2401 1079 2471 1125
rect 2517 1079 2587 1125
rect 2633 1079 2703 1125
rect 2749 1079 2819 1125
rect 2865 1079 2884 1125
rect -2884 1009 2884 1079
rect -2884 963 -2865 1009
rect -2819 963 -2749 1009
rect -2703 963 -2633 1009
rect -2587 963 -2517 1009
rect -2471 963 -2401 1009
rect -2355 963 -2285 1009
rect -2239 963 -2169 1009
rect -2123 963 -2053 1009
rect -2007 963 -1937 1009
rect -1891 963 -1821 1009
rect -1775 963 -1705 1009
rect -1659 963 -1589 1009
rect -1543 963 -1473 1009
rect -1427 963 -1357 1009
rect -1311 963 -1241 1009
rect -1195 963 -1125 1009
rect -1079 963 -1009 1009
rect -963 963 -893 1009
rect -847 963 -777 1009
rect -731 963 -661 1009
rect -615 963 -545 1009
rect -499 963 -429 1009
rect -383 963 -313 1009
rect -267 963 -197 1009
rect -151 963 -81 1009
rect -35 963 35 1009
rect 81 963 151 1009
rect 197 963 267 1009
rect 313 963 383 1009
rect 429 963 499 1009
rect 545 963 615 1009
rect 661 963 731 1009
rect 777 963 847 1009
rect 893 963 963 1009
rect 1009 963 1079 1009
rect 1125 963 1195 1009
rect 1241 963 1311 1009
rect 1357 963 1427 1009
rect 1473 963 1543 1009
rect 1589 963 1659 1009
rect 1705 963 1775 1009
rect 1821 963 1891 1009
rect 1937 963 2007 1009
rect 2053 963 2123 1009
rect 2169 963 2239 1009
rect 2285 963 2355 1009
rect 2401 963 2471 1009
rect 2517 963 2587 1009
rect 2633 963 2703 1009
rect 2749 963 2819 1009
rect 2865 963 2884 1009
rect -2884 893 2884 963
rect -2884 847 -2865 893
rect -2819 847 -2749 893
rect -2703 847 -2633 893
rect -2587 847 -2517 893
rect -2471 847 -2401 893
rect -2355 847 -2285 893
rect -2239 847 -2169 893
rect -2123 847 -2053 893
rect -2007 847 -1937 893
rect -1891 847 -1821 893
rect -1775 847 -1705 893
rect -1659 847 -1589 893
rect -1543 847 -1473 893
rect -1427 847 -1357 893
rect -1311 847 -1241 893
rect -1195 847 -1125 893
rect -1079 847 -1009 893
rect -963 847 -893 893
rect -847 847 -777 893
rect -731 847 -661 893
rect -615 847 -545 893
rect -499 847 -429 893
rect -383 847 -313 893
rect -267 847 -197 893
rect -151 847 -81 893
rect -35 847 35 893
rect 81 847 151 893
rect 197 847 267 893
rect 313 847 383 893
rect 429 847 499 893
rect 545 847 615 893
rect 661 847 731 893
rect 777 847 847 893
rect 893 847 963 893
rect 1009 847 1079 893
rect 1125 847 1195 893
rect 1241 847 1311 893
rect 1357 847 1427 893
rect 1473 847 1543 893
rect 1589 847 1659 893
rect 1705 847 1775 893
rect 1821 847 1891 893
rect 1937 847 2007 893
rect 2053 847 2123 893
rect 2169 847 2239 893
rect 2285 847 2355 893
rect 2401 847 2471 893
rect 2517 847 2587 893
rect 2633 847 2703 893
rect 2749 847 2819 893
rect 2865 847 2884 893
rect -2884 777 2884 847
rect -2884 731 -2865 777
rect -2819 731 -2749 777
rect -2703 731 -2633 777
rect -2587 731 -2517 777
rect -2471 731 -2401 777
rect -2355 731 -2285 777
rect -2239 731 -2169 777
rect -2123 731 -2053 777
rect -2007 731 -1937 777
rect -1891 731 -1821 777
rect -1775 731 -1705 777
rect -1659 731 -1589 777
rect -1543 731 -1473 777
rect -1427 731 -1357 777
rect -1311 731 -1241 777
rect -1195 731 -1125 777
rect -1079 731 -1009 777
rect -963 731 -893 777
rect -847 731 -777 777
rect -731 731 -661 777
rect -615 731 -545 777
rect -499 731 -429 777
rect -383 731 -313 777
rect -267 731 -197 777
rect -151 731 -81 777
rect -35 731 35 777
rect 81 731 151 777
rect 197 731 267 777
rect 313 731 383 777
rect 429 731 499 777
rect 545 731 615 777
rect 661 731 731 777
rect 777 731 847 777
rect 893 731 963 777
rect 1009 731 1079 777
rect 1125 731 1195 777
rect 1241 731 1311 777
rect 1357 731 1427 777
rect 1473 731 1543 777
rect 1589 731 1659 777
rect 1705 731 1775 777
rect 1821 731 1891 777
rect 1937 731 2007 777
rect 2053 731 2123 777
rect 2169 731 2239 777
rect 2285 731 2355 777
rect 2401 731 2471 777
rect 2517 731 2587 777
rect 2633 731 2703 777
rect 2749 731 2819 777
rect 2865 731 2884 777
rect -2884 661 2884 731
rect -2884 615 -2865 661
rect -2819 615 -2749 661
rect -2703 615 -2633 661
rect -2587 615 -2517 661
rect -2471 615 -2401 661
rect -2355 615 -2285 661
rect -2239 615 -2169 661
rect -2123 615 -2053 661
rect -2007 615 -1937 661
rect -1891 615 -1821 661
rect -1775 615 -1705 661
rect -1659 615 -1589 661
rect -1543 615 -1473 661
rect -1427 615 -1357 661
rect -1311 615 -1241 661
rect -1195 615 -1125 661
rect -1079 615 -1009 661
rect -963 615 -893 661
rect -847 615 -777 661
rect -731 615 -661 661
rect -615 615 -545 661
rect -499 615 -429 661
rect -383 615 -313 661
rect -267 615 -197 661
rect -151 615 -81 661
rect -35 615 35 661
rect 81 615 151 661
rect 197 615 267 661
rect 313 615 383 661
rect 429 615 499 661
rect 545 615 615 661
rect 661 615 731 661
rect 777 615 847 661
rect 893 615 963 661
rect 1009 615 1079 661
rect 1125 615 1195 661
rect 1241 615 1311 661
rect 1357 615 1427 661
rect 1473 615 1543 661
rect 1589 615 1659 661
rect 1705 615 1775 661
rect 1821 615 1891 661
rect 1937 615 2007 661
rect 2053 615 2123 661
rect 2169 615 2239 661
rect 2285 615 2355 661
rect 2401 615 2471 661
rect 2517 615 2587 661
rect 2633 615 2703 661
rect 2749 615 2819 661
rect 2865 615 2884 661
rect -2884 545 2884 615
rect -2884 499 -2865 545
rect -2819 499 -2749 545
rect -2703 499 -2633 545
rect -2587 499 -2517 545
rect -2471 499 -2401 545
rect -2355 499 -2285 545
rect -2239 499 -2169 545
rect -2123 499 -2053 545
rect -2007 499 -1937 545
rect -1891 499 -1821 545
rect -1775 499 -1705 545
rect -1659 499 -1589 545
rect -1543 499 -1473 545
rect -1427 499 -1357 545
rect -1311 499 -1241 545
rect -1195 499 -1125 545
rect -1079 499 -1009 545
rect -963 499 -893 545
rect -847 499 -777 545
rect -731 499 -661 545
rect -615 499 -545 545
rect -499 499 -429 545
rect -383 499 -313 545
rect -267 499 -197 545
rect -151 499 -81 545
rect -35 499 35 545
rect 81 499 151 545
rect 197 499 267 545
rect 313 499 383 545
rect 429 499 499 545
rect 545 499 615 545
rect 661 499 731 545
rect 777 499 847 545
rect 893 499 963 545
rect 1009 499 1079 545
rect 1125 499 1195 545
rect 1241 499 1311 545
rect 1357 499 1427 545
rect 1473 499 1543 545
rect 1589 499 1659 545
rect 1705 499 1775 545
rect 1821 499 1891 545
rect 1937 499 2007 545
rect 2053 499 2123 545
rect 2169 499 2239 545
rect 2285 499 2355 545
rect 2401 499 2471 545
rect 2517 499 2587 545
rect 2633 499 2703 545
rect 2749 499 2819 545
rect 2865 499 2884 545
rect -2884 429 2884 499
rect -2884 383 -2865 429
rect -2819 383 -2749 429
rect -2703 383 -2633 429
rect -2587 383 -2517 429
rect -2471 383 -2401 429
rect -2355 383 -2285 429
rect -2239 383 -2169 429
rect -2123 383 -2053 429
rect -2007 383 -1937 429
rect -1891 383 -1821 429
rect -1775 383 -1705 429
rect -1659 383 -1589 429
rect -1543 383 -1473 429
rect -1427 383 -1357 429
rect -1311 383 -1241 429
rect -1195 383 -1125 429
rect -1079 383 -1009 429
rect -963 383 -893 429
rect -847 383 -777 429
rect -731 383 -661 429
rect -615 383 -545 429
rect -499 383 -429 429
rect -383 383 -313 429
rect -267 383 -197 429
rect -151 383 -81 429
rect -35 383 35 429
rect 81 383 151 429
rect 197 383 267 429
rect 313 383 383 429
rect 429 383 499 429
rect 545 383 615 429
rect 661 383 731 429
rect 777 383 847 429
rect 893 383 963 429
rect 1009 383 1079 429
rect 1125 383 1195 429
rect 1241 383 1311 429
rect 1357 383 1427 429
rect 1473 383 1543 429
rect 1589 383 1659 429
rect 1705 383 1775 429
rect 1821 383 1891 429
rect 1937 383 2007 429
rect 2053 383 2123 429
rect 2169 383 2239 429
rect 2285 383 2355 429
rect 2401 383 2471 429
rect 2517 383 2587 429
rect 2633 383 2703 429
rect 2749 383 2819 429
rect 2865 383 2884 429
rect -2884 313 2884 383
rect -2884 267 -2865 313
rect -2819 267 -2749 313
rect -2703 267 -2633 313
rect -2587 267 -2517 313
rect -2471 267 -2401 313
rect -2355 267 -2285 313
rect -2239 267 -2169 313
rect -2123 267 -2053 313
rect -2007 267 -1937 313
rect -1891 267 -1821 313
rect -1775 267 -1705 313
rect -1659 267 -1589 313
rect -1543 267 -1473 313
rect -1427 267 -1357 313
rect -1311 267 -1241 313
rect -1195 267 -1125 313
rect -1079 267 -1009 313
rect -963 267 -893 313
rect -847 267 -777 313
rect -731 267 -661 313
rect -615 267 -545 313
rect -499 267 -429 313
rect -383 267 -313 313
rect -267 267 -197 313
rect -151 267 -81 313
rect -35 267 35 313
rect 81 267 151 313
rect 197 267 267 313
rect 313 267 383 313
rect 429 267 499 313
rect 545 267 615 313
rect 661 267 731 313
rect 777 267 847 313
rect 893 267 963 313
rect 1009 267 1079 313
rect 1125 267 1195 313
rect 1241 267 1311 313
rect 1357 267 1427 313
rect 1473 267 1543 313
rect 1589 267 1659 313
rect 1705 267 1775 313
rect 1821 267 1891 313
rect 1937 267 2007 313
rect 2053 267 2123 313
rect 2169 267 2239 313
rect 2285 267 2355 313
rect 2401 267 2471 313
rect 2517 267 2587 313
rect 2633 267 2703 313
rect 2749 267 2819 313
rect 2865 267 2884 313
rect -2884 197 2884 267
rect -2884 151 -2865 197
rect -2819 151 -2749 197
rect -2703 151 -2633 197
rect -2587 151 -2517 197
rect -2471 151 -2401 197
rect -2355 151 -2285 197
rect -2239 151 -2169 197
rect -2123 151 -2053 197
rect -2007 151 -1937 197
rect -1891 151 -1821 197
rect -1775 151 -1705 197
rect -1659 151 -1589 197
rect -1543 151 -1473 197
rect -1427 151 -1357 197
rect -1311 151 -1241 197
rect -1195 151 -1125 197
rect -1079 151 -1009 197
rect -963 151 -893 197
rect -847 151 -777 197
rect -731 151 -661 197
rect -615 151 -545 197
rect -499 151 -429 197
rect -383 151 -313 197
rect -267 151 -197 197
rect -151 151 -81 197
rect -35 151 35 197
rect 81 151 151 197
rect 197 151 267 197
rect 313 151 383 197
rect 429 151 499 197
rect 545 151 615 197
rect 661 151 731 197
rect 777 151 847 197
rect 893 151 963 197
rect 1009 151 1079 197
rect 1125 151 1195 197
rect 1241 151 1311 197
rect 1357 151 1427 197
rect 1473 151 1543 197
rect 1589 151 1659 197
rect 1705 151 1775 197
rect 1821 151 1891 197
rect 1937 151 2007 197
rect 2053 151 2123 197
rect 2169 151 2239 197
rect 2285 151 2355 197
rect 2401 151 2471 197
rect 2517 151 2587 197
rect 2633 151 2703 197
rect 2749 151 2819 197
rect 2865 151 2884 197
rect -2884 81 2884 151
rect -2884 35 -2865 81
rect -2819 35 -2749 81
rect -2703 35 -2633 81
rect -2587 35 -2517 81
rect -2471 35 -2401 81
rect -2355 35 -2285 81
rect -2239 35 -2169 81
rect -2123 35 -2053 81
rect -2007 35 -1937 81
rect -1891 35 -1821 81
rect -1775 35 -1705 81
rect -1659 35 -1589 81
rect -1543 35 -1473 81
rect -1427 35 -1357 81
rect -1311 35 -1241 81
rect -1195 35 -1125 81
rect -1079 35 -1009 81
rect -963 35 -893 81
rect -847 35 -777 81
rect -731 35 -661 81
rect -615 35 -545 81
rect -499 35 -429 81
rect -383 35 -313 81
rect -267 35 -197 81
rect -151 35 -81 81
rect -35 35 35 81
rect 81 35 151 81
rect 197 35 267 81
rect 313 35 383 81
rect 429 35 499 81
rect 545 35 615 81
rect 661 35 731 81
rect 777 35 847 81
rect 893 35 963 81
rect 1009 35 1079 81
rect 1125 35 1195 81
rect 1241 35 1311 81
rect 1357 35 1427 81
rect 1473 35 1543 81
rect 1589 35 1659 81
rect 1705 35 1775 81
rect 1821 35 1891 81
rect 1937 35 2007 81
rect 2053 35 2123 81
rect 2169 35 2239 81
rect 2285 35 2355 81
rect 2401 35 2471 81
rect 2517 35 2587 81
rect 2633 35 2703 81
rect 2749 35 2819 81
rect 2865 35 2884 81
rect -2884 -35 2884 35
rect -2884 -81 -2865 -35
rect -2819 -81 -2749 -35
rect -2703 -81 -2633 -35
rect -2587 -81 -2517 -35
rect -2471 -81 -2401 -35
rect -2355 -81 -2285 -35
rect -2239 -81 -2169 -35
rect -2123 -81 -2053 -35
rect -2007 -81 -1937 -35
rect -1891 -81 -1821 -35
rect -1775 -81 -1705 -35
rect -1659 -81 -1589 -35
rect -1543 -81 -1473 -35
rect -1427 -81 -1357 -35
rect -1311 -81 -1241 -35
rect -1195 -81 -1125 -35
rect -1079 -81 -1009 -35
rect -963 -81 -893 -35
rect -847 -81 -777 -35
rect -731 -81 -661 -35
rect -615 -81 -545 -35
rect -499 -81 -429 -35
rect -383 -81 -313 -35
rect -267 -81 -197 -35
rect -151 -81 -81 -35
rect -35 -81 35 -35
rect 81 -81 151 -35
rect 197 -81 267 -35
rect 313 -81 383 -35
rect 429 -81 499 -35
rect 545 -81 615 -35
rect 661 -81 731 -35
rect 777 -81 847 -35
rect 893 -81 963 -35
rect 1009 -81 1079 -35
rect 1125 -81 1195 -35
rect 1241 -81 1311 -35
rect 1357 -81 1427 -35
rect 1473 -81 1543 -35
rect 1589 -81 1659 -35
rect 1705 -81 1775 -35
rect 1821 -81 1891 -35
rect 1937 -81 2007 -35
rect 2053 -81 2123 -35
rect 2169 -81 2239 -35
rect 2285 -81 2355 -35
rect 2401 -81 2471 -35
rect 2517 -81 2587 -35
rect 2633 -81 2703 -35
rect 2749 -81 2819 -35
rect 2865 -81 2884 -35
rect -2884 -151 2884 -81
rect -2884 -197 -2865 -151
rect -2819 -197 -2749 -151
rect -2703 -197 -2633 -151
rect -2587 -197 -2517 -151
rect -2471 -197 -2401 -151
rect -2355 -197 -2285 -151
rect -2239 -197 -2169 -151
rect -2123 -197 -2053 -151
rect -2007 -197 -1937 -151
rect -1891 -197 -1821 -151
rect -1775 -197 -1705 -151
rect -1659 -197 -1589 -151
rect -1543 -197 -1473 -151
rect -1427 -197 -1357 -151
rect -1311 -197 -1241 -151
rect -1195 -197 -1125 -151
rect -1079 -197 -1009 -151
rect -963 -197 -893 -151
rect -847 -197 -777 -151
rect -731 -197 -661 -151
rect -615 -197 -545 -151
rect -499 -197 -429 -151
rect -383 -197 -313 -151
rect -267 -197 -197 -151
rect -151 -197 -81 -151
rect -35 -197 35 -151
rect 81 -197 151 -151
rect 197 -197 267 -151
rect 313 -197 383 -151
rect 429 -197 499 -151
rect 545 -197 615 -151
rect 661 -197 731 -151
rect 777 -197 847 -151
rect 893 -197 963 -151
rect 1009 -197 1079 -151
rect 1125 -197 1195 -151
rect 1241 -197 1311 -151
rect 1357 -197 1427 -151
rect 1473 -197 1543 -151
rect 1589 -197 1659 -151
rect 1705 -197 1775 -151
rect 1821 -197 1891 -151
rect 1937 -197 2007 -151
rect 2053 -197 2123 -151
rect 2169 -197 2239 -151
rect 2285 -197 2355 -151
rect 2401 -197 2471 -151
rect 2517 -197 2587 -151
rect 2633 -197 2703 -151
rect 2749 -197 2819 -151
rect 2865 -197 2884 -151
rect -2884 -267 2884 -197
rect -2884 -313 -2865 -267
rect -2819 -313 -2749 -267
rect -2703 -313 -2633 -267
rect -2587 -313 -2517 -267
rect -2471 -313 -2401 -267
rect -2355 -313 -2285 -267
rect -2239 -313 -2169 -267
rect -2123 -313 -2053 -267
rect -2007 -313 -1937 -267
rect -1891 -313 -1821 -267
rect -1775 -313 -1705 -267
rect -1659 -313 -1589 -267
rect -1543 -313 -1473 -267
rect -1427 -313 -1357 -267
rect -1311 -313 -1241 -267
rect -1195 -313 -1125 -267
rect -1079 -313 -1009 -267
rect -963 -313 -893 -267
rect -847 -313 -777 -267
rect -731 -313 -661 -267
rect -615 -313 -545 -267
rect -499 -313 -429 -267
rect -383 -313 -313 -267
rect -267 -313 -197 -267
rect -151 -313 -81 -267
rect -35 -313 35 -267
rect 81 -313 151 -267
rect 197 -313 267 -267
rect 313 -313 383 -267
rect 429 -313 499 -267
rect 545 -313 615 -267
rect 661 -313 731 -267
rect 777 -313 847 -267
rect 893 -313 963 -267
rect 1009 -313 1079 -267
rect 1125 -313 1195 -267
rect 1241 -313 1311 -267
rect 1357 -313 1427 -267
rect 1473 -313 1543 -267
rect 1589 -313 1659 -267
rect 1705 -313 1775 -267
rect 1821 -313 1891 -267
rect 1937 -313 2007 -267
rect 2053 -313 2123 -267
rect 2169 -313 2239 -267
rect 2285 -313 2355 -267
rect 2401 -313 2471 -267
rect 2517 -313 2587 -267
rect 2633 -313 2703 -267
rect 2749 -313 2819 -267
rect 2865 -313 2884 -267
rect -2884 -383 2884 -313
rect -2884 -429 -2865 -383
rect -2819 -429 -2749 -383
rect -2703 -429 -2633 -383
rect -2587 -429 -2517 -383
rect -2471 -429 -2401 -383
rect -2355 -429 -2285 -383
rect -2239 -429 -2169 -383
rect -2123 -429 -2053 -383
rect -2007 -429 -1937 -383
rect -1891 -429 -1821 -383
rect -1775 -429 -1705 -383
rect -1659 -429 -1589 -383
rect -1543 -429 -1473 -383
rect -1427 -429 -1357 -383
rect -1311 -429 -1241 -383
rect -1195 -429 -1125 -383
rect -1079 -429 -1009 -383
rect -963 -429 -893 -383
rect -847 -429 -777 -383
rect -731 -429 -661 -383
rect -615 -429 -545 -383
rect -499 -429 -429 -383
rect -383 -429 -313 -383
rect -267 -429 -197 -383
rect -151 -429 -81 -383
rect -35 -429 35 -383
rect 81 -429 151 -383
rect 197 -429 267 -383
rect 313 -429 383 -383
rect 429 -429 499 -383
rect 545 -429 615 -383
rect 661 -429 731 -383
rect 777 -429 847 -383
rect 893 -429 963 -383
rect 1009 -429 1079 -383
rect 1125 -429 1195 -383
rect 1241 -429 1311 -383
rect 1357 -429 1427 -383
rect 1473 -429 1543 -383
rect 1589 -429 1659 -383
rect 1705 -429 1775 -383
rect 1821 -429 1891 -383
rect 1937 -429 2007 -383
rect 2053 -429 2123 -383
rect 2169 -429 2239 -383
rect 2285 -429 2355 -383
rect 2401 -429 2471 -383
rect 2517 -429 2587 -383
rect 2633 -429 2703 -383
rect 2749 -429 2819 -383
rect 2865 -429 2884 -383
rect -2884 -499 2884 -429
rect -2884 -545 -2865 -499
rect -2819 -545 -2749 -499
rect -2703 -545 -2633 -499
rect -2587 -545 -2517 -499
rect -2471 -545 -2401 -499
rect -2355 -545 -2285 -499
rect -2239 -545 -2169 -499
rect -2123 -545 -2053 -499
rect -2007 -545 -1937 -499
rect -1891 -545 -1821 -499
rect -1775 -545 -1705 -499
rect -1659 -545 -1589 -499
rect -1543 -545 -1473 -499
rect -1427 -545 -1357 -499
rect -1311 -545 -1241 -499
rect -1195 -545 -1125 -499
rect -1079 -545 -1009 -499
rect -963 -545 -893 -499
rect -847 -545 -777 -499
rect -731 -545 -661 -499
rect -615 -545 -545 -499
rect -499 -545 -429 -499
rect -383 -545 -313 -499
rect -267 -545 -197 -499
rect -151 -545 -81 -499
rect -35 -545 35 -499
rect 81 -545 151 -499
rect 197 -545 267 -499
rect 313 -545 383 -499
rect 429 -545 499 -499
rect 545 -545 615 -499
rect 661 -545 731 -499
rect 777 -545 847 -499
rect 893 -545 963 -499
rect 1009 -545 1079 -499
rect 1125 -545 1195 -499
rect 1241 -545 1311 -499
rect 1357 -545 1427 -499
rect 1473 -545 1543 -499
rect 1589 -545 1659 -499
rect 1705 -545 1775 -499
rect 1821 -545 1891 -499
rect 1937 -545 2007 -499
rect 2053 -545 2123 -499
rect 2169 -545 2239 -499
rect 2285 -545 2355 -499
rect 2401 -545 2471 -499
rect 2517 -545 2587 -499
rect 2633 -545 2703 -499
rect 2749 -545 2819 -499
rect 2865 -545 2884 -499
rect -2884 -615 2884 -545
rect -2884 -661 -2865 -615
rect -2819 -661 -2749 -615
rect -2703 -661 -2633 -615
rect -2587 -661 -2517 -615
rect -2471 -661 -2401 -615
rect -2355 -661 -2285 -615
rect -2239 -661 -2169 -615
rect -2123 -661 -2053 -615
rect -2007 -661 -1937 -615
rect -1891 -661 -1821 -615
rect -1775 -661 -1705 -615
rect -1659 -661 -1589 -615
rect -1543 -661 -1473 -615
rect -1427 -661 -1357 -615
rect -1311 -661 -1241 -615
rect -1195 -661 -1125 -615
rect -1079 -661 -1009 -615
rect -963 -661 -893 -615
rect -847 -661 -777 -615
rect -731 -661 -661 -615
rect -615 -661 -545 -615
rect -499 -661 -429 -615
rect -383 -661 -313 -615
rect -267 -661 -197 -615
rect -151 -661 -81 -615
rect -35 -661 35 -615
rect 81 -661 151 -615
rect 197 -661 267 -615
rect 313 -661 383 -615
rect 429 -661 499 -615
rect 545 -661 615 -615
rect 661 -661 731 -615
rect 777 -661 847 -615
rect 893 -661 963 -615
rect 1009 -661 1079 -615
rect 1125 -661 1195 -615
rect 1241 -661 1311 -615
rect 1357 -661 1427 -615
rect 1473 -661 1543 -615
rect 1589 -661 1659 -615
rect 1705 -661 1775 -615
rect 1821 -661 1891 -615
rect 1937 -661 2007 -615
rect 2053 -661 2123 -615
rect 2169 -661 2239 -615
rect 2285 -661 2355 -615
rect 2401 -661 2471 -615
rect 2517 -661 2587 -615
rect 2633 -661 2703 -615
rect 2749 -661 2819 -615
rect 2865 -661 2884 -615
rect -2884 -731 2884 -661
rect -2884 -777 -2865 -731
rect -2819 -777 -2749 -731
rect -2703 -777 -2633 -731
rect -2587 -777 -2517 -731
rect -2471 -777 -2401 -731
rect -2355 -777 -2285 -731
rect -2239 -777 -2169 -731
rect -2123 -777 -2053 -731
rect -2007 -777 -1937 -731
rect -1891 -777 -1821 -731
rect -1775 -777 -1705 -731
rect -1659 -777 -1589 -731
rect -1543 -777 -1473 -731
rect -1427 -777 -1357 -731
rect -1311 -777 -1241 -731
rect -1195 -777 -1125 -731
rect -1079 -777 -1009 -731
rect -963 -777 -893 -731
rect -847 -777 -777 -731
rect -731 -777 -661 -731
rect -615 -777 -545 -731
rect -499 -777 -429 -731
rect -383 -777 -313 -731
rect -267 -777 -197 -731
rect -151 -777 -81 -731
rect -35 -777 35 -731
rect 81 -777 151 -731
rect 197 -777 267 -731
rect 313 -777 383 -731
rect 429 -777 499 -731
rect 545 -777 615 -731
rect 661 -777 731 -731
rect 777 -777 847 -731
rect 893 -777 963 -731
rect 1009 -777 1079 -731
rect 1125 -777 1195 -731
rect 1241 -777 1311 -731
rect 1357 -777 1427 -731
rect 1473 -777 1543 -731
rect 1589 -777 1659 -731
rect 1705 -777 1775 -731
rect 1821 -777 1891 -731
rect 1937 -777 2007 -731
rect 2053 -777 2123 -731
rect 2169 -777 2239 -731
rect 2285 -777 2355 -731
rect 2401 -777 2471 -731
rect 2517 -777 2587 -731
rect 2633 -777 2703 -731
rect 2749 -777 2819 -731
rect 2865 -777 2884 -731
rect -2884 -847 2884 -777
rect -2884 -893 -2865 -847
rect -2819 -893 -2749 -847
rect -2703 -893 -2633 -847
rect -2587 -893 -2517 -847
rect -2471 -893 -2401 -847
rect -2355 -893 -2285 -847
rect -2239 -893 -2169 -847
rect -2123 -893 -2053 -847
rect -2007 -893 -1937 -847
rect -1891 -893 -1821 -847
rect -1775 -893 -1705 -847
rect -1659 -893 -1589 -847
rect -1543 -893 -1473 -847
rect -1427 -893 -1357 -847
rect -1311 -893 -1241 -847
rect -1195 -893 -1125 -847
rect -1079 -893 -1009 -847
rect -963 -893 -893 -847
rect -847 -893 -777 -847
rect -731 -893 -661 -847
rect -615 -893 -545 -847
rect -499 -893 -429 -847
rect -383 -893 -313 -847
rect -267 -893 -197 -847
rect -151 -893 -81 -847
rect -35 -893 35 -847
rect 81 -893 151 -847
rect 197 -893 267 -847
rect 313 -893 383 -847
rect 429 -893 499 -847
rect 545 -893 615 -847
rect 661 -893 731 -847
rect 777 -893 847 -847
rect 893 -893 963 -847
rect 1009 -893 1079 -847
rect 1125 -893 1195 -847
rect 1241 -893 1311 -847
rect 1357 -893 1427 -847
rect 1473 -893 1543 -847
rect 1589 -893 1659 -847
rect 1705 -893 1775 -847
rect 1821 -893 1891 -847
rect 1937 -893 2007 -847
rect 2053 -893 2123 -847
rect 2169 -893 2239 -847
rect 2285 -893 2355 -847
rect 2401 -893 2471 -847
rect 2517 -893 2587 -847
rect 2633 -893 2703 -847
rect 2749 -893 2819 -847
rect 2865 -893 2884 -847
rect -2884 -963 2884 -893
rect -2884 -1009 -2865 -963
rect -2819 -1009 -2749 -963
rect -2703 -1009 -2633 -963
rect -2587 -1009 -2517 -963
rect -2471 -1009 -2401 -963
rect -2355 -1009 -2285 -963
rect -2239 -1009 -2169 -963
rect -2123 -1009 -2053 -963
rect -2007 -1009 -1937 -963
rect -1891 -1009 -1821 -963
rect -1775 -1009 -1705 -963
rect -1659 -1009 -1589 -963
rect -1543 -1009 -1473 -963
rect -1427 -1009 -1357 -963
rect -1311 -1009 -1241 -963
rect -1195 -1009 -1125 -963
rect -1079 -1009 -1009 -963
rect -963 -1009 -893 -963
rect -847 -1009 -777 -963
rect -731 -1009 -661 -963
rect -615 -1009 -545 -963
rect -499 -1009 -429 -963
rect -383 -1009 -313 -963
rect -267 -1009 -197 -963
rect -151 -1009 -81 -963
rect -35 -1009 35 -963
rect 81 -1009 151 -963
rect 197 -1009 267 -963
rect 313 -1009 383 -963
rect 429 -1009 499 -963
rect 545 -1009 615 -963
rect 661 -1009 731 -963
rect 777 -1009 847 -963
rect 893 -1009 963 -963
rect 1009 -1009 1079 -963
rect 1125 -1009 1195 -963
rect 1241 -1009 1311 -963
rect 1357 -1009 1427 -963
rect 1473 -1009 1543 -963
rect 1589 -1009 1659 -963
rect 1705 -1009 1775 -963
rect 1821 -1009 1891 -963
rect 1937 -1009 2007 -963
rect 2053 -1009 2123 -963
rect 2169 -1009 2239 -963
rect 2285 -1009 2355 -963
rect 2401 -1009 2471 -963
rect 2517 -1009 2587 -963
rect 2633 -1009 2703 -963
rect 2749 -1009 2819 -963
rect 2865 -1009 2884 -963
rect -2884 -1079 2884 -1009
rect -2884 -1125 -2865 -1079
rect -2819 -1125 -2749 -1079
rect -2703 -1125 -2633 -1079
rect -2587 -1125 -2517 -1079
rect -2471 -1125 -2401 -1079
rect -2355 -1125 -2285 -1079
rect -2239 -1125 -2169 -1079
rect -2123 -1125 -2053 -1079
rect -2007 -1125 -1937 -1079
rect -1891 -1125 -1821 -1079
rect -1775 -1125 -1705 -1079
rect -1659 -1125 -1589 -1079
rect -1543 -1125 -1473 -1079
rect -1427 -1125 -1357 -1079
rect -1311 -1125 -1241 -1079
rect -1195 -1125 -1125 -1079
rect -1079 -1125 -1009 -1079
rect -963 -1125 -893 -1079
rect -847 -1125 -777 -1079
rect -731 -1125 -661 -1079
rect -615 -1125 -545 -1079
rect -499 -1125 -429 -1079
rect -383 -1125 -313 -1079
rect -267 -1125 -197 -1079
rect -151 -1125 -81 -1079
rect -35 -1125 35 -1079
rect 81 -1125 151 -1079
rect 197 -1125 267 -1079
rect 313 -1125 383 -1079
rect 429 -1125 499 -1079
rect 545 -1125 615 -1079
rect 661 -1125 731 -1079
rect 777 -1125 847 -1079
rect 893 -1125 963 -1079
rect 1009 -1125 1079 -1079
rect 1125 -1125 1195 -1079
rect 1241 -1125 1311 -1079
rect 1357 -1125 1427 -1079
rect 1473 -1125 1543 -1079
rect 1589 -1125 1659 -1079
rect 1705 -1125 1775 -1079
rect 1821 -1125 1891 -1079
rect 1937 -1125 2007 -1079
rect 2053 -1125 2123 -1079
rect 2169 -1125 2239 -1079
rect 2285 -1125 2355 -1079
rect 2401 -1125 2471 -1079
rect 2517 -1125 2587 -1079
rect 2633 -1125 2703 -1079
rect 2749 -1125 2819 -1079
rect 2865 -1125 2884 -1079
rect -2884 -1144 2884 -1125
<< psubdiffcont >>
rect -2865 1079 -2819 1125
rect -2749 1079 -2703 1125
rect -2633 1079 -2587 1125
rect -2517 1079 -2471 1125
rect -2401 1079 -2355 1125
rect -2285 1079 -2239 1125
rect -2169 1079 -2123 1125
rect -2053 1079 -2007 1125
rect -1937 1079 -1891 1125
rect -1821 1079 -1775 1125
rect -1705 1079 -1659 1125
rect -1589 1079 -1543 1125
rect -1473 1079 -1427 1125
rect -1357 1079 -1311 1125
rect -1241 1079 -1195 1125
rect -1125 1079 -1079 1125
rect -1009 1079 -963 1125
rect -893 1079 -847 1125
rect -777 1079 -731 1125
rect -661 1079 -615 1125
rect -545 1079 -499 1125
rect -429 1079 -383 1125
rect -313 1079 -267 1125
rect -197 1079 -151 1125
rect -81 1079 -35 1125
rect 35 1079 81 1125
rect 151 1079 197 1125
rect 267 1079 313 1125
rect 383 1079 429 1125
rect 499 1079 545 1125
rect 615 1079 661 1125
rect 731 1079 777 1125
rect 847 1079 893 1125
rect 963 1079 1009 1125
rect 1079 1079 1125 1125
rect 1195 1079 1241 1125
rect 1311 1079 1357 1125
rect 1427 1079 1473 1125
rect 1543 1079 1589 1125
rect 1659 1079 1705 1125
rect 1775 1079 1821 1125
rect 1891 1079 1937 1125
rect 2007 1079 2053 1125
rect 2123 1079 2169 1125
rect 2239 1079 2285 1125
rect 2355 1079 2401 1125
rect 2471 1079 2517 1125
rect 2587 1079 2633 1125
rect 2703 1079 2749 1125
rect 2819 1079 2865 1125
rect -2865 963 -2819 1009
rect -2749 963 -2703 1009
rect -2633 963 -2587 1009
rect -2517 963 -2471 1009
rect -2401 963 -2355 1009
rect -2285 963 -2239 1009
rect -2169 963 -2123 1009
rect -2053 963 -2007 1009
rect -1937 963 -1891 1009
rect -1821 963 -1775 1009
rect -1705 963 -1659 1009
rect -1589 963 -1543 1009
rect -1473 963 -1427 1009
rect -1357 963 -1311 1009
rect -1241 963 -1195 1009
rect -1125 963 -1079 1009
rect -1009 963 -963 1009
rect -893 963 -847 1009
rect -777 963 -731 1009
rect -661 963 -615 1009
rect -545 963 -499 1009
rect -429 963 -383 1009
rect -313 963 -267 1009
rect -197 963 -151 1009
rect -81 963 -35 1009
rect 35 963 81 1009
rect 151 963 197 1009
rect 267 963 313 1009
rect 383 963 429 1009
rect 499 963 545 1009
rect 615 963 661 1009
rect 731 963 777 1009
rect 847 963 893 1009
rect 963 963 1009 1009
rect 1079 963 1125 1009
rect 1195 963 1241 1009
rect 1311 963 1357 1009
rect 1427 963 1473 1009
rect 1543 963 1589 1009
rect 1659 963 1705 1009
rect 1775 963 1821 1009
rect 1891 963 1937 1009
rect 2007 963 2053 1009
rect 2123 963 2169 1009
rect 2239 963 2285 1009
rect 2355 963 2401 1009
rect 2471 963 2517 1009
rect 2587 963 2633 1009
rect 2703 963 2749 1009
rect 2819 963 2865 1009
rect -2865 847 -2819 893
rect -2749 847 -2703 893
rect -2633 847 -2587 893
rect -2517 847 -2471 893
rect -2401 847 -2355 893
rect -2285 847 -2239 893
rect -2169 847 -2123 893
rect -2053 847 -2007 893
rect -1937 847 -1891 893
rect -1821 847 -1775 893
rect -1705 847 -1659 893
rect -1589 847 -1543 893
rect -1473 847 -1427 893
rect -1357 847 -1311 893
rect -1241 847 -1195 893
rect -1125 847 -1079 893
rect -1009 847 -963 893
rect -893 847 -847 893
rect -777 847 -731 893
rect -661 847 -615 893
rect -545 847 -499 893
rect -429 847 -383 893
rect -313 847 -267 893
rect -197 847 -151 893
rect -81 847 -35 893
rect 35 847 81 893
rect 151 847 197 893
rect 267 847 313 893
rect 383 847 429 893
rect 499 847 545 893
rect 615 847 661 893
rect 731 847 777 893
rect 847 847 893 893
rect 963 847 1009 893
rect 1079 847 1125 893
rect 1195 847 1241 893
rect 1311 847 1357 893
rect 1427 847 1473 893
rect 1543 847 1589 893
rect 1659 847 1705 893
rect 1775 847 1821 893
rect 1891 847 1937 893
rect 2007 847 2053 893
rect 2123 847 2169 893
rect 2239 847 2285 893
rect 2355 847 2401 893
rect 2471 847 2517 893
rect 2587 847 2633 893
rect 2703 847 2749 893
rect 2819 847 2865 893
rect -2865 731 -2819 777
rect -2749 731 -2703 777
rect -2633 731 -2587 777
rect -2517 731 -2471 777
rect -2401 731 -2355 777
rect -2285 731 -2239 777
rect -2169 731 -2123 777
rect -2053 731 -2007 777
rect -1937 731 -1891 777
rect -1821 731 -1775 777
rect -1705 731 -1659 777
rect -1589 731 -1543 777
rect -1473 731 -1427 777
rect -1357 731 -1311 777
rect -1241 731 -1195 777
rect -1125 731 -1079 777
rect -1009 731 -963 777
rect -893 731 -847 777
rect -777 731 -731 777
rect -661 731 -615 777
rect -545 731 -499 777
rect -429 731 -383 777
rect -313 731 -267 777
rect -197 731 -151 777
rect -81 731 -35 777
rect 35 731 81 777
rect 151 731 197 777
rect 267 731 313 777
rect 383 731 429 777
rect 499 731 545 777
rect 615 731 661 777
rect 731 731 777 777
rect 847 731 893 777
rect 963 731 1009 777
rect 1079 731 1125 777
rect 1195 731 1241 777
rect 1311 731 1357 777
rect 1427 731 1473 777
rect 1543 731 1589 777
rect 1659 731 1705 777
rect 1775 731 1821 777
rect 1891 731 1937 777
rect 2007 731 2053 777
rect 2123 731 2169 777
rect 2239 731 2285 777
rect 2355 731 2401 777
rect 2471 731 2517 777
rect 2587 731 2633 777
rect 2703 731 2749 777
rect 2819 731 2865 777
rect -2865 615 -2819 661
rect -2749 615 -2703 661
rect -2633 615 -2587 661
rect -2517 615 -2471 661
rect -2401 615 -2355 661
rect -2285 615 -2239 661
rect -2169 615 -2123 661
rect -2053 615 -2007 661
rect -1937 615 -1891 661
rect -1821 615 -1775 661
rect -1705 615 -1659 661
rect -1589 615 -1543 661
rect -1473 615 -1427 661
rect -1357 615 -1311 661
rect -1241 615 -1195 661
rect -1125 615 -1079 661
rect -1009 615 -963 661
rect -893 615 -847 661
rect -777 615 -731 661
rect -661 615 -615 661
rect -545 615 -499 661
rect -429 615 -383 661
rect -313 615 -267 661
rect -197 615 -151 661
rect -81 615 -35 661
rect 35 615 81 661
rect 151 615 197 661
rect 267 615 313 661
rect 383 615 429 661
rect 499 615 545 661
rect 615 615 661 661
rect 731 615 777 661
rect 847 615 893 661
rect 963 615 1009 661
rect 1079 615 1125 661
rect 1195 615 1241 661
rect 1311 615 1357 661
rect 1427 615 1473 661
rect 1543 615 1589 661
rect 1659 615 1705 661
rect 1775 615 1821 661
rect 1891 615 1937 661
rect 2007 615 2053 661
rect 2123 615 2169 661
rect 2239 615 2285 661
rect 2355 615 2401 661
rect 2471 615 2517 661
rect 2587 615 2633 661
rect 2703 615 2749 661
rect 2819 615 2865 661
rect -2865 499 -2819 545
rect -2749 499 -2703 545
rect -2633 499 -2587 545
rect -2517 499 -2471 545
rect -2401 499 -2355 545
rect -2285 499 -2239 545
rect -2169 499 -2123 545
rect -2053 499 -2007 545
rect -1937 499 -1891 545
rect -1821 499 -1775 545
rect -1705 499 -1659 545
rect -1589 499 -1543 545
rect -1473 499 -1427 545
rect -1357 499 -1311 545
rect -1241 499 -1195 545
rect -1125 499 -1079 545
rect -1009 499 -963 545
rect -893 499 -847 545
rect -777 499 -731 545
rect -661 499 -615 545
rect -545 499 -499 545
rect -429 499 -383 545
rect -313 499 -267 545
rect -197 499 -151 545
rect -81 499 -35 545
rect 35 499 81 545
rect 151 499 197 545
rect 267 499 313 545
rect 383 499 429 545
rect 499 499 545 545
rect 615 499 661 545
rect 731 499 777 545
rect 847 499 893 545
rect 963 499 1009 545
rect 1079 499 1125 545
rect 1195 499 1241 545
rect 1311 499 1357 545
rect 1427 499 1473 545
rect 1543 499 1589 545
rect 1659 499 1705 545
rect 1775 499 1821 545
rect 1891 499 1937 545
rect 2007 499 2053 545
rect 2123 499 2169 545
rect 2239 499 2285 545
rect 2355 499 2401 545
rect 2471 499 2517 545
rect 2587 499 2633 545
rect 2703 499 2749 545
rect 2819 499 2865 545
rect -2865 383 -2819 429
rect -2749 383 -2703 429
rect -2633 383 -2587 429
rect -2517 383 -2471 429
rect -2401 383 -2355 429
rect -2285 383 -2239 429
rect -2169 383 -2123 429
rect -2053 383 -2007 429
rect -1937 383 -1891 429
rect -1821 383 -1775 429
rect -1705 383 -1659 429
rect -1589 383 -1543 429
rect -1473 383 -1427 429
rect -1357 383 -1311 429
rect -1241 383 -1195 429
rect -1125 383 -1079 429
rect -1009 383 -963 429
rect -893 383 -847 429
rect -777 383 -731 429
rect -661 383 -615 429
rect -545 383 -499 429
rect -429 383 -383 429
rect -313 383 -267 429
rect -197 383 -151 429
rect -81 383 -35 429
rect 35 383 81 429
rect 151 383 197 429
rect 267 383 313 429
rect 383 383 429 429
rect 499 383 545 429
rect 615 383 661 429
rect 731 383 777 429
rect 847 383 893 429
rect 963 383 1009 429
rect 1079 383 1125 429
rect 1195 383 1241 429
rect 1311 383 1357 429
rect 1427 383 1473 429
rect 1543 383 1589 429
rect 1659 383 1705 429
rect 1775 383 1821 429
rect 1891 383 1937 429
rect 2007 383 2053 429
rect 2123 383 2169 429
rect 2239 383 2285 429
rect 2355 383 2401 429
rect 2471 383 2517 429
rect 2587 383 2633 429
rect 2703 383 2749 429
rect 2819 383 2865 429
rect -2865 267 -2819 313
rect -2749 267 -2703 313
rect -2633 267 -2587 313
rect -2517 267 -2471 313
rect -2401 267 -2355 313
rect -2285 267 -2239 313
rect -2169 267 -2123 313
rect -2053 267 -2007 313
rect -1937 267 -1891 313
rect -1821 267 -1775 313
rect -1705 267 -1659 313
rect -1589 267 -1543 313
rect -1473 267 -1427 313
rect -1357 267 -1311 313
rect -1241 267 -1195 313
rect -1125 267 -1079 313
rect -1009 267 -963 313
rect -893 267 -847 313
rect -777 267 -731 313
rect -661 267 -615 313
rect -545 267 -499 313
rect -429 267 -383 313
rect -313 267 -267 313
rect -197 267 -151 313
rect -81 267 -35 313
rect 35 267 81 313
rect 151 267 197 313
rect 267 267 313 313
rect 383 267 429 313
rect 499 267 545 313
rect 615 267 661 313
rect 731 267 777 313
rect 847 267 893 313
rect 963 267 1009 313
rect 1079 267 1125 313
rect 1195 267 1241 313
rect 1311 267 1357 313
rect 1427 267 1473 313
rect 1543 267 1589 313
rect 1659 267 1705 313
rect 1775 267 1821 313
rect 1891 267 1937 313
rect 2007 267 2053 313
rect 2123 267 2169 313
rect 2239 267 2285 313
rect 2355 267 2401 313
rect 2471 267 2517 313
rect 2587 267 2633 313
rect 2703 267 2749 313
rect 2819 267 2865 313
rect -2865 151 -2819 197
rect -2749 151 -2703 197
rect -2633 151 -2587 197
rect -2517 151 -2471 197
rect -2401 151 -2355 197
rect -2285 151 -2239 197
rect -2169 151 -2123 197
rect -2053 151 -2007 197
rect -1937 151 -1891 197
rect -1821 151 -1775 197
rect -1705 151 -1659 197
rect -1589 151 -1543 197
rect -1473 151 -1427 197
rect -1357 151 -1311 197
rect -1241 151 -1195 197
rect -1125 151 -1079 197
rect -1009 151 -963 197
rect -893 151 -847 197
rect -777 151 -731 197
rect -661 151 -615 197
rect -545 151 -499 197
rect -429 151 -383 197
rect -313 151 -267 197
rect -197 151 -151 197
rect -81 151 -35 197
rect 35 151 81 197
rect 151 151 197 197
rect 267 151 313 197
rect 383 151 429 197
rect 499 151 545 197
rect 615 151 661 197
rect 731 151 777 197
rect 847 151 893 197
rect 963 151 1009 197
rect 1079 151 1125 197
rect 1195 151 1241 197
rect 1311 151 1357 197
rect 1427 151 1473 197
rect 1543 151 1589 197
rect 1659 151 1705 197
rect 1775 151 1821 197
rect 1891 151 1937 197
rect 2007 151 2053 197
rect 2123 151 2169 197
rect 2239 151 2285 197
rect 2355 151 2401 197
rect 2471 151 2517 197
rect 2587 151 2633 197
rect 2703 151 2749 197
rect 2819 151 2865 197
rect -2865 35 -2819 81
rect -2749 35 -2703 81
rect -2633 35 -2587 81
rect -2517 35 -2471 81
rect -2401 35 -2355 81
rect -2285 35 -2239 81
rect -2169 35 -2123 81
rect -2053 35 -2007 81
rect -1937 35 -1891 81
rect -1821 35 -1775 81
rect -1705 35 -1659 81
rect -1589 35 -1543 81
rect -1473 35 -1427 81
rect -1357 35 -1311 81
rect -1241 35 -1195 81
rect -1125 35 -1079 81
rect -1009 35 -963 81
rect -893 35 -847 81
rect -777 35 -731 81
rect -661 35 -615 81
rect -545 35 -499 81
rect -429 35 -383 81
rect -313 35 -267 81
rect -197 35 -151 81
rect -81 35 -35 81
rect 35 35 81 81
rect 151 35 197 81
rect 267 35 313 81
rect 383 35 429 81
rect 499 35 545 81
rect 615 35 661 81
rect 731 35 777 81
rect 847 35 893 81
rect 963 35 1009 81
rect 1079 35 1125 81
rect 1195 35 1241 81
rect 1311 35 1357 81
rect 1427 35 1473 81
rect 1543 35 1589 81
rect 1659 35 1705 81
rect 1775 35 1821 81
rect 1891 35 1937 81
rect 2007 35 2053 81
rect 2123 35 2169 81
rect 2239 35 2285 81
rect 2355 35 2401 81
rect 2471 35 2517 81
rect 2587 35 2633 81
rect 2703 35 2749 81
rect 2819 35 2865 81
rect -2865 -81 -2819 -35
rect -2749 -81 -2703 -35
rect -2633 -81 -2587 -35
rect -2517 -81 -2471 -35
rect -2401 -81 -2355 -35
rect -2285 -81 -2239 -35
rect -2169 -81 -2123 -35
rect -2053 -81 -2007 -35
rect -1937 -81 -1891 -35
rect -1821 -81 -1775 -35
rect -1705 -81 -1659 -35
rect -1589 -81 -1543 -35
rect -1473 -81 -1427 -35
rect -1357 -81 -1311 -35
rect -1241 -81 -1195 -35
rect -1125 -81 -1079 -35
rect -1009 -81 -963 -35
rect -893 -81 -847 -35
rect -777 -81 -731 -35
rect -661 -81 -615 -35
rect -545 -81 -499 -35
rect -429 -81 -383 -35
rect -313 -81 -267 -35
rect -197 -81 -151 -35
rect -81 -81 -35 -35
rect 35 -81 81 -35
rect 151 -81 197 -35
rect 267 -81 313 -35
rect 383 -81 429 -35
rect 499 -81 545 -35
rect 615 -81 661 -35
rect 731 -81 777 -35
rect 847 -81 893 -35
rect 963 -81 1009 -35
rect 1079 -81 1125 -35
rect 1195 -81 1241 -35
rect 1311 -81 1357 -35
rect 1427 -81 1473 -35
rect 1543 -81 1589 -35
rect 1659 -81 1705 -35
rect 1775 -81 1821 -35
rect 1891 -81 1937 -35
rect 2007 -81 2053 -35
rect 2123 -81 2169 -35
rect 2239 -81 2285 -35
rect 2355 -81 2401 -35
rect 2471 -81 2517 -35
rect 2587 -81 2633 -35
rect 2703 -81 2749 -35
rect 2819 -81 2865 -35
rect -2865 -197 -2819 -151
rect -2749 -197 -2703 -151
rect -2633 -197 -2587 -151
rect -2517 -197 -2471 -151
rect -2401 -197 -2355 -151
rect -2285 -197 -2239 -151
rect -2169 -197 -2123 -151
rect -2053 -197 -2007 -151
rect -1937 -197 -1891 -151
rect -1821 -197 -1775 -151
rect -1705 -197 -1659 -151
rect -1589 -197 -1543 -151
rect -1473 -197 -1427 -151
rect -1357 -197 -1311 -151
rect -1241 -197 -1195 -151
rect -1125 -197 -1079 -151
rect -1009 -197 -963 -151
rect -893 -197 -847 -151
rect -777 -197 -731 -151
rect -661 -197 -615 -151
rect -545 -197 -499 -151
rect -429 -197 -383 -151
rect -313 -197 -267 -151
rect -197 -197 -151 -151
rect -81 -197 -35 -151
rect 35 -197 81 -151
rect 151 -197 197 -151
rect 267 -197 313 -151
rect 383 -197 429 -151
rect 499 -197 545 -151
rect 615 -197 661 -151
rect 731 -197 777 -151
rect 847 -197 893 -151
rect 963 -197 1009 -151
rect 1079 -197 1125 -151
rect 1195 -197 1241 -151
rect 1311 -197 1357 -151
rect 1427 -197 1473 -151
rect 1543 -197 1589 -151
rect 1659 -197 1705 -151
rect 1775 -197 1821 -151
rect 1891 -197 1937 -151
rect 2007 -197 2053 -151
rect 2123 -197 2169 -151
rect 2239 -197 2285 -151
rect 2355 -197 2401 -151
rect 2471 -197 2517 -151
rect 2587 -197 2633 -151
rect 2703 -197 2749 -151
rect 2819 -197 2865 -151
rect -2865 -313 -2819 -267
rect -2749 -313 -2703 -267
rect -2633 -313 -2587 -267
rect -2517 -313 -2471 -267
rect -2401 -313 -2355 -267
rect -2285 -313 -2239 -267
rect -2169 -313 -2123 -267
rect -2053 -313 -2007 -267
rect -1937 -313 -1891 -267
rect -1821 -313 -1775 -267
rect -1705 -313 -1659 -267
rect -1589 -313 -1543 -267
rect -1473 -313 -1427 -267
rect -1357 -313 -1311 -267
rect -1241 -313 -1195 -267
rect -1125 -313 -1079 -267
rect -1009 -313 -963 -267
rect -893 -313 -847 -267
rect -777 -313 -731 -267
rect -661 -313 -615 -267
rect -545 -313 -499 -267
rect -429 -313 -383 -267
rect -313 -313 -267 -267
rect -197 -313 -151 -267
rect -81 -313 -35 -267
rect 35 -313 81 -267
rect 151 -313 197 -267
rect 267 -313 313 -267
rect 383 -313 429 -267
rect 499 -313 545 -267
rect 615 -313 661 -267
rect 731 -313 777 -267
rect 847 -313 893 -267
rect 963 -313 1009 -267
rect 1079 -313 1125 -267
rect 1195 -313 1241 -267
rect 1311 -313 1357 -267
rect 1427 -313 1473 -267
rect 1543 -313 1589 -267
rect 1659 -313 1705 -267
rect 1775 -313 1821 -267
rect 1891 -313 1937 -267
rect 2007 -313 2053 -267
rect 2123 -313 2169 -267
rect 2239 -313 2285 -267
rect 2355 -313 2401 -267
rect 2471 -313 2517 -267
rect 2587 -313 2633 -267
rect 2703 -313 2749 -267
rect 2819 -313 2865 -267
rect -2865 -429 -2819 -383
rect -2749 -429 -2703 -383
rect -2633 -429 -2587 -383
rect -2517 -429 -2471 -383
rect -2401 -429 -2355 -383
rect -2285 -429 -2239 -383
rect -2169 -429 -2123 -383
rect -2053 -429 -2007 -383
rect -1937 -429 -1891 -383
rect -1821 -429 -1775 -383
rect -1705 -429 -1659 -383
rect -1589 -429 -1543 -383
rect -1473 -429 -1427 -383
rect -1357 -429 -1311 -383
rect -1241 -429 -1195 -383
rect -1125 -429 -1079 -383
rect -1009 -429 -963 -383
rect -893 -429 -847 -383
rect -777 -429 -731 -383
rect -661 -429 -615 -383
rect -545 -429 -499 -383
rect -429 -429 -383 -383
rect -313 -429 -267 -383
rect -197 -429 -151 -383
rect -81 -429 -35 -383
rect 35 -429 81 -383
rect 151 -429 197 -383
rect 267 -429 313 -383
rect 383 -429 429 -383
rect 499 -429 545 -383
rect 615 -429 661 -383
rect 731 -429 777 -383
rect 847 -429 893 -383
rect 963 -429 1009 -383
rect 1079 -429 1125 -383
rect 1195 -429 1241 -383
rect 1311 -429 1357 -383
rect 1427 -429 1473 -383
rect 1543 -429 1589 -383
rect 1659 -429 1705 -383
rect 1775 -429 1821 -383
rect 1891 -429 1937 -383
rect 2007 -429 2053 -383
rect 2123 -429 2169 -383
rect 2239 -429 2285 -383
rect 2355 -429 2401 -383
rect 2471 -429 2517 -383
rect 2587 -429 2633 -383
rect 2703 -429 2749 -383
rect 2819 -429 2865 -383
rect -2865 -545 -2819 -499
rect -2749 -545 -2703 -499
rect -2633 -545 -2587 -499
rect -2517 -545 -2471 -499
rect -2401 -545 -2355 -499
rect -2285 -545 -2239 -499
rect -2169 -545 -2123 -499
rect -2053 -545 -2007 -499
rect -1937 -545 -1891 -499
rect -1821 -545 -1775 -499
rect -1705 -545 -1659 -499
rect -1589 -545 -1543 -499
rect -1473 -545 -1427 -499
rect -1357 -545 -1311 -499
rect -1241 -545 -1195 -499
rect -1125 -545 -1079 -499
rect -1009 -545 -963 -499
rect -893 -545 -847 -499
rect -777 -545 -731 -499
rect -661 -545 -615 -499
rect -545 -545 -499 -499
rect -429 -545 -383 -499
rect -313 -545 -267 -499
rect -197 -545 -151 -499
rect -81 -545 -35 -499
rect 35 -545 81 -499
rect 151 -545 197 -499
rect 267 -545 313 -499
rect 383 -545 429 -499
rect 499 -545 545 -499
rect 615 -545 661 -499
rect 731 -545 777 -499
rect 847 -545 893 -499
rect 963 -545 1009 -499
rect 1079 -545 1125 -499
rect 1195 -545 1241 -499
rect 1311 -545 1357 -499
rect 1427 -545 1473 -499
rect 1543 -545 1589 -499
rect 1659 -545 1705 -499
rect 1775 -545 1821 -499
rect 1891 -545 1937 -499
rect 2007 -545 2053 -499
rect 2123 -545 2169 -499
rect 2239 -545 2285 -499
rect 2355 -545 2401 -499
rect 2471 -545 2517 -499
rect 2587 -545 2633 -499
rect 2703 -545 2749 -499
rect 2819 -545 2865 -499
rect -2865 -661 -2819 -615
rect -2749 -661 -2703 -615
rect -2633 -661 -2587 -615
rect -2517 -661 -2471 -615
rect -2401 -661 -2355 -615
rect -2285 -661 -2239 -615
rect -2169 -661 -2123 -615
rect -2053 -661 -2007 -615
rect -1937 -661 -1891 -615
rect -1821 -661 -1775 -615
rect -1705 -661 -1659 -615
rect -1589 -661 -1543 -615
rect -1473 -661 -1427 -615
rect -1357 -661 -1311 -615
rect -1241 -661 -1195 -615
rect -1125 -661 -1079 -615
rect -1009 -661 -963 -615
rect -893 -661 -847 -615
rect -777 -661 -731 -615
rect -661 -661 -615 -615
rect -545 -661 -499 -615
rect -429 -661 -383 -615
rect -313 -661 -267 -615
rect -197 -661 -151 -615
rect -81 -661 -35 -615
rect 35 -661 81 -615
rect 151 -661 197 -615
rect 267 -661 313 -615
rect 383 -661 429 -615
rect 499 -661 545 -615
rect 615 -661 661 -615
rect 731 -661 777 -615
rect 847 -661 893 -615
rect 963 -661 1009 -615
rect 1079 -661 1125 -615
rect 1195 -661 1241 -615
rect 1311 -661 1357 -615
rect 1427 -661 1473 -615
rect 1543 -661 1589 -615
rect 1659 -661 1705 -615
rect 1775 -661 1821 -615
rect 1891 -661 1937 -615
rect 2007 -661 2053 -615
rect 2123 -661 2169 -615
rect 2239 -661 2285 -615
rect 2355 -661 2401 -615
rect 2471 -661 2517 -615
rect 2587 -661 2633 -615
rect 2703 -661 2749 -615
rect 2819 -661 2865 -615
rect -2865 -777 -2819 -731
rect -2749 -777 -2703 -731
rect -2633 -777 -2587 -731
rect -2517 -777 -2471 -731
rect -2401 -777 -2355 -731
rect -2285 -777 -2239 -731
rect -2169 -777 -2123 -731
rect -2053 -777 -2007 -731
rect -1937 -777 -1891 -731
rect -1821 -777 -1775 -731
rect -1705 -777 -1659 -731
rect -1589 -777 -1543 -731
rect -1473 -777 -1427 -731
rect -1357 -777 -1311 -731
rect -1241 -777 -1195 -731
rect -1125 -777 -1079 -731
rect -1009 -777 -963 -731
rect -893 -777 -847 -731
rect -777 -777 -731 -731
rect -661 -777 -615 -731
rect -545 -777 -499 -731
rect -429 -777 -383 -731
rect -313 -777 -267 -731
rect -197 -777 -151 -731
rect -81 -777 -35 -731
rect 35 -777 81 -731
rect 151 -777 197 -731
rect 267 -777 313 -731
rect 383 -777 429 -731
rect 499 -777 545 -731
rect 615 -777 661 -731
rect 731 -777 777 -731
rect 847 -777 893 -731
rect 963 -777 1009 -731
rect 1079 -777 1125 -731
rect 1195 -777 1241 -731
rect 1311 -777 1357 -731
rect 1427 -777 1473 -731
rect 1543 -777 1589 -731
rect 1659 -777 1705 -731
rect 1775 -777 1821 -731
rect 1891 -777 1937 -731
rect 2007 -777 2053 -731
rect 2123 -777 2169 -731
rect 2239 -777 2285 -731
rect 2355 -777 2401 -731
rect 2471 -777 2517 -731
rect 2587 -777 2633 -731
rect 2703 -777 2749 -731
rect 2819 -777 2865 -731
rect -2865 -893 -2819 -847
rect -2749 -893 -2703 -847
rect -2633 -893 -2587 -847
rect -2517 -893 -2471 -847
rect -2401 -893 -2355 -847
rect -2285 -893 -2239 -847
rect -2169 -893 -2123 -847
rect -2053 -893 -2007 -847
rect -1937 -893 -1891 -847
rect -1821 -893 -1775 -847
rect -1705 -893 -1659 -847
rect -1589 -893 -1543 -847
rect -1473 -893 -1427 -847
rect -1357 -893 -1311 -847
rect -1241 -893 -1195 -847
rect -1125 -893 -1079 -847
rect -1009 -893 -963 -847
rect -893 -893 -847 -847
rect -777 -893 -731 -847
rect -661 -893 -615 -847
rect -545 -893 -499 -847
rect -429 -893 -383 -847
rect -313 -893 -267 -847
rect -197 -893 -151 -847
rect -81 -893 -35 -847
rect 35 -893 81 -847
rect 151 -893 197 -847
rect 267 -893 313 -847
rect 383 -893 429 -847
rect 499 -893 545 -847
rect 615 -893 661 -847
rect 731 -893 777 -847
rect 847 -893 893 -847
rect 963 -893 1009 -847
rect 1079 -893 1125 -847
rect 1195 -893 1241 -847
rect 1311 -893 1357 -847
rect 1427 -893 1473 -847
rect 1543 -893 1589 -847
rect 1659 -893 1705 -847
rect 1775 -893 1821 -847
rect 1891 -893 1937 -847
rect 2007 -893 2053 -847
rect 2123 -893 2169 -847
rect 2239 -893 2285 -847
rect 2355 -893 2401 -847
rect 2471 -893 2517 -847
rect 2587 -893 2633 -847
rect 2703 -893 2749 -847
rect 2819 -893 2865 -847
rect -2865 -1009 -2819 -963
rect -2749 -1009 -2703 -963
rect -2633 -1009 -2587 -963
rect -2517 -1009 -2471 -963
rect -2401 -1009 -2355 -963
rect -2285 -1009 -2239 -963
rect -2169 -1009 -2123 -963
rect -2053 -1009 -2007 -963
rect -1937 -1009 -1891 -963
rect -1821 -1009 -1775 -963
rect -1705 -1009 -1659 -963
rect -1589 -1009 -1543 -963
rect -1473 -1009 -1427 -963
rect -1357 -1009 -1311 -963
rect -1241 -1009 -1195 -963
rect -1125 -1009 -1079 -963
rect -1009 -1009 -963 -963
rect -893 -1009 -847 -963
rect -777 -1009 -731 -963
rect -661 -1009 -615 -963
rect -545 -1009 -499 -963
rect -429 -1009 -383 -963
rect -313 -1009 -267 -963
rect -197 -1009 -151 -963
rect -81 -1009 -35 -963
rect 35 -1009 81 -963
rect 151 -1009 197 -963
rect 267 -1009 313 -963
rect 383 -1009 429 -963
rect 499 -1009 545 -963
rect 615 -1009 661 -963
rect 731 -1009 777 -963
rect 847 -1009 893 -963
rect 963 -1009 1009 -963
rect 1079 -1009 1125 -963
rect 1195 -1009 1241 -963
rect 1311 -1009 1357 -963
rect 1427 -1009 1473 -963
rect 1543 -1009 1589 -963
rect 1659 -1009 1705 -963
rect 1775 -1009 1821 -963
rect 1891 -1009 1937 -963
rect 2007 -1009 2053 -963
rect 2123 -1009 2169 -963
rect 2239 -1009 2285 -963
rect 2355 -1009 2401 -963
rect 2471 -1009 2517 -963
rect 2587 -1009 2633 -963
rect 2703 -1009 2749 -963
rect 2819 -1009 2865 -963
rect -2865 -1125 -2819 -1079
rect -2749 -1125 -2703 -1079
rect -2633 -1125 -2587 -1079
rect -2517 -1125 -2471 -1079
rect -2401 -1125 -2355 -1079
rect -2285 -1125 -2239 -1079
rect -2169 -1125 -2123 -1079
rect -2053 -1125 -2007 -1079
rect -1937 -1125 -1891 -1079
rect -1821 -1125 -1775 -1079
rect -1705 -1125 -1659 -1079
rect -1589 -1125 -1543 -1079
rect -1473 -1125 -1427 -1079
rect -1357 -1125 -1311 -1079
rect -1241 -1125 -1195 -1079
rect -1125 -1125 -1079 -1079
rect -1009 -1125 -963 -1079
rect -893 -1125 -847 -1079
rect -777 -1125 -731 -1079
rect -661 -1125 -615 -1079
rect -545 -1125 -499 -1079
rect -429 -1125 -383 -1079
rect -313 -1125 -267 -1079
rect -197 -1125 -151 -1079
rect -81 -1125 -35 -1079
rect 35 -1125 81 -1079
rect 151 -1125 197 -1079
rect 267 -1125 313 -1079
rect 383 -1125 429 -1079
rect 499 -1125 545 -1079
rect 615 -1125 661 -1079
rect 731 -1125 777 -1079
rect 847 -1125 893 -1079
rect 963 -1125 1009 -1079
rect 1079 -1125 1125 -1079
rect 1195 -1125 1241 -1079
rect 1311 -1125 1357 -1079
rect 1427 -1125 1473 -1079
rect 1543 -1125 1589 -1079
rect 1659 -1125 1705 -1079
rect 1775 -1125 1821 -1079
rect 1891 -1125 1937 -1079
rect 2007 -1125 2053 -1079
rect 2123 -1125 2169 -1079
rect 2239 -1125 2285 -1079
rect 2355 -1125 2401 -1079
rect 2471 -1125 2517 -1079
rect 2587 -1125 2633 -1079
rect 2703 -1125 2749 -1079
rect 2819 -1125 2865 -1079
<< metal1 >>
rect -2876 1125 2876 1136
rect -2876 1079 -2865 1125
rect -2819 1079 -2749 1125
rect -2703 1079 -2633 1125
rect -2587 1079 -2517 1125
rect -2471 1079 -2401 1125
rect -2355 1079 -2285 1125
rect -2239 1079 -2169 1125
rect -2123 1079 -2053 1125
rect -2007 1079 -1937 1125
rect -1891 1079 -1821 1125
rect -1775 1079 -1705 1125
rect -1659 1079 -1589 1125
rect -1543 1079 -1473 1125
rect -1427 1079 -1357 1125
rect -1311 1079 -1241 1125
rect -1195 1079 -1125 1125
rect -1079 1079 -1009 1125
rect -963 1079 -893 1125
rect -847 1079 -777 1125
rect -731 1079 -661 1125
rect -615 1079 -545 1125
rect -499 1079 -429 1125
rect -383 1079 -313 1125
rect -267 1079 -197 1125
rect -151 1079 -81 1125
rect -35 1079 35 1125
rect 81 1079 151 1125
rect 197 1079 267 1125
rect 313 1079 383 1125
rect 429 1079 499 1125
rect 545 1079 615 1125
rect 661 1079 731 1125
rect 777 1079 847 1125
rect 893 1079 963 1125
rect 1009 1079 1079 1125
rect 1125 1079 1195 1125
rect 1241 1079 1311 1125
rect 1357 1079 1427 1125
rect 1473 1079 1543 1125
rect 1589 1079 1659 1125
rect 1705 1079 1775 1125
rect 1821 1079 1891 1125
rect 1937 1079 2007 1125
rect 2053 1079 2123 1125
rect 2169 1079 2239 1125
rect 2285 1079 2355 1125
rect 2401 1079 2471 1125
rect 2517 1079 2587 1125
rect 2633 1079 2703 1125
rect 2749 1079 2819 1125
rect 2865 1079 2876 1125
rect -2876 1009 2876 1079
rect -2876 963 -2865 1009
rect -2819 963 -2749 1009
rect -2703 963 -2633 1009
rect -2587 963 -2517 1009
rect -2471 963 -2401 1009
rect -2355 963 -2285 1009
rect -2239 963 -2169 1009
rect -2123 963 -2053 1009
rect -2007 963 -1937 1009
rect -1891 963 -1821 1009
rect -1775 963 -1705 1009
rect -1659 963 -1589 1009
rect -1543 963 -1473 1009
rect -1427 963 -1357 1009
rect -1311 963 -1241 1009
rect -1195 963 -1125 1009
rect -1079 963 -1009 1009
rect -963 963 -893 1009
rect -847 963 -777 1009
rect -731 963 -661 1009
rect -615 963 -545 1009
rect -499 963 -429 1009
rect -383 963 -313 1009
rect -267 963 -197 1009
rect -151 963 -81 1009
rect -35 963 35 1009
rect 81 963 151 1009
rect 197 963 267 1009
rect 313 963 383 1009
rect 429 963 499 1009
rect 545 963 615 1009
rect 661 963 731 1009
rect 777 963 847 1009
rect 893 963 963 1009
rect 1009 963 1079 1009
rect 1125 963 1195 1009
rect 1241 963 1311 1009
rect 1357 963 1427 1009
rect 1473 963 1543 1009
rect 1589 963 1659 1009
rect 1705 963 1775 1009
rect 1821 963 1891 1009
rect 1937 963 2007 1009
rect 2053 963 2123 1009
rect 2169 963 2239 1009
rect 2285 963 2355 1009
rect 2401 963 2471 1009
rect 2517 963 2587 1009
rect 2633 963 2703 1009
rect 2749 963 2819 1009
rect 2865 963 2876 1009
rect -2876 893 2876 963
rect -2876 847 -2865 893
rect -2819 847 -2749 893
rect -2703 847 -2633 893
rect -2587 847 -2517 893
rect -2471 847 -2401 893
rect -2355 847 -2285 893
rect -2239 847 -2169 893
rect -2123 847 -2053 893
rect -2007 847 -1937 893
rect -1891 847 -1821 893
rect -1775 847 -1705 893
rect -1659 847 -1589 893
rect -1543 847 -1473 893
rect -1427 847 -1357 893
rect -1311 847 -1241 893
rect -1195 847 -1125 893
rect -1079 847 -1009 893
rect -963 847 -893 893
rect -847 847 -777 893
rect -731 847 -661 893
rect -615 847 -545 893
rect -499 847 -429 893
rect -383 847 -313 893
rect -267 847 -197 893
rect -151 847 -81 893
rect -35 847 35 893
rect 81 847 151 893
rect 197 847 267 893
rect 313 847 383 893
rect 429 847 499 893
rect 545 847 615 893
rect 661 847 731 893
rect 777 847 847 893
rect 893 847 963 893
rect 1009 847 1079 893
rect 1125 847 1195 893
rect 1241 847 1311 893
rect 1357 847 1427 893
rect 1473 847 1543 893
rect 1589 847 1659 893
rect 1705 847 1775 893
rect 1821 847 1891 893
rect 1937 847 2007 893
rect 2053 847 2123 893
rect 2169 847 2239 893
rect 2285 847 2355 893
rect 2401 847 2471 893
rect 2517 847 2587 893
rect 2633 847 2703 893
rect 2749 847 2819 893
rect 2865 847 2876 893
rect -2876 777 2876 847
rect -2876 731 -2865 777
rect -2819 731 -2749 777
rect -2703 731 -2633 777
rect -2587 731 -2517 777
rect -2471 731 -2401 777
rect -2355 731 -2285 777
rect -2239 731 -2169 777
rect -2123 731 -2053 777
rect -2007 731 -1937 777
rect -1891 731 -1821 777
rect -1775 731 -1705 777
rect -1659 731 -1589 777
rect -1543 731 -1473 777
rect -1427 731 -1357 777
rect -1311 731 -1241 777
rect -1195 731 -1125 777
rect -1079 731 -1009 777
rect -963 731 -893 777
rect -847 731 -777 777
rect -731 731 -661 777
rect -615 731 -545 777
rect -499 731 -429 777
rect -383 731 -313 777
rect -267 731 -197 777
rect -151 731 -81 777
rect -35 731 35 777
rect 81 731 151 777
rect 197 731 267 777
rect 313 731 383 777
rect 429 731 499 777
rect 545 731 615 777
rect 661 731 731 777
rect 777 731 847 777
rect 893 731 963 777
rect 1009 731 1079 777
rect 1125 731 1195 777
rect 1241 731 1311 777
rect 1357 731 1427 777
rect 1473 731 1543 777
rect 1589 731 1659 777
rect 1705 731 1775 777
rect 1821 731 1891 777
rect 1937 731 2007 777
rect 2053 731 2123 777
rect 2169 731 2239 777
rect 2285 731 2355 777
rect 2401 731 2471 777
rect 2517 731 2587 777
rect 2633 731 2703 777
rect 2749 731 2819 777
rect 2865 731 2876 777
rect -2876 661 2876 731
rect -2876 615 -2865 661
rect -2819 615 -2749 661
rect -2703 615 -2633 661
rect -2587 615 -2517 661
rect -2471 615 -2401 661
rect -2355 615 -2285 661
rect -2239 615 -2169 661
rect -2123 615 -2053 661
rect -2007 615 -1937 661
rect -1891 615 -1821 661
rect -1775 615 -1705 661
rect -1659 615 -1589 661
rect -1543 615 -1473 661
rect -1427 615 -1357 661
rect -1311 615 -1241 661
rect -1195 615 -1125 661
rect -1079 615 -1009 661
rect -963 615 -893 661
rect -847 615 -777 661
rect -731 615 -661 661
rect -615 615 -545 661
rect -499 615 -429 661
rect -383 615 -313 661
rect -267 615 -197 661
rect -151 615 -81 661
rect -35 615 35 661
rect 81 615 151 661
rect 197 615 267 661
rect 313 615 383 661
rect 429 615 499 661
rect 545 615 615 661
rect 661 615 731 661
rect 777 615 847 661
rect 893 615 963 661
rect 1009 615 1079 661
rect 1125 615 1195 661
rect 1241 615 1311 661
rect 1357 615 1427 661
rect 1473 615 1543 661
rect 1589 615 1659 661
rect 1705 615 1775 661
rect 1821 615 1891 661
rect 1937 615 2007 661
rect 2053 615 2123 661
rect 2169 615 2239 661
rect 2285 615 2355 661
rect 2401 615 2471 661
rect 2517 615 2587 661
rect 2633 615 2703 661
rect 2749 615 2819 661
rect 2865 615 2876 661
rect -2876 545 2876 615
rect -2876 499 -2865 545
rect -2819 499 -2749 545
rect -2703 499 -2633 545
rect -2587 499 -2517 545
rect -2471 499 -2401 545
rect -2355 499 -2285 545
rect -2239 499 -2169 545
rect -2123 499 -2053 545
rect -2007 499 -1937 545
rect -1891 499 -1821 545
rect -1775 499 -1705 545
rect -1659 499 -1589 545
rect -1543 499 -1473 545
rect -1427 499 -1357 545
rect -1311 499 -1241 545
rect -1195 499 -1125 545
rect -1079 499 -1009 545
rect -963 499 -893 545
rect -847 499 -777 545
rect -731 499 -661 545
rect -615 499 -545 545
rect -499 499 -429 545
rect -383 499 -313 545
rect -267 499 -197 545
rect -151 499 -81 545
rect -35 499 35 545
rect 81 499 151 545
rect 197 499 267 545
rect 313 499 383 545
rect 429 499 499 545
rect 545 499 615 545
rect 661 499 731 545
rect 777 499 847 545
rect 893 499 963 545
rect 1009 499 1079 545
rect 1125 499 1195 545
rect 1241 499 1311 545
rect 1357 499 1427 545
rect 1473 499 1543 545
rect 1589 499 1659 545
rect 1705 499 1775 545
rect 1821 499 1891 545
rect 1937 499 2007 545
rect 2053 499 2123 545
rect 2169 499 2239 545
rect 2285 499 2355 545
rect 2401 499 2471 545
rect 2517 499 2587 545
rect 2633 499 2703 545
rect 2749 499 2819 545
rect 2865 499 2876 545
rect -2876 429 2876 499
rect -2876 383 -2865 429
rect -2819 383 -2749 429
rect -2703 383 -2633 429
rect -2587 383 -2517 429
rect -2471 383 -2401 429
rect -2355 383 -2285 429
rect -2239 383 -2169 429
rect -2123 383 -2053 429
rect -2007 383 -1937 429
rect -1891 383 -1821 429
rect -1775 383 -1705 429
rect -1659 383 -1589 429
rect -1543 383 -1473 429
rect -1427 383 -1357 429
rect -1311 383 -1241 429
rect -1195 383 -1125 429
rect -1079 383 -1009 429
rect -963 383 -893 429
rect -847 383 -777 429
rect -731 383 -661 429
rect -615 383 -545 429
rect -499 383 -429 429
rect -383 383 -313 429
rect -267 383 -197 429
rect -151 383 -81 429
rect -35 383 35 429
rect 81 383 151 429
rect 197 383 267 429
rect 313 383 383 429
rect 429 383 499 429
rect 545 383 615 429
rect 661 383 731 429
rect 777 383 847 429
rect 893 383 963 429
rect 1009 383 1079 429
rect 1125 383 1195 429
rect 1241 383 1311 429
rect 1357 383 1427 429
rect 1473 383 1543 429
rect 1589 383 1659 429
rect 1705 383 1775 429
rect 1821 383 1891 429
rect 1937 383 2007 429
rect 2053 383 2123 429
rect 2169 383 2239 429
rect 2285 383 2355 429
rect 2401 383 2471 429
rect 2517 383 2587 429
rect 2633 383 2703 429
rect 2749 383 2819 429
rect 2865 383 2876 429
rect -2876 313 2876 383
rect -2876 267 -2865 313
rect -2819 267 -2749 313
rect -2703 267 -2633 313
rect -2587 267 -2517 313
rect -2471 267 -2401 313
rect -2355 267 -2285 313
rect -2239 267 -2169 313
rect -2123 267 -2053 313
rect -2007 267 -1937 313
rect -1891 267 -1821 313
rect -1775 267 -1705 313
rect -1659 267 -1589 313
rect -1543 267 -1473 313
rect -1427 267 -1357 313
rect -1311 267 -1241 313
rect -1195 267 -1125 313
rect -1079 267 -1009 313
rect -963 267 -893 313
rect -847 267 -777 313
rect -731 267 -661 313
rect -615 267 -545 313
rect -499 267 -429 313
rect -383 267 -313 313
rect -267 267 -197 313
rect -151 267 -81 313
rect -35 267 35 313
rect 81 267 151 313
rect 197 267 267 313
rect 313 267 383 313
rect 429 267 499 313
rect 545 267 615 313
rect 661 267 731 313
rect 777 267 847 313
rect 893 267 963 313
rect 1009 267 1079 313
rect 1125 267 1195 313
rect 1241 267 1311 313
rect 1357 267 1427 313
rect 1473 267 1543 313
rect 1589 267 1659 313
rect 1705 267 1775 313
rect 1821 267 1891 313
rect 1937 267 2007 313
rect 2053 267 2123 313
rect 2169 267 2239 313
rect 2285 267 2355 313
rect 2401 267 2471 313
rect 2517 267 2587 313
rect 2633 267 2703 313
rect 2749 267 2819 313
rect 2865 267 2876 313
rect -2876 197 2876 267
rect -2876 151 -2865 197
rect -2819 151 -2749 197
rect -2703 151 -2633 197
rect -2587 151 -2517 197
rect -2471 151 -2401 197
rect -2355 151 -2285 197
rect -2239 151 -2169 197
rect -2123 151 -2053 197
rect -2007 151 -1937 197
rect -1891 151 -1821 197
rect -1775 151 -1705 197
rect -1659 151 -1589 197
rect -1543 151 -1473 197
rect -1427 151 -1357 197
rect -1311 151 -1241 197
rect -1195 151 -1125 197
rect -1079 151 -1009 197
rect -963 151 -893 197
rect -847 151 -777 197
rect -731 151 -661 197
rect -615 151 -545 197
rect -499 151 -429 197
rect -383 151 -313 197
rect -267 151 -197 197
rect -151 151 -81 197
rect -35 151 35 197
rect 81 151 151 197
rect 197 151 267 197
rect 313 151 383 197
rect 429 151 499 197
rect 545 151 615 197
rect 661 151 731 197
rect 777 151 847 197
rect 893 151 963 197
rect 1009 151 1079 197
rect 1125 151 1195 197
rect 1241 151 1311 197
rect 1357 151 1427 197
rect 1473 151 1543 197
rect 1589 151 1659 197
rect 1705 151 1775 197
rect 1821 151 1891 197
rect 1937 151 2007 197
rect 2053 151 2123 197
rect 2169 151 2239 197
rect 2285 151 2355 197
rect 2401 151 2471 197
rect 2517 151 2587 197
rect 2633 151 2703 197
rect 2749 151 2819 197
rect 2865 151 2876 197
rect -2876 81 2876 151
rect -2876 35 -2865 81
rect -2819 35 -2749 81
rect -2703 35 -2633 81
rect -2587 35 -2517 81
rect -2471 35 -2401 81
rect -2355 35 -2285 81
rect -2239 35 -2169 81
rect -2123 35 -2053 81
rect -2007 35 -1937 81
rect -1891 35 -1821 81
rect -1775 35 -1705 81
rect -1659 35 -1589 81
rect -1543 35 -1473 81
rect -1427 35 -1357 81
rect -1311 35 -1241 81
rect -1195 35 -1125 81
rect -1079 35 -1009 81
rect -963 35 -893 81
rect -847 35 -777 81
rect -731 35 -661 81
rect -615 35 -545 81
rect -499 35 -429 81
rect -383 35 -313 81
rect -267 35 -197 81
rect -151 35 -81 81
rect -35 35 35 81
rect 81 35 151 81
rect 197 35 267 81
rect 313 35 383 81
rect 429 35 499 81
rect 545 35 615 81
rect 661 35 731 81
rect 777 35 847 81
rect 893 35 963 81
rect 1009 35 1079 81
rect 1125 35 1195 81
rect 1241 35 1311 81
rect 1357 35 1427 81
rect 1473 35 1543 81
rect 1589 35 1659 81
rect 1705 35 1775 81
rect 1821 35 1891 81
rect 1937 35 2007 81
rect 2053 35 2123 81
rect 2169 35 2239 81
rect 2285 35 2355 81
rect 2401 35 2471 81
rect 2517 35 2587 81
rect 2633 35 2703 81
rect 2749 35 2819 81
rect 2865 35 2876 81
rect -2876 -35 2876 35
rect -2876 -81 -2865 -35
rect -2819 -81 -2749 -35
rect -2703 -81 -2633 -35
rect -2587 -81 -2517 -35
rect -2471 -81 -2401 -35
rect -2355 -81 -2285 -35
rect -2239 -81 -2169 -35
rect -2123 -81 -2053 -35
rect -2007 -81 -1937 -35
rect -1891 -81 -1821 -35
rect -1775 -81 -1705 -35
rect -1659 -81 -1589 -35
rect -1543 -81 -1473 -35
rect -1427 -81 -1357 -35
rect -1311 -81 -1241 -35
rect -1195 -81 -1125 -35
rect -1079 -81 -1009 -35
rect -963 -81 -893 -35
rect -847 -81 -777 -35
rect -731 -81 -661 -35
rect -615 -81 -545 -35
rect -499 -81 -429 -35
rect -383 -81 -313 -35
rect -267 -81 -197 -35
rect -151 -81 -81 -35
rect -35 -81 35 -35
rect 81 -81 151 -35
rect 197 -81 267 -35
rect 313 -81 383 -35
rect 429 -81 499 -35
rect 545 -81 615 -35
rect 661 -81 731 -35
rect 777 -81 847 -35
rect 893 -81 963 -35
rect 1009 -81 1079 -35
rect 1125 -81 1195 -35
rect 1241 -81 1311 -35
rect 1357 -81 1427 -35
rect 1473 -81 1543 -35
rect 1589 -81 1659 -35
rect 1705 -81 1775 -35
rect 1821 -81 1891 -35
rect 1937 -81 2007 -35
rect 2053 -81 2123 -35
rect 2169 -81 2239 -35
rect 2285 -81 2355 -35
rect 2401 -81 2471 -35
rect 2517 -81 2587 -35
rect 2633 -81 2703 -35
rect 2749 -81 2819 -35
rect 2865 -81 2876 -35
rect -2876 -151 2876 -81
rect -2876 -197 -2865 -151
rect -2819 -197 -2749 -151
rect -2703 -197 -2633 -151
rect -2587 -197 -2517 -151
rect -2471 -197 -2401 -151
rect -2355 -197 -2285 -151
rect -2239 -197 -2169 -151
rect -2123 -197 -2053 -151
rect -2007 -197 -1937 -151
rect -1891 -197 -1821 -151
rect -1775 -197 -1705 -151
rect -1659 -197 -1589 -151
rect -1543 -197 -1473 -151
rect -1427 -197 -1357 -151
rect -1311 -197 -1241 -151
rect -1195 -197 -1125 -151
rect -1079 -197 -1009 -151
rect -963 -197 -893 -151
rect -847 -197 -777 -151
rect -731 -197 -661 -151
rect -615 -197 -545 -151
rect -499 -197 -429 -151
rect -383 -197 -313 -151
rect -267 -197 -197 -151
rect -151 -197 -81 -151
rect -35 -197 35 -151
rect 81 -197 151 -151
rect 197 -197 267 -151
rect 313 -197 383 -151
rect 429 -197 499 -151
rect 545 -197 615 -151
rect 661 -197 731 -151
rect 777 -197 847 -151
rect 893 -197 963 -151
rect 1009 -197 1079 -151
rect 1125 -197 1195 -151
rect 1241 -197 1311 -151
rect 1357 -197 1427 -151
rect 1473 -197 1543 -151
rect 1589 -197 1659 -151
rect 1705 -197 1775 -151
rect 1821 -197 1891 -151
rect 1937 -197 2007 -151
rect 2053 -197 2123 -151
rect 2169 -197 2239 -151
rect 2285 -197 2355 -151
rect 2401 -197 2471 -151
rect 2517 -197 2587 -151
rect 2633 -197 2703 -151
rect 2749 -197 2819 -151
rect 2865 -197 2876 -151
rect -2876 -267 2876 -197
rect -2876 -313 -2865 -267
rect -2819 -313 -2749 -267
rect -2703 -313 -2633 -267
rect -2587 -313 -2517 -267
rect -2471 -313 -2401 -267
rect -2355 -313 -2285 -267
rect -2239 -313 -2169 -267
rect -2123 -313 -2053 -267
rect -2007 -313 -1937 -267
rect -1891 -313 -1821 -267
rect -1775 -313 -1705 -267
rect -1659 -313 -1589 -267
rect -1543 -313 -1473 -267
rect -1427 -313 -1357 -267
rect -1311 -313 -1241 -267
rect -1195 -313 -1125 -267
rect -1079 -313 -1009 -267
rect -963 -313 -893 -267
rect -847 -313 -777 -267
rect -731 -313 -661 -267
rect -615 -313 -545 -267
rect -499 -313 -429 -267
rect -383 -313 -313 -267
rect -267 -313 -197 -267
rect -151 -313 -81 -267
rect -35 -313 35 -267
rect 81 -313 151 -267
rect 197 -313 267 -267
rect 313 -313 383 -267
rect 429 -313 499 -267
rect 545 -313 615 -267
rect 661 -313 731 -267
rect 777 -313 847 -267
rect 893 -313 963 -267
rect 1009 -313 1079 -267
rect 1125 -313 1195 -267
rect 1241 -313 1311 -267
rect 1357 -313 1427 -267
rect 1473 -313 1543 -267
rect 1589 -313 1659 -267
rect 1705 -313 1775 -267
rect 1821 -313 1891 -267
rect 1937 -313 2007 -267
rect 2053 -313 2123 -267
rect 2169 -313 2239 -267
rect 2285 -313 2355 -267
rect 2401 -313 2471 -267
rect 2517 -313 2587 -267
rect 2633 -313 2703 -267
rect 2749 -313 2819 -267
rect 2865 -313 2876 -267
rect -2876 -383 2876 -313
rect -2876 -429 -2865 -383
rect -2819 -429 -2749 -383
rect -2703 -429 -2633 -383
rect -2587 -429 -2517 -383
rect -2471 -429 -2401 -383
rect -2355 -429 -2285 -383
rect -2239 -429 -2169 -383
rect -2123 -429 -2053 -383
rect -2007 -429 -1937 -383
rect -1891 -429 -1821 -383
rect -1775 -429 -1705 -383
rect -1659 -429 -1589 -383
rect -1543 -429 -1473 -383
rect -1427 -429 -1357 -383
rect -1311 -429 -1241 -383
rect -1195 -429 -1125 -383
rect -1079 -429 -1009 -383
rect -963 -429 -893 -383
rect -847 -429 -777 -383
rect -731 -429 -661 -383
rect -615 -429 -545 -383
rect -499 -429 -429 -383
rect -383 -429 -313 -383
rect -267 -429 -197 -383
rect -151 -429 -81 -383
rect -35 -429 35 -383
rect 81 -429 151 -383
rect 197 -429 267 -383
rect 313 -429 383 -383
rect 429 -429 499 -383
rect 545 -429 615 -383
rect 661 -429 731 -383
rect 777 -429 847 -383
rect 893 -429 963 -383
rect 1009 -429 1079 -383
rect 1125 -429 1195 -383
rect 1241 -429 1311 -383
rect 1357 -429 1427 -383
rect 1473 -429 1543 -383
rect 1589 -429 1659 -383
rect 1705 -429 1775 -383
rect 1821 -429 1891 -383
rect 1937 -429 2007 -383
rect 2053 -429 2123 -383
rect 2169 -429 2239 -383
rect 2285 -429 2355 -383
rect 2401 -429 2471 -383
rect 2517 -429 2587 -383
rect 2633 -429 2703 -383
rect 2749 -429 2819 -383
rect 2865 -429 2876 -383
rect -2876 -499 2876 -429
rect -2876 -545 -2865 -499
rect -2819 -545 -2749 -499
rect -2703 -545 -2633 -499
rect -2587 -545 -2517 -499
rect -2471 -545 -2401 -499
rect -2355 -545 -2285 -499
rect -2239 -545 -2169 -499
rect -2123 -545 -2053 -499
rect -2007 -545 -1937 -499
rect -1891 -545 -1821 -499
rect -1775 -545 -1705 -499
rect -1659 -545 -1589 -499
rect -1543 -545 -1473 -499
rect -1427 -545 -1357 -499
rect -1311 -545 -1241 -499
rect -1195 -545 -1125 -499
rect -1079 -545 -1009 -499
rect -963 -545 -893 -499
rect -847 -545 -777 -499
rect -731 -545 -661 -499
rect -615 -545 -545 -499
rect -499 -545 -429 -499
rect -383 -545 -313 -499
rect -267 -545 -197 -499
rect -151 -545 -81 -499
rect -35 -545 35 -499
rect 81 -545 151 -499
rect 197 -545 267 -499
rect 313 -545 383 -499
rect 429 -545 499 -499
rect 545 -545 615 -499
rect 661 -545 731 -499
rect 777 -545 847 -499
rect 893 -545 963 -499
rect 1009 -545 1079 -499
rect 1125 -545 1195 -499
rect 1241 -545 1311 -499
rect 1357 -545 1427 -499
rect 1473 -545 1543 -499
rect 1589 -545 1659 -499
rect 1705 -545 1775 -499
rect 1821 -545 1891 -499
rect 1937 -545 2007 -499
rect 2053 -545 2123 -499
rect 2169 -545 2239 -499
rect 2285 -545 2355 -499
rect 2401 -545 2471 -499
rect 2517 -545 2587 -499
rect 2633 -545 2703 -499
rect 2749 -545 2819 -499
rect 2865 -545 2876 -499
rect -2876 -615 2876 -545
rect -2876 -661 -2865 -615
rect -2819 -661 -2749 -615
rect -2703 -661 -2633 -615
rect -2587 -661 -2517 -615
rect -2471 -661 -2401 -615
rect -2355 -661 -2285 -615
rect -2239 -661 -2169 -615
rect -2123 -661 -2053 -615
rect -2007 -661 -1937 -615
rect -1891 -661 -1821 -615
rect -1775 -661 -1705 -615
rect -1659 -661 -1589 -615
rect -1543 -661 -1473 -615
rect -1427 -661 -1357 -615
rect -1311 -661 -1241 -615
rect -1195 -661 -1125 -615
rect -1079 -661 -1009 -615
rect -963 -661 -893 -615
rect -847 -661 -777 -615
rect -731 -661 -661 -615
rect -615 -661 -545 -615
rect -499 -661 -429 -615
rect -383 -661 -313 -615
rect -267 -661 -197 -615
rect -151 -661 -81 -615
rect -35 -661 35 -615
rect 81 -661 151 -615
rect 197 -661 267 -615
rect 313 -661 383 -615
rect 429 -661 499 -615
rect 545 -661 615 -615
rect 661 -661 731 -615
rect 777 -661 847 -615
rect 893 -661 963 -615
rect 1009 -661 1079 -615
rect 1125 -661 1195 -615
rect 1241 -661 1311 -615
rect 1357 -661 1427 -615
rect 1473 -661 1543 -615
rect 1589 -661 1659 -615
rect 1705 -661 1775 -615
rect 1821 -661 1891 -615
rect 1937 -661 2007 -615
rect 2053 -661 2123 -615
rect 2169 -661 2239 -615
rect 2285 -661 2355 -615
rect 2401 -661 2471 -615
rect 2517 -661 2587 -615
rect 2633 -661 2703 -615
rect 2749 -661 2819 -615
rect 2865 -661 2876 -615
rect -2876 -731 2876 -661
rect -2876 -777 -2865 -731
rect -2819 -777 -2749 -731
rect -2703 -777 -2633 -731
rect -2587 -777 -2517 -731
rect -2471 -777 -2401 -731
rect -2355 -777 -2285 -731
rect -2239 -777 -2169 -731
rect -2123 -777 -2053 -731
rect -2007 -777 -1937 -731
rect -1891 -777 -1821 -731
rect -1775 -777 -1705 -731
rect -1659 -777 -1589 -731
rect -1543 -777 -1473 -731
rect -1427 -777 -1357 -731
rect -1311 -777 -1241 -731
rect -1195 -777 -1125 -731
rect -1079 -777 -1009 -731
rect -963 -777 -893 -731
rect -847 -777 -777 -731
rect -731 -777 -661 -731
rect -615 -777 -545 -731
rect -499 -777 -429 -731
rect -383 -777 -313 -731
rect -267 -777 -197 -731
rect -151 -777 -81 -731
rect -35 -777 35 -731
rect 81 -777 151 -731
rect 197 -777 267 -731
rect 313 -777 383 -731
rect 429 -777 499 -731
rect 545 -777 615 -731
rect 661 -777 731 -731
rect 777 -777 847 -731
rect 893 -777 963 -731
rect 1009 -777 1079 -731
rect 1125 -777 1195 -731
rect 1241 -777 1311 -731
rect 1357 -777 1427 -731
rect 1473 -777 1543 -731
rect 1589 -777 1659 -731
rect 1705 -777 1775 -731
rect 1821 -777 1891 -731
rect 1937 -777 2007 -731
rect 2053 -777 2123 -731
rect 2169 -777 2239 -731
rect 2285 -777 2355 -731
rect 2401 -777 2471 -731
rect 2517 -777 2587 -731
rect 2633 -777 2703 -731
rect 2749 -777 2819 -731
rect 2865 -777 2876 -731
rect -2876 -847 2876 -777
rect -2876 -893 -2865 -847
rect -2819 -893 -2749 -847
rect -2703 -893 -2633 -847
rect -2587 -893 -2517 -847
rect -2471 -893 -2401 -847
rect -2355 -893 -2285 -847
rect -2239 -893 -2169 -847
rect -2123 -893 -2053 -847
rect -2007 -893 -1937 -847
rect -1891 -893 -1821 -847
rect -1775 -893 -1705 -847
rect -1659 -893 -1589 -847
rect -1543 -893 -1473 -847
rect -1427 -893 -1357 -847
rect -1311 -893 -1241 -847
rect -1195 -893 -1125 -847
rect -1079 -893 -1009 -847
rect -963 -893 -893 -847
rect -847 -893 -777 -847
rect -731 -893 -661 -847
rect -615 -893 -545 -847
rect -499 -893 -429 -847
rect -383 -893 -313 -847
rect -267 -893 -197 -847
rect -151 -893 -81 -847
rect -35 -893 35 -847
rect 81 -893 151 -847
rect 197 -893 267 -847
rect 313 -893 383 -847
rect 429 -893 499 -847
rect 545 -893 615 -847
rect 661 -893 731 -847
rect 777 -893 847 -847
rect 893 -893 963 -847
rect 1009 -893 1079 -847
rect 1125 -893 1195 -847
rect 1241 -893 1311 -847
rect 1357 -893 1427 -847
rect 1473 -893 1543 -847
rect 1589 -893 1659 -847
rect 1705 -893 1775 -847
rect 1821 -893 1891 -847
rect 1937 -893 2007 -847
rect 2053 -893 2123 -847
rect 2169 -893 2239 -847
rect 2285 -893 2355 -847
rect 2401 -893 2471 -847
rect 2517 -893 2587 -847
rect 2633 -893 2703 -847
rect 2749 -893 2819 -847
rect 2865 -893 2876 -847
rect -2876 -963 2876 -893
rect -2876 -1009 -2865 -963
rect -2819 -1009 -2749 -963
rect -2703 -1009 -2633 -963
rect -2587 -1009 -2517 -963
rect -2471 -1009 -2401 -963
rect -2355 -1009 -2285 -963
rect -2239 -1009 -2169 -963
rect -2123 -1009 -2053 -963
rect -2007 -1009 -1937 -963
rect -1891 -1009 -1821 -963
rect -1775 -1009 -1705 -963
rect -1659 -1009 -1589 -963
rect -1543 -1009 -1473 -963
rect -1427 -1009 -1357 -963
rect -1311 -1009 -1241 -963
rect -1195 -1009 -1125 -963
rect -1079 -1009 -1009 -963
rect -963 -1009 -893 -963
rect -847 -1009 -777 -963
rect -731 -1009 -661 -963
rect -615 -1009 -545 -963
rect -499 -1009 -429 -963
rect -383 -1009 -313 -963
rect -267 -1009 -197 -963
rect -151 -1009 -81 -963
rect -35 -1009 35 -963
rect 81 -1009 151 -963
rect 197 -1009 267 -963
rect 313 -1009 383 -963
rect 429 -1009 499 -963
rect 545 -1009 615 -963
rect 661 -1009 731 -963
rect 777 -1009 847 -963
rect 893 -1009 963 -963
rect 1009 -1009 1079 -963
rect 1125 -1009 1195 -963
rect 1241 -1009 1311 -963
rect 1357 -1009 1427 -963
rect 1473 -1009 1543 -963
rect 1589 -1009 1659 -963
rect 1705 -1009 1775 -963
rect 1821 -1009 1891 -963
rect 1937 -1009 2007 -963
rect 2053 -1009 2123 -963
rect 2169 -1009 2239 -963
rect 2285 -1009 2355 -963
rect 2401 -1009 2471 -963
rect 2517 -1009 2587 -963
rect 2633 -1009 2703 -963
rect 2749 -1009 2819 -963
rect 2865 -1009 2876 -963
rect -2876 -1079 2876 -1009
rect -2876 -1125 -2865 -1079
rect -2819 -1125 -2749 -1079
rect -2703 -1125 -2633 -1079
rect -2587 -1125 -2517 -1079
rect -2471 -1125 -2401 -1079
rect -2355 -1125 -2285 -1079
rect -2239 -1125 -2169 -1079
rect -2123 -1125 -2053 -1079
rect -2007 -1125 -1937 -1079
rect -1891 -1125 -1821 -1079
rect -1775 -1125 -1705 -1079
rect -1659 -1125 -1589 -1079
rect -1543 -1125 -1473 -1079
rect -1427 -1125 -1357 -1079
rect -1311 -1125 -1241 -1079
rect -1195 -1125 -1125 -1079
rect -1079 -1125 -1009 -1079
rect -963 -1125 -893 -1079
rect -847 -1125 -777 -1079
rect -731 -1125 -661 -1079
rect -615 -1125 -545 -1079
rect -499 -1125 -429 -1079
rect -383 -1125 -313 -1079
rect -267 -1125 -197 -1079
rect -151 -1125 -81 -1079
rect -35 -1125 35 -1079
rect 81 -1125 151 -1079
rect 197 -1125 267 -1079
rect 313 -1125 383 -1079
rect 429 -1125 499 -1079
rect 545 -1125 615 -1079
rect 661 -1125 731 -1079
rect 777 -1125 847 -1079
rect 893 -1125 963 -1079
rect 1009 -1125 1079 -1079
rect 1125 -1125 1195 -1079
rect 1241 -1125 1311 -1079
rect 1357 -1125 1427 -1079
rect 1473 -1125 1543 -1079
rect 1589 -1125 1659 -1079
rect 1705 -1125 1775 -1079
rect 1821 -1125 1891 -1079
rect 1937 -1125 2007 -1079
rect 2053 -1125 2123 -1079
rect 2169 -1125 2239 -1079
rect 2285 -1125 2355 -1079
rect 2401 -1125 2471 -1079
rect 2517 -1125 2587 -1079
rect 2633 -1125 2703 -1079
rect 2749 -1125 2819 -1079
rect 2865 -1125 2876 -1079
rect -2876 -1136 2876 -1125
<< properties >>
string GDS_END 2138856
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2074660
<< end >>
