magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 760 1620
<< nmos >>
rect 160 190 220 360
rect 330 190 390 360
rect 500 190 560 360
<< pmos >>
rect 190 1090 250 1430
rect 300 1090 360 1430
rect 500 1090 560 1430
<< ndiff >>
rect 60 298 160 360
rect 60 252 82 298
rect 128 252 160 298
rect 60 190 160 252
rect 220 298 330 360
rect 220 252 252 298
rect 298 252 330 298
rect 220 190 330 252
rect 390 298 500 360
rect 390 252 422 298
rect 468 252 500 298
rect 390 190 500 252
rect 560 298 660 360
rect 560 252 592 298
rect 638 252 660 298
rect 560 190 660 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1090 300 1430
rect 360 1377 500 1430
rect 360 1143 407 1377
rect 453 1143 500 1377
rect 360 1090 500 1143
rect 560 1377 660 1430
rect 560 1143 592 1377
rect 638 1143 660 1377
rect 560 1090 660 1143
<< ndiffc >>
rect 82 252 128 298
rect 252 252 298 298
rect 422 252 468 298
rect 592 252 638 298
<< pdiffc >>
rect 112 1143 158 1377
rect 407 1143 453 1377
rect 592 1143 638 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 300 1430 360 1480
rect 500 1430 560 1480
rect 190 1050 250 1090
rect 160 1000 250 1050
rect 300 1060 360 1090
rect 300 1000 390 1060
rect 160 780 220 1000
rect 160 753 280 780
rect 160 707 207 753
rect 253 707 280 753
rect 160 680 280 707
rect 160 360 220 680
rect 330 650 390 1000
rect 500 910 560 1090
rect 440 883 560 910
rect 440 837 467 883
rect 513 837 560 883
rect 440 810 560 837
rect 330 623 430 650
rect 330 577 357 623
rect 403 577 430 623
rect 330 550 430 577
rect 330 360 390 550
rect 500 360 560 810
rect 160 140 220 190
rect 330 140 390 190
rect 500 140 560 190
<< polycontact >>
rect 207 707 253 753
rect 467 837 513 883
rect 357 577 403 623
<< metal1 >>
rect 0 1568 760 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 760 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 760 1566
rect 0 1470 760 1514
rect 110 1377 160 1430
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1100 160 1143
rect 80 1050 160 1100
rect 390 1377 470 1470
rect 390 1143 407 1377
rect 453 1143 470 1377
rect 390 1060 470 1143
rect 590 1377 640 1430
rect 590 1143 592 1377
rect 638 1143 640 1377
rect 80 890 130 1050
rect 590 1020 640 1143
rect 590 1016 690 1020
rect 590 964 614 1016
rect 666 964 690 1016
rect 590 930 690 964
rect 80 886 540 890
rect 80 834 464 886
rect 516 834 540 886
rect 80 830 540 834
rect 80 490 130 830
rect 180 756 280 760
rect 180 704 204 756
rect 256 704 280 756
rect 180 670 280 704
rect 330 626 430 630
rect 330 574 354 626
rect 406 574 430 626
rect 330 540 430 574
rect 80 440 300 490
rect 80 298 130 360
rect 80 252 82 298
rect 128 252 130 298
rect 80 120 130 252
rect 250 298 300 440
rect 250 252 252 298
rect 298 252 300 298
rect 250 190 300 252
rect 420 298 470 360
rect 420 252 422 298
rect 468 252 470 298
rect 420 120 470 252
rect 590 298 640 930
rect 590 252 592 298
rect 638 252 640 298
rect 590 160 640 252
rect 0 106 760 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 760 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 760 54
rect 0 -30 760 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 614 964 666 1016
rect 464 883 516 886
rect 464 837 467 883
rect 467 837 513 883
rect 513 837 516 883
rect 464 834 516 837
rect 204 753 256 756
rect 204 707 207 753
rect 207 707 253 753
rect 253 707 256 753
rect 204 704 256 707
rect 354 623 406 626
rect 354 577 357 623
rect 357 577 403 623
rect 403 577 406 623
rect 354 574 406 577
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
<< metal2 >>
rect 90 1566 190 1580
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1470 190 1514
rect 330 1566 430 1580
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1470 430 1514
rect 570 1566 670 1580
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1470 670 1514
rect 590 1016 690 1030
rect 590 964 614 1016
rect 666 964 690 1016
rect 590 920 690 964
rect 440 886 540 900
rect 440 834 464 886
rect 516 834 540 886
rect 440 820 540 834
rect 180 756 280 770
rect 180 704 204 756
rect 256 704 280 756
rect 180 660 280 704
rect 330 626 430 640
rect 330 574 354 626
rect 406 574 430 626
rect 330 530 430 574
rect 90 106 190 120
rect 90 54 114 106
rect 166 54 190 106
rect 90 10 190 54
rect 330 106 430 120
rect 330 54 354 106
rect 406 54 430 106
rect 330 10 430 54
rect 570 106 670 120
rect 570 54 594 106
rect 646 54 670 106
rect 570 10 670 54
<< labels >>
rlabel metal2 s 90 10 190 90 4 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 90 1470 190 1550 4 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 530 430 610 4 B
port 1 nsew signal input
rlabel metal2 s 180 660 280 740 4 A
port 2 nsew signal input
rlabel metal2 s 590 920 690 1000 4 Y
port 3 nsew signal output
rlabel metal1 s 180 670 280 730 1 A
port 2 nsew signal input
rlabel metal1 s 330 540 430 600 1 B
port 1 nsew signal input
rlabel metal2 s 330 1470 430 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 570 1470 670 1550 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 390 1060 470 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 0 1470 760 1590 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal2 s 330 10 430 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal2 s 570 10 670 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 80 -30 130 330 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 420 -30 470 330 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 0 -30 760 90 1 VSS
port 9 nsew ground bidirectional
rlabel metal1 s 590 160 640 1400 1 Y
port 3 nsew signal output
rlabel metal1 s 590 930 690 990 1 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 760 1590
string GDS_END 425518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 419176
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
