magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect 85432 578 85816 53502
<< metal1 >>
rect 0 403 1000 53494
<< metal2 >>
rect 424 403 1424 52949
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105905487112_128x8m81  M1_PSUB43105905487112_128x8m81_0
timestamp 1669390400
transform -1 0 85672 0 1 53088
box -42 -42 85602 414
use M1_PSUB43105905487112_128x8m81  M1_PSUB43105905487112_128x8m81_1
timestamp 1669390400
transform -1 0 85672 0 1 620
box -42 -42 85602 414
use M1_PSUB43105905487113_128x8m81  M1_PSUB43105905487113_128x8m81_0
timestamp 1669390400
transform 1 0 85474 0 1 1140
box -42 -42 342 51842
use M1_PSUB43105905487113_128x8m81  M1_PSUB43105905487113_128x8m81_1
timestamp 1669390400
transform 1 0 112 0 1 1140
box -42 -42 342 51842
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2235368
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2234712
string path 4.620 11.160 4.620 0.000 
<< end >>
