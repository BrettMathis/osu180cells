magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1680 844
rect 69 590 115 724
rect 132 232 204 542
rect 356 304 428 664
rect 474 430 538 664
rect 611 594 1013 652
rect 1089 640 1135 724
rect 1207 594 1620 652
rect 611 580 1620 594
rect 951 548 1620 580
rect 474 354 872 430
rect 918 354 1096 430
rect 1032 212 1096 354
rect 1144 354 1322 430
rect 1144 212 1208 354
rect 1368 244 1414 548
rect 1302 198 1414 244
rect 1460 354 1654 430
rect 1460 212 1544 354
rect 49 60 95 152
rect 497 60 543 152
rect 0 -60 1680 60
<< obsm1 >>
rect 273 198 922 244
rect 273 106 319 198
rect 630 106 1640 152
<< labels >>
rlabel metal1 s 1460 354 1654 430 6 A1
port 1 nsew default input
rlabel metal1 s 1460 212 1544 354 6 A1
port 1 nsew default input
rlabel metal1 s 1144 354 1322 430 6 A2
port 2 nsew default input
rlabel metal1 s 1144 212 1208 354 6 A2
port 2 nsew default input
rlabel metal1 s 474 430 538 664 6 B1
port 3 nsew default input
rlabel metal1 s 474 354 872 430 6 B1
port 3 nsew default input
rlabel metal1 s 918 354 1096 430 6 B2
port 4 nsew default input
rlabel metal1 s 1032 212 1096 354 6 B2
port 4 nsew default input
rlabel metal1 s 356 304 428 664 6 C1
port 5 nsew default input
rlabel metal1 s 132 232 204 542 6 C2
port 6 nsew default input
rlabel metal1 s 1207 594 1620 652 6 ZN
port 7 nsew default output
rlabel metal1 s 611 594 1013 652 6 ZN
port 7 nsew default output
rlabel metal1 s 611 580 1620 594 6 ZN
port 7 nsew default output
rlabel metal1 s 951 548 1620 580 6 ZN
port 7 nsew default output
rlabel metal1 s 1368 244 1414 548 6 ZN
port 7 nsew default output
rlabel metal1 s 1302 198 1414 244 6 ZN
port 7 nsew default output
rlabel metal1 s 0 724 1680 844 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1089 640 1135 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 69 640 115 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 69 590 115 640 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 497 60 543 152 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 152 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1680 60 8 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1680 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 124588
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 120322
<< end >>
