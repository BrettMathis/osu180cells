magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 274
<< mvndiff >>
rect -88 261 0 274
rect -88 13 -75 261
rect -29 13 0 261
rect -88 0 0 13
rect 120 261 208 274
rect 120 13 149 261
rect 195 13 208 261
rect 120 0 208 13
<< mvndiffc >>
rect -75 13 -29 261
rect 149 13 195 261
<< polysilicon >>
rect 0 274 120 318
rect 0 -44 120 0
<< metal1 >>
rect -75 261 -29 274
rect -75 0 -29 13
rect 149 261 195 274
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 137 -52 137 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 137 172 137 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 89676
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 88396
<< end >>
