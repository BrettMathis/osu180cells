magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -586 453 310 1094
<< pwell >>
rect -586 -86 310 453
<< mvpsubdiff >>
rect 72 276 144 289
rect 72 136 85 276
rect 131 136 144 276
rect 72 82 144 136
<< mvnsubdiff >>
rect 72 638 144 651
rect 72 498 85 638
rect 131 498 144 638
rect 72 485 144 498
<< mvpsubdiffcont >>
rect 85 136 131 276
<< mvnsubdiffcont >>
rect 85 498 131 638
<< metal1 >>
rect 0 918 224 1098
rect 46 638 170 918
rect 46 498 85 638
rect 131 498 170 638
rect 46 468 170 498
rect 46 276 170 306
rect 46 136 85 276
rect 131 136 170 276
rect 46 90 170 136
rect 0 -90 224 90
<< labels >>
flabel metal1 s 46 90 170 306 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel metal1 s 0 918 224 1098 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 46 468 170 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -90 224 90 1 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 1008
string GDS_END 750844
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 749194
string LEFclass gf180mcu_fd_sc_mcu9t5v0__endcap PRE
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
