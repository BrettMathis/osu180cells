magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 1654 1094
<< pwell >>
rect -86 -86 1654 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
<< mvpmos >>
rect 144 610 244 939
rect 348 610 448 939
rect 592 573 692 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1244 573 1344 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 287 348 333
rect 244 147 273 287
rect 319 147 348 287
rect 244 69 348 147
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 285 796 333
rect 692 239 721 285
rect 767 239 796 285
rect 692 69 796 239
rect 916 287 1020 333
rect 916 147 945 287
rect 991 147 1020 287
rect 916 69 1020 147
rect 1140 285 1244 333
rect 1140 239 1169 285
rect 1215 239 1244 285
rect 1140 69 1244 239
rect 1364 287 1452 333
rect 1364 147 1393 287
rect 1439 147 1452 287
rect 1364 69 1452 147
<< mvpdiff >>
rect 56 884 144 939
rect 56 744 69 884
rect 115 744 144 884
rect 56 610 144 744
rect 244 853 348 939
rect 244 713 273 853
rect 319 713 348 853
rect 244 610 348 713
rect 448 923 592 939
rect 448 783 477 923
rect 523 783 592 923
rect 448 610 592 783
rect 512 573 592 610
rect 692 573 806 939
rect 906 861 1030 939
rect 906 721 935 861
rect 981 721 1030 861
rect 906 573 1030 721
rect 1130 573 1244 939
rect 1344 923 1432 939
rect 1344 783 1373 923
rect 1419 783 1432 923
rect 1344 573 1432 783
<< mvndiffc >>
rect 49 147 95 287
rect 273 147 319 287
rect 497 147 543 287
rect 721 239 767 285
rect 945 147 991 287
rect 1169 239 1215 285
rect 1393 147 1439 287
<< mvpdiffc >>
rect 69 744 115 884
rect 273 713 319 853
rect 477 783 523 923
rect 935 721 981 861
rect 1373 783 1419 923
<< polysilicon >>
rect 144 939 244 983
rect 348 939 448 983
rect 592 939 692 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1244 939 1344 983
rect 144 513 244 610
rect 348 513 448 610
rect 144 500 448 513
rect 144 454 157 500
rect 203 454 448 500
rect 144 441 448 454
rect 144 377 244 441
rect 124 333 244 377
rect 348 377 448 441
rect 592 500 692 573
rect 592 454 605 500
rect 651 454 692 500
rect 592 377 692 454
rect 806 513 906 573
rect 1030 513 1130 573
rect 806 500 1130 513
rect 806 454 819 500
rect 865 454 1130 500
rect 806 441 1130 454
rect 806 377 916 441
rect 348 333 468 377
rect 572 333 692 377
rect 796 333 916 377
rect 1020 377 1130 441
rect 1244 500 1344 573
rect 1244 454 1257 500
rect 1303 454 1344 500
rect 1244 377 1344 454
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
<< polycontact >>
rect 157 454 203 500
rect 605 454 651 500
rect 819 454 865 500
rect 1257 454 1303 500
<< metal1 >>
rect 0 923 1568 1098
rect 0 918 477 923
rect 69 884 115 918
rect 69 733 115 744
rect 273 853 319 864
rect 523 918 1373 923
rect 477 772 523 783
rect 935 861 981 872
rect 319 721 935 726
rect 1419 918 1568 923
rect 1373 772 1419 783
rect 981 721 1395 726
rect 319 713 1395 721
rect 273 680 1395 713
rect 590 588 1303 634
rect 130 500 214 530
rect 130 454 157 500
rect 203 454 214 500
rect 590 500 662 588
rect 590 454 605 500
rect 651 454 662 500
rect 807 500 866 542
rect 807 454 819 500
rect 865 454 866 500
rect 807 443 866 454
rect 1257 500 1303 588
rect 1257 443 1303 454
rect 1349 390 1395 680
rect 49 344 543 390
rect 49 287 95 344
rect 49 136 95 147
rect 273 287 319 298
rect 273 90 319 147
rect 497 287 543 344
rect 721 344 1395 390
rect 721 285 767 344
rect 721 228 767 239
rect 945 287 991 298
rect 543 147 945 182
rect 1038 285 1215 344
rect 1038 239 1169 285
rect 1038 228 1215 239
rect 1393 287 1439 298
rect 991 147 1393 182
rect 497 136 1439 147
rect 0 -90 1568 90
<< labels >>
flabel metal1 s 807 443 866 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 590 588 1303 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 130 454 214 530 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 0 918 1568 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 273 90 319 298 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 935 864 981 872 0 FreeSans 200 0 0 0 ZN
port 4 nsew default output
rlabel metal1 s 1257 454 1303 588 1 A2
port 2 nsew default input
rlabel metal1 s 590 454 662 588 1 A2
port 2 nsew default input
rlabel metal1 s 1257 443 1303 454 1 A2
port 2 nsew default input
rlabel metal1 s 935 726 981 864 1 ZN
port 4 nsew default output
rlabel metal1 s 273 726 319 864 1 ZN
port 4 nsew default output
rlabel metal1 s 273 680 1395 726 1 ZN
port 4 nsew default output
rlabel metal1 s 1349 390 1395 680 1 ZN
port 4 nsew default output
rlabel metal1 s 721 344 1395 390 1 ZN
port 4 nsew default output
rlabel metal1 s 1038 228 1215 344 1 ZN
port 4 nsew default output
rlabel metal1 s 721 228 767 344 1 ZN
port 4 nsew default output
rlabel metal1 s 1373 772 1419 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 477 772 523 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 772 115 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 733 115 772 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 -90 1568 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1568 1008
string GDS_END 118816
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 114542
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
