magic
tech gf180mcuB
timestamp 1669390400
<< metal1 >>
rect 0 147 78 159
rect 11 106 16 147
rect 45 106 50 147
rect 62 101 67 140
rect 62 100 69 101
rect 62 94 72 100
rect 62 93 70 94
rect 12 67 22 73
rect 38 54 48 60
rect 42 9 50 33
rect 62 16 67 93
rect 0 -3 78 9
<< obsm1 >>
rect 28 86 33 140
rect 26 80 57 86
rect 28 40 33 80
rect 14 35 33 40
rect 14 16 19 35
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 9 148 19 154
rect 33 148 43 154
rect 57 148 67 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 62 93 72 101
rect 12 66 22 74
rect 38 53 48 61
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 9 2 19 8
rect 33 2 43 8
rect 57 2 67 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
<< obsm2 >>
rect 26 79 36 87
rect 47 79 57 87
<< labels >>
rlabel metal2 s 12 66 22 74 6 A
port 1 nsew signal input
rlabel metal1 s 12 67 22 73 6 A
port 1 nsew signal input
rlabel metal2 s 38 53 48 61 6 B
port 2 nsew signal input
rlabel metal1 s 38 54 48 60 6 B
port 2 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 34 147 42 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 33 148 43 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 58 147 66 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 57 148 67 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 45 106 50 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 147 78 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 34 1 42 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 33 2 43 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 58 1 66 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 57 2 67 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 42 -3 50 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 0 -3 78 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 62 93 72 101 6 Y
port 3 nsew signal output
rlabel metal1 s 62 16 67 140 6 Y
port 3 nsew signal output
rlabel metal1 s 62 93 69 101 6 Y
port 3 nsew signal output
rlabel metal1 s 62 93 70 100 6 Y
port 3 nsew signal output
rlabel metal1 s 62 94 72 100 6 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 78 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 47360
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 39994
<< end >>
