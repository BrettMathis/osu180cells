magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 3000 1230
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
rect 1550 190 1610 360
rect 1720 190 1780 360
rect 1890 190 1950 360
rect 2060 190 2120 360
rect 2230 190 2290 360
rect 2400 190 2460 360
rect 2570 190 2630 360
rect 2740 190 2800 360
<< pmos >>
rect 190 700 250 1040
rect 360 700 420 1040
rect 530 700 590 1040
rect 700 700 760 1040
rect 870 700 930 1040
rect 1040 700 1100 1040
rect 1210 700 1270 1040
rect 1380 700 1440 1040
rect 1550 700 1610 1040
rect 1720 700 1780 1040
rect 1890 700 1950 1040
rect 2060 700 2120 1040
rect 2230 700 2290 1040
rect 2400 700 2460 1040
rect 2570 700 2630 1040
rect 2740 700 2800 1040
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 870 360
rect 760 252 792 298
rect 838 252 870 298
rect 760 190 870 252
rect 930 298 1040 360
rect 930 252 962 298
rect 1008 252 1040 298
rect 930 190 1040 252
rect 1100 298 1210 360
rect 1100 252 1132 298
rect 1178 252 1210 298
rect 1100 190 1210 252
rect 1270 298 1380 360
rect 1270 252 1302 298
rect 1348 252 1380 298
rect 1270 190 1380 252
rect 1440 298 1550 360
rect 1440 252 1472 298
rect 1518 252 1550 298
rect 1440 190 1550 252
rect 1610 298 1720 360
rect 1610 252 1642 298
rect 1688 252 1720 298
rect 1610 190 1720 252
rect 1780 298 1890 360
rect 1780 252 1812 298
rect 1858 252 1890 298
rect 1780 190 1890 252
rect 1950 298 2060 360
rect 1950 252 1982 298
rect 2028 252 2060 298
rect 1950 190 2060 252
rect 2120 298 2230 360
rect 2120 252 2152 298
rect 2198 252 2230 298
rect 2120 190 2230 252
rect 2290 298 2400 360
rect 2290 252 2322 298
rect 2368 252 2400 298
rect 2290 190 2400 252
rect 2460 298 2570 360
rect 2460 252 2492 298
rect 2538 252 2570 298
rect 2460 190 2570 252
rect 2630 298 2740 360
rect 2630 252 2662 298
rect 2708 252 2740 298
rect 2630 190 2740 252
rect 2800 298 2900 360
rect 2800 252 2832 298
rect 2878 252 2900 298
rect 2800 190 2900 252
<< pdiff >>
rect 90 987 190 1040
rect 90 753 112 987
rect 158 753 190 987
rect 90 700 190 753
rect 250 987 360 1040
rect 250 753 282 987
rect 328 753 360 987
rect 250 700 360 753
rect 420 987 530 1040
rect 420 753 452 987
rect 498 753 530 987
rect 420 700 530 753
rect 590 987 700 1040
rect 590 753 622 987
rect 668 753 700 987
rect 590 700 700 753
rect 760 987 870 1040
rect 760 753 792 987
rect 838 753 870 987
rect 760 700 870 753
rect 930 987 1040 1040
rect 930 753 962 987
rect 1008 753 1040 987
rect 930 700 1040 753
rect 1100 987 1210 1040
rect 1100 753 1132 987
rect 1178 753 1210 987
rect 1100 700 1210 753
rect 1270 987 1380 1040
rect 1270 753 1302 987
rect 1348 753 1380 987
rect 1270 700 1380 753
rect 1440 987 1550 1040
rect 1440 753 1472 987
rect 1518 753 1550 987
rect 1440 700 1550 753
rect 1610 987 1720 1040
rect 1610 753 1642 987
rect 1688 753 1720 987
rect 1610 700 1720 753
rect 1780 987 1890 1040
rect 1780 753 1812 987
rect 1858 753 1890 987
rect 1780 700 1890 753
rect 1950 987 2060 1040
rect 1950 753 1982 987
rect 2028 753 2060 987
rect 1950 700 2060 753
rect 2120 987 2230 1040
rect 2120 753 2152 987
rect 2198 753 2230 987
rect 2120 700 2230 753
rect 2290 987 2400 1040
rect 2290 753 2322 987
rect 2368 753 2400 987
rect 2290 700 2400 753
rect 2460 987 2570 1040
rect 2460 753 2492 987
rect 2538 753 2570 987
rect 2460 700 2570 753
rect 2630 987 2740 1040
rect 2630 753 2662 987
rect 2708 753 2740 987
rect 2630 700 2740 753
rect 2800 987 2910 1040
rect 2800 753 2832 987
rect 2878 753 2910 987
rect 2800 700 2910 753
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
rect 962 252 1008 298
rect 1132 252 1178 298
rect 1302 252 1348 298
rect 1472 252 1518 298
rect 1642 252 1688 298
rect 1812 252 1858 298
rect 1982 252 2028 298
rect 2152 252 2198 298
rect 2322 252 2368 298
rect 2492 252 2538 298
rect 2662 252 2708 298
rect 2832 252 2878 298
<< pdiffc >>
rect 112 753 158 987
rect 282 753 328 987
rect 452 753 498 987
rect 622 753 668 987
rect 792 753 838 987
rect 962 753 1008 987
rect 1132 753 1178 987
rect 1302 753 1348 987
rect 1472 753 1518 987
rect 1642 753 1688 987
rect 1812 753 1858 987
rect 1982 753 2028 987
rect 2152 753 2198 987
rect 2322 753 2368 987
rect 2492 753 2538 987
rect 2662 753 2708 987
rect 2832 753 2878 987
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
rect 1530 98 1620 120
rect 1530 52 1552 98
rect 1598 52 1620 98
rect 1530 30 1620 52
rect 1770 98 1860 120
rect 1770 52 1792 98
rect 1838 52 1860 98
rect 1770 30 1860 52
rect 2010 98 2100 120
rect 2010 52 2032 98
rect 2078 52 2100 98
rect 2010 30 2100 52
rect 2250 98 2340 120
rect 2250 52 2272 98
rect 2318 52 2340 98
rect 2250 30 2340 52
rect 2490 98 2580 120
rect 2490 52 2512 98
rect 2558 52 2580 98
rect 2490 30 2580 52
rect 2730 98 2820 120
rect 2730 52 2752 98
rect 2798 52 2820 98
rect 2730 30 2820 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
rect 810 1178 900 1200
rect 810 1132 832 1178
rect 878 1132 900 1178
rect 810 1110 900 1132
rect 1050 1178 1140 1200
rect 1050 1132 1072 1178
rect 1118 1132 1140 1178
rect 1050 1110 1140 1132
rect 1290 1178 1380 1200
rect 1290 1132 1312 1178
rect 1358 1132 1380 1178
rect 1290 1110 1380 1132
rect 1530 1178 1620 1200
rect 1530 1132 1552 1178
rect 1598 1132 1620 1178
rect 1530 1110 1620 1132
rect 1770 1178 1860 1200
rect 1770 1132 1792 1178
rect 1838 1132 1860 1178
rect 1770 1110 1860 1132
rect 2010 1178 2100 1200
rect 2010 1132 2032 1178
rect 2078 1132 2100 1178
rect 2010 1110 2100 1132
rect 2250 1178 2340 1200
rect 2250 1132 2272 1178
rect 2318 1132 2340 1178
rect 2250 1110 2340 1132
rect 2490 1178 2580 1200
rect 2490 1132 2512 1178
rect 2558 1132 2580 1178
rect 2490 1110 2580 1132
rect 2730 1178 2820 1200
rect 2730 1132 2752 1178
rect 2798 1132 2820 1178
rect 2730 1110 2820 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
rect 1552 52 1598 98
rect 1792 52 1838 98
rect 2032 52 2078 98
rect 2272 52 2318 98
rect 2512 52 2558 98
rect 2752 52 2798 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
rect 832 1132 878 1178
rect 1072 1132 1118 1178
rect 1312 1132 1358 1178
rect 1552 1132 1598 1178
rect 1792 1132 1838 1178
rect 2032 1132 2078 1178
rect 2272 1132 2318 1178
rect 2512 1132 2558 1178
rect 2752 1132 2798 1178
<< polysilicon >>
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 870 1040 930 1090
rect 1040 1040 1100 1090
rect 1210 1040 1270 1090
rect 1380 1040 1440 1090
rect 1550 1040 1610 1090
rect 1720 1040 1780 1090
rect 1890 1040 1950 1090
rect 2060 1040 2120 1090
rect 2230 1040 2290 1090
rect 2400 1040 2460 1090
rect 2570 1040 2630 1090
rect 2740 1040 2800 1090
rect 190 650 250 700
rect 360 650 420 700
rect 530 650 590 700
rect 700 650 760 700
rect 870 650 930 700
rect 1040 650 1100 700
rect 1210 650 1270 700
rect 1380 650 1440 700
rect 1550 650 1610 700
rect 1720 650 1780 700
rect 1890 650 1950 700
rect 2060 650 2120 700
rect 2230 650 2290 700
rect 2400 650 2460 700
rect 2570 650 2630 700
rect 2740 650 2800 700
rect 190 600 2800 650
rect 190 520 250 600
rect 90 498 250 520
rect 90 452 112 498
rect 158 460 250 498
rect 158 452 2800 460
rect 90 430 2800 452
rect 190 400 2800 430
rect 190 360 250 400
rect 360 360 420 400
rect 530 360 590 400
rect 700 360 760 400
rect 870 360 930 400
rect 1040 360 1100 400
rect 1210 360 1270 400
rect 1380 360 1440 400
rect 1550 360 1610 400
rect 1720 360 1780 400
rect 1890 360 1950 400
rect 2060 360 2120 400
rect 2230 360 2290 400
rect 2400 360 2460 400
rect 2570 360 2630 400
rect 2740 360 2800 400
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
rect 1550 140 1610 190
rect 1720 140 1780 190
rect 1890 140 1950 190
rect 2060 140 2120 190
rect 2230 140 2290 190
rect 2400 140 2460 190
rect 2570 140 2630 190
rect 2740 140 2800 190
<< polycontact >>
rect 112 452 158 498
<< metal1 >>
rect 0 1178 3000 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 832 1178
rect 878 1176 1072 1178
rect 1118 1176 1312 1178
rect 1358 1176 1552 1178
rect 1598 1176 1792 1178
rect 1838 1176 2032 1178
rect 2078 1176 2272 1178
rect 2318 1176 2512 1178
rect 2558 1176 2752 1178
rect 2798 1176 3000 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 646 1132 832 1176
rect 886 1132 1072 1176
rect 1126 1132 1312 1176
rect 1366 1132 1552 1176
rect 1606 1132 1792 1176
rect 1846 1132 2032 1176
rect 2086 1132 2272 1176
rect 2326 1132 2512 1176
rect 2566 1132 2752 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 834 1132
rect 886 1124 1074 1132
rect 1126 1124 1314 1132
rect 1366 1124 1554 1132
rect 1606 1124 1794 1132
rect 1846 1124 2034 1132
rect 2086 1124 2274 1132
rect 2326 1124 2514 1132
rect 2566 1124 2754 1132
rect 2806 1124 3000 1176
rect 0 1110 3000 1124
rect 110 987 160 1110
rect 110 753 112 987
rect 158 753 160 987
rect 110 700 160 753
rect 280 987 330 1040
rect 280 753 282 987
rect 328 753 330 987
rect 280 650 330 753
rect 450 987 500 1110
rect 450 753 452 987
rect 498 753 500 987
rect 450 700 500 753
rect 620 987 670 1040
rect 620 753 622 987
rect 668 753 670 987
rect 620 650 670 753
rect 790 987 840 1110
rect 790 753 792 987
rect 838 753 840 987
rect 790 700 840 753
rect 960 987 1010 1040
rect 960 753 962 987
rect 1008 753 1010 987
rect 960 650 1010 753
rect 1130 987 1180 1110
rect 1130 753 1132 987
rect 1178 753 1180 987
rect 1130 700 1180 753
rect 1300 987 1350 1040
rect 1300 753 1302 987
rect 1348 753 1350 987
rect 1300 650 1350 753
rect 1470 987 1520 1110
rect 1470 753 1472 987
rect 1518 753 1520 987
rect 1470 700 1520 753
rect 1640 987 1690 1040
rect 1640 753 1642 987
rect 1688 753 1690 987
rect 1640 650 1690 753
rect 1810 987 1860 1110
rect 1810 753 1812 987
rect 1858 753 1860 987
rect 1810 700 1860 753
rect 1980 987 2030 1040
rect 1980 753 1982 987
rect 2028 753 2030 987
rect 1980 650 2030 753
rect 2150 987 2200 1110
rect 2150 753 2152 987
rect 2198 753 2200 987
rect 2150 700 2200 753
rect 2320 987 2370 1040
rect 2320 753 2322 987
rect 2368 753 2370 987
rect 2320 650 2370 753
rect 2490 987 2540 1110
rect 2490 753 2492 987
rect 2538 753 2540 987
rect 2490 700 2540 753
rect 2660 987 2710 1040
rect 2660 753 2662 987
rect 2708 760 2710 987
rect 2830 987 2880 1110
rect 2708 756 2770 760
rect 2660 704 2694 753
rect 2746 704 2770 756
rect 2660 700 2770 704
rect 2830 753 2832 987
rect 2878 753 2880 987
rect 2830 700 2880 753
rect 2660 650 2710 700
rect 280 600 2710 650
rect 80 498 180 500
rect 80 496 112 498
rect 80 444 104 496
rect 158 452 180 498
rect 156 444 180 452
rect 80 440 180 444
rect 280 460 330 600
rect 620 460 670 600
rect 960 460 1010 600
rect 1300 460 1350 600
rect 1640 460 1690 600
rect 1980 460 2030 600
rect 2320 460 2370 600
rect 2660 460 2710 600
rect 280 410 2710 460
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 410
rect 280 252 282 298
rect 328 252 330 298
rect 280 190 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 410
rect 620 252 622 298
rect 668 252 670 298
rect 620 190 670 252
rect 790 298 840 360
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 960 298 1010 410
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 190 1010 252
rect 1130 298 1180 360
rect 1130 252 1132 298
rect 1178 252 1180 298
rect 1130 120 1180 252
rect 1300 298 1350 410
rect 1300 252 1302 298
rect 1348 252 1350 298
rect 1300 190 1350 252
rect 1470 298 1520 360
rect 1470 252 1472 298
rect 1518 252 1520 298
rect 1470 120 1520 252
rect 1640 298 1690 410
rect 1640 252 1642 298
rect 1688 252 1690 298
rect 1640 190 1690 252
rect 1810 298 1860 360
rect 1810 252 1812 298
rect 1858 252 1860 298
rect 1810 120 1860 252
rect 1980 298 2030 410
rect 1980 252 1982 298
rect 2028 252 2030 298
rect 1980 190 2030 252
rect 2150 298 2200 360
rect 2150 252 2152 298
rect 2198 252 2200 298
rect 2150 120 2200 252
rect 2320 298 2370 410
rect 2320 252 2322 298
rect 2368 252 2370 298
rect 2320 190 2370 252
rect 2490 298 2540 360
rect 2490 252 2492 298
rect 2538 252 2540 298
rect 2490 120 2540 252
rect 2660 298 2710 410
rect 2660 252 2662 298
rect 2708 252 2710 298
rect 2660 190 2710 252
rect 2830 298 2880 360
rect 2830 252 2832 298
rect 2878 252 2880 298
rect 2830 120 2880 252
rect 0 106 3000 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 1366 98 1554 106
rect 1606 98 1794 106
rect 1846 98 2034 106
rect 2086 98 2274 106
rect 2326 98 2514 106
rect 2566 98 2754 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1552 98
rect 1606 54 1792 98
rect 1846 54 2032 98
rect 2086 54 2272 98
rect 2326 54 2512 98
rect 2566 54 2752 98
rect 2806 54 3000 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1552 54
rect 1598 52 1792 54
rect 1838 52 2032 54
rect 2078 52 2272 54
rect 2318 52 2512 54
rect 2558 52 2752 54
rect 2798 52 3000 54
rect 0 0 3000 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 834 1132 878 1176
rect 878 1132 886 1176
rect 1074 1132 1118 1176
rect 1118 1132 1126 1176
rect 1314 1132 1358 1176
rect 1358 1132 1366 1176
rect 1554 1132 1598 1176
rect 1598 1132 1606 1176
rect 1794 1132 1838 1176
rect 1838 1132 1846 1176
rect 2034 1132 2078 1176
rect 2078 1132 2086 1176
rect 2274 1132 2318 1176
rect 2318 1132 2326 1176
rect 2514 1132 2558 1176
rect 2558 1132 2566 1176
rect 2754 1132 2798 1176
rect 2798 1132 2806 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 834 1124 886 1132
rect 1074 1124 1126 1132
rect 1314 1124 1366 1132
rect 1554 1124 1606 1132
rect 1794 1124 1846 1132
rect 2034 1124 2086 1132
rect 2274 1124 2326 1132
rect 2514 1124 2566 1132
rect 2754 1124 2806 1132
rect 2694 753 2708 756
rect 2708 753 2746 756
rect 2694 704 2746 753
rect 104 452 112 496
rect 112 452 156 496
rect 104 444 156 452
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 1554 98 1606 106
rect 1794 98 1846 106
rect 2034 98 2086 106
rect 2274 98 2326 106
rect 2514 98 2566 106
rect 2754 98 2806 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
rect 1554 54 1598 98
rect 1598 54 1606 98
rect 1794 54 1838 98
rect 1838 54 1846 98
rect 2034 54 2078 98
rect 2078 54 2086 98
rect 2274 54 2318 98
rect 2318 54 2326 98
rect 2514 54 2558 98
rect 2558 54 2566 98
rect 2754 54 2798 98
rect 2798 54 2806 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 820 1180 900 1190
rect 1060 1180 1140 1190
rect 1300 1180 1380 1190
rect 1540 1180 1620 1190
rect 1780 1180 1860 1190
rect 2020 1180 2100 1190
rect 2260 1180 2340 1190
rect 2500 1180 2580 1190
rect 2740 1180 2820 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 810 1176 910 1180
rect 810 1124 834 1176
rect 886 1124 910 1176
rect 810 1120 910 1124
rect 1050 1176 1150 1180
rect 1050 1124 1074 1176
rect 1126 1124 1150 1176
rect 1050 1120 1150 1124
rect 1290 1176 1390 1180
rect 1290 1124 1314 1176
rect 1366 1124 1390 1176
rect 1290 1120 1390 1124
rect 1530 1176 1630 1180
rect 1530 1124 1554 1176
rect 1606 1124 1630 1176
rect 1530 1120 1630 1124
rect 1770 1176 1870 1180
rect 1770 1124 1794 1176
rect 1846 1124 1870 1176
rect 1770 1120 1870 1124
rect 2010 1176 2110 1180
rect 2010 1124 2034 1176
rect 2086 1124 2110 1176
rect 2010 1120 2110 1124
rect 2250 1176 2350 1180
rect 2250 1124 2274 1176
rect 2326 1124 2350 1176
rect 2250 1120 2350 1124
rect 2490 1176 2590 1180
rect 2490 1124 2514 1176
rect 2566 1124 2590 1176
rect 2490 1120 2590 1124
rect 2730 1176 2830 1180
rect 2730 1124 2754 1176
rect 2806 1124 2830 1176
rect 2730 1120 2830 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 820 1110 900 1120
rect 1060 1110 1140 1120
rect 1300 1110 1380 1120
rect 1540 1110 1620 1120
rect 1780 1110 1860 1120
rect 2020 1110 2100 1120
rect 2260 1110 2340 1120
rect 2500 1110 2580 1120
rect 2740 1110 2820 1120
rect 2680 760 2760 770
rect 2670 756 2770 760
rect 2670 704 2694 756
rect 2746 704 2770 756
rect 2670 700 2770 704
rect 2680 690 2760 700
rect 80 496 180 510
rect 80 444 104 496
rect 156 444 180 496
rect 80 430 180 444
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 1540 110 1620 120
rect 1780 110 1860 120
rect 2020 110 2100 120
rect 2260 110 2340 120
rect 2500 110 2580 120
rect 2740 110 2820 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 1530 106 1630 110
rect 1530 54 1554 106
rect 1606 54 1630 106
rect 1530 50 1630 54
rect 1770 106 1870 110
rect 1770 54 1794 106
rect 1846 54 1870 106
rect 1770 50 1870 54
rect 2010 106 2110 110
rect 2010 54 2034 106
rect 2086 54 2110 106
rect 2010 50 2110 54
rect 2250 106 2350 110
rect 2250 54 2274 106
rect 2326 54 2350 106
rect 2250 50 2350 54
rect 2490 106 2590 110
rect 2490 54 2514 106
rect 2566 54 2590 106
rect 2490 50 2590 54
rect 2730 106 2830 110
rect 2730 54 2754 106
rect 2806 54 2830 106
rect 2730 50 2830 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
rect 1540 40 1620 50
rect 1780 40 1860 50
rect 2020 40 2100 50
rect 2260 40 2340 50
rect 2500 40 2580 50
rect 2740 40 2820 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 80 430 180 510 4 A
port 1 nsew signal input
rlabel metal2 s 2680 690 2760 770 4 Y
port 2 nsew signal output
rlabel metal1 s 80 440 180 500 1 A
port 1 nsew signal input
rlabel metal2 s 90 1120 190 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 820 1110 900 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 810 1120 910 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1060 1110 1140 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1050 1120 1150 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1300 1110 1380 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1290 1120 1390 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1540 1110 1620 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1530 1120 1630 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1780 1110 1860 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1770 1120 1870 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2020 1110 2100 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2010 1120 2110 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2260 1110 2340 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2250 1120 2350 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2500 1110 2580 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2490 1120 2590 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2740 1110 2820 1190 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 2730 1120 2830 1180 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 700 160 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 700 500 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 700 840 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1130 700 1180 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1470 700 1520 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1810 700 1860 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2150 700 2200 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2490 700 2540 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2830 700 2880 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1110 3000 1230 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1540 40 1620 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1530 50 1630 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1780 40 1860 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1770 50 1870 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2020 40 2100 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2010 50 2110 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2260 40 2340 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2250 50 2350 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2500 40 2580 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2490 50 2590 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2740 40 2820 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2730 50 2830 110 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 0 160 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 0 500 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 0 840 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1130 0 1180 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1470 0 1520 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1810 0 1860 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2150 0 2200 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2490 0 2540 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 2830 0 2880 360 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 3000 120 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 2670 700 2770 760 1 Y
port 2 nsew signal output
rlabel metal1 s 280 190 330 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 620 190 670 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 960 190 1010 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 190 1350 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 1640 190 1690 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 1980 190 2030 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 2320 190 2370 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 280 410 2710 460 1 Y
port 2 nsew signal output
rlabel metal1 s 280 600 2710 650 1 Y
port 2 nsew signal output
rlabel metal1 s 2660 190 2710 1040 1 Y
port 2 nsew signal output
rlabel metal1 s 2660 700 2770 760 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3000 1230
string GDS_END 221814
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 199254
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
