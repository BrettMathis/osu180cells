magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 320
<< mvndiff >>
rect -88 307 0 320
rect -88 261 -75 307
rect -29 261 0 307
rect -88 183 0 261
rect -88 137 -75 183
rect -29 137 0 183
rect -88 59 0 137
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 307 208 320
rect 120 261 149 307
rect 195 261 208 307
rect 120 183 208 261
rect 120 137 149 183
rect 195 137 208 183
rect 120 59 208 137
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 261 -29 307
rect -75 137 -29 183
rect -75 13 -29 59
rect 149 261 195 307
rect 149 137 195 183
rect 149 13 195 59
<< polysilicon >>
rect 0 320 120 364
rect 0 -44 120 0
<< metal1 >>
rect -75 307 -29 320
rect -75 183 -29 261
rect -75 59 -29 137
rect -75 0 -29 13
rect 149 307 195 320
rect 149 183 195 261
rect 149 59 195 137
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 160 -52 160 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 160 172 160 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 374180
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 372900
<< end >>
