magic
tech gf180mcuA
timestamp 1669390400
<< metal1 >>
rect 0 111 290 123
rect 28 95 33 111
rect 100 82 105 111
rect 172 95 177 111
rect 208 70 213 111
rect 50 65 179 66
rect 50 63 188 65
rect 35 57 45 63
rect 50 60 190 63
rect 78 46 84 60
rect 76 40 86 46
rect 121 45 127 60
rect 180 57 190 60
rect 119 39 129 45
rect 28 12 33 30
rect 100 12 105 28
rect 172 12 177 30
rect 240 76 245 104
rect 257 81 262 111
rect 274 90 279 104
rect 274 83 285 90
rect 274 82 284 83
rect 240 70 269 76
rect 208 12 213 28
rect 261 42 267 70
rect 240 37 267 42
rect 240 19 245 37
rect 257 12 262 32
rect 274 19 279 82
rect 0 0 290 12
<< obsm1 >>
rect 11 47 16 104
rect 66 90 77 104
rect 10 46 16 47
rect 8 40 16 46
rect 10 38 16 40
rect 11 19 16 38
rect 21 84 77 90
rect 21 66 27 84
rect 128 84 139 104
rect 161 84 171 90
rect 128 82 134 84
rect 163 82 169 84
rect 189 75 194 104
rect 189 70 200 75
rect 21 60 29 66
rect 21 41 27 60
rect 94 46 100 47
rect 21 36 45 41
rect 54 40 64 46
rect 92 40 102 46
rect 195 50 200 70
rect 139 46 145 48
rect 138 40 151 46
rect 161 44 171 50
rect 189 44 200 50
rect 139 38 151 40
rect 40 33 45 36
rect 40 28 77 33
rect 126 28 139 33
rect 145 29 151 38
rect 66 19 77 28
rect 128 19 139 28
rect 189 29 195 44
rect 212 39 218 59
rect 225 57 230 104
rect 225 51 253 57
rect 210 33 220 39
rect 189 19 194 29
rect 225 19 230 51
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 177 112 187 118
rect 201 112 211 118
rect 225 112 235 118
rect 249 112 259 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 35 63 45 64
rect 34 57 46 63
rect 35 56 45 57
rect 276 89 284 90
rect 181 63 189 64
rect 180 57 190 63
rect 275 83 285 89
rect 276 82 284 83
rect 260 76 268 77
rect 259 70 269 76
rect 260 69 268 70
rect 181 56 189 57
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< obsm2 >>
rect 56 98 151 104
rect 56 47 62 98
rect 128 91 134 92
rect 127 83 135 91
rect 9 46 17 47
rect 55 46 64 47
rect 93 46 101 47
rect 8 40 18 46
rect 54 40 64 46
rect 92 40 102 46
rect 9 39 17 40
rect 55 39 64 40
rect 93 39 101 40
rect 10 27 16 39
rect 94 27 100 39
rect 128 34 134 83
rect 145 38 151 98
rect 162 90 170 91
rect 161 84 229 90
rect 162 83 170 84
rect 163 51 169 83
rect 223 57 229 84
rect 244 57 252 58
rect 223 51 253 57
rect 162 50 170 51
rect 244 50 252 51
rect 161 44 171 50
rect 162 43 170 44
rect 211 39 219 40
rect 144 37 152 38
rect 188 37 196 38
rect 127 33 135 34
rect 126 27 135 33
rect 143 31 198 37
rect 204 33 220 39
rect 204 32 219 33
rect 144 30 152 31
rect 188 30 196 31
rect 10 21 100 27
rect 127 26 135 27
rect 128 24 135 26
rect 204 24 210 32
rect 128 18 210 24
<< labels >>
rlabel metal2 s 181 56 189 64 6 CLK
port 4 nsew clock input
rlabel metal2 s 180 57 190 63 6 CLK
port 4 nsew clock input
rlabel metal1 s 78 40 84 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 76 40 86 46 6 CLK
port 4 nsew clock input
rlabel metal1 s 121 39 127 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 119 39 129 45 6 CLK
port 4 nsew clock input
rlabel metal1 s 50 60 179 66 6 CLK
port 4 nsew clock input
rlabel metal1 s 50 60 188 65 6 CLK
port 4 nsew clock input
rlabel metal1 s 180 57 190 63 6 CLK
port 4 nsew clock input
rlabel metal2 s 35 56 45 64 6 D
port 1 nsew signal input
rlabel metal2 s 34 57 46 63 6 D
port 1 nsew signal input
rlabel metal1 s 35 57 45 63 6 D
port 1 nsew signal input
rlabel metal2 s 276 82 284 90 6 Q
port 2 nsew signal output
rlabel metal2 s 275 83 285 89 6 Q
port 2 nsew signal output
rlabel metal1 s 274 19 279 104 6 Q
port 2 nsew signal output
rlabel metal1 s 274 82 284 90 6 Q
port 2 nsew signal output
rlabel metal1 s 274 83 285 90 6 Q
port 2 nsew signal output
rlabel metal2 s 260 69 268 77 6 QN
port 3 nsew signal output
rlabel metal2 s 259 70 269 76 6 QN
port 3 nsew signal output
rlabel metal1 s 240 19 245 42 6 QN
port 3 nsew signal output
rlabel metal1 s 240 70 245 104 6 QN
port 3 nsew signal output
rlabel metal1 s 240 37 267 42 6 QN
port 3 nsew signal output
rlabel metal1 s 261 37 267 76 6 QN
port 3 nsew signal output
rlabel metal1 s 240 70 269 76 6 QN
port 3 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 178 111 186 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 177 112 187 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 202 111 210 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 201 112 211 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 226 111 234 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 225 112 235 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 250 111 258 119 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 249 112 259 118 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 28 95 33 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 100 82 105 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 172 95 177 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 208 70 213 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 257 81 262 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 111 290 123 6 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 28 0 33 30 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 100 0 105 28 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 172 0 177 30 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 208 0 213 28 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 257 0 262 32 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 290 12 6 VSS
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 290 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 249564
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 221870
<< end >>
