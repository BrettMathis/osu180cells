magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -384 16828 1102 16875
rect -384 16776 39 16828
rect 91 16776 147 16828
rect 199 16776 255 16828
rect 307 16776 363 16828
rect 415 16776 471 16828
rect 523 16776 579 16828
rect 631 16776 687 16828
rect 739 16776 795 16828
rect 847 16776 903 16828
rect 955 16776 1011 16828
rect 1063 16776 1102 16828
rect -384 16720 1102 16776
rect -384 16668 39 16720
rect 91 16668 147 16720
rect 199 16668 255 16720
rect 307 16668 363 16720
rect 415 16668 471 16720
rect 523 16668 579 16720
rect 631 16668 687 16720
rect 739 16668 795 16720
rect 847 16668 903 16720
rect 955 16668 1011 16720
rect 1063 16668 1102 16720
rect -384 16623 1102 16668
rect 1450 16118 3254 16130
rect 1450 16066 1462 16118
rect 1514 16066 1570 16118
rect 1622 16066 1678 16118
rect 1730 16066 1786 16118
rect 1838 16066 1894 16118
rect 1946 16066 2002 16118
rect 2054 16066 2110 16118
rect 2162 16066 2218 16118
rect 2270 16066 2326 16118
rect 2378 16066 2434 16118
rect 2486 16066 2542 16118
rect 2594 16066 2650 16118
rect 2702 16066 2758 16118
rect 2810 16066 2866 16118
rect 2918 16066 2974 16118
rect 3026 16066 3082 16118
rect 3134 16066 3190 16118
rect 3242 16066 3254 16118
rect 1450 16010 3254 16066
rect 1450 15958 1462 16010
rect 1514 15958 1570 16010
rect 1622 15958 1678 16010
rect 1730 15958 1786 16010
rect 1838 15958 1894 16010
rect 1946 15958 2002 16010
rect 2054 15958 2110 16010
rect 2162 15958 2218 16010
rect 2270 15958 2326 16010
rect 2378 15958 2434 16010
rect 2486 15958 2542 16010
rect 2594 15958 2650 16010
rect 2702 15958 2758 16010
rect 2810 15958 2866 16010
rect 2918 15958 2974 16010
rect 3026 15958 3082 16010
rect 3134 15958 3190 16010
rect 3242 15958 3254 16010
rect 1450 15946 3254 15958
rect 5317 16118 6365 16130
rect 5317 16066 5329 16118
rect 5381 16066 5437 16118
rect 5489 16066 5545 16118
rect 5597 16066 5653 16118
rect 5705 16066 5761 16118
rect 5813 16066 5869 16118
rect 5921 16066 5977 16118
rect 6029 16066 6085 16118
rect 6137 16066 6193 16118
rect 6245 16066 6301 16118
rect 6353 16066 6365 16118
rect 5317 16010 6365 16066
rect 5317 15958 5329 16010
rect 5381 15958 5437 16010
rect 5489 15958 5545 16010
rect 5597 15958 5653 16010
rect 5705 15958 5761 16010
rect 5813 15958 5869 16010
rect 5921 15958 5977 16010
rect 6029 15958 6085 16010
rect 6137 15958 6193 16010
rect 6245 15958 6301 16010
rect 6353 15958 6365 16010
rect 5317 15946 6365 15958
rect 7694 16118 9498 16130
rect 7694 16066 7706 16118
rect 7758 16066 7814 16118
rect 7866 16066 7922 16118
rect 7974 16066 8030 16118
rect 8082 16066 8138 16118
rect 8190 16066 8246 16118
rect 8298 16066 8354 16118
rect 8406 16066 8462 16118
rect 8514 16066 8570 16118
rect 8622 16066 8678 16118
rect 8730 16066 8786 16118
rect 8838 16066 8894 16118
rect 8946 16066 9002 16118
rect 9054 16066 9110 16118
rect 9162 16066 9218 16118
rect 9270 16066 9326 16118
rect 9378 16066 9434 16118
rect 9486 16066 9498 16118
rect 7694 16010 9498 16066
rect 7694 15958 7706 16010
rect 7758 15958 7814 16010
rect 7866 15958 7922 16010
rect 7974 15958 8030 16010
rect 8082 15958 8138 16010
rect 8190 15958 8246 16010
rect 8298 15958 8354 16010
rect 8406 15958 8462 16010
rect 8514 15958 8570 16010
rect 8622 15958 8678 16010
rect 8730 15958 8786 16010
rect 8838 15958 8894 16010
rect 8946 15958 9002 16010
rect 9054 15958 9110 16010
rect 9162 15958 9218 16010
rect 9270 15958 9326 16010
rect 9378 15958 9434 16010
rect 9486 15958 9498 16010
rect 7694 15946 9498 15958
rect 1446 10381 3258 10393
rect 1446 10329 1458 10381
rect 1510 10329 1582 10381
rect 1634 10329 1706 10381
rect 1758 10329 1830 10381
rect 1882 10329 1954 10381
rect 2006 10329 2078 10381
rect 2130 10329 2202 10381
rect 2254 10329 2326 10381
rect 2378 10329 2450 10381
rect 2502 10329 2574 10381
rect 2626 10329 2698 10381
rect 2750 10329 2822 10381
rect 2874 10329 2946 10381
rect 2998 10329 3070 10381
rect 3122 10329 3194 10381
rect 3246 10329 3258 10381
rect 1446 10257 3258 10329
rect 1446 10205 1458 10257
rect 1510 10205 1582 10257
rect 1634 10205 1706 10257
rect 1758 10205 1830 10257
rect 1882 10205 1954 10257
rect 2006 10205 2078 10257
rect 2130 10205 2202 10257
rect 2254 10205 2326 10257
rect 2378 10205 2450 10257
rect 2502 10205 2574 10257
rect 2626 10205 2698 10257
rect 2750 10205 2822 10257
rect 2874 10205 2946 10257
rect 2998 10205 3070 10257
rect 3122 10205 3194 10257
rect 3246 10205 3258 10257
rect 1446 10133 3258 10205
rect 1446 10081 1458 10133
rect 1510 10081 1582 10133
rect 1634 10081 1706 10133
rect 1758 10081 1830 10133
rect 1882 10081 1954 10133
rect 2006 10081 2078 10133
rect 2130 10081 2202 10133
rect 2254 10081 2326 10133
rect 2378 10081 2450 10133
rect 2502 10081 2574 10133
rect 2626 10081 2698 10133
rect 2750 10081 2822 10133
rect 2874 10081 2946 10133
rect 2998 10081 3070 10133
rect 3122 10081 3194 10133
rect 3246 10081 3258 10133
rect 1446 10009 3258 10081
rect 1446 9957 1458 10009
rect 1510 9957 1582 10009
rect 1634 9957 1706 10009
rect 1758 9957 1830 10009
rect 1882 9957 1954 10009
rect 2006 9957 2078 10009
rect 2130 9957 2202 10009
rect 2254 9957 2326 10009
rect 2378 9957 2450 10009
rect 2502 9957 2574 10009
rect 2626 9957 2698 10009
rect 2750 9957 2822 10009
rect 2874 9957 2946 10009
rect 2998 9957 3070 10009
rect 3122 9957 3194 10009
rect 3246 9957 3258 10009
rect 1446 9885 3258 9957
rect 1446 9833 1458 9885
rect 1510 9833 1582 9885
rect 1634 9833 1706 9885
rect 1758 9833 1830 9885
rect 1882 9833 1954 9885
rect 2006 9833 2078 9885
rect 2130 9833 2202 9885
rect 2254 9833 2326 9885
rect 2378 9833 2450 9885
rect 2502 9833 2574 9885
rect 2626 9833 2698 9885
rect 2750 9833 2822 9885
rect 2874 9833 2946 9885
rect 2998 9833 3070 9885
rect 3122 9833 3194 9885
rect 3246 9833 3258 9885
rect 1446 9761 3258 9833
rect 1446 9709 1458 9761
rect 1510 9709 1582 9761
rect 1634 9709 1706 9761
rect 1758 9709 1830 9761
rect 1882 9709 1954 9761
rect 2006 9709 2078 9761
rect 2130 9709 2202 9761
rect 2254 9709 2326 9761
rect 2378 9709 2450 9761
rect 2502 9709 2574 9761
rect 2626 9709 2698 9761
rect 2750 9709 2822 9761
rect 2874 9709 2946 9761
rect 2998 9709 3070 9761
rect 3122 9709 3194 9761
rect 3246 9709 3258 9761
rect 1446 9697 3258 9709
rect 5307 10381 6375 10393
rect 5307 10329 5319 10381
rect 5371 10329 5443 10381
rect 5495 10329 5567 10381
rect 5619 10329 5691 10381
rect 5743 10329 5815 10381
rect 5867 10329 5939 10381
rect 5991 10329 6063 10381
rect 6115 10329 6187 10381
rect 6239 10329 6311 10381
rect 6363 10329 6375 10381
rect 5307 10257 6375 10329
rect 5307 10205 5319 10257
rect 5371 10205 5443 10257
rect 5495 10205 5567 10257
rect 5619 10205 5691 10257
rect 5743 10205 5815 10257
rect 5867 10205 5939 10257
rect 5991 10205 6063 10257
rect 6115 10205 6187 10257
rect 6239 10205 6311 10257
rect 6363 10205 6375 10257
rect 5307 10133 6375 10205
rect 5307 10081 5319 10133
rect 5371 10081 5443 10133
rect 5495 10081 5567 10133
rect 5619 10081 5691 10133
rect 5743 10081 5815 10133
rect 5867 10081 5939 10133
rect 5991 10081 6063 10133
rect 6115 10081 6187 10133
rect 6239 10081 6311 10133
rect 6363 10081 6375 10133
rect 5307 10009 6375 10081
rect 5307 9957 5319 10009
rect 5371 9957 5443 10009
rect 5495 9957 5567 10009
rect 5619 9957 5691 10009
rect 5743 9957 5815 10009
rect 5867 9957 5939 10009
rect 5991 9957 6063 10009
rect 6115 9957 6187 10009
rect 6239 9957 6311 10009
rect 6363 9957 6375 10009
rect 5307 9885 6375 9957
rect 5307 9833 5319 9885
rect 5371 9833 5443 9885
rect 5495 9833 5567 9885
rect 5619 9833 5691 9885
rect 5743 9833 5815 9885
rect 5867 9833 5939 9885
rect 5991 9833 6063 9885
rect 6115 9833 6187 9885
rect 6239 9833 6311 9885
rect 6363 9833 6375 9885
rect 5307 9761 6375 9833
rect 5307 9709 5319 9761
rect 5371 9709 5443 9761
rect 5495 9709 5567 9761
rect 5619 9709 5691 9761
rect 5743 9709 5815 9761
rect 5867 9709 5939 9761
rect 5991 9709 6063 9761
rect 6115 9709 6187 9761
rect 6239 9709 6311 9761
rect 6363 9709 6375 9761
rect 5307 9697 6375 9709
rect 7690 10381 9502 10393
rect 7690 10329 7702 10381
rect 7754 10329 7826 10381
rect 7878 10329 7950 10381
rect 8002 10329 8074 10381
rect 8126 10329 8198 10381
rect 8250 10329 8322 10381
rect 8374 10329 8446 10381
rect 8498 10329 8570 10381
rect 8622 10329 8694 10381
rect 8746 10329 8818 10381
rect 8870 10329 8942 10381
rect 8994 10329 9066 10381
rect 9118 10329 9190 10381
rect 9242 10329 9314 10381
rect 9366 10329 9438 10381
rect 9490 10329 9502 10381
rect 7690 10257 9502 10329
rect 7690 10205 7702 10257
rect 7754 10205 7826 10257
rect 7878 10205 7950 10257
rect 8002 10205 8074 10257
rect 8126 10205 8198 10257
rect 8250 10205 8322 10257
rect 8374 10205 8446 10257
rect 8498 10205 8570 10257
rect 8622 10205 8694 10257
rect 8746 10205 8818 10257
rect 8870 10205 8942 10257
rect 8994 10205 9066 10257
rect 9118 10205 9190 10257
rect 9242 10205 9314 10257
rect 9366 10205 9438 10257
rect 9490 10205 9502 10257
rect 7690 10133 9502 10205
rect 7690 10081 7702 10133
rect 7754 10081 7826 10133
rect 7878 10081 7950 10133
rect 8002 10081 8074 10133
rect 8126 10081 8198 10133
rect 8250 10081 8322 10133
rect 8374 10081 8446 10133
rect 8498 10081 8570 10133
rect 8622 10081 8694 10133
rect 8746 10081 8818 10133
rect 8870 10081 8942 10133
rect 8994 10081 9066 10133
rect 9118 10081 9190 10133
rect 9242 10081 9314 10133
rect 9366 10081 9438 10133
rect 9490 10081 9502 10133
rect 7690 10009 9502 10081
rect 7690 9957 7702 10009
rect 7754 9957 7826 10009
rect 7878 9957 7950 10009
rect 8002 9957 8074 10009
rect 8126 9957 8198 10009
rect 8250 9957 8322 10009
rect 8374 9957 8446 10009
rect 8498 9957 8570 10009
rect 8622 9957 8694 10009
rect 8746 9957 8818 10009
rect 8870 9957 8942 10009
rect 8994 9957 9066 10009
rect 9118 9957 9190 10009
rect 9242 9957 9314 10009
rect 9366 9957 9438 10009
rect 9490 9957 9502 10009
rect 7690 9885 9502 9957
rect 7690 9833 7702 9885
rect 7754 9833 7826 9885
rect 7878 9833 7950 9885
rect 8002 9833 8074 9885
rect 8126 9833 8198 9885
rect 8250 9833 8322 9885
rect 8374 9833 8446 9885
rect 8498 9833 8570 9885
rect 8622 9833 8694 9885
rect 8746 9833 8818 9885
rect 8870 9833 8942 9885
rect 8994 9833 9066 9885
rect 9118 9833 9190 9885
rect 9242 9833 9314 9885
rect 9366 9833 9438 9885
rect 9490 9833 9502 9885
rect 7690 9761 9502 9833
rect 7690 9709 7702 9761
rect 7754 9709 7826 9761
rect 7878 9709 7950 9761
rect 8002 9709 8074 9761
rect 8126 9709 8198 9761
rect 8250 9709 8322 9761
rect 8374 9709 8446 9761
rect 8498 9709 8570 9761
rect 8622 9709 8694 9761
rect 8746 9709 8818 9761
rect 8870 9709 8942 9761
rect 8994 9709 9066 9761
rect 9118 9709 9190 9761
rect 9242 9709 9314 9761
rect 9366 9709 9438 9761
rect 9490 9709 9502 9761
rect 7690 9697 9502 9709
rect 1450 4034 3254 4046
rect 1450 3982 1462 4034
rect 1514 3982 1570 4034
rect 1622 3982 1678 4034
rect 1730 3982 1786 4034
rect 1838 3982 1894 4034
rect 1946 3982 2002 4034
rect 2054 3982 2110 4034
rect 2162 3982 2218 4034
rect 2270 3982 2326 4034
rect 2378 3982 2434 4034
rect 2486 3982 2542 4034
rect 2594 3982 2650 4034
rect 2702 3982 2758 4034
rect 2810 3982 2866 4034
rect 2918 3982 2974 4034
rect 3026 3982 3082 4034
rect 3134 3982 3190 4034
rect 3242 3982 3254 4034
rect 1450 3926 3254 3982
rect 1450 3874 1462 3926
rect 1514 3874 1570 3926
rect 1622 3874 1678 3926
rect 1730 3874 1786 3926
rect 1838 3874 1894 3926
rect 1946 3874 2002 3926
rect 2054 3874 2110 3926
rect 2162 3874 2218 3926
rect 2270 3874 2326 3926
rect 2378 3874 2434 3926
rect 2486 3874 2542 3926
rect 2594 3874 2650 3926
rect 2702 3874 2758 3926
rect 2810 3874 2866 3926
rect 2918 3874 2974 3926
rect 3026 3874 3082 3926
rect 3134 3874 3190 3926
rect 3242 3874 3254 3926
rect 1450 3862 3254 3874
rect 5317 4034 6365 4046
rect 5317 3982 5329 4034
rect 5381 3982 5437 4034
rect 5489 3982 5545 4034
rect 5597 3982 5653 4034
rect 5705 3982 5761 4034
rect 5813 3982 5869 4034
rect 5921 3982 5977 4034
rect 6029 3982 6085 4034
rect 6137 3982 6193 4034
rect 6245 3982 6301 4034
rect 6353 3982 6365 4034
rect 5317 3926 6365 3982
rect 5317 3874 5329 3926
rect 5381 3874 5437 3926
rect 5489 3874 5545 3926
rect 5597 3874 5653 3926
rect 5705 3874 5761 3926
rect 5813 3874 5869 3926
rect 5921 3874 5977 3926
rect 6029 3874 6085 3926
rect 6137 3874 6193 3926
rect 6245 3874 6301 3926
rect 6353 3874 6365 3926
rect 5317 3862 6365 3874
rect 7694 4034 9498 4046
rect 7694 3982 7706 4034
rect 7758 3982 7814 4034
rect 7866 3982 7922 4034
rect 7974 3982 8030 4034
rect 8082 3982 8138 4034
rect 8190 3982 8246 4034
rect 8298 3982 8354 4034
rect 8406 3982 8462 4034
rect 8514 3982 8570 4034
rect 8622 3982 8678 4034
rect 8730 3982 8786 4034
rect 8838 3982 8894 4034
rect 8946 3982 9002 4034
rect 9054 3982 9110 4034
rect 9162 3982 9218 4034
rect 9270 3982 9326 4034
rect 9378 3982 9434 4034
rect 9486 3982 9498 4034
rect 7694 3926 9498 3982
rect 7694 3874 7706 3926
rect 7758 3874 7814 3926
rect 7866 3874 7922 3926
rect 7974 3874 8030 3926
rect 8082 3874 8138 3926
rect 8190 3874 8246 3926
rect 8298 3874 8354 3926
rect 8406 3874 8462 3926
rect 8514 3874 8570 3926
rect 8622 3874 8678 3926
rect 8730 3874 8786 3926
rect 8838 3874 8894 3926
rect 8946 3874 9002 3926
rect 9054 3874 9110 3926
rect 9162 3874 9218 3926
rect 9270 3874 9326 3926
rect 9378 3874 9434 3926
rect 9486 3874 9498 3926
rect 7694 3862 9498 3874
rect 124 3566 12876 3586
rect 124 3514 150 3566
rect 202 3514 258 3566
rect 310 3514 366 3566
rect 418 3514 474 3566
rect 526 3514 582 3566
rect 634 3514 690 3566
rect 742 3514 798 3566
rect 850 3514 906 3566
rect 958 3514 1014 3566
rect 1066 3514 3390 3566
rect 3442 3514 3498 3566
rect 3550 3514 3606 3566
rect 3658 3514 3714 3566
rect 3766 3514 3822 3566
rect 3874 3514 3930 3566
rect 3982 3514 4038 3566
rect 4090 3514 4146 3566
rect 4198 3514 4254 3566
rect 4306 3514 4362 3566
rect 4414 3514 4470 3566
rect 4522 3514 4578 3566
rect 4630 3514 4686 3566
rect 4738 3514 4794 3566
rect 4846 3514 4902 3566
rect 4954 3514 5010 3566
rect 5062 3514 5118 3566
rect 5170 3514 6523 3566
rect 6575 3514 6631 3566
rect 6683 3514 6739 3566
rect 6791 3514 6847 3566
rect 6899 3514 6955 3566
rect 7007 3514 7063 3566
rect 7115 3514 7171 3566
rect 7223 3514 7279 3566
rect 7331 3514 7387 3566
rect 7439 3514 7495 3566
rect 7547 3514 9634 3566
rect 9686 3514 9742 3566
rect 9794 3514 9850 3566
rect 9902 3514 9958 3566
rect 10010 3514 10066 3566
rect 10118 3514 10174 3566
rect 10226 3514 10282 3566
rect 10334 3514 10390 3566
rect 10442 3514 10498 3566
rect 10550 3514 10606 3566
rect 10658 3514 10714 3566
rect 10766 3514 10822 3566
rect 10874 3514 10930 3566
rect 10982 3514 11038 3566
rect 11090 3514 11146 3566
rect 11198 3514 11254 3566
rect 11306 3514 11362 3566
rect 11414 3514 12876 3566
rect 124 3458 12876 3514
rect 124 3406 150 3458
rect 202 3406 258 3458
rect 310 3406 366 3458
rect 418 3406 474 3458
rect 526 3406 582 3458
rect 634 3406 690 3458
rect 742 3406 798 3458
rect 850 3406 906 3458
rect 958 3406 1014 3458
rect 1066 3406 3390 3458
rect 3442 3406 3498 3458
rect 3550 3406 3606 3458
rect 3658 3406 3714 3458
rect 3766 3406 3822 3458
rect 3874 3406 3930 3458
rect 3982 3406 4038 3458
rect 4090 3406 4146 3458
rect 4198 3406 4254 3458
rect 4306 3406 4362 3458
rect 4414 3406 4470 3458
rect 4522 3406 4578 3458
rect 4630 3406 4686 3458
rect 4738 3406 4794 3458
rect 4846 3406 4902 3458
rect 4954 3406 5010 3458
rect 5062 3406 5118 3458
rect 5170 3406 6523 3458
rect 6575 3406 6631 3458
rect 6683 3406 6739 3458
rect 6791 3406 6847 3458
rect 6899 3406 6955 3458
rect 7007 3406 7063 3458
rect 7115 3406 7171 3458
rect 7223 3406 7279 3458
rect 7331 3406 7387 3458
rect 7439 3406 7495 3458
rect 7547 3406 9634 3458
rect 9686 3406 9742 3458
rect 9794 3406 9850 3458
rect 9902 3406 9958 3458
rect 10010 3406 10066 3458
rect 10118 3406 10174 3458
rect 10226 3406 10282 3458
rect 10334 3406 10390 3458
rect 10442 3406 10498 3458
rect 10550 3406 10606 3458
rect 10658 3406 10714 3458
rect 10766 3406 10822 3458
rect 10874 3406 10930 3458
rect 10982 3406 11038 3458
rect 11090 3406 11146 3458
rect 11198 3406 11254 3458
rect 11306 3406 11362 3458
rect 11414 3406 12876 3458
rect 124 3386 12876 3406
rect 0 286 6716 306
rect 0 234 1462 286
rect 1514 234 1570 286
rect 1622 234 1678 286
rect 1730 234 1786 286
rect 1838 234 1894 286
rect 1946 234 2002 286
rect 2054 234 2110 286
rect 2162 234 2218 286
rect 2270 234 2326 286
rect 2378 234 2434 286
rect 2486 234 2542 286
rect 2594 234 2650 286
rect 2702 234 2758 286
rect 2810 234 2866 286
rect 2918 234 2974 286
rect 3026 234 3082 286
rect 3134 234 3190 286
rect 3242 234 5329 286
rect 5381 234 5437 286
rect 5489 234 5545 286
rect 5597 234 5653 286
rect 5705 234 5761 286
rect 5813 234 5869 286
rect 5921 234 5977 286
rect 6029 234 6085 286
rect 6137 234 6193 286
rect 6245 234 6301 286
rect 6353 234 6716 286
rect 0 178 6716 234
rect 0 126 1462 178
rect 1514 126 1570 178
rect 1622 126 1678 178
rect 1730 126 1786 178
rect 1838 126 1894 178
rect 1946 126 2002 178
rect 2054 126 2110 178
rect 2162 126 2218 178
rect 2270 126 2326 178
rect 2378 126 2434 178
rect 2486 126 2542 178
rect 2594 126 2650 178
rect 2702 126 2758 178
rect 2810 126 2866 178
rect 2918 126 2974 178
rect 3026 126 3082 178
rect 3134 126 3190 178
rect 3242 126 5329 178
rect 5381 126 5437 178
rect 5489 126 5545 178
rect 5597 126 5653 178
rect 5705 126 5761 178
rect 5813 126 5869 178
rect 5921 126 5977 178
rect 6029 126 6085 178
rect 6137 126 6193 178
rect 6245 126 6301 178
rect 6353 126 6716 178
rect 0 106 6716 126
rect 6892 286 12876 306
rect 6892 234 7904 286
rect 7956 234 8012 286
rect 8064 234 8120 286
rect 8172 234 8228 286
rect 8280 234 8336 286
rect 8388 234 8444 286
rect 8496 234 8552 286
rect 8604 234 8660 286
rect 8712 234 8768 286
rect 8820 234 8876 286
rect 8928 234 8984 286
rect 9036 234 9092 286
rect 9144 234 9200 286
rect 9252 234 9308 286
rect 9360 234 9416 286
rect 9468 234 11813 286
rect 11865 234 11921 286
rect 11973 234 12029 286
rect 12081 234 12137 286
rect 12189 234 12245 286
rect 12297 234 12353 286
rect 12405 234 12461 286
rect 12513 234 12569 286
rect 12621 234 12677 286
rect 12729 234 12785 286
rect 12837 234 12876 286
rect 6892 178 12876 234
rect 6892 126 7904 178
rect 7956 126 8012 178
rect 8064 126 8120 178
rect 8172 126 8228 178
rect 8280 126 8336 178
rect 8388 126 8444 178
rect 8496 126 8552 178
rect 8604 126 8660 178
rect 8712 126 8768 178
rect 8820 126 8876 178
rect 8928 126 8984 178
rect 9036 126 9092 178
rect 9144 126 9200 178
rect 9252 126 9308 178
rect 9360 126 9416 178
rect 9468 126 11813 178
rect 11865 126 11921 178
rect 11973 126 12029 178
rect 12081 126 12137 178
rect 12189 126 12245 178
rect 12297 126 12353 178
rect 12405 126 12461 178
rect 12513 126 12569 178
rect 12621 126 12677 178
rect 12729 126 12785 178
rect 12837 126 12876 178
rect 6892 106 12876 126
<< via1 >>
rect 39 16776 91 16828
rect 147 16776 199 16828
rect 255 16776 307 16828
rect 363 16776 415 16828
rect 471 16776 523 16828
rect 579 16776 631 16828
rect 687 16776 739 16828
rect 795 16776 847 16828
rect 903 16776 955 16828
rect 1011 16776 1063 16828
rect 39 16668 91 16720
rect 147 16668 199 16720
rect 255 16668 307 16720
rect 363 16668 415 16720
rect 471 16668 523 16720
rect 579 16668 631 16720
rect 687 16668 739 16720
rect 795 16668 847 16720
rect 903 16668 955 16720
rect 1011 16668 1063 16720
rect 1462 16066 1514 16118
rect 1570 16066 1622 16118
rect 1678 16066 1730 16118
rect 1786 16066 1838 16118
rect 1894 16066 1946 16118
rect 2002 16066 2054 16118
rect 2110 16066 2162 16118
rect 2218 16066 2270 16118
rect 2326 16066 2378 16118
rect 2434 16066 2486 16118
rect 2542 16066 2594 16118
rect 2650 16066 2702 16118
rect 2758 16066 2810 16118
rect 2866 16066 2918 16118
rect 2974 16066 3026 16118
rect 3082 16066 3134 16118
rect 3190 16066 3242 16118
rect 1462 15958 1514 16010
rect 1570 15958 1622 16010
rect 1678 15958 1730 16010
rect 1786 15958 1838 16010
rect 1894 15958 1946 16010
rect 2002 15958 2054 16010
rect 2110 15958 2162 16010
rect 2218 15958 2270 16010
rect 2326 15958 2378 16010
rect 2434 15958 2486 16010
rect 2542 15958 2594 16010
rect 2650 15958 2702 16010
rect 2758 15958 2810 16010
rect 2866 15958 2918 16010
rect 2974 15958 3026 16010
rect 3082 15958 3134 16010
rect 3190 15958 3242 16010
rect 5329 16066 5381 16118
rect 5437 16066 5489 16118
rect 5545 16066 5597 16118
rect 5653 16066 5705 16118
rect 5761 16066 5813 16118
rect 5869 16066 5921 16118
rect 5977 16066 6029 16118
rect 6085 16066 6137 16118
rect 6193 16066 6245 16118
rect 6301 16066 6353 16118
rect 5329 15958 5381 16010
rect 5437 15958 5489 16010
rect 5545 15958 5597 16010
rect 5653 15958 5705 16010
rect 5761 15958 5813 16010
rect 5869 15958 5921 16010
rect 5977 15958 6029 16010
rect 6085 15958 6137 16010
rect 6193 15958 6245 16010
rect 6301 15958 6353 16010
rect 7706 16066 7758 16118
rect 7814 16066 7866 16118
rect 7922 16066 7974 16118
rect 8030 16066 8082 16118
rect 8138 16066 8190 16118
rect 8246 16066 8298 16118
rect 8354 16066 8406 16118
rect 8462 16066 8514 16118
rect 8570 16066 8622 16118
rect 8678 16066 8730 16118
rect 8786 16066 8838 16118
rect 8894 16066 8946 16118
rect 9002 16066 9054 16118
rect 9110 16066 9162 16118
rect 9218 16066 9270 16118
rect 9326 16066 9378 16118
rect 9434 16066 9486 16118
rect 7706 15958 7758 16010
rect 7814 15958 7866 16010
rect 7922 15958 7974 16010
rect 8030 15958 8082 16010
rect 8138 15958 8190 16010
rect 8246 15958 8298 16010
rect 8354 15958 8406 16010
rect 8462 15958 8514 16010
rect 8570 15958 8622 16010
rect 8678 15958 8730 16010
rect 8786 15958 8838 16010
rect 8894 15958 8946 16010
rect 9002 15958 9054 16010
rect 9110 15958 9162 16010
rect 9218 15958 9270 16010
rect 9326 15958 9378 16010
rect 9434 15958 9486 16010
rect 1458 10329 1510 10381
rect 1582 10329 1634 10381
rect 1706 10329 1758 10381
rect 1830 10329 1882 10381
rect 1954 10329 2006 10381
rect 2078 10329 2130 10381
rect 2202 10329 2254 10381
rect 2326 10329 2378 10381
rect 2450 10329 2502 10381
rect 2574 10329 2626 10381
rect 2698 10329 2750 10381
rect 2822 10329 2874 10381
rect 2946 10329 2998 10381
rect 3070 10329 3122 10381
rect 3194 10329 3246 10381
rect 1458 10205 1510 10257
rect 1582 10205 1634 10257
rect 1706 10205 1758 10257
rect 1830 10205 1882 10257
rect 1954 10205 2006 10257
rect 2078 10205 2130 10257
rect 2202 10205 2254 10257
rect 2326 10205 2378 10257
rect 2450 10205 2502 10257
rect 2574 10205 2626 10257
rect 2698 10205 2750 10257
rect 2822 10205 2874 10257
rect 2946 10205 2998 10257
rect 3070 10205 3122 10257
rect 3194 10205 3246 10257
rect 1458 10081 1510 10133
rect 1582 10081 1634 10133
rect 1706 10081 1758 10133
rect 1830 10081 1882 10133
rect 1954 10081 2006 10133
rect 2078 10081 2130 10133
rect 2202 10081 2254 10133
rect 2326 10081 2378 10133
rect 2450 10081 2502 10133
rect 2574 10081 2626 10133
rect 2698 10081 2750 10133
rect 2822 10081 2874 10133
rect 2946 10081 2998 10133
rect 3070 10081 3122 10133
rect 3194 10081 3246 10133
rect 1458 9957 1510 10009
rect 1582 9957 1634 10009
rect 1706 9957 1758 10009
rect 1830 9957 1882 10009
rect 1954 9957 2006 10009
rect 2078 9957 2130 10009
rect 2202 9957 2254 10009
rect 2326 9957 2378 10009
rect 2450 9957 2502 10009
rect 2574 9957 2626 10009
rect 2698 9957 2750 10009
rect 2822 9957 2874 10009
rect 2946 9957 2998 10009
rect 3070 9957 3122 10009
rect 3194 9957 3246 10009
rect 1458 9833 1510 9885
rect 1582 9833 1634 9885
rect 1706 9833 1758 9885
rect 1830 9833 1882 9885
rect 1954 9833 2006 9885
rect 2078 9833 2130 9885
rect 2202 9833 2254 9885
rect 2326 9833 2378 9885
rect 2450 9833 2502 9885
rect 2574 9833 2626 9885
rect 2698 9833 2750 9885
rect 2822 9833 2874 9885
rect 2946 9833 2998 9885
rect 3070 9833 3122 9885
rect 3194 9833 3246 9885
rect 1458 9709 1510 9761
rect 1582 9709 1634 9761
rect 1706 9709 1758 9761
rect 1830 9709 1882 9761
rect 1954 9709 2006 9761
rect 2078 9709 2130 9761
rect 2202 9709 2254 9761
rect 2326 9709 2378 9761
rect 2450 9709 2502 9761
rect 2574 9709 2626 9761
rect 2698 9709 2750 9761
rect 2822 9709 2874 9761
rect 2946 9709 2998 9761
rect 3070 9709 3122 9761
rect 3194 9709 3246 9761
rect 5319 10329 5371 10381
rect 5443 10329 5495 10381
rect 5567 10329 5619 10381
rect 5691 10329 5743 10381
rect 5815 10329 5867 10381
rect 5939 10329 5991 10381
rect 6063 10329 6115 10381
rect 6187 10329 6239 10381
rect 6311 10329 6363 10381
rect 5319 10205 5371 10257
rect 5443 10205 5495 10257
rect 5567 10205 5619 10257
rect 5691 10205 5743 10257
rect 5815 10205 5867 10257
rect 5939 10205 5991 10257
rect 6063 10205 6115 10257
rect 6187 10205 6239 10257
rect 6311 10205 6363 10257
rect 5319 10081 5371 10133
rect 5443 10081 5495 10133
rect 5567 10081 5619 10133
rect 5691 10081 5743 10133
rect 5815 10081 5867 10133
rect 5939 10081 5991 10133
rect 6063 10081 6115 10133
rect 6187 10081 6239 10133
rect 6311 10081 6363 10133
rect 5319 9957 5371 10009
rect 5443 9957 5495 10009
rect 5567 9957 5619 10009
rect 5691 9957 5743 10009
rect 5815 9957 5867 10009
rect 5939 9957 5991 10009
rect 6063 9957 6115 10009
rect 6187 9957 6239 10009
rect 6311 9957 6363 10009
rect 5319 9833 5371 9885
rect 5443 9833 5495 9885
rect 5567 9833 5619 9885
rect 5691 9833 5743 9885
rect 5815 9833 5867 9885
rect 5939 9833 5991 9885
rect 6063 9833 6115 9885
rect 6187 9833 6239 9885
rect 6311 9833 6363 9885
rect 5319 9709 5371 9761
rect 5443 9709 5495 9761
rect 5567 9709 5619 9761
rect 5691 9709 5743 9761
rect 5815 9709 5867 9761
rect 5939 9709 5991 9761
rect 6063 9709 6115 9761
rect 6187 9709 6239 9761
rect 6311 9709 6363 9761
rect 7702 10329 7754 10381
rect 7826 10329 7878 10381
rect 7950 10329 8002 10381
rect 8074 10329 8126 10381
rect 8198 10329 8250 10381
rect 8322 10329 8374 10381
rect 8446 10329 8498 10381
rect 8570 10329 8622 10381
rect 8694 10329 8746 10381
rect 8818 10329 8870 10381
rect 8942 10329 8994 10381
rect 9066 10329 9118 10381
rect 9190 10329 9242 10381
rect 9314 10329 9366 10381
rect 9438 10329 9490 10381
rect 7702 10205 7754 10257
rect 7826 10205 7878 10257
rect 7950 10205 8002 10257
rect 8074 10205 8126 10257
rect 8198 10205 8250 10257
rect 8322 10205 8374 10257
rect 8446 10205 8498 10257
rect 8570 10205 8622 10257
rect 8694 10205 8746 10257
rect 8818 10205 8870 10257
rect 8942 10205 8994 10257
rect 9066 10205 9118 10257
rect 9190 10205 9242 10257
rect 9314 10205 9366 10257
rect 9438 10205 9490 10257
rect 7702 10081 7754 10133
rect 7826 10081 7878 10133
rect 7950 10081 8002 10133
rect 8074 10081 8126 10133
rect 8198 10081 8250 10133
rect 8322 10081 8374 10133
rect 8446 10081 8498 10133
rect 8570 10081 8622 10133
rect 8694 10081 8746 10133
rect 8818 10081 8870 10133
rect 8942 10081 8994 10133
rect 9066 10081 9118 10133
rect 9190 10081 9242 10133
rect 9314 10081 9366 10133
rect 9438 10081 9490 10133
rect 7702 9957 7754 10009
rect 7826 9957 7878 10009
rect 7950 9957 8002 10009
rect 8074 9957 8126 10009
rect 8198 9957 8250 10009
rect 8322 9957 8374 10009
rect 8446 9957 8498 10009
rect 8570 9957 8622 10009
rect 8694 9957 8746 10009
rect 8818 9957 8870 10009
rect 8942 9957 8994 10009
rect 9066 9957 9118 10009
rect 9190 9957 9242 10009
rect 9314 9957 9366 10009
rect 9438 9957 9490 10009
rect 7702 9833 7754 9885
rect 7826 9833 7878 9885
rect 7950 9833 8002 9885
rect 8074 9833 8126 9885
rect 8198 9833 8250 9885
rect 8322 9833 8374 9885
rect 8446 9833 8498 9885
rect 8570 9833 8622 9885
rect 8694 9833 8746 9885
rect 8818 9833 8870 9885
rect 8942 9833 8994 9885
rect 9066 9833 9118 9885
rect 9190 9833 9242 9885
rect 9314 9833 9366 9885
rect 9438 9833 9490 9885
rect 7702 9709 7754 9761
rect 7826 9709 7878 9761
rect 7950 9709 8002 9761
rect 8074 9709 8126 9761
rect 8198 9709 8250 9761
rect 8322 9709 8374 9761
rect 8446 9709 8498 9761
rect 8570 9709 8622 9761
rect 8694 9709 8746 9761
rect 8818 9709 8870 9761
rect 8942 9709 8994 9761
rect 9066 9709 9118 9761
rect 9190 9709 9242 9761
rect 9314 9709 9366 9761
rect 9438 9709 9490 9761
rect 1462 3982 1514 4034
rect 1570 3982 1622 4034
rect 1678 3982 1730 4034
rect 1786 3982 1838 4034
rect 1894 3982 1946 4034
rect 2002 3982 2054 4034
rect 2110 3982 2162 4034
rect 2218 3982 2270 4034
rect 2326 3982 2378 4034
rect 2434 3982 2486 4034
rect 2542 3982 2594 4034
rect 2650 3982 2702 4034
rect 2758 3982 2810 4034
rect 2866 3982 2918 4034
rect 2974 3982 3026 4034
rect 3082 3982 3134 4034
rect 3190 3982 3242 4034
rect 1462 3874 1514 3926
rect 1570 3874 1622 3926
rect 1678 3874 1730 3926
rect 1786 3874 1838 3926
rect 1894 3874 1946 3926
rect 2002 3874 2054 3926
rect 2110 3874 2162 3926
rect 2218 3874 2270 3926
rect 2326 3874 2378 3926
rect 2434 3874 2486 3926
rect 2542 3874 2594 3926
rect 2650 3874 2702 3926
rect 2758 3874 2810 3926
rect 2866 3874 2918 3926
rect 2974 3874 3026 3926
rect 3082 3874 3134 3926
rect 3190 3874 3242 3926
rect 5329 3982 5381 4034
rect 5437 3982 5489 4034
rect 5545 3982 5597 4034
rect 5653 3982 5705 4034
rect 5761 3982 5813 4034
rect 5869 3982 5921 4034
rect 5977 3982 6029 4034
rect 6085 3982 6137 4034
rect 6193 3982 6245 4034
rect 6301 3982 6353 4034
rect 5329 3874 5381 3926
rect 5437 3874 5489 3926
rect 5545 3874 5597 3926
rect 5653 3874 5705 3926
rect 5761 3874 5813 3926
rect 5869 3874 5921 3926
rect 5977 3874 6029 3926
rect 6085 3874 6137 3926
rect 6193 3874 6245 3926
rect 6301 3874 6353 3926
rect 7706 3982 7758 4034
rect 7814 3982 7866 4034
rect 7922 3982 7974 4034
rect 8030 3982 8082 4034
rect 8138 3982 8190 4034
rect 8246 3982 8298 4034
rect 8354 3982 8406 4034
rect 8462 3982 8514 4034
rect 8570 3982 8622 4034
rect 8678 3982 8730 4034
rect 8786 3982 8838 4034
rect 8894 3982 8946 4034
rect 9002 3982 9054 4034
rect 9110 3982 9162 4034
rect 9218 3982 9270 4034
rect 9326 3982 9378 4034
rect 9434 3982 9486 4034
rect 7706 3874 7758 3926
rect 7814 3874 7866 3926
rect 7922 3874 7974 3926
rect 8030 3874 8082 3926
rect 8138 3874 8190 3926
rect 8246 3874 8298 3926
rect 8354 3874 8406 3926
rect 8462 3874 8514 3926
rect 8570 3874 8622 3926
rect 8678 3874 8730 3926
rect 8786 3874 8838 3926
rect 8894 3874 8946 3926
rect 9002 3874 9054 3926
rect 9110 3874 9162 3926
rect 9218 3874 9270 3926
rect 9326 3874 9378 3926
rect 9434 3874 9486 3926
rect 150 3514 202 3566
rect 258 3514 310 3566
rect 366 3514 418 3566
rect 474 3514 526 3566
rect 582 3514 634 3566
rect 690 3514 742 3566
rect 798 3514 850 3566
rect 906 3514 958 3566
rect 1014 3514 1066 3566
rect 3390 3514 3442 3566
rect 3498 3514 3550 3566
rect 3606 3514 3658 3566
rect 3714 3514 3766 3566
rect 3822 3514 3874 3566
rect 3930 3514 3982 3566
rect 4038 3514 4090 3566
rect 4146 3514 4198 3566
rect 4254 3514 4306 3566
rect 4362 3514 4414 3566
rect 4470 3514 4522 3566
rect 4578 3514 4630 3566
rect 4686 3514 4738 3566
rect 4794 3514 4846 3566
rect 4902 3514 4954 3566
rect 5010 3514 5062 3566
rect 5118 3514 5170 3566
rect 6523 3514 6575 3566
rect 6631 3514 6683 3566
rect 6739 3514 6791 3566
rect 6847 3514 6899 3566
rect 6955 3514 7007 3566
rect 7063 3514 7115 3566
rect 7171 3514 7223 3566
rect 7279 3514 7331 3566
rect 7387 3514 7439 3566
rect 7495 3514 7547 3566
rect 9634 3514 9686 3566
rect 9742 3514 9794 3566
rect 9850 3514 9902 3566
rect 9958 3514 10010 3566
rect 10066 3514 10118 3566
rect 10174 3514 10226 3566
rect 10282 3514 10334 3566
rect 10390 3514 10442 3566
rect 10498 3514 10550 3566
rect 10606 3514 10658 3566
rect 10714 3514 10766 3566
rect 10822 3514 10874 3566
rect 10930 3514 10982 3566
rect 11038 3514 11090 3566
rect 11146 3514 11198 3566
rect 11254 3514 11306 3566
rect 11362 3514 11414 3566
rect 150 3406 202 3458
rect 258 3406 310 3458
rect 366 3406 418 3458
rect 474 3406 526 3458
rect 582 3406 634 3458
rect 690 3406 742 3458
rect 798 3406 850 3458
rect 906 3406 958 3458
rect 1014 3406 1066 3458
rect 3390 3406 3442 3458
rect 3498 3406 3550 3458
rect 3606 3406 3658 3458
rect 3714 3406 3766 3458
rect 3822 3406 3874 3458
rect 3930 3406 3982 3458
rect 4038 3406 4090 3458
rect 4146 3406 4198 3458
rect 4254 3406 4306 3458
rect 4362 3406 4414 3458
rect 4470 3406 4522 3458
rect 4578 3406 4630 3458
rect 4686 3406 4738 3458
rect 4794 3406 4846 3458
rect 4902 3406 4954 3458
rect 5010 3406 5062 3458
rect 5118 3406 5170 3458
rect 6523 3406 6575 3458
rect 6631 3406 6683 3458
rect 6739 3406 6791 3458
rect 6847 3406 6899 3458
rect 6955 3406 7007 3458
rect 7063 3406 7115 3458
rect 7171 3406 7223 3458
rect 7279 3406 7331 3458
rect 7387 3406 7439 3458
rect 7495 3406 7547 3458
rect 9634 3406 9686 3458
rect 9742 3406 9794 3458
rect 9850 3406 9902 3458
rect 9958 3406 10010 3458
rect 10066 3406 10118 3458
rect 10174 3406 10226 3458
rect 10282 3406 10334 3458
rect 10390 3406 10442 3458
rect 10498 3406 10550 3458
rect 10606 3406 10658 3458
rect 10714 3406 10766 3458
rect 10822 3406 10874 3458
rect 10930 3406 10982 3458
rect 11038 3406 11090 3458
rect 11146 3406 11198 3458
rect 11254 3406 11306 3458
rect 11362 3406 11414 3458
rect 1462 234 1514 286
rect 1570 234 1622 286
rect 1678 234 1730 286
rect 1786 234 1838 286
rect 1894 234 1946 286
rect 2002 234 2054 286
rect 2110 234 2162 286
rect 2218 234 2270 286
rect 2326 234 2378 286
rect 2434 234 2486 286
rect 2542 234 2594 286
rect 2650 234 2702 286
rect 2758 234 2810 286
rect 2866 234 2918 286
rect 2974 234 3026 286
rect 3082 234 3134 286
rect 3190 234 3242 286
rect 5329 234 5381 286
rect 5437 234 5489 286
rect 5545 234 5597 286
rect 5653 234 5705 286
rect 5761 234 5813 286
rect 5869 234 5921 286
rect 5977 234 6029 286
rect 6085 234 6137 286
rect 6193 234 6245 286
rect 6301 234 6353 286
rect 1462 126 1514 178
rect 1570 126 1622 178
rect 1678 126 1730 178
rect 1786 126 1838 178
rect 1894 126 1946 178
rect 2002 126 2054 178
rect 2110 126 2162 178
rect 2218 126 2270 178
rect 2326 126 2378 178
rect 2434 126 2486 178
rect 2542 126 2594 178
rect 2650 126 2702 178
rect 2758 126 2810 178
rect 2866 126 2918 178
rect 2974 126 3026 178
rect 3082 126 3134 178
rect 3190 126 3242 178
rect 5329 126 5381 178
rect 5437 126 5489 178
rect 5545 126 5597 178
rect 5653 126 5705 178
rect 5761 126 5813 178
rect 5869 126 5921 178
rect 5977 126 6029 178
rect 6085 126 6137 178
rect 6193 126 6245 178
rect 6301 126 6353 178
rect 7904 234 7956 286
rect 8012 234 8064 286
rect 8120 234 8172 286
rect 8228 234 8280 286
rect 8336 234 8388 286
rect 8444 234 8496 286
rect 8552 234 8604 286
rect 8660 234 8712 286
rect 8768 234 8820 286
rect 8876 234 8928 286
rect 8984 234 9036 286
rect 9092 234 9144 286
rect 9200 234 9252 286
rect 9308 234 9360 286
rect 9416 234 9468 286
rect 11813 234 11865 286
rect 11921 234 11973 286
rect 12029 234 12081 286
rect 12137 234 12189 286
rect 12245 234 12297 286
rect 12353 234 12405 286
rect 12461 234 12513 286
rect 12569 234 12621 286
rect 12677 234 12729 286
rect 12785 234 12837 286
rect 7904 126 7956 178
rect 8012 126 8064 178
rect 8120 126 8172 178
rect 8228 126 8280 178
rect 8336 126 8388 178
rect 8444 126 8496 178
rect 8552 126 8604 178
rect 8660 126 8712 178
rect 8768 126 8820 178
rect 8876 126 8928 178
rect 8984 126 9036 178
rect 9092 126 9144 178
rect 9200 126 9252 178
rect 9308 126 9360 178
rect 9416 126 9468 178
rect 11813 126 11865 178
rect 11921 126 11973 178
rect 12029 126 12081 178
rect 12137 126 12189 178
rect 12245 126 12297 178
rect 12353 126 12405 178
rect 12461 126 12513 178
rect 12569 126 12621 178
rect 12677 126 12729 178
rect 12785 126 12837 178
<< metal2 >>
rect 4891 29422 6125 31350
rect 3963 28014 6125 29422
rect 3963 22978 5194 28014
rect 6307 27877 7506 31333
rect 0 16828 1102 17740
rect 0 16776 39 16828
rect 91 16776 147 16828
rect 199 16776 255 16828
rect 307 16776 363 16828
rect 415 16776 471 16828
rect 523 16776 579 16828
rect 631 16776 687 16828
rect 739 16776 795 16828
rect 847 16776 903 16828
rect 955 16776 1011 16828
rect 1063 16776 1102 16828
rect 0 16720 1102 16776
rect 0 16668 39 16720
rect 91 16668 147 16720
rect 199 16668 255 16720
rect 307 16668 363 16720
rect 415 16668 471 16720
rect 523 16668 579 16720
rect 631 16668 687 16720
rect 739 16668 795 16720
rect 847 16668 903 16720
rect 955 16668 1011 16720
rect 1063 16668 1102 16720
rect 0 3566 1102 16668
rect 0 3514 150 3566
rect 202 3514 258 3566
rect 310 3514 366 3566
rect 418 3514 474 3566
rect 526 3514 582 3566
rect 634 3514 690 3566
rect 742 3514 798 3566
rect 850 3514 906 3566
rect 958 3514 1014 3566
rect 1066 3514 1102 3566
rect 0 3458 1102 3514
rect 0 3406 150 3458
rect 202 3406 258 3458
rect 310 3406 366 3458
rect 418 3406 474 3458
rect 526 3406 582 3458
rect 634 3406 690 3458
rect 742 3406 798 3458
rect 850 3406 906 3458
rect 958 3406 1014 3458
rect 1066 3406 1102 3458
rect 0 0 1102 3406
rect 1438 16118 3266 16554
rect 1438 16066 1462 16118
rect 1514 16066 1570 16118
rect 1622 16066 1678 16118
rect 1730 16066 1786 16118
rect 1838 16066 1894 16118
rect 1946 16066 2002 16118
rect 2054 16066 2110 16118
rect 2162 16066 2218 16118
rect 2270 16066 2326 16118
rect 2378 16066 2434 16118
rect 2486 16066 2542 16118
rect 2594 16066 2650 16118
rect 2702 16066 2758 16118
rect 2810 16066 2866 16118
rect 2918 16066 2974 16118
rect 3026 16066 3082 16118
rect 3134 16066 3190 16118
rect 3242 16066 3266 16118
rect 1438 16010 3266 16066
rect 1438 15958 1462 16010
rect 1514 15958 1570 16010
rect 1622 15958 1678 16010
rect 1730 15958 1786 16010
rect 1838 15958 1894 16010
rect 1946 15958 2002 16010
rect 2054 15958 2110 16010
rect 2162 15958 2218 16010
rect 2270 15958 2326 16010
rect 2378 15958 2434 16010
rect 2486 15958 2542 16010
rect 2594 15958 2650 16010
rect 2702 15958 2758 16010
rect 2810 15958 2866 16010
rect 2918 15958 2974 16010
rect 3026 15958 3082 16010
rect 3134 15958 3190 16010
rect 3242 15958 3266 16010
rect 1438 10381 3266 15958
rect 1438 10329 1458 10381
rect 1510 10329 1582 10381
rect 1634 10329 1706 10381
rect 1758 10329 1830 10381
rect 1882 10329 1954 10381
rect 2006 10329 2078 10381
rect 2130 10329 2202 10381
rect 2254 10329 2326 10381
rect 2378 10329 2450 10381
rect 2502 10329 2574 10381
rect 2626 10329 2698 10381
rect 2750 10329 2822 10381
rect 2874 10329 2946 10381
rect 2998 10329 3070 10381
rect 3122 10329 3194 10381
rect 3246 10329 3266 10381
rect 1438 10257 3266 10329
rect 1438 10205 1458 10257
rect 1510 10205 1582 10257
rect 1634 10205 1706 10257
rect 1758 10205 1830 10257
rect 1882 10205 1954 10257
rect 2006 10205 2078 10257
rect 2130 10205 2202 10257
rect 2254 10205 2326 10257
rect 2378 10205 2450 10257
rect 2502 10205 2574 10257
rect 2626 10205 2698 10257
rect 2750 10205 2822 10257
rect 2874 10205 2946 10257
rect 2998 10205 3070 10257
rect 3122 10205 3194 10257
rect 3246 10205 3266 10257
rect 1438 10133 3266 10205
rect 1438 10081 1458 10133
rect 1510 10081 1582 10133
rect 1634 10081 1706 10133
rect 1758 10081 1830 10133
rect 1882 10081 1954 10133
rect 2006 10081 2078 10133
rect 2130 10081 2202 10133
rect 2254 10081 2326 10133
rect 2378 10081 2450 10133
rect 2502 10081 2574 10133
rect 2626 10081 2698 10133
rect 2750 10081 2822 10133
rect 2874 10081 2946 10133
rect 2998 10081 3070 10133
rect 3122 10081 3194 10133
rect 3246 10081 3266 10133
rect 1438 10009 3266 10081
rect 1438 9957 1458 10009
rect 1510 9957 1582 10009
rect 1634 9957 1706 10009
rect 1758 9957 1830 10009
rect 1882 9957 1954 10009
rect 2006 9957 2078 10009
rect 2130 9957 2202 10009
rect 2254 9957 2326 10009
rect 2378 9957 2450 10009
rect 2502 9957 2574 10009
rect 2626 9957 2698 10009
rect 2750 9957 2822 10009
rect 2874 9957 2946 10009
rect 2998 9957 3070 10009
rect 3122 9957 3194 10009
rect 3246 9957 3266 10009
rect 1438 9885 3266 9957
rect 1438 9833 1458 9885
rect 1510 9833 1582 9885
rect 1634 9833 1706 9885
rect 1758 9833 1830 9885
rect 1882 9833 1954 9885
rect 2006 9833 2078 9885
rect 2130 9833 2202 9885
rect 2254 9833 2326 9885
rect 2378 9833 2450 9885
rect 2502 9833 2574 9885
rect 2626 9833 2698 9885
rect 2750 9833 2822 9885
rect 2874 9833 2946 9885
rect 2998 9833 3070 9885
rect 3122 9833 3194 9885
rect 3246 9833 3266 9885
rect 1438 9761 3266 9833
rect 1438 9709 1458 9761
rect 1510 9709 1582 9761
rect 1634 9709 1706 9761
rect 1758 9709 1830 9761
rect 1882 9709 1954 9761
rect 2006 9709 2078 9761
rect 2130 9709 2202 9761
rect 2254 9709 2326 9761
rect 2378 9709 2450 9761
rect 2502 9709 2574 9761
rect 2626 9709 2698 9761
rect 2750 9709 2822 9761
rect 2874 9709 2946 9761
rect 2998 9709 3070 9761
rect 3122 9709 3194 9761
rect 3246 9709 3266 9761
rect 1438 4034 3266 9709
rect 1438 3982 1462 4034
rect 1514 3982 1570 4034
rect 1622 3982 1678 4034
rect 1730 3982 1786 4034
rect 1838 3982 1894 4034
rect 1946 3982 2002 4034
rect 2054 3982 2110 4034
rect 2162 3982 2218 4034
rect 2270 3982 2326 4034
rect 2378 3982 2434 4034
rect 2486 3982 2542 4034
rect 2594 3982 2650 4034
rect 2702 3982 2758 4034
rect 2810 3982 2866 4034
rect 2918 3982 2974 4034
rect 3026 3982 3082 4034
rect 3134 3982 3190 4034
rect 3242 3982 3266 4034
rect 1438 3926 3266 3982
rect 1438 3874 1462 3926
rect 1514 3874 1570 3926
rect 1622 3874 1678 3926
rect 1730 3874 1786 3926
rect 1838 3874 1894 3926
rect 1946 3874 2002 3926
rect 2054 3874 2110 3926
rect 2162 3874 2218 3926
rect 2270 3874 2326 3926
rect 2378 3874 2434 3926
rect 2486 3874 2542 3926
rect 2594 3874 2650 3926
rect 2702 3874 2758 3926
rect 2810 3874 2866 3926
rect 2918 3874 2974 3926
rect 3026 3874 3082 3926
rect 3134 3874 3190 3926
rect 3242 3874 3266 3926
rect 1438 286 3266 3874
rect 1438 234 1462 286
rect 1514 234 1570 286
rect 1622 234 1678 286
rect 1730 234 1786 286
rect 1838 234 1894 286
rect 1946 234 2002 286
rect 2054 234 2110 286
rect 2162 234 2218 286
rect 2270 234 2326 286
rect 2378 234 2434 286
rect 2486 234 2542 286
rect 2594 234 2650 286
rect 2702 234 2758 286
rect 2810 234 2866 286
rect 2918 234 2974 286
rect 3026 234 3082 286
rect 3134 234 3190 286
rect 3242 234 3266 286
rect 1438 178 3266 234
rect 1438 126 1462 178
rect 1514 126 1570 178
rect 1622 126 1678 178
rect 1730 126 1786 178
rect 1838 126 1894 178
rect 1946 126 2002 178
rect 2054 126 2110 178
rect 2162 126 2218 178
rect 2270 126 2326 178
rect 2378 126 2434 178
rect 2486 126 2542 178
rect 2594 126 2650 178
rect 2702 126 2758 178
rect 2810 126 2866 178
rect 2918 126 2974 178
rect 3026 126 3082 178
rect 3134 126 3190 178
rect 3242 126 3266 178
rect 1438 0 3266 126
rect 3366 3566 5194 22978
rect 3366 3514 3390 3566
rect 3442 3514 3498 3566
rect 3550 3514 3606 3566
rect 3658 3514 3714 3566
rect 3766 3514 3822 3566
rect 3874 3514 3930 3566
rect 3982 3514 4038 3566
rect 4090 3514 4146 3566
rect 4198 3514 4254 3566
rect 4306 3514 4362 3566
rect 4414 3514 4470 3566
rect 4522 3514 4578 3566
rect 4630 3514 4686 3566
rect 4738 3514 4794 3566
rect 4846 3514 4902 3566
rect 4954 3514 5010 3566
rect 5062 3514 5118 3566
rect 5170 3514 5194 3566
rect 3366 3458 5194 3514
rect 3366 3406 3390 3458
rect 3442 3406 3498 3458
rect 3550 3406 3606 3458
rect 3658 3406 3714 3458
rect 3766 3406 3822 3458
rect 3874 3406 3930 3458
rect 3982 3406 4038 3458
rect 4090 3406 4146 3458
rect 4198 3406 4254 3458
rect 4306 3406 4362 3458
rect 4414 3406 4470 3458
rect 4522 3406 4578 3458
rect 4630 3406 4686 3458
rect 4738 3406 4794 3458
rect 4846 3406 4902 3458
rect 4954 3406 5010 3458
rect 5062 3406 5118 3458
rect 5170 3406 5194 3458
rect 3366 0 5194 3406
rect 5294 26749 7506 27877
rect 5294 16118 6388 26749
rect 5294 16066 5329 16118
rect 5381 16066 5437 16118
rect 5489 16066 5545 16118
rect 5597 16066 5653 16118
rect 5705 16066 5761 16118
rect 5813 16066 5869 16118
rect 5921 16066 5977 16118
rect 6029 16066 6085 16118
rect 6137 16066 6193 16118
rect 6245 16066 6301 16118
rect 6353 16066 6388 16118
rect 5294 16010 6388 16066
rect 5294 15958 5329 16010
rect 5381 15958 5437 16010
rect 5489 15958 5545 16010
rect 5597 15958 5653 16010
rect 5705 15958 5761 16010
rect 5813 15958 5869 16010
rect 5921 15958 5977 16010
rect 6029 15958 6085 16010
rect 6137 15958 6193 16010
rect 6245 15958 6301 16010
rect 6353 15958 6388 16010
rect 5294 10381 6388 15958
rect 5294 10329 5319 10381
rect 5371 10329 5443 10381
rect 5495 10329 5567 10381
rect 5619 10329 5691 10381
rect 5743 10329 5815 10381
rect 5867 10329 5939 10381
rect 5991 10329 6063 10381
rect 6115 10329 6187 10381
rect 6239 10329 6311 10381
rect 6363 10329 6388 10381
rect 5294 10257 6388 10329
rect 5294 10205 5319 10257
rect 5371 10205 5443 10257
rect 5495 10205 5567 10257
rect 5619 10205 5691 10257
rect 5743 10205 5815 10257
rect 5867 10205 5939 10257
rect 5991 10205 6063 10257
rect 6115 10205 6187 10257
rect 6239 10205 6311 10257
rect 6363 10205 6388 10257
rect 5294 10133 6388 10205
rect 5294 10081 5319 10133
rect 5371 10081 5443 10133
rect 5495 10081 5567 10133
rect 5619 10081 5691 10133
rect 5743 10081 5815 10133
rect 5867 10081 5939 10133
rect 5991 10081 6063 10133
rect 6115 10081 6187 10133
rect 6239 10081 6311 10133
rect 6363 10081 6388 10133
rect 5294 10009 6388 10081
rect 5294 9957 5319 10009
rect 5371 9957 5443 10009
rect 5495 9957 5567 10009
rect 5619 9957 5691 10009
rect 5743 9957 5815 10009
rect 5867 9957 5939 10009
rect 5991 9957 6063 10009
rect 6115 9957 6187 10009
rect 6239 9957 6311 10009
rect 6363 9957 6388 10009
rect 5294 9885 6388 9957
rect 5294 9833 5319 9885
rect 5371 9833 5443 9885
rect 5495 9833 5567 9885
rect 5619 9833 5691 9885
rect 5743 9833 5815 9885
rect 5867 9833 5939 9885
rect 5991 9833 6063 9885
rect 6115 9833 6187 9885
rect 6239 9833 6311 9885
rect 6363 9833 6388 9885
rect 5294 9761 6388 9833
rect 5294 9709 5319 9761
rect 5371 9709 5443 9761
rect 5495 9709 5567 9761
rect 5619 9709 5691 9761
rect 5743 9709 5815 9761
rect 5867 9709 5939 9761
rect 5991 9709 6063 9761
rect 6115 9709 6187 9761
rect 6239 9709 6311 9761
rect 6363 9709 6388 9761
rect 5294 4034 6388 9709
rect 5294 3982 5329 4034
rect 5381 3982 5437 4034
rect 5489 3982 5545 4034
rect 5597 3982 5653 4034
rect 5705 3982 5761 4034
rect 5813 3982 5869 4034
rect 5921 3982 5977 4034
rect 6029 3982 6085 4034
rect 6137 3982 6193 4034
rect 6245 3982 6301 4034
rect 6353 3982 6388 4034
rect 5294 3926 6388 3982
rect 5294 3874 5329 3926
rect 5381 3874 5437 3926
rect 5489 3874 5545 3926
rect 5597 3874 5653 3926
rect 5705 3874 5761 3926
rect 5813 3874 5869 3926
rect 5921 3874 5977 3926
rect 6029 3874 6085 3926
rect 6137 3874 6193 3926
rect 6245 3874 6301 3926
rect 6353 3874 6388 3926
rect 5294 286 6388 3874
rect 5294 234 5329 286
rect 5381 234 5437 286
rect 5489 234 5545 286
rect 5597 234 5653 286
rect 5705 234 5761 286
rect 5813 234 5869 286
rect 5921 234 5977 286
rect 6029 234 6085 286
rect 6137 234 6193 286
rect 6245 234 6301 286
rect 6353 234 6388 286
rect 5294 178 6388 234
rect 5294 126 5329 178
rect 5381 126 5437 178
rect 5489 126 5545 178
rect 5597 126 5653 178
rect 5705 126 5761 178
rect 5813 126 5869 178
rect 5921 126 5977 178
rect 6029 126 6085 178
rect 6137 126 6193 178
rect 6245 126 6301 178
rect 6353 126 6388 178
rect 5294 0 6388 126
rect 6488 3566 7582 26448
rect 9945 16554 11438 24232
rect 6488 3514 6523 3566
rect 6575 3514 6631 3566
rect 6683 3514 6739 3566
rect 6791 3514 6847 3566
rect 6899 3514 6955 3566
rect 7007 3514 7063 3566
rect 7115 3514 7171 3566
rect 7223 3514 7279 3566
rect 7331 3514 7387 3566
rect 7439 3514 7495 3566
rect 7547 3514 7582 3566
rect 6488 3458 7582 3514
rect 6488 3406 6523 3458
rect 6575 3406 6631 3458
rect 6683 3406 6739 3458
rect 6791 3406 6847 3458
rect 6899 3406 6955 3458
rect 7007 3406 7063 3458
rect 7115 3406 7171 3458
rect 7223 3406 7279 3458
rect 7331 3406 7387 3458
rect 7439 3406 7495 3458
rect 7547 3406 7582 3458
rect 6488 0 7582 3406
rect 7682 16118 9510 16554
rect 7682 16066 7706 16118
rect 7758 16066 7814 16118
rect 7866 16066 7922 16118
rect 7974 16066 8030 16118
rect 8082 16066 8138 16118
rect 8190 16066 8246 16118
rect 8298 16066 8354 16118
rect 8406 16066 8462 16118
rect 8514 16066 8570 16118
rect 8622 16066 8678 16118
rect 8730 16066 8786 16118
rect 8838 16066 8894 16118
rect 8946 16066 9002 16118
rect 9054 16066 9110 16118
rect 9162 16066 9218 16118
rect 9270 16066 9326 16118
rect 9378 16066 9434 16118
rect 9486 16066 9510 16118
rect 7682 16010 9510 16066
rect 7682 15958 7706 16010
rect 7758 15958 7814 16010
rect 7866 15958 7922 16010
rect 7974 15958 8030 16010
rect 8082 15958 8138 16010
rect 8190 15958 8246 16010
rect 8298 15958 8354 16010
rect 8406 15958 8462 16010
rect 8514 15958 8570 16010
rect 8622 15958 8678 16010
rect 8730 15958 8786 16010
rect 8838 15958 8894 16010
rect 8946 15958 9002 16010
rect 9054 15958 9110 16010
rect 9162 15958 9218 16010
rect 9270 15958 9326 16010
rect 9378 15958 9434 16010
rect 9486 15958 9510 16010
rect 7682 10381 9510 15958
rect 7682 10329 7702 10381
rect 7754 10329 7826 10381
rect 7878 10329 7950 10381
rect 8002 10329 8074 10381
rect 8126 10329 8198 10381
rect 8250 10329 8322 10381
rect 8374 10329 8446 10381
rect 8498 10329 8570 10381
rect 8622 10329 8694 10381
rect 8746 10329 8818 10381
rect 8870 10329 8942 10381
rect 8994 10329 9066 10381
rect 9118 10329 9190 10381
rect 9242 10329 9314 10381
rect 9366 10329 9438 10381
rect 9490 10329 9510 10381
rect 7682 10257 9510 10329
rect 7682 10205 7702 10257
rect 7754 10205 7826 10257
rect 7878 10205 7950 10257
rect 8002 10205 8074 10257
rect 8126 10205 8198 10257
rect 8250 10205 8322 10257
rect 8374 10205 8446 10257
rect 8498 10205 8570 10257
rect 8622 10205 8694 10257
rect 8746 10205 8818 10257
rect 8870 10205 8942 10257
rect 8994 10205 9066 10257
rect 9118 10205 9190 10257
rect 9242 10205 9314 10257
rect 9366 10205 9438 10257
rect 9490 10205 9510 10257
rect 7682 10133 9510 10205
rect 7682 10081 7702 10133
rect 7754 10081 7826 10133
rect 7878 10081 7950 10133
rect 8002 10081 8074 10133
rect 8126 10081 8198 10133
rect 8250 10081 8322 10133
rect 8374 10081 8446 10133
rect 8498 10081 8570 10133
rect 8622 10081 8694 10133
rect 8746 10081 8818 10133
rect 8870 10081 8942 10133
rect 8994 10081 9066 10133
rect 9118 10081 9190 10133
rect 9242 10081 9314 10133
rect 9366 10081 9438 10133
rect 9490 10081 9510 10133
rect 7682 10009 9510 10081
rect 7682 9957 7702 10009
rect 7754 9957 7826 10009
rect 7878 9957 7950 10009
rect 8002 9957 8074 10009
rect 8126 9957 8198 10009
rect 8250 9957 8322 10009
rect 8374 9957 8446 10009
rect 8498 9957 8570 10009
rect 8622 9957 8694 10009
rect 8746 9957 8818 10009
rect 8870 9957 8942 10009
rect 8994 9957 9066 10009
rect 9118 9957 9190 10009
rect 9242 9957 9314 10009
rect 9366 9957 9438 10009
rect 9490 9957 9510 10009
rect 7682 9885 9510 9957
rect 7682 9833 7702 9885
rect 7754 9833 7826 9885
rect 7878 9833 7950 9885
rect 8002 9833 8074 9885
rect 8126 9833 8198 9885
rect 8250 9833 8322 9885
rect 8374 9833 8446 9885
rect 8498 9833 8570 9885
rect 8622 9833 8694 9885
rect 8746 9833 8818 9885
rect 8870 9833 8942 9885
rect 8994 9833 9066 9885
rect 9118 9833 9190 9885
rect 9242 9833 9314 9885
rect 9366 9833 9438 9885
rect 9490 9833 9510 9885
rect 7682 9761 9510 9833
rect 7682 9709 7702 9761
rect 7754 9709 7826 9761
rect 7878 9709 7950 9761
rect 8002 9709 8074 9761
rect 8126 9709 8198 9761
rect 8250 9709 8322 9761
rect 8374 9709 8446 9761
rect 8498 9709 8570 9761
rect 8622 9709 8694 9761
rect 8746 9709 8818 9761
rect 8870 9709 8942 9761
rect 8994 9709 9066 9761
rect 9118 9709 9190 9761
rect 9242 9709 9314 9761
rect 9366 9709 9438 9761
rect 9490 9709 9510 9761
rect 7682 4034 9510 9709
rect 7682 3982 7706 4034
rect 7758 3982 7814 4034
rect 7866 3982 7922 4034
rect 7974 3982 8030 4034
rect 8082 3982 8138 4034
rect 8190 3982 8246 4034
rect 8298 3982 8354 4034
rect 8406 3982 8462 4034
rect 8514 3982 8570 4034
rect 8622 3982 8678 4034
rect 8730 3982 8786 4034
rect 8838 3982 8894 4034
rect 8946 3982 9002 4034
rect 9054 3982 9110 4034
rect 9162 3982 9218 4034
rect 9270 3982 9326 4034
rect 9378 3982 9434 4034
rect 9486 3982 9510 4034
rect 7682 3926 9510 3982
rect 7682 3874 7706 3926
rect 7758 3874 7814 3926
rect 7866 3874 7922 3926
rect 7974 3874 8030 3926
rect 8082 3874 8138 3926
rect 8190 3874 8246 3926
rect 8298 3874 8354 3926
rect 8406 3874 8462 3926
rect 8514 3874 8570 3926
rect 8622 3874 8678 3926
rect 8730 3874 8786 3926
rect 8838 3874 8894 3926
rect 8946 3874 9002 3926
rect 9054 3874 9110 3926
rect 9162 3874 9218 3926
rect 9270 3874 9326 3926
rect 9378 3874 9434 3926
rect 9486 3874 9510 3926
rect 7682 286 9510 3874
rect 7682 234 7904 286
rect 7956 234 8012 286
rect 8064 234 8120 286
rect 8172 234 8228 286
rect 8280 234 8336 286
rect 8388 234 8444 286
rect 8496 234 8552 286
rect 8604 234 8660 286
rect 8712 234 8768 286
rect 8820 234 8876 286
rect 8928 234 8984 286
rect 9036 234 9092 286
rect 9144 234 9200 286
rect 9252 234 9308 286
rect 9360 234 9416 286
rect 9468 234 9510 286
rect 7682 178 9510 234
rect 7682 126 7904 178
rect 7956 126 8012 178
rect 8064 126 8120 178
rect 8172 126 8228 178
rect 8280 126 8336 178
rect 8388 126 8444 178
rect 8496 126 8552 178
rect 8604 126 8660 178
rect 8712 126 8768 178
rect 8820 126 8876 178
rect 8928 126 8984 178
rect 9036 126 9092 178
rect 9144 126 9200 178
rect 9252 126 9308 178
rect 9360 126 9416 178
rect 9468 126 9510 178
rect 7682 0 9510 126
rect 9610 3566 11438 16554
rect 9610 3514 9634 3566
rect 9686 3514 9742 3566
rect 9794 3514 9850 3566
rect 9902 3514 9958 3566
rect 10010 3514 10066 3566
rect 10118 3514 10174 3566
rect 10226 3514 10282 3566
rect 10334 3514 10390 3566
rect 10442 3514 10498 3566
rect 10550 3514 10606 3566
rect 10658 3514 10714 3566
rect 10766 3514 10822 3566
rect 10874 3514 10930 3566
rect 10982 3514 11038 3566
rect 11090 3514 11146 3566
rect 11198 3514 11254 3566
rect 11306 3514 11362 3566
rect 11414 3514 11438 3566
rect 9610 3458 11438 3514
rect 9610 3406 9634 3458
rect 9686 3406 9742 3458
rect 9794 3406 9850 3458
rect 9902 3406 9958 3458
rect 10010 3406 10066 3458
rect 10118 3406 10174 3458
rect 10226 3406 10282 3458
rect 10334 3406 10390 3458
rect 10442 3406 10498 3458
rect 10550 3406 10606 3458
rect 10658 3406 10714 3458
rect 10766 3406 10822 3458
rect 10874 3406 10930 3458
rect 10982 3406 11038 3458
rect 11090 3406 11146 3458
rect 11198 3406 11254 3458
rect 11306 3406 11362 3458
rect 11414 3406 11438 3458
rect 9610 0 11438 3406
rect 11774 16554 12656 25832
rect 11774 286 12876 16554
rect 11774 234 11813 286
rect 11865 234 11921 286
rect 11973 234 12029 286
rect 12081 234 12137 286
rect 12189 234 12245 286
rect 12297 234 12353 286
rect 12405 234 12461 286
rect 12513 234 12569 286
rect 12621 234 12677 286
rect 12729 234 12785 286
rect 12837 234 12876 286
rect 11774 178 12876 234
rect 11774 126 11813 178
rect 11865 126 11921 178
rect 11973 126 12029 178
rect 12081 126 12137 178
rect 12189 126 12245 178
rect 12297 126 12353 178
rect 12405 126 12461 178
rect 12513 126 12569 178
rect 12621 126 12677 178
rect 12729 126 12785 178
rect 12837 126 12876 178
rect 11774 0 12876 126
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_0
timestamp 1669390400
transform 1 0 10524 0 1 3486
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_1
timestamp 1669390400
transform 1 0 8596 0 1 16038
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_2
timestamp 1669390400
transform 1 0 8596 0 1 3954
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_3
timestamp 1669390400
transform 1 0 4280 0 1 3486
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_4
timestamp 1669390400
transform 1 0 2352 0 1 16038
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_5
timestamp 1669390400
transform 1 0 2352 0 1 3954
box 0 0 1 1
use M2_M1_CDNS_40661956134143  M2_M1_CDNS_40661956134143_6
timestamp 1669390400
transform 1 0 2352 0 1 206
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_0
timestamp 1669390400
transform 1 0 551 0 1 16748
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_1
timestamp 1669390400
transform 1 0 5841 0 1 206
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_2
timestamp 1669390400
transform 1 0 5841 0 1 3954
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_3
timestamp 1669390400
transform 1 0 5841 0 1 16038
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_4
timestamp 1669390400
transform 1 0 12325 0 1 206
box 0 0 1 1
use M2_M1_CDNS_40661956134147  M2_M1_CDNS_40661956134147_5
timestamp 1669390400
transform 1 0 7035 0 1 3486
box 0 0 1 1
use M2_M1_CDNS_40661956134149  M2_M1_CDNS_40661956134149_0
timestamp 1669390400
transform 1 0 608 0 1 3486
box 0 0 1 1
use M2_M1_CDNS_40661956134150  M2_M1_CDNS_40661956134150_0
timestamp 1669390400
transform 1 0 8596 0 1 10045
box 0 0 1 1
use M2_M1_CDNS_40661956134150  M2_M1_CDNS_40661956134150_1
timestamp 1669390400
transform 1 0 2352 0 1 10045
box 0 0 1 1
use M2_M1_CDNS_40661956134151  M2_M1_CDNS_40661956134151_0
timestamp 1669390400
transform 1 0 5841 0 1 10045
box 0 0 1 1
use M2_M1_CDNS_40661956134152  M2_M1_CDNS_40661956134152_0
timestamp 1669390400
transform 1 0 8686 0 1 206
box 0 0 1 1
<< properties >>
string GDS_END 4724986
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4722588
string path 308.125 0.000 308.125 413.850 
<< end >>
