magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 960 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 860 360
rect 760 252 792 298
rect 838 252 860 298
rect 760 190 860 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 860 1430
rect 760 1143 792 1377
rect 838 1143 860 1377
rect 760 1090 860 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 190 990 760 1040
rect 190 800 250 990
rect 160 780 250 800
rect 90 758 250 780
rect 90 712 112 758
rect 158 712 250 758
rect 90 690 250 712
rect 160 680 250 690
rect 190 450 250 680
rect 190 400 760 450
rect 190 360 250 400
rect 360 360 420 400
rect 530 360 590 400
rect 700 360 760 400
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
<< polycontact >>
rect 112 712 158 758
<< metal1 >>
rect 0 1568 960 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 960 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 960 1566
rect 0 1470 960 1514
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1060 160 1143
rect 280 1377 330 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 940 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1060 500 1143
rect 620 1377 670 1430
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 940 670 1143
rect 790 1377 840 1470
rect 790 1143 792 1377
rect 838 1143 840 1377
rect 790 1060 840 1143
rect 280 936 670 940
rect 280 884 614 936
rect 666 884 670 936
rect 280 860 670 884
rect 80 758 180 760
rect 80 756 112 758
rect 80 704 104 756
rect 158 712 180 758
rect 156 704 180 712
rect 80 670 180 704
rect 280 460 330 860
rect 590 840 670 860
rect 620 460 670 840
rect 280 380 670 460
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 380
rect 280 252 282 298
rect 328 252 330 298
rect 280 160 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 380
rect 620 252 622 298
rect 668 252 670 298
rect 620 160 670 252
rect 790 298 840 360
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 0 106 960 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 960 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 960 54
rect 0 -30 960 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 614 884 666 936
rect 104 712 112 756
rect 112 712 156 756
rect 104 704 156 712
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1480 670 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 580 1470 660 1480
rect 590 936 690 950
rect 590 884 614 936
rect 666 884 690 936
rect 590 840 690 884
rect 80 756 180 770
rect 80 704 104 756
rect 156 704 180 756
rect 80 660 180 704
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 20 670 54
rect 100 10 180 20
rect 340 10 420 20
rect 580 10 660 20
<< labels >>
rlabel metal2 s 100 1470 180 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 100 10 180 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 80 660 180 740 4 A
port 1 nsew signal input
rlabel metal2 s 590 840 690 920 4 Y
port 2 nsew signal output
rlabel metal1 s 80 670 180 730 1 A
port 1 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 580 1470 660 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 570 1480 670 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 1060 840 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1470 960 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 580 10 660 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 570 20 670 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 -30 840 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 -30 960 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 380 670 430 1 Y
port 2 nsew signal output
rlabel metal1 s 590 840 670 910 1 Y
port 2 nsew signal output
rlabel metal1 s 280 860 670 910 1 Y
port 2 nsew signal output
rlabel metal1 s 620 160 670 1400 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 960 1590
string GDS_END 357800
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 350472
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
