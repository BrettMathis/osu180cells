magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -64 1007 64 1045
rect -64 951 -28 1007
rect 28 951 64 1007
rect -64 790 64 951
rect -64 734 -28 790
rect 28 734 64 790
rect -64 572 64 734
rect -64 516 -28 572
rect 28 516 64 572
rect -64 355 64 516
rect -64 299 -28 355
rect 28 299 64 355
rect -64 137 64 299
rect -64 81 -28 137
rect 28 81 64 137
rect -64 -81 64 81
rect -64 -137 -28 -81
rect 28 -137 64 -81
rect -64 -299 64 -137
rect -64 -355 -28 -299
rect 28 -355 64 -299
rect -64 -516 64 -355
rect -64 -572 -28 -516
rect 28 -572 64 -516
rect -64 -734 64 -572
rect -64 -790 -28 -734
rect 28 -790 64 -734
rect -64 -951 64 -790
rect -64 -1007 -28 -951
rect 28 -1007 64 -951
rect -64 -1046 64 -1007
<< via2 >>
rect -28 951 28 1007
rect -28 734 28 790
rect -28 516 28 572
rect -28 299 28 355
rect -28 81 28 137
rect -28 -137 28 -81
rect -28 -355 28 -299
rect -28 -572 28 -516
rect -28 -790 28 -734
rect -28 -1007 28 -951
<< metal3 >>
rect -65 1007 65 1046
rect -65 951 -28 1007
rect 28 951 65 1007
rect -65 790 65 951
rect -65 734 -28 790
rect 28 734 65 790
rect -65 572 65 734
rect -65 516 -28 572
rect 28 516 65 572
rect -65 355 65 516
rect -65 299 -28 355
rect 28 299 65 355
rect -65 137 65 299
rect -65 81 -28 137
rect 28 81 65 137
rect -65 -81 65 81
rect -65 -137 -28 -81
rect 28 -137 65 -81
rect -65 -299 65 -137
rect -65 -355 -28 -299
rect 28 -355 65 -299
rect -65 -516 65 -355
rect -65 -572 -28 -516
rect 28 -572 65 -516
rect -65 -734 65 -572
rect -65 -790 -28 -734
rect 28 -790 65 -734
rect -65 -951 65 -790
rect -65 -1007 -28 -951
rect 28 -1007 65 -951
rect -65 -1046 65 -1007
<< properties >>
string GDS_END 253596
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 252824
<< end >>
