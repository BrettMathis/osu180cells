magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect -17 147 299 159
rect 11 106 16 147
rect 28 100 33 140
rect 45 106 50 147
rect 62 100 67 140
rect 79 106 84 147
rect 96 100 101 140
rect 113 106 118 147
rect 130 100 135 140
rect 147 106 152 147
rect 164 100 169 140
rect 181 106 186 147
rect 198 100 203 140
rect 215 106 220 147
rect 232 100 237 140
rect 249 106 254 147
rect 266 100 271 140
rect 283 106 288 147
rect 28 94 274 100
rect 4 80 14 86
rect 28 43 33 94
rect 62 43 67 94
rect 96 43 101 94
rect 130 43 135 94
rect 164 43 169 94
rect 198 43 203 94
rect 232 43 237 94
rect 266 43 271 94
rect 28 38 271 43
rect 11 9 16 33
rect 28 16 33 38
rect 45 9 50 33
rect 62 16 67 38
rect 79 9 84 33
rect 96 16 101 38
rect 113 9 118 33
rect 130 16 135 38
rect 147 9 152 33
rect 164 16 169 38
rect 181 9 186 33
rect 198 16 203 38
rect 215 9 220 33
rect 232 16 237 38
rect 249 9 254 33
rect 266 16 271 38
rect 283 9 288 33
rect -17 -3 299 9
<< obsm1 >>
rect -6 61 -1 140
rect -6 55 23 61
rect -6 16 -1 55
<< metal2 >>
rect -7 154 1 155
rect 17 154 25 155
rect 41 154 49 155
rect 65 154 73 155
rect 89 154 97 155
rect 113 154 121 155
rect 137 154 145 155
rect 161 154 169 155
rect 185 154 193 155
rect 209 154 217 155
rect 233 154 241 155
rect 257 154 265 155
rect -8 148 2 154
rect 16 148 26 154
rect 40 148 50 154
rect 64 148 74 154
rect 88 148 98 154
rect 112 148 122 154
rect 136 148 146 154
rect 160 148 170 154
rect 184 148 194 154
rect 208 148 218 154
rect 232 148 242 154
rect 256 148 266 154
rect -7 147 1 148
rect 17 147 25 148
rect 41 147 49 148
rect 65 147 73 148
rect 89 147 97 148
rect 113 147 121 148
rect 137 147 145 148
rect 161 147 169 148
rect 185 147 193 148
rect 209 147 217 148
rect 233 147 241 148
rect 257 147 265 148
rect 264 100 274 101
rect 263 94 274 100
rect 264 93 274 94
rect 5 86 13 87
rect 4 80 14 86
rect 5 79 13 80
rect -7 8 1 9
rect 17 8 25 9
rect 41 8 49 9
rect 65 8 73 9
rect 89 8 97 9
rect 113 8 121 9
rect 137 8 145 9
rect 161 8 169 9
rect 185 8 193 9
rect 209 8 217 9
rect 233 8 241 9
rect 257 8 265 9
rect -8 2 2 8
rect 16 2 26 8
rect 40 2 50 8
rect 64 2 74 8
rect 88 2 98 8
rect 112 2 122 8
rect 136 2 146 8
rect 160 2 170 8
rect 184 2 194 8
rect 208 2 218 8
rect 232 2 242 8
rect 256 2 266 8
rect -7 1 1 2
rect 17 1 25 2
rect 41 1 49 2
rect 65 1 73 2
rect 89 1 97 2
rect 113 1 121 2
rect 137 1 145 2
rect 161 1 169 2
rect 185 1 193 2
rect 209 1 217 2
rect 233 1 241 2
rect 257 1 265 2
<< labels >>
rlabel metal2 s 5 79 13 87 6 A
port 1 nsew signal input
rlabel metal2 s 4 80 14 86 6 A
port 1 nsew signal input
rlabel metal1 s 4 80 14 86 6 A
port 1 nsew signal input
rlabel metal2 s -7 147 1 155 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s -8 148 2 154 4 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 17 147 25 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 16 148 26 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 41 147 49 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 40 148 50 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 65 147 73 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 64 148 74 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 89 147 97 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 88 148 98 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 113 147 121 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 112 148 122 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 137 147 145 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 136 148 146 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 161 147 169 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 160 148 170 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 185 147 193 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 184 148 194 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 209 147 217 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 208 148 218 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 233 147 241 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 232 148 242 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 257 147 265 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 256 148 266 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 45 106 50 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 79 106 84 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 113 106 118 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 147 106 152 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 181 106 186 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 215 106 220 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 249 106 254 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 283 106 288 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s -17 147 299 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s -7 1 1 9 4 VSS
port 6 nsew ground bidirectional
rlabel metal2 s -8 2 2 8 4 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 17 1 25 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 16 2 26 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 41 1 49 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 40 2 50 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 65 1 73 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 64 2 74 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 89 1 97 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 88 2 98 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 113 1 121 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 112 2 122 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 137 1 145 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 136 2 146 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 161 1 169 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 160 2 170 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 185 1 193 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 184 2 194 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 209 1 217 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 208 2 218 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 233 1 241 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 232 2 242 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 257 1 265 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 256 2 266 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 45 -3 50 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 79 -3 84 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 113 -3 118 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 147 -3 152 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 181 -3 186 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 215 -3 220 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 249 -3 254 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 283 -3 288 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s -17 -3 299 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 263 94 274 100 6 Y
port 2 nsew signal output
rlabel metal2 s 264 93 274 101 6 Y
port 2 nsew signal output
rlabel metal1 s 28 16 33 140 6 Y
port 2 nsew signal output
rlabel metal1 s 62 16 67 140 6 Y
port 2 nsew signal output
rlabel metal1 s 96 16 101 140 6 Y
port 2 nsew signal output
rlabel metal1 s 130 16 135 140 6 Y
port 2 nsew signal output
rlabel metal1 s 164 16 169 140 6 Y
port 2 nsew signal output
rlabel metal1 s 198 16 203 140 6 Y
port 2 nsew signal output
rlabel metal1 s 232 16 237 140 6 Y
port 2 nsew signal output
rlabel metal1 s 28 38 271 43 6 Y
port 2 nsew signal output
rlabel metal1 s 266 16 271 140 6 Y
port 2 nsew signal output
rlabel metal1 s 28 94 274 100 6 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX -17 -3 299 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 166456
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 143448
<< end >>
