magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 322 23861 5755 29123
rect 1448 9376 1506 9429
rect 2252 9374 2303 9400
rect 3186 2694 3236 2701
<< mvpmos >>
rect 5069 27944 5189 28626
rect 5294 27944 5414 28626
rect 5069 27169 5189 27851
rect 5294 27169 5414 27851
<< mvpdiff >>
rect 4963 27944 5069 28626
rect 5189 27944 5294 28626
rect 5414 27944 5520 28626
rect 4963 27169 5069 27851
rect 5189 27169 5294 27851
rect 5414 27169 5520 27851
<< metal1 >>
rect 412 27097 540 27118
rect 412 27045 448 27097
rect 500 27045 540 27097
rect 412 27025 540 27045
rect 698 18380 826 18401
rect 698 18328 734 18380
rect 786 18328 826 18380
rect 698 18308 826 18328
rect 1717 18380 2025 18400
rect 1717 18328 1747 18380
rect 1799 18328 1933 18380
rect 1985 18328 2025 18380
rect 1717 18308 2025 18328
rect 2955 18380 3263 18400
rect 2955 18328 2985 18380
rect 3037 18328 3171 18380
rect 3223 18328 3263 18380
rect 2955 18308 3263 18328
rect 4194 18380 4502 18400
rect 4194 18328 4224 18380
rect 4276 18328 4410 18380
rect 4462 18328 4502 18380
rect 4194 18308 4502 18328
rect 5389 18380 5517 18401
rect 5389 18328 5429 18380
rect 5481 18328 5517 18380
rect 5389 18308 5517 18328
rect 4824 16408 5132 16428
rect 4824 16356 4854 16408
rect 4906 16356 5040 16408
rect 5092 16356 5132 16408
rect 4824 16336 5132 16356
rect 3720 16180 4482 16220
rect 3720 16128 3758 16180
rect 3810 16128 3969 16180
rect 4021 16128 4181 16180
rect 4233 16128 4392 16180
rect 4444 16128 4482 16180
rect 3720 16087 4482 16128
rect 500 15946 628 15967
rect 500 15894 536 15946
rect 588 15894 628 15946
rect 500 15874 628 15894
rect 2258 15929 2350 15970
rect 2258 15877 2278 15929
rect 2330 15877 2350 15929
rect 2258 15743 2350 15877
rect 2258 15691 2278 15743
rect 2330 15691 2350 15743
rect 2258 15651 2350 15691
rect 5344 10239 5438 11046
rect 5344 10187 5365 10239
rect 5417 10187 5438 10239
rect 5344 10069 5438 10187
rect 5345 10053 5437 10069
rect 5345 10001 5365 10053
rect 5417 10001 5437 10053
rect 5345 9960 5437 10001
rect 617 8863 925 8883
rect 617 8811 647 8863
rect 699 8811 833 8863
rect 885 8811 925 8863
rect 617 8791 925 8811
rect 2741 8732 2824 9040
rect 461 8523 553 8563
rect 461 8471 481 8523
rect 533 8471 553 8523
rect 461 8337 553 8471
rect 461 8285 481 8337
rect 533 8285 553 8337
rect 461 8244 553 8285
rect 3416 7513 3620 7821
rect 1485 6634 1577 6675
rect 1485 6582 1505 6634
rect 1557 6582 1577 6634
rect 1485 6448 1577 6582
rect 1485 6396 1505 6448
rect 1557 6396 1577 6448
rect 1485 6356 1577 6396
rect 4639 5591 4715 5603
rect 4639 5435 4651 5591
rect 4703 5435 4715 5591
rect 4639 5423 4715 5435
rect 5125 5591 5201 5603
rect 5125 5435 5137 5591
rect 5189 5435 5201 5591
rect 5125 5423 5201 5435
rect 2257 3604 2349 3644
rect 2257 3552 2277 3604
rect 2329 3552 2349 3604
rect 2257 3418 2349 3552
rect 2257 3366 2277 3418
rect 2329 3366 2349 3418
rect 2257 3325 2349 3366
rect 1813 1020 1929 1178
rect 2397 907 2480 1027
rect 2621 979 2677 1001
rect 2621 907 2698 979
rect 3346 907 3413 1001
rect 2621 370 2741 559
rect 3366 370 3466 559
rect 866 -101 1046 -89
rect 866 -153 878 -101
rect 1034 -153 1046 -101
rect 866 -165 1046 -153
rect 3000 -2266 3076 -2254
rect 3000 -2422 3012 -2266
rect 3064 -2422 3076 -2266
rect 3000 -2434 3076 -2422
<< via1 >>
rect 448 27045 500 27097
rect 734 18328 786 18380
rect 1747 18328 1799 18380
rect 1933 18328 1985 18380
rect 2985 18328 3037 18380
rect 3171 18328 3223 18380
rect 4224 18328 4276 18380
rect 4410 18328 4462 18380
rect 5429 18328 5481 18380
rect 4854 16356 4906 16408
rect 5040 16356 5092 16408
rect 3758 16128 3810 16180
rect 3969 16128 4021 16180
rect 4181 16128 4233 16180
rect 4392 16128 4444 16180
rect 536 15894 588 15946
rect 2278 15877 2330 15929
rect 2278 15691 2330 15743
rect 5365 10187 5417 10239
rect 5365 10001 5417 10053
rect 647 8811 699 8863
rect 833 8811 885 8863
rect 481 8471 533 8523
rect 481 8285 533 8337
rect 1505 6582 1557 6634
rect 1505 6396 1557 6448
rect 4651 5435 4703 5591
rect 5137 5435 5189 5591
rect 2277 3552 2329 3604
rect 2277 3366 2329 3418
rect 878 -153 1034 -101
rect 3012 -2422 3064 -2266
<< metal2 >>
rect 271 27118 478 27121
rect 271 27097 540 27118
rect 271 27045 448 27097
rect 500 27045 540 27097
rect 271 27025 540 27045
rect 271 27024 478 27025
rect 80 22626 174 26890
rect 80 22570 99 22626
rect 155 22570 174 22626
rect 80 22440 174 22570
rect 80 22384 99 22440
rect 155 22384 174 22440
rect 80 16131 174 22384
rect 271 15970 366 27024
rect 473 22626 568 26890
rect 473 22570 492 22626
rect 548 22570 568 22626
rect 473 22440 568 22570
rect 473 22384 492 22440
rect 548 22384 568 22440
rect 473 16131 568 22384
rect 5448 21179 5542 21217
rect 5448 21123 5467 21179
rect 5523 21123 5542 21179
rect 5448 21084 5542 21123
rect 4393 20860 4487 20898
rect 4393 20804 4412 20860
rect 4468 20804 4487 20860
rect 4393 20765 4487 20804
rect 4209 20531 4303 20569
rect 4209 20475 4228 20531
rect 4284 20475 4303 20531
rect 4209 20436 4303 20475
rect 3155 20218 3249 20256
rect 3155 20162 3174 20218
rect 3230 20162 3249 20218
rect 3155 20123 3249 20162
rect 2970 19558 3064 19596
rect 2970 19502 2989 19558
rect 3045 19502 3064 19558
rect 2970 19463 3064 19502
rect 1916 19246 2010 19284
rect 1916 19190 1935 19246
rect 1991 19190 2010 19246
rect 1916 19151 2010 19190
rect 1732 18919 1826 18957
rect 1732 18863 1751 18919
rect 1807 18863 1826 18919
rect 1732 18824 1826 18863
rect 678 18604 772 18642
rect 678 18548 697 18604
rect 753 18548 772 18604
rect 678 18509 772 18548
rect 699 18400 826 18401
rect 697 18380 826 18400
rect 697 18328 734 18380
rect 786 18328 826 18380
rect 697 18308 826 18328
rect 1717 18380 2025 18400
rect 1717 18328 1747 18380
rect 1799 18328 1933 18380
rect 1985 18328 2025 18380
rect 1717 18308 2025 18328
rect 2955 18380 3263 18400
rect 2955 18328 2985 18380
rect 3037 18328 3171 18380
rect 3223 18328 3263 18380
rect 2955 18308 3263 18328
rect 4194 18380 4502 18400
rect 4194 18328 4224 18380
rect 4276 18328 4410 18380
rect 4462 18328 4502 18380
rect 4194 18308 4502 18328
rect 5389 18380 5522 18401
rect 5389 18328 5429 18380
rect 5481 18328 5522 18380
rect 5389 18308 5522 18328
rect 697 16544 787 18308
rect 1826 16639 1916 18308
rect 3065 16639 3154 18308
rect 4303 16639 4393 18308
rect 5432 16432 5522 18308
rect 5045 16428 5522 16432
rect 4824 16408 5522 16428
rect 4824 16356 4854 16408
rect 4906 16356 5040 16408
rect 5092 16356 5522 16408
rect 4824 16336 5522 16356
rect 5045 16335 5522 16336
rect 3720 16182 4482 16220
rect 3720 16126 3756 16182
rect 3812 16126 3967 16182
rect 4023 16126 4179 16182
rect 4235 16126 4390 16182
rect 4446 16126 4482 16182
rect 3720 16087 4482 16126
rect 271 15946 628 15970
rect 271 15894 536 15946
rect 588 15894 628 15946
rect 271 15873 628 15894
rect 2072 10257 2166 15972
rect 2256 15929 2351 15970
rect 2256 15877 2278 15929
rect 2330 15877 2351 15929
rect 2256 15743 2351 15877
rect 2256 15691 2278 15743
rect 2330 15691 2351 15743
rect 1004 10192 1913 10248
rect 617 8863 926 8883
rect 617 8811 647 8863
rect 699 8811 833 8863
rect 885 8811 926 8863
rect 617 8791 926 8811
rect 461 8523 553 8563
rect 461 8471 481 8523
rect 533 8471 553 8523
rect 461 8427 553 8471
rect 460 8337 554 8427
rect 460 8285 481 8337
rect 533 8285 554 8337
rect 460 -1 554 8285
rect 831 7768 926 8791
rect 831 7634 1158 7768
rect 1063 5917 1158 7634
rect 1857 7689 1913 10192
rect 2256 7803 2351 15691
rect 2441 12624 2535 15972
rect 2441 12568 2460 12624
rect 2516 12568 2535 12624
rect 2441 12438 2535 12568
rect 2441 12382 2460 12438
rect 2516 12382 2535 12438
rect 2441 11849 2535 12382
rect 2441 11793 2460 11849
rect 2516 11793 2535 11849
rect 2441 11663 2535 11793
rect 2441 11607 2460 11663
rect 2516 11607 2535 11663
rect 2441 10933 2535 11607
rect 2441 10877 2460 10933
rect 2516 10877 2535 10933
rect 2441 10747 2535 10877
rect 2441 10691 2460 10747
rect 2516 10691 2535 10747
rect 2441 10257 2535 10691
rect 5345 10239 5437 10279
rect 5345 10187 5365 10239
rect 5417 10187 5437 10239
rect 5345 10100 5437 10187
rect 5344 10053 5438 10100
rect 5344 10001 5365 10053
rect 5417 10001 5438 10053
rect 4233 8339 4327 8518
rect 4692 8470 4786 8518
rect 4692 8373 5050 8470
rect 4233 8242 4435 8339
rect 4956 8158 5050 8373
rect 1857 7633 2004 7689
rect 2256 7687 2863 7803
rect 1497 6674 1591 6675
rect 1485 6634 1591 6674
rect 1485 6582 1505 6634
rect 1557 6582 1591 6634
rect 1485 6448 1591 6582
rect 1485 6396 1505 6448
rect 1557 6396 1591 6448
rect 1485 6356 1591 6396
rect 845 5811 1158 5917
rect 845 1505 940 5811
rect 1497 5738 1591 6356
rect 1948 6076 2004 7633
rect 1308 5625 1591 5738
rect 1877 6020 2004 6076
rect 911 -89 1006 1366
rect 1308 1 1402 5625
rect 1877 1853 1933 6020
rect 2298 4999 2354 5859
rect 2768 5039 2863 7687
rect 5344 6043 5438 10001
rect 4370 5909 4715 6043
rect 4639 5591 4715 5909
rect 4639 5435 4651 5591
rect 4703 5435 4715 5591
rect 4639 5423 4715 5435
rect 5125 5909 5438 6043
rect 5125 5591 5201 5909
rect 5125 5435 5137 5591
rect 5189 5435 5201 5591
rect 5125 5423 5201 5435
rect 2131 4989 2354 4999
rect 2131 4933 2141 4989
rect 2301 4933 2354 4989
rect 2466 4948 2863 5039
rect 2131 4923 2311 4933
rect 2466 4680 2577 4948
rect 2256 4594 2577 4680
rect 2256 3604 2351 4594
rect 2256 3552 2277 3604
rect 2329 3552 2351 3604
rect 2256 3418 2351 3552
rect 2256 3366 2277 3418
rect 2329 3366 2351 3418
rect 2256 3325 2351 3366
rect 1877 1797 1984 1853
rect 1928 986 1984 1797
rect 1928 910 2054 986
rect 866 -101 1046 -89
rect 866 -153 878 -101
rect 1034 -153 1046 -101
rect 866 -165 1046 -153
rect 1998 -1907 2054 910
rect 1998 -1963 3066 -1907
rect 3010 -2254 3066 -1963
rect 3000 -2266 3076 -2254
rect 3000 -2422 3012 -2266
rect 3064 -2422 3076 -2266
rect 3000 -2434 3076 -2422
<< via2 >>
rect 99 22570 155 22626
rect 99 22384 155 22440
rect 492 22570 548 22626
rect 492 22384 548 22440
rect 5467 21123 5523 21179
rect 4412 20804 4468 20860
rect 4228 20475 4284 20531
rect 3174 20162 3230 20218
rect 2989 19502 3045 19558
rect 1935 19190 1991 19246
rect 1751 18863 1807 18919
rect 697 18548 753 18604
rect 3756 16180 3812 16182
rect 3756 16128 3758 16180
rect 3758 16128 3810 16180
rect 3810 16128 3812 16180
rect 3756 16126 3812 16128
rect 3967 16180 4023 16182
rect 3967 16128 3969 16180
rect 3969 16128 4021 16180
rect 4021 16128 4023 16180
rect 3967 16126 4023 16128
rect 4179 16180 4235 16182
rect 4179 16128 4181 16180
rect 4181 16128 4233 16180
rect 4233 16128 4235 16180
rect 4179 16126 4235 16128
rect 4390 16180 4446 16182
rect 4390 16128 4392 16180
rect 4392 16128 4444 16180
rect 4444 16128 4446 16180
rect 4390 16126 4446 16128
rect 2460 12568 2516 12624
rect 2460 12382 2516 12438
rect 2460 11793 2516 11849
rect 2460 11607 2516 11663
rect 2460 10877 2516 10933
rect 2460 10691 2516 10747
rect 2141 4933 2301 4989
<< metal3 >>
rect -1 22626 324 23409
rect -1 22570 99 22626
rect 155 22570 324 22626
rect -1 22440 324 22570
rect -1 22384 99 22440
rect 155 22384 324 22440
rect -1 21410 324 22384
rect 474 22626 567 22664
rect 474 22570 492 22626
rect 548 22570 567 22626
rect 474 22440 567 22570
rect 474 22384 492 22440
rect 548 22384 567 22440
rect 474 22345 567 22384
rect 5448 21179 5542 21217
rect 5448 21123 5467 21179
rect 5523 21123 5542 21179
rect 5448 21084 5542 21123
rect 4393 20860 4487 20898
rect 4393 20804 4412 20860
rect 4468 20804 4487 20860
rect 4393 20765 4487 20804
rect 4209 20531 4303 20569
rect 4209 20475 4228 20531
rect 4284 20475 4303 20531
rect 4209 20436 4303 20475
rect 3155 20218 3249 20256
rect 3155 20162 3174 20218
rect 3230 20162 3249 20218
rect 3155 20123 3249 20162
rect 2970 19558 3064 19596
rect 2970 19502 2989 19558
rect 3045 19502 3064 19558
rect 2970 19463 3064 19502
rect 1916 19246 2010 19284
rect 1916 19190 1935 19246
rect 1991 19190 2010 19246
rect 1916 19151 2010 19190
rect 1732 18919 1826 18957
rect 1732 18863 1751 18919
rect 1807 18863 1826 18919
rect 1732 18824 1826 18863
rect 678 18604 772 18642
rect 678 18548 697 18604
rect 753 18548 772 18604
rect 678 18509 772 18548
rect 368 16182 5517 16228
rect 368 16126 3756 16182
rect 3812 16126 3967 16182
rect 4023 16126 4179 16182
rect 4235 16126 4390 16182
rect 4446 16126 5517 16182
rect 368 16000 5517 16126
rect 5493 12991 5794 15714
rect 2442 12624 2535 12662
rect 2442 12568 2460 12624
rect 2516 12568 2535 12624
rect 2442 12438 2535 12568
rect 2442 12382 2460 12438
rect 2516 12382 2535 12438
rect 2442 12343 2535 12382
rect 2442 11849 2535 11887
rect 2442 11793 2460 11849
rect 2516 11793 2535 11849
rect 2442 11663 2535 11793
rect 2442 11607 2460 11663
rect 2516 11607 2535 11663
rect 2442 11568 2535 11607
rect 2442 10933 2535 10971
rect 2442 10877 2460 10933
rect 2516 10877 2535 10933
rect 2442 10747 2535 10877
rect 2442 10691 2460 10747
rect 2516 10691 2535 10747
rect 2442 10652 2535 10691
rect 318 4989 2311 5005
rect 318 4933 2141 4989
rect 2301 4933 2311 4989
rect 318 4917 2311 4933
rect 5627 3128 5794 4490
rect 5636 149 5794 604
use M2_M1$$45012012_256x8m81  M2_M1$$45012012_256x8m81_0
timestamp 1669390400
transform 1 0 2570 0 1 16154
box -803 -67 803 66
use M2_M1$$45013036_256x8m81  M2_M1$$45013036_256x8m81_0
timestamp 1669390400
transform 1 0 4101 0 1 16154
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1669390400
transform 0 -1 5163 1 0 5513
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_1
timestamp 1669390400
transform 0 -1 4677 1 0 5513
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_2
timestamp 1669390400
transform 1 0 956 0 1 -127
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_0
timestamp 1669390400
transform 1 0 3038 0 1 -2344
box 0 0 1 1
use M3_M2$$43370540_256x8m81  M3_M2$$43370540_256x8m81_0
timestamp 1669390400
transform 1 0 4101 0 1 16154
box 0 0 1 1
use M3_M2$$44741676_256x8m81  M3_M2$$44741676_256x8m81_0
timestamp 1669390400
transform 1 0 2570 0 1 16154
box -803 -67 803 67
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_0
timestamp 1669390400
transform 1 0 2221 0 1 4961
box 0 0 1 1
use din_256x8m81  din_256x8m81_0
timestamp 1669390400
transform 1 0 323 0 1 7805
box -223 -57 2607 8999
use m2_saout01_256x8m81  m2_saout01_256x8m81_0
timestamp 1669390400
transform 1 0 686 0 1 28980
box -89 -63 4849 2153
use mux821_256x8m81  mux821_256x8m81_0
timestamp 1669390400
transform 1 0 553 0 1 16662
box -822 81 7080 12461
use outbuf_oe_256x8m81  outbuf_oe_256x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 5509
box -532 -359 5177 3324
use sa_256x8m81  sa_256x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 8608
box -357 -196 5034 8146
use sacntl_2_256x8m81  sacntl_2_256x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 23
box -530 -24 5176 5655
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1669390400
transform 1 0 2073 0 1 12344
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1669390400
transform 1 0 2073 0 1 11569
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1669390400
transform 1 0 2073 0 1 10653
box 0 -1 93 308
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1669390400
transform 0 1 5389 1 0 18308
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_1
timestamp 1669390400
transform 0 -1 628 1 0 15874
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_2
timestamp 1669390400
transform 0 -1 540 1 0 27025
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_3
timestamp 1669390400
transform 0 -1 826 1 0 18308
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1669390400
transform -1 0 2350 0 -1 15969
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1669390400
transform -1 0 1577 0 -1 6674
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1669390400
transform 1 0 2257 0 1 3326
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1669390400
transform 1 0 5345 0 1 9961
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1669390400
transform 1 0 461 0 1 8245
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1669390400
transform 0 -1 5132 1 0 16336
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1669390400
transform 0 -1 2025 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1669390400
transform 0 -1 3263 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_3
timestamp 1669390400
transform 0 -1 4502 1 0 18308
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_4
timestamp 1669390400
transform 0 -1 925 1 0 8791
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_0
timestamp 1669390400
transform -1 0 771 0 1 18510
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_1
timestamp 1669390400
transform -1 0 1825 0 1 18825
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_2
timestamp 1669390400
transform -1 0 2009 0 1 19152
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_3
timestamp 1669390400
transform -1 0 4302 0 1 20437
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_4
timestamp 1669390400
transform -1 0 4486 0 1 20766
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_5
timestamp 1669390400
transform -1 0 5541 0 1 21085
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_6
timestamp 1669390400
transform 1 0 2971 0 1 19464
box 0 0 1 1
use via2_256x8m81  via2_256x8m81_7
timestamp 1669390400
transform 1 0 3156 0 1 20124
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_0
timestamp 1669390400
transform 1 0 474 0 1 22346
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_1
timestamp 1669390400
transform 1 0 81 0 1 22346
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_2
timestamp 1669390400
transform 1 0 2442 0 1 12344
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_3
timestamp 1669390400
transform 1 0 2442 0 1 11569
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_4
timestamp 1669390400
transform 1 0 2442 0 1 10653
box 0 0 1 1
use wen_wm1_256x8m81  wen_wm1_256x8m81_0
timestamp 1669390400
transform 1 0 322 0 1 -3376
box -156 -24 4946 3287
<< labels >>
rlabel metal1 s 993 27075 993 27075 4 pcb
port 1 nsew
rlabel metal1 s 698 8313 698 8313 4 datain
port 2 nsew
rlabel metal1 s 993 27073 993 27073 4 pcb
port 1 nsew
rlabel metal1 s 933 18156 933 18156 4 vdd
port 3 nsew
flabel metal1 s 709 -3344 709 -3344 0 FreeSans 600 0 0 0 WEN
port 4 nsew
rlabel metal3 s 810 18907 810 18907 4 ypass[1]
port 5 nsew
rlabel metal3 s 810 19224 810 19224 4 ypass[2]
port 6 nsew
rlabel metal3 s 810 19542 810 19542 4 ypass[3]
port 7 nsew
rlabel metal3 s 810 20197 810 20197 4 ypass[4]
port 8 nsew
rlabel metal3 s 810 20521 810 20521 4 ypass[5]
port 9 nsew
rlabel metal3 s 810 20838 810 20838 4 ypass[6]
port 10 nsew
rlabel metal3 s 810 21156 810 21156 4 ypass[7]
port 11 nsew
rlabel metal3 s 881 1460 881 1460 4 men
port 12 nsew
rlabel metal3 s 373 1086 373 1086 4 vss
port 13 nsew
rlabel metal3 s 440 2179 440 2179 4 vss
port 13 nsew
rlabel metal3 s 810 20197 810 20197 4 ypass[4]
port 8 nsew
rlabel metal3 s 545 3843 545 3843 4 vdd
port 3 nsew
rlabel metal3 s 393 399 393 399 4 vdd
port 3 nsew
rlabel metal3 s 454 6155 454 6155 4 vss
port 13 nsew
rlabel metal3 s 439 11029 439 11029 4 vss
port 13 nsew
rlabel metal3 s 810 21156 810 21156 4 ypass[7]
port 11 nsew
rlabel metal3 s 810 20838 810 20838 4 ypass[6]
port 10 nsew
rlabel metal3 s 810 20521 810 20521 4 ypass[5]
port 9 nsew
rlabel metal3 s 810 19542 810 19542 4 ypass[3]
port 7 nsew
rlabel metal3 s 810 19224 810 19224 4 ypass[2]
port 6 nsew
rlabel metal3 s 810 18907 810 18907 4 ypass[1]
port 5 nsew
rlabel metal3 s 810 18585 810 18585 4 ypass[0]
port 14 nsew
rlabel metal3 s 398 1458 398 1458 4 men
port 12 nsew
rlabel metal3 s 933 28895 933 28895 4 vdd
port 3 nsew
rlabel metal3 s 949 22008 949 22008 4 vss
port 13 nsew
rlabel metal3 s 477 17166 477 17166 4 vss
port 13 nsew
rlabel metal3 s 466 13763 466 13763 4 vdd
port 3 nsew
rlabel metal3 s 401 8726 401 8726 4 vdd
port 3 nsew
rlabel metal3 s 335 7368 335 7368 4 vdd
port 3 nsew
rlabel metal3 s 810 18585 810 18585 4 ypass[0]
port 14 nsew
flabel metal3 s 644 4959 644 4959 0 FreeSans 600 0 0 0 GWE
port 15 nsew
rlabel metal3 s 393 -592 393 -592 4 vdd
port 3 nsew
rlabel metal3 s 373 -1762 373 -1762 4 vss
port 13 nsew
rlabel metal3 s 373 -2331 373 -2331 4 vss
port 13 nsew
rlabel metal3 s 393 -2997 393 -2997 4 vdd
port 3 nsew
rlabel metal3 s 373 -1375 373 -1375 4 vss
port 13 nsew
flabel metal3 s 705 -2005 705 -2005 0 FreeSans 600 0 0 0 GWEN
port 16 nsew
rlabel metal2 s 501 1625 501 1625 4 datain
port 2 nsew
rlabel metal2 s 5501 28725 5501 28725 4 b[7]
port 17 nsew
rlabel metal2 s 4464 28725 4464 28725 4 b[6]
port 18 nsew
rlabel metal2 s 4256 28725 4256 28725 4 b[5]
port 19 nsew
rlabel metal2 s 3228 28725 3228 28725 4 b[4]
port 20 nsew
rlabel metal2 s 3024 28725 3024 28725 4 b[3]
port 21 nsew
rlabel metal2 s 1983 28725 1983 28725 4 b[2]
port 22 nsew
rlabel metal2 s 1781 28725 1781 28725 4 b[1]
port 23 nsew
rlabel metal2 s 736 28727 736 28727 4 b[0]
port 24 nsew
rlabel metal2 s 4880 28727 4880 28727 4 bb[6]
port 25 nsew
rlabel metal2 s 5082 28734 5082 28734 4 bb[7]
port 26 nsew
rlabel metal2 s 3841 28727 3841 28727 4 bb[5]
port 27 nsew
rlabel metal2 s 1351 1158 1351 1158 4 q
port 28 nsew
rlabel metal2 s 3641 28727 3641 28727 4 bb[4]
port 29 nsew
rlabel metal2 s 2604 28734 2604 28734 4 bb[3]
port 30 nsew
rlabel metal2 s 2405 28730 2405 28730 4 bb[2]
port 31 nsew
rlabel metal2 s 1162 28725 1162 28725 4 bb[0]
port 32 nsew
rlabel metal2 s 1368 28725 1368 28725 4 bb[1]
port 33 nsew
rlabel metal2 s 1351 1124 1351 1124 4 q
port 28 nsew
<< properties >>
string GDS_END 819028
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 810674
string path 10.130 4.930 10.130 -9.675 15.190 -9.675 15.190 -12.125 
<< end >>
