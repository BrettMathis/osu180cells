magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1008 844
rect 49 312 115 579
rect 645 507 691 724
rect 49 231 790 312
rect 49 113 95 231
rect 645 60 691 185
rect 0 -60 1008 60
<< obsm1 >>
rect 849 437 915 636
rect 490 377 915 437
rect 869 115 915 377
<< labels >>
rlabel metal1 s 49 312 115 579 6 Z
port 1 nsew default bidirectional
rlabel metal1 s 49 231 790 312 6 Z
port 1 nsew default bidirectional
rlabel metal1 s 49 113 95 231 6 Z
port 1 nsew default bidirectional
rlabel metal1 s 0 724 1008 844 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 645 507 691 724 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 645 60 691 185 6 VSS
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1008 60 8 VSS
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1008 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 418222
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 415896
<< end >>
