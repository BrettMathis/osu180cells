magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -27 702 7407 2956
<< ndiff >>
rect 79 484 233 541
rect 79 438 133 484
rect 179 438 233 484
rect 79 320 233 438
rect 79 274 133 320
rect 179 274 233 320
rect 79 218 233 274
<< pdiff >>
rect 1938 843 1987 1035
rect 2212 843 2335 1035
rect 4378 1105 4435 1297
<< ndiffc >>
rect 133 438 179 484
rect 133 274 179 320
<< psubdiff >>
rect 4372 3525 4456 3544
rect 4372 3291 4391 3525
rect 4437 3291 4456 3525
rect 7032 3525 7210 3544
rect 4372 3272 4456 3291
rect 7032 3291 7051 3525
rect 7191 3291 7210 3525
rect 7032 3272 7210 3291
rect 7032 490 7210 509
rect 7032 256 7051 490
rect 7191 256 7210 490
rect 7032 237 7210 256
<< nsubdiff >>
rect 1706 2249 1790 2268
rect 1706 2015 1725 2249
rect 1771 2015 1790 2249
rect 1706 1996 1790 2015
rect 4372 2249 4456 2268
rect 4372 2015 4391 2249
rect 4437 2015 4456 2249
rect 4372 1996 4456 2015
rect 7032 2249 7210 2268
rect 7032 2015 7051 2249
rect 7191 2015 7210 2249
rect 7032 1996 7210 2015
rect 79 1186 233 1243
rect 79 1140 133 1186
rect 179 1140 233 1186
rect 79 1022 233 1140
rect 79 976 133 1022
rect 179 976 233 1022
rect 79 920 233 976
rect 7047 1186 7201 1243
rect 7047 1140 7101 1186
rect 7147 1140 7201 1186
rect 7047 1022 7201 1140
rect 7047 976 7101 1022
rect 7147 976 7201 1022
rect 7047 920 7201 976
<< psubdiffcont >>
rect 4391 3291 4437 3525
rect 7051 3291 7191 3525
rect 7051 256 7191 490
<< nsubdiffcont >>
rect 1725 2015 1771 2249
rect 4391 2015 4437 2249
rect 7051 2015 7191 2249
rect 133 1140 179 1186
rect 133 976 179 1022
rect 7101 1140 7147 1186
rect 7101 976 7147 1022
<< polysilicon >>
rect 252 1705 372 3369
rect 476 1705 596 3369
rect 700 1705 820 3369
rect 2023 3004 2143 3484
rect 2247 3004 2367 3484
rect 2471 3004 2591 3484
rect 2695 3004 2815 3484
rect 2919 3004 3039 3484
rect 3143 3004 3263 3484
rect 3367 3004 3487 3484
rect 3591 3004 3711 3484
rect 3815 3004 3935 3484
rect 4039 3004 4159 3484
rect 1607 2920 4159 3004
rect 1607 2870 1785 2920
rect 1607 2824 1626 2870
rect 1766 2824 1785 2870
rect 1607 2805 1785 2824
rect 2023 2737 2143 2920
rect 2247 2737 2367 2920
rect 2471 2737 2591 2920
rect 2695 2737 2815 2920
rect 2919 2737 3039 2920
rect 3143 2737 3263 2920
rect 3367 2737 3487 2920
rect 3591 2737 3711 2920
rect 3815 2737 3935 2920
rect 4039 2737 4159 2920
rect 924 1705 1044 2490
rect 1148 1705 1268 2490
rect 1372 1705 1492 2490
rect 252 1686 1492 1705
rect 252 1640 470 1686
rect 610 1640 1492 1686
rect 252 1621 1492 1640
rect 4669 1698 4789 3369
rect 4893 1698 5013 3369
rect 5117 1698 5237 3369
rect 5341 1698 5461 3369
rect 5565 1698 5685 3369
rect 5789 1698 5909 3369
rect 6013 1698 6133 3369
rect 6237 1698 6357 3369
rect 6461 1698 6581 3369
rect 6685 1698 6805 3369
rect 4669 1679 6805 1698
rect 4669 1633 5407 1679
rect 5547 1633 5849 1679
rect 5989 1633 6303 1679
rect 6443 1633 6646 1679
rect 6786 1633 6805 1679
rect 4669 1614 6805 1633
rect 1181 1459 2156 1520
rect 451 1429 629 1448
rect 451 1383 470 1429
rect 610 1383 629 1429
rect 451 1364 629 1383
rect 509 1297 629 1364
rect 733 1297 853 1370
rect 1181 1324 1301 1459
rect 1181 1297 1300 1324
rect 2036 1036 2156 1459
rect 4510 1469 4767 1488
rect 3950 1430 4426 1449
rect 3950 1384 4267 1430
rect 4407 1384 4426 1430
rect 3950 1365 4426 1384
rect 4510 1423 4608 1469
rect 4748 1423 4767 1469
rect 4510 1404 4767 1423
rect 509 827 628 843
rect 733 827 852 843
rect 509 441 629 827
rect 509 140 629 213
rect 733 103 853 827
rect 1181 819 1300 843
rect 1181 677 1301 819
rect 1011 658 1301 677
rect 1011 612 1030 658
rect 1170 612 1301 658
rect 1011 593 1301 612
rect 1364 764 1974 783
rect 1364 624 1383 764
rect 1429 722 1974 764
rect 1429 624 1448 722
rect 1883 685 1974 722
rect 2374 753 2494 819
rect 2374 734 2668 753
rect 2374 688 2509 734
rect 2649 688 2668 734
rect 1364 605 1448 624
rect 733 84 911 103
rect 733 38 752 84
rect 892 38 911 84
rect 733 19 911 38
rect 1181 32 1301 593
rect 1688 563 1808 636
rect 1883 624 2270 685
rect 2374 669 2668 688
rect 2374 583 2494 669
rect 1688 32 1808 108
rect 2822 89 2942 1341
rect 3950 1297 4070 1365
rect 4174 1297 4294 1365
rect 4510 1077 4630 1404
rect 4842 1217 4962 1614
rect 5307 1297 5426 1370
rect 5531 1297 5650 1370
rect 5755 1297 5874 1370
rect 5979 1297 6098 1370
rect 6203 1297 6322 1370
rect 6427 1297 6546 1370
rect 6651 1297 6770 1370
rect 1181 -73 1808 32
rect 2439 70 2942 89
rect 2439 24 2458 70
rect 2598 24 2942 70
rect 2439 5 2942 24
rect 3293 89 3413 816
rect 3517 89 3637 816
rect 3950 769 4070 843
rect 4174 769 4294 843
rect 3950 563 4069 636
rect 4174 563 4293 636
rect 4842 327 4962 1105
rect 5307 751 5427 908
rect 5531 751 5651 908
rect 5755 751 5875 908
rect 5979 751 6099 908
rect 6203 751 6323 908
rect 6427 751 6547 908
rect 6651 751 6771 908
rect 5154 732 6771 751
rect 5154 686 5173 732
rect 5313 686 6771 732
rect 5154 667 6771 686
rect 5307 563 5427 667
rect 5531 563 5651 667
rect 5755 563 5875 667
rect 5979 563 6099 667
rect 6203 563 6323 667
rect 6427 563 6547 667
rect 6651 563 6771 667
rect 5307 308 5426 380
rect 5531 308 5650 380
rect 5755 308 5874 380
rect 5979 308 6098 380
rect 6203 308 6322 380
rect 3293 70 3637 89
rect 3293 24 3312 70
rect 3452 24 3637 70
rect 3293 5 3637 24
rect 3950 8 4070 108
rect 4174 8 4294 108
rect 4618 83 4738 225
rect 1688 -182 1808 -73
rect 3950 -18 4294 8
rect 4560 64 4738 83
rect 4560 18 4579 64
rect 4719 18 4738 64
rect 4560 -1 4738 18
rect 3950 -64 3969 -18
rect 4109 -58 4294 -18
rect 4109 -64 4128 -58
rect 3950 -83 4128 -64
rect 1688 -201 1866 -182
rect 1688 -247 1707 -201
rect 1847 -247 1866 -201
rect 1688 -266 1866 -247
<< polycontact >>
rect 1626 2824 1766 2870
rect 470 1640 610 1686
rect 5407 1633 5547 1679
rect 5849 1633 5989 1679
rect 6303 1633 6443 1679
rect 6646 1633 6786 1679
rect 470 1383 610 1429
rect 4267 1384 4407 1430
rect 4608 1423 4748 1469
rect 1030 612 1170 658
rect 1383 624 1429 764
rect 2509 688 2649 734
rect 752 38 892 84
rect 2458 24 2598 70
rect 5173 686 5313 732
rect 3312 24 3452 70
rect 4579 18 4719 64
rect 3969 -64 4109 -18
rect 1707 -247 1847 -201
<< metal1 >>
rect 162 3543 238 3555
rect 162 3283 174 3543
rect 226 3283 238 3543
rect 610 3543 686 3555
rect 162 3271 238 3283
rect 401 2881 447 3360
rect 610 3283 622 3543
rect 674 3283 686 3543
rect 1933 3543 2009 3555
rect 610 3271 686 3283
rect 849 2881 895 3360
rect 1933 3283 1945 3543
rect 1997 3283 2009 3543
rect 2381 3543 2457 3555
rect 1933 3271 2009 3283
rect 2172 3052 2218 3360
rect 2381 3283 2393 3543
rect 2445 3283 2457 3543
rect 2829 3543 2905 3555
rect 2381 3271 2457 3283
rect 2003 3040 2391 3052
rect 2003 3037 2015 3040
rect 1397 2991 2015 3037
rect 2003 2988 2015 2991
rect 2379 3037 2391 3040
rect 2620 3037 2666 3360
rect 2829 3283 2841 3543
rect 2893 3283 2905 3543
rect 3277 3543 3353 3555
rect 2829 3271 2905 3283
rect 3068 3037 3114 3360
rect 3277 3283 3289 3543
rect 3341 3283 3353 3543
rect 3725 3543 3801 3555
rect 3277 3271 3353 3283
rect 3516 3037 3562 3360
rect 3725 3283 3737 3543
rect 3789 3283 3801 3543
rect 4173 3543 4249 3555
rect 3725 3271 3801 3283
rect 3964 3037 4010 3360
rect 4173 3283 4185 3543
rect 4237 3283 4249 3543
rect 4173 3271 4249 3283
rect 4376 3543 4452 3555
rect 4376 3283 4388 3543
rect 4440 3283 4452 3543
rect 4376 3271 4452 3283
rect 4579 3543 4655 3555
rect 4579 3283 4591 3543
rect 4643 3283 4655 3543
rect 5027 3543 5103 3555
rect 4579 3271 4655 3283
rect 2379 2991 4010 3037
rect 2379 2988 2391 2991
rect 2003 2976 2391 2988
rect 401 2870 1777 2881
rect 401 2824 1626 2870
rect 1766 2824 1777 2870
rect 401 2813 1777 2824
rect 162 2267 238 2279
rect 162 2007 174 2267
rect 226 2007 238 2267
rect 401 2260 447 2813
rect 610 2267 686 2279
rect 162 1995 238 2007
rect 610 2007 622 2267
rect 674 2007 686 2267
rect 849 2260 895 2813
rect 1058 2267 1134 2279
rect 610 1995 686 2007
rect 1058 2007 1070 2267
rect 1122 2007 1134 2267
rect 1297 2260 1343 2813
rect 1506 2267 1582 2279
rect 1058 1995 1134 2007
rect 1506 2007 1518 2267
rect 1570 2007 1582 2267
rect 1506 1995 1582 2007
rect 1710 2267 1786 2279
rect 1710 2007 1722 2267
rect 1774 2007 1786 2267
rect 1710 1995 1786 2007
rect 1933 2267 2009 2279
rect 1933 2007 1945 2267
rect 1997 2007 2009 2267
rect 2172 2260 2218 2976
rect 2381 2267 2457 2279
rect 1933 1995 2009 2007
rect 2381 2007 2393 2267
rect 2445 2007 2457 2267
rect 2620 2260 2666 2991
rect 2829 2267 2905 2279
rect 2381 1995 2457 2007
rect 2829 2007 2841 2267
rect 2893 2007 2905 2267
rect 3068 2260 3114 2991
rect 3277 2267 3353 2279
rect 2829 1995 2905 2007
rect 3277 2007 3289 2267
rect 3341 2007 3353 2267
rect 3516 2260 3562 2991
rect 3725 2267 3801 2279
rect 3277 1995 3353 2007
rect 3725 2007 3737 2267
rect 3789 2007 3801 2267
rect 3964 2260 4010 2991
rect 4818 3025 4864 3360
rect 5027 3283 5039 3543
rect 5091 3283 5103 3543
rect 5475 3543 5551 3555
rect 5027 3271 5103 3283
rect 5266 3025 5312 3360
rect 5475 3283 5487 3543
rect 5539 3283 5551 3543
rect 5923 3543 5999 3555
rect 5475 3271 5551 3283
rect 5714 3025 5760 3360
rect 5923 3283 5935 3543
rect 5987 3283 5999 3543
rect 6371 3543 6447 3555
rect 5923 3271 5999 3283
rect 6162 3025 6208 3360
rect 6371 3283 6383 3543
rect 6435 3283 6447 3543
rect 6819 3543 6895 3555
rect 6371 3271 6447 3283
rect 6610 3025 6656 3360
rect 6819 3283 6831 3543
rect 6883 3283 6895 3543
rect 6819 3271 6895 3283
rect 7038 3543 7218 3555
rect 7038 3283 7050 3543
rect 7206 3283 7218 3543
rect 7038 3271 7218 3283
rect 4818 2979 6656 3025
rect 4173 2267 4249 2279
rect 3725 1995 3801 2007
rect 4173 2007 4185 2267
rect 4237 2007 4249 2267
rect 4173 1995 4249 2007
rect 4376 2267 4452 2279
rect 4376 2007 4388 2267
rect 4440 2007 4452 2267
rect 4376 1995 4452 2007
rect 4579 2267 4655 2279
rect 4579 2007 4591 2267
rect 4643 2007 4655 2267
rect 4818 2260 4864 2979
rect 5027 2267 5103 2279
rect 4579 1995 4655 2007
rect 5027 2007 5039 2267
rect 5091 2007 5103 2267
rect 5266 2260 5312 2979
rect 5475 2267 5551 2279
rect 5027 1995 5103 2007
rect 5475 2007 5487 2267
rect 5539 2007 5551 2267
rect 5714 2260 5760 2979
rect 5923 2267 5999 2279
rect 5475 1995 5551 2007
rect 5923 2007 5935 2267
rect 5987 2007 5999 2267
rect 6162 2260 6208 2979
rect 6371 2267 6447 2279
rect 5923 1995 5999 2007
rect 6371 2007 6383 2267
rect 6435 2007 6447 2267
rect 6610 2260 6656 2979
rect 6819 2267 6895 2279
rect 6371 1995 6447 2007
rect 6819 2007 6831 2267
rect 6883 2007 6895 2267
rect 6819 1995 6895 2007
rect 7032 2267 7212 2279
rect 7032 2007 7044 2267
rect 7200 2007 7212 2267
rect 7032 1995 7212 2007
rect 459 1686 621 1697
rect 459 1640 470 1686
rect 610 1640 621 1686
rect 459 1429 621 1640
rect 5396 1679 5558 1690
rect 5396 1633 5407 1679
rect 5547 1633 5558 1679
rect 5396 1622 5558 1633
rect 5838 1679 6000 1690
rect 5838 1633 5849 1679
rect 5989 1633 6000 1679
rect 5838 1622 6000 1633
rect 6292 1679 6454 1690
rect 6292 1633 6303 1679
rect 6443 1633 6454 1679
rect 6292 1622 6454 1633
rect 6635 1679 6846 1690
rect 6635 1633 6646 1679
rect 6786 1633 6846 1679
rect 6635 1622 6846 1633
rect 459 1383 470 1429
rect 610 1383 621 1429
rect 459 1372 621 1383
rect 882 1563 4327 1609
rect 882 1261 928 1563
rect 1262 1476 1442 1488
rect 1262 1424 1274 1476
rect 1430 1424 1442 1476
rect 1262 1412 1442 1424
rect 3442 1457 4145 1512
rect 91 1216 221 1257
rect 1064 1246 1193 1289
rect 91 1164 130 1216
rect 182 1164 221 1216
rect 91 1140 133 1164
rect 179 1140 221 1164
rect 91 1022 221 1140
rect 91 998 133 1022
rect 179 998 221 1022
rect 91 946 130 998
rect 182 946 221 998
rect 91 906 221 946
rect 616 1205 746 1246
rect 616 1153 655 1205
rect 707 1153 746 1205
rect 616 987 746 1153
rect 616 935 655 987
rect 707 935 746 987
rect 91 514 221 555
rect 91 462 130 514
rect 182 462 221 514
rect 91 438 133 462
rect 179 438 221 462
rect 91 320 221 438
rect 91 296 133 320
rect 179 296 221 320
rect 91 244 130 296
rect 182 244 221 296
rect 91 204 221 244
rect 434 -85 480 902
rect 616 895 746 935
rect 1064 1205 1194 1246
rect 1064 1153 1103 1205
rect 1155 1153 1194 1205
rect 1064 987 1194 1153
rect 1064 935 1103 987
rect 1155 935 1194 987
rect 882 669 928 902
rect 1064 895 1194 935
rect 1064 852 1193 895
rect 1330 775 1376 1412
rect 1572 1164 1700 1289
rect 1572 1112 1610 1164
rect 1662 1112 1700 1164
rect 1572 947 1700 1112
rect 1572 895 1610 947
rect 1662 895 1700 947
rect 1330 764 1440 775
rect 882 658 1181 669
rect 882 612 1030 658
rect 1170 612 1181 658
rect 882 601 1181 612
rect 1330 624 1383 764
rect 1429 624 1440 764
rect 1330 613 1440 624
rect 1572 729 1700 895
rect 1572 677 1610 729
rect 1662 677 1700 729
rect 616 514 746 555
rect 616 462 655 514
rect 707 462 746 514
rect 616 296 746 462
rect 616 244 655 296
rect 707 244 746 296
rect 616 204 746 244
rect 882 221 928 601
rect 1065 513 1193 554
rect 1065 461 1103 513
rect 1155 461 1193 513
rect 1065 327 1193 461
rect 1065 275 1103 327
rect 1155 275 1193 327
rect 1065 235 1193 275
rect 632 84 972 95
rect 632 55 752 84
rect 892 55 972 84
rect 632 3 670 55
rect 722 38 752 55
rect 722 3 882 38
rect 934 3 972 55
rect 632 -38 972 3
rect 1330 -76 1376 613
rect 1572 511 1700 677
rect 1572 459 1610 511
rect 1662 459 1700 511
rect 1572 294 1700 459
rect 1572 242 1610 294
rect 1662 242 1700 294
rect 1572 201 1700 242
rect 1796 1035 1924 1289
rect 2299 1036 2345 1289
rect 2481 1246 2609 1289
rect 1796 843 2005 1035
rect 2190 843 2345 1036
rect 2480 1205 2610 1246
rect 2480 1153 2519 1205
rect 2571 1153 2610 1205
rect 2480 987 2610 1153
rect 2480 935 2519 987
rect 2571 935 2610 987
rect 2480 895 2610 935
rect 2481 852 2609 895
rect 1796 554 1924 843
rect 1796 380 2155 554
rect 2299 380 2345 843
rect 2734 745 2806 1289
rect 2929 1246 3057 1289
rect 2928 1205 3058 1246
rect 2928 1153 2967 1205
rect 3019 1153 3058 1205
rect 2928 987 3058 1153
rect 2928 935 2967 987
rect 3019 935 3058 987
rect 3203 1219 3279 1231
rect 3203 959 3215 1219
rect 3267 959 3279 1219
rect 3203 947 3279 959
rect 2928 895 3058 935
rect 2929 852 3057 895
rect 2498 734 2806 745
rect 2498 688 2509 734
rect 2649 688 2806 734
rect 2498 677 2806 688
rect 2481 513 2609 554
rect 2481 461 2519 513
rect 2571 461 2609 513
rect 1796 81 1924 380
rect 2481 327 2609 461
rect 2481 275 2519 327
rect 2571 275 2609 327
rect 2481 235 2609 275
rect 2734 81 2806 677
rect 2929 513 3057 554
rect 2929 461 2967 513
rect 3019 461 3057 513
rect 2929 327 3057 461
rect 2929 275 2967 327
rect 3019 275 3057 327
rect 2929 235 3057 275
rect 3203 490 3279 502
rect 3203 230 3215 490
rect 3267 230 3279 490
rect 3442 382 3488 1457
rect 3651 1219 3727 1231
rect 3651 959 3663 1219
rect 3715 959 3727 1219
rect 3651 947 3727 959
rect 3833 763 3961 1289
rect 4099 1246 4145 1457
rect 4281 1441 4327 1563
rect 4590 1476 4770 1488
rect 4256 1430 4418 1441
rect 4256 1384 4267 1430
rect 4407 1384 4418 1430
rect 4590 1424 4602 1476
rect 4758 1424 4770 1476
rect 4590 1423 4608 1424
rect 4748 1423 4770 1424
rect 4590 1412 4770 1423
rect 4256 1373 4418 1384
rect 4056 1205 4186 1246
rect 4056 1153 4095 1205
rect 4147 1153 4186 1205
rect 4056 987 4186 1153
rect 4056 935 4095 987
rect 4147 935 4186 987
rect 4056 895 4186 935
rect 4323 1105 4475 1297
rect 4659 1205 4855 1298
rect 4950 1246 5078 1289
rect 5191 1254 5319 1289
rect 4659 1153 4764 1205
rect 4816 1153 4855 1205
rect 4659 1105 4855 1153
rect 4099 852 4145 895
rect 4323 763 4409 1105
rect 4725 987 4855 1105
rect 4725 935 4764 987
rect 4816 935 4855 987
rect 4725 895 4855 935
rect 4949 1205 5079 1246
rect 4949 1153 4988 1205
rect 5040 1153 5079 1205
rect 4949 987 5079 1153
rect 4949 935 4988 987
rect 5040 935 5079 987
rect 4949 895 5079 935
rect 5190 1214 5320 1254
rect 5190 1162 5229 1214
rect 5281 1162 5320 1214
rect 5190 996 5320 1162
rect 5190 944 5229 996
rect 5281 944 5320 996
rect 5190 903 5320 944
rect 4950 852 5078 895
rect 5191 852 5319 903
rect 3833 743 4409 763
rect 5418 763 5534 1622
rect 5638 1254 5767 1289
rect 5638 1214 5768 1254
rect 5638 1162 5677 1214
rect 5729 1162 5768 1214
rect 5638 996 5768 1162
rect 5638 944 5677 996
rect 5729 944 5768 996
rect 5638 903 5768 944
rect 5638 852 5767 903
rect 5866 763 5981 1622
rect 6086 1254 6215 1289
rect 6086 1214 6216 1254
rect 6086 1162 6125 1214
rect 6177 1162 6216 1214
rect 6086 996 6216 1162
rect 6086 944 6125 996
rect 6177 944 6216 996
rect 6086 903 6216 944
rect 6086 852 6215 903
rect 6314 763 6429 1622
rect 6534 1254 6663 1289
rect 6534 1214 6664 1254
rect 6534 1162 6573 1214
rect 6625 1162 6664 1214
rect 6534 996 6664 1162
rect 6534 944 6573 996
rect 6625 944 6664 996
rect 6534 903 6664 944
rect 6534 852 6663 903
rect 6762 763 6846 1622
rect 7059 1216 7189 1257
rect 7059 1164 7098 1216
rect 7150 1164 7189 1216
rect 7059 1140 7101 1164
rect 7147 1140 7189 1164
rect 7059 1022 7189 1140
rect 7059 998 7101 1022
rect 7147 998 7189 1022
rect 7059 946 7098 998
rect 7150 946 7189 998
rect 7059 906 7189 946
rect 3833 732 5324 743
rect 3833 686 5173 732
rect 5313 686 5324 732
rect 3833 675 5324 686
rect 3833 667 5275 675
rect 3833 643 4409 667
rect 3651 490 3727 502
rect 3203 218 3279 230
rect 3651 230 3663 490
rect 3715 230 3727 490
rect 3651 218 3727 230
rect 3833 117 3961 643
rect 4057 512 4185 554
rect 4056 471 4186 512
rect 4056 419 4095 471
rect 4147 419 4186 471
rect 4056 253 4186 419
rect 4056 201 4095 253
rect 4147 201 4186 253
rect 4056 161 4186 201
rect 4057 117 4185 161
rect 4281 117 4409 643
rect 4543 398 4589 667
rect 5418 643 6846 763
rect 4950 513 5078 554
rect 4725 471 4855 512
rect 4725 419 4764 471
rect 4816 419 4855 471
rect 4725 253 4855 419
rect 4725 201 4764 253
rect 4816 201 4855 253
rect 4950 461 4988 513
rect 5040 461 5078 513
rect 4950 327 5078 461
rect 4950 275 4988 327
rect 5040 275 5078 327
rect 4950 235 5078 275
rect 5190 514 5320 555
rect 5190 462 5229 514
rect 5281 462 5320 514
rect 5190 296 5320 462
rect 5418 389 5534 643
rect 5638 514 5768 555
rect 5638 462 5677 514
rect 5729 462 5768 514
rect 5190 244 5229 296
rect 5281 244 5320 296
rect 5190 204 5320 244
rect 5638 296 5768 462
rect 5866 389 5981 643
rect 6086 514 6216 555
rect 6086 462 6125 514
rect 6177 462 6216 514
rect 5638 244 5677 296
rect 5729 244 5768 296
rect 5638 204 5768 244
rect 6086 296 6216 462
rect 6314 389 6429 643
rect 6534 514 6664 555
rect 6534 462 6573 514
rect 6625 462 6664 514
rect 6086 244 6125 296
rect 6177 244 6216 296
rect 6086 204 6216 244
rect 6534 296 6664 462
rect 6800 381 6846 643
rect 7038 508 7218 520
rect 6534 244 6573 296
rect 6625 244 6664 296
rect 6534 204 6664 244
rect 7038 248 7050 508
rect 7206 248 7218 508
rect 7038 236 7218 248
rect 4725 161 4855 201
rect 1796 70 2609 81
rect 1796 24 2458 70
rect 2598 24 2609 70
rect 1796 13 2609 24
rect 2734 70 3463 81
rect 2734 24 3312 70
rect 3452 24 3463 70
rect 2734 13 3463 24
rect 4568 64 4730 75
rect 4568 18 4579 64
rect 4719 18 4730 64
rect 4568 7 4730 18
rect 3958 -18 4120 -7
rect 3958 -64 3969 -18
rect 4109 -64 4120 -18
rect 3958 -76 4120 -64
rect 366 -97 546 -85
rect 366 -149 378 -97
rect 534 -149 546 -97
rect 1330 -122 4120 -76
rect 366 -161 546 -149
rect 1696 -201 1858 -190
rect 4633 -201 4679 7
rect 1696 -247 1707 -201
rect 1847 -247 4679 -201
rect 1696 -258 1858 -247
<< via1 >>
rect 174 3283 226 3543
rect 622 3283 674 3543
rect 1945 3283 1997 3543
rect 2393 3283 2445 3543
rect 2015 2988 2379 3040
rect 2841 3283 2893 3543
rect 3289 3283 3341 3543
rect 3737 3283 3789 3543
rect 4185 3283 4237 3543
rect 4388 3525 4440 3543
rect 4388 3291 4391 3525
rect 4391 3291 4437 3525
rect 4437 3291 4440 3525
rect 4388 3283 4440 3291
rect 4591 3283 4643 3543
rect 174 2007 226 2267
rect 622 2007 674 2267
rect 1070 2007 1122 2267
rect 1518 2007 1570 2267
rect 1722 2249 1774 2267
rect 1722 2015 1725 2249
rect 1725 2015 1771 2249
rect 1771 2015 1774 2249
rect 1722 2007 1774 2015
rect 1945 2007 1997 2267
rect 2393 2007 2445 2267
rect 2841 2007 2893 2267
rect 3289 2007 3341 2267
rect 3737 2007 3789 2267
rect 5039 3283 5091 3543
rect 5487 3283 5539 3543
rect 5935 3283 5987 3543
rect 6383 3283 6435 3543
rect 6831 3283 6883 3543
rect 7050 3525 7206 3543
rect 7050 3291 7051 3525
rect 7051 3291 7191 3525
rect 7191 3291 7206 3525
rect 7050 3283 7206 3291
rect 4185 2007 4237 2267
rect 4388 2249 4440 2267
rect 4388 2015 4391 2249
rect 4391 2015 4437 2249
rect 4437 2015 4440 2249
rect 4388 2007 4440 2015
rect 4591 2007 4643 2267
rect 5039 2007 5091 2267
rect 5487 2007 5539 2267
rect 5935 2007 5987 2267
rect 6383 2007 6435 2267
rect 6831 2007 6883 2267
rect 7044 2249 7200 2267
rect 7044 2015 7051 2249
rect 7051 2015 7191 2249
rect 7191 2015 7200 2249
rect 7044 2007 7200 2015
rect 1274 1424 1430 1476
rect 130 1186 182 1216
rect 130 1164 133 1186
rect 133 1164 179 1186
rect 179 1164 182 1186
rect 130 976 133 998
rect 133 976 179 998
rect 179 976 182 998
rect 130 946 182 976
rect 655 1153 707 1205
rect 655 935 707 987
rect 130 484 182 514
rect 130 462 133 484
rect 133 462 179 484
rect 179 462 182 484
rect 130 274 133 296
rect 133 274 179 296
rect 179 274 182 296
rect 130 244 182 274
rect 1103 1153 1155 1205
rect 1103 935 1155 987
rect 1610 1112 1662 1164
rect 1610 895 1662 947
rect 1610 677 1662 729
rect 655 462 707 514
rect 655 244 707 296
rect 1103 461 1155 513
rect 1103 275 1155 327
rect 670 3 722 55
rect 882 38 892 55
rect 892 38 934 55
rect 882 3 934 38
rect 1610 459 1662 511
rect 1610 242 1662 294
rect 2519 1153 2571 1205
rect 2519 935 2571 987
rect 2967 1153 3019 1205
rect 2967 935 3019 987
rect 3215 959 3267 1219
rect 2519 461 2571 513
rect 2519 275 2571 327
rect 2967 461 3019 513
rect 2967 275 3019 327
rect 3215 230 3267 490
rect 3663 959 3715 1219
rect 4602 1469 4758 1476
rect 4602 1424 4608 1469
rect 4608 1424 4748 1469
rect 4748 1424 4758 1469
rect 4095 1153 4147 1205
rect 4095 935 4147 987
rect 4764 1153 4816 1205
rect 4764 935 4816 987
rect 4988 1153 5040 1205
rect 4988 935 5040 987
rect 5229 1162 5281 1214
rect 5229 944 5281 996
rect 5677 1162 5729 1214
rect 5677 944 5729 996
rect 6125 1162 6177 1214
rect 6125 944 6177 996
rect 6573 1162 6625 1214
rect 6573 944 6625 996
rect 7098 1186 7150 1216
rect 7098 1164 7101 1186
rect 7101 1164 7147 1186
rect 7147 1164 7150 1186
rect 7098 976 7101 998
rect 7101 976 7147 998
rect 7147 976 7150 998
rect 7098 946 7150 976
rect 3663 230 3715 490
rect 4095 419 4147 471
rect 4095 201 4147 253
rect 4764 419 4816 471
rect 4764 201 4816 253
rect 4988 461 5040 513
rect 4988 275 5040 327
rect 5229 462 5281 514
rect 5677 462 5729 514
rect 5229 244 5281 296
rect 6125 462 6177 514
rect 5677 244 5729 296
rect 6573 462 6625 514
rect 6125 244 6177 296
rect 6573 244 6625 296
rect 7050 490 7206 508
rect 7050 256 7051 490
rect 7051 256 7191 490
rect 7191 256 7206 490
rect 7050 248 7206 256
rect 378 -149 534 -97
<< metal2 >>
rect 162 3545 238 3555
rect 162 3281 172 3545
rect 228 3281 238 3545
rect 162 3271 238 3281
rect 610 3545 686 3555
rect 610 3281 620 3545
rect 676 3281 686 3545
rect 610 3271 686 3281
rect 1933 3545 2009 3555
rect 1933 3281 1943 3545
rect 1999 3281 2009 3545
rect 1933 3271 2009 3281
rect 2381 3545 2457 3555
rect 2381 3281 2391 3545
rect 2447 3281 2457 3545
rect 2381 3271 2457 3281
rect 2829 3545 2905 3555
rect 2829 3281 2839 3545
rect 2895 3281 2905 3545
rect 2829 3271 2905 3281
rect 3277 3545 3353 3555
rect 3277 3281 3287 3545
rect 3343 3281 3353 3545
rect 3277 3271 3353 3281
rect 3725 3545 3801 3555
rect 3725 3281 3735 3545
rect 3791 3281 3801 3545
rect 3725 3271 3801 3281
rect 4173 3545 4249 3555
rect 4173 3281 4183 3545
rect 4239 3281 4249 3545
rect 4173 3271 4249 3281
rect 4376 3545 4452 3555
rect 4376 3281 4386 3545
rect 4442 3281 4452 3545
rect 4376 3271 4452 3281
rect 4579 3545 4655 3555
rect 4579 3281 4589 3545
rect 4645 3281 4655 3545
rect 4579 3271 4655 3281
rect 5027 3545 5103 3555
rect 5027 3281 5037 3545
rect 5093 3281 5103 3545
rect 5027 3271 5103 3281
rect 5475 3545 5551 3555
rect 5475 3281 5485 3545
rect 5541 3281 5551 3545
rect 5475 3271 5551 3281
rect 5923 3545 5999 3555
rect 5923 3281 5933 3545
rect 5989 3281 5999 3545
rect 5923 3271 5999 3281
rect 6371 3545 6447 3555
rect 6371 3281 6381 3545
rect 6437 3281 6447 3545
rect 6371 3271 6447 3281
rect 6819 3545 6895 3555
rect 6819 3281 6829 3545
rect 6885 3281 6895 3545
rect 6819 3271 6895 3281
rect 7038 3545 7218 3555
rect 7038 3281 7048 3545
rect 7208 3281 7218 3545
rect 7038 3271 7218 3281
rect 2003 3042 2391 3052
rect 2003 2986 2013 3042
rect 2381 2986 2391 3042
rect 2003 2976 2391 2986
rect 162 2269 238 2279
rect 162 2005 172 2269
rect 228 2005 238 2269
rect 162 1995 238 2005
rect 610 2269 686 2279
rect 610 2005 620 2269
rect 676 2005 686 2269
rect 610 1995 686 2005
rect 1058 2269 1134 2279
rect 1058 2005 1068 2269
rect 1124 2005 1134 2269
rect 1058 1995 1134 2005
rect 1506 2269 1582 2279
rect 1506 2005 1516 2269
rect 1572 2005 1582 2269
rect 1506 1995 1582 2005
rect 1710 2269 1786 2279
rect 1710 2005 1720 2269
rect 1776 2005 1786 2269
rect 1710 1995 1786 2005
rect 1933 2269 2009 2279
rect 1933 2005 1943 2269
rect 1999 2005 2009 2269
rect 1933 1995 2009 2005
rect 2381 2269 2457 2279
rect 2381 2005 2391 2269
rect 2447 2005 2457 2269
rect 2381 1995 2457 2005
rect 2829 2269 2905 2279
rect 2829 2005 2839 2269
rect 2895 2005 2905 2269
rect 2829 1995 2905 2005
rect 3277 2269 3353 2279
rect 3277 2005 3287 2269
rect 3343 2005 3353 2269
rect 3277 1995 3353 2005
rect 3725 2269 3801 2279
rect 3725 2005 3735 2269
rect 3791 2005 3801 2269
rect 3725 1995 3801 2005
rect 4173 2269 4249 2279
rect 4173 2005 4183 2269
rect 4239 2005 4249 2269
rect 4173 1995 4249 2005
rect 4376 2269 4452 2279
rect 4376 2005 4386 2269
rect 4442 2005 4452 2269
rect 4376 1995 4452 2005
rect 4579 2269 4655 2279
rect 4579 2005 4589 2269
rect 4645 2005 4655 2269
rect 4579 1995 4655 2005
rect 5027 2269 5103 2279
rect 5027 2005 5037 2269
rect 5093 2005 5103 2269
rect 5027 1995 5103 2005
rect 5475 2269 5551 2279
rect 5475 2005 5485 2269
rect 5541 2005 5551 2269
rect 5475 1995 5551 2005
rect 5923 2269 5999 2279
rect 5923 2005 5933 2269
rect 5989 2005 5999 2269
rect 5923 1995 5999 2005
rect 6371 2269 6447 2279
rect 6371 2005 6381 2269
rect 6437 2005 6447 2269
rect 6371 1995 6447 2005
rect 6819 2269 6895 2279
rect 6819 2005 6829 2269
rect 6885 2005 6895 2269
rect 6819 1995 6895 2005
rect 7032 2269 7212 2279
rect 7032 2005 7042 2269
rect 7202 2005 7212 2269
rect 7032 1995 7212 2005
rect 1262 1478 1442 1488
rect 1262 1422 1272 1478
rect 1432 1422 1442 1478
rect 1262 1412 1442 1422
rect 4590 1478 4770 1488
rect 4590 1422 4600 1478
rect 4760 1422 4770 1478
rect 4590 1412 4770 1422
rect 91 1218 221 1257
rect 91 1162 128 1218
rect 184 1162 221 1218
rect 91 1000 221 1162
rect 91 944 128 1000
rect 184 944 221 1000
rect 91 906 221 944
rect 616 1207 746 1246
rect 616 1151 653 1207
rect 709 1151 746 1207
rect 616 989 746 1151
rect 616 933 653 989
rect 709 933 746 989
rect 616 895 746 933
rect 1064 1207 1194 1246
rect 1064 1151 1101 1207
rect 1157 1151 1194 1207
rect 1064 989 1194 1151
rect 1064 933 1101 989
rect 1157 933 1194 989
rect 1064 895 1194 933
rect 1572 1164 1700 1289
rect 4057 1246 4185 1289
rect 4726 1246 4854 1289
rect 1572 1112 1610 1164
rect 1662 1112 1700 1164
rect 1572 947 1700 1112
rect 1572 895 1610 947
rect 1662 895 1700 947
rect 2480 1207 2610 1246
rect 2480 1151 2517 1207
rect 2573 1151 2610 1207
rect 2480 989 2610 1151
rect 2480 933 2517 989
rect 2573 933 2610 989
rect 2480 895 2610 933
rect 2928 1207 3058 1246
rect 2928 1151 2965 1207
rect 3021 1151 3058 1207
rect 2928 989 3058 1151
rect 2928 933 2965 989
rect 3021 933 3058 989
rect 3203 1221 3279 1231
rect 3203 957 3213 1221
rect 3269 957 3279 1221
rect 3203 947 3279 957
rect 3651 1221 3727 1231
rect 3651 957 3661 1221
rect 3717 957 3727 1221
rect 3651 947 3727 957
rect 4056 1205 4186 1246
rect 4056 1153 4095 1205
rect 4147 1153 4186 1205
rect 4056 987 4186 1153
rect 2928 895 3058 933
rect 4056 935 4095 987
rect 4147 935 4186 987
rect 4056 895 4186 935
rect 4725 1205 4855 1246
rect 4725 1153 4764 1205
rect 4816 1153 4855 1205
rect 4725 987 4855 1153
rect 4725 935 4764 987
rect 4816 935 4855 987
rect 4725 895 4855 935
rect 4949 1207 5079 1246
rect 4949 1151 4986 1207
rect 5042 1151 5079 1207
rect 4949 989 5079 1151
rect 4949 933 4986 989
rect 5042 933 5079 989
rect 4949 895 5079 933
rect 5190 1216 5320 1254
rect 5190 1160 5227 1216
rect 5283 1160 5320 1216
rect 5190 998 5320 1160
rect 5190 942 5227 998
rect 5283 942 5320 998
rect 5190 903 5320 942
rect 5638 1216 5768 1254
rect 5638 1160 5675 1216
rect 5731 1160 5768 1216
rect 5638 998 5768 1160
rect 5638 942 5675 998
rect 5731 942 5768 998
rect 5638 903 5768 942
rect 6086 1216 6216 1254
rect 6086 1160 6123 1216
rect 6179 1160 6216 1216
rect 6086 998 6216 1160
rect 6086 942 6123 998
rect 6179 942 6216 998
rect 6086 903 6216 942
rect 6534 1216 6664 1254
rect 6534 1160 6571 1216
rect 6627 1160 6664 1216
rect 6534 998 6664 1160
rect 6534 942 6571 998
rect 6627 942 6664 998
rect 6534 903 6664 942
rect 7059 1218 7189 1257
rect 7059 1162 7096 1218
rect 7152 1162 7189 1218
rect 7059 1000 7189 1162
rect 7059 944 7096 1000
rect 7152 944 7189 1000
rect 7059 906 7189 944
rect 1572 729 1700 895
rect 1572 677 1610 729
rect 1662 677 1700 729
rect 91 516 221 555
rect 91 460 128 516
rect 184 460 221 516
rect 91 298 221 460
rect 91 242 128 298
rect 184 242 221 298
rect 91 204 221 242
rect 616 516 746 555
rect 616 460 653 516
rect 709 460 746 516
rect 616 298 746 460
rect 616 242 653 298
rect 709 242 746 298
rect 616 204 746 242
rect 1065 515 1193 554
rect 1065 459 1101 515
rect 1157 459 1193 515
rect 1065 329 1193 459
rect 1065 273 1101 329
rect 1157 273 1193 329
rect 1065 235 1193 273
rect 1572 511 1700 677
rect 1572 459 1610 511
rect 1662 459 1700 511
rect 1572 294 1700 459
rect 1572 242 1610 294
rect 1662 242 1700 294
rect 1572 201 1700 242
rect 2481 515 2609 554
rect 2481 459 2517 515
rect 2573 459 2609 515
rect 2481 329 2609 459
rect 2481 273 2517 329
rect 2573 273 2609 329
rect 2481 235 2609 273
rect 2929 515 3057 554
rect 2929 459 2965 515
rect 3021 459 3057 515
rect 4057 512 4185 895
rect 4726 512 4854 895
rect 4950 515 5078 554
rect 2929 329 3057 459
rect 2929 273 2965 329
rect 3021 273 3057 329
rect 2929 235 3057 273
rect 3203 492 3279 502
rect 3203 228 3213 492
rect 3269 228 3279 492
rect 3203 218 3279 228
rect 3651 492 3727 502
rect 3651 228 3661 492
rect 3717 228 3727 492
rect 3651 218 3727 228
rect 4056 471 4186 512
rect 4056 419 4095 471
rect 4147 419 4186 471
rect 4056 253 4186 419
rect 4056 201 4095 253
rect 4147 201 4186 253
rect 632 56 972 96
rect 632 0 668 56
rect 724 0 880 56
rect 936 0 972 56
rect 632 -38 972 0
rect 366 -94 546 -85
rect 1608 -94 1664 201
rect 4056 161 4186 201
rect 4725 471 4855 512
rect 4725 419 4764 471
rect 4816 419 4855 471
rect 4725 253 4855 419
rect 4725 201 4764 253
rect 4816 201 4855 253
rect 4950 459 4986 515
rect 5042 459 5078 515
rect 4950 329 5078 459
rect 4950 273 4986 329
rect 5042 273 5078 329
rect 4950 235 5078 273
rect 5190 516 5320 555
rect 5190 460 5227 516
rect 5283 460 5320 516
rect 5190 298 5320 460
rect 5190 242 5227 298
rect 5283 242 5320 298
rect 5190 204 5320 242
rect 5638 516 5768 555
rect 5638 460 5675 516
rect 5731 460 5768 516
rect 5638 298 5768 460
rect 5638 242 5675 298
rect 5731 242 5768 298
rect 5638 204 5768 242
rect 6086 516 6216 555
rect 6086 460 6123 516
rect 6179 460 6216 516
rect 6086 298 6216 460
rect 6086 242 6123 298
rect 6179 242 6216 298
rect 6086 204 6216 242
rect 6534 516 6664 555
rect 6534 460 6571 516
rect 6627 460 6664 516
rect 6534 298 6664 460
rect 6534 242 6571 298
rect 6627 242 6664 298
rect 6534 204 6664 242
rect 7038 510 7218 520
rect 7038 246 7048 510
rect 7208 246 7218 510
rect 7038 236 7218 246
rect 4725 161 4855 201
rect 4057 117 4185 161
rect 4726 117 4854 161
rect 366 -97 1664 -94
rect 366 -149 378 -97
rect 534 -149 1664 -97
rect 366 -150 1664 -149
rect 366 -161 546 -150
<< via2 >>
rect 172 3543 228 3545
rect 172 3283 174 3543
rect 174 3283 226 3543
rect 226 3283 228 3543
rect 172 3281 228 3283
rect 620 3543 676 3545
rect 620 3283 622 3543
rect 622 3283 674 3543
rect 674 3283 676 3543
rect 620 3281 676 3283
rect 1943 3543 1999 3545
rect 1943 3283 1945 3543
rect 1945 3283 1997 3543
rect 1997 3283 1999 3543
rect 1943 3281 1999 3283
rect 2391 3543 2447 3545
rect 2391 3283 2393 3543
rect 2393 3283 2445 3543
rect 2445 3283 2447 3543
rect 2391 3281 2447 3283
rect 2839 3543 2895 3545
rect 2839 3283 2841 3543
rect 2841 3283 2893 3543
rect 2893 3283 2895 3543
rect 2839 3281 2895 3283
rect 3287 3543 3343 3545
rect 3287 3283 3289 3543
rect 3289 3283 3341 3543
rect 3341 3283 3343 3543
rect 3287 3281 3343 3283
rect 3735 3543 3791 3545
rect 3735 3283 3737 3543
rect 3737 3283 3789 3543
rect 3789 3283 3791 3543
rect 3735 3281 3791 3283
rect 4183 3543 4239 3545
rect 4183 3283 4185 3543
rect 4185 3283 4237 3543
rect 4237 3283 4239 3543
rect 4183 3281 4239 3283
rect 4386 3543 4442 3545
rect 4386 3283 4388 3543
rect 4388 3283 4440 3543
rect 4440 3283 4442 3543
rect 4386 3281 4442 3283
rect 4589 3543 4645 3545
rect 4589 3283 4591 3543
rect 4591 3283 4643 3543
rect 4643 3283 4645 3543
rect 4589 3281 4645 3283
rect 5037 3543 5093 3545
rect 5037 3283 5039 3543
rect 5039 3283 5091 3543
rect 5091 3283 5093 3543
rect 5037 3281 5093 3283
rect 5485 3543 5541 3545
rect 5485 3283 5487 3543
rect 5487 3283 5539 3543
rect 5539 3283 5541 3543
rect 5485 3281 5541 3283
rect 5933 3543 5989 3545
rect 5933 3283 5935 3543
rect 5935 3283 5987 3543
rect 5987 3283 5989 3543
rect 5933 3281 5989 3283
rect 6381 3543 6437 3545
rect 6381 3283 6383 3543
rect 6383 3283 6435 3543
rect 6435 3283 6437 3543
rect 6381 3281 6437 3283
rect 6829 3543 6885 3545
rect 6829 3283 6831 3543
rect 6831 3283 6883 3543
rect 6883 3283 6885 3543
rect 6829 3281 6885 3283
rect 7048 3543 7208 3545
rect 7048 3283 7050 3543
rect 7050 3283 7206 3543
rect 7206 3283 7208 3543
rect 7048 3281 7208 3283
rect 2013 3040 2381 3042
rect 2013 2988 2015 3040
rect 2015 2988 2379 3040
rect 2379 2988 2381 3040
rect 2013 2986 2381 2988
rect 172 2267 228 2269
rect 172 2007 174 2267
rect 174 2007 226 2267
rect 226 2007 228 2267
rect 172 2005 228 2007
rect 620 2267 676 2269
rect 620 2007 622 2267
rect 622 2007 674 2267
rect 674 2007 676 2267
rect 620 2005 676 2007
rect 1068 2267 1124 2269
rect 1068 2007 1070 2267
rect 1070 2007 1122 2267
rect 1122 2007 1124 2267
rect 1068 2005 1124 2007
rect 1516 2267 1572 2269
rect 1516 2007 1518 2267
rect 1518 2007 1570 2267
rect 1570 2007 1572 2267
rect 1516 2005 1572 2007
rect 1720 2267 1776 2269
rect 1720 2007 1722 2267
rect 1722 2007 1774 2267
rect 1774 2007 1776 2267
rect 1720 2005 1776 2007
rect 1943 2267 1999 2269
rect 1943 2007 1945 2267
rect 1945 2007 1997 2267
rect 1997 2007 1999 2267
rect 1943 2005 1999 2007
rect 2391 2267 2447 2269
rect 2391 2007 2393 2267
rect 2393 2007 2445 2267
rect 2445 2007 2447 2267
rect 2391 2005 2447 2007
rect 2839 2267 2895 2269
rect 2839 2007 2841 2267
rect 2841 2007 2893 2267
rect 2893 2007 2895 2267
rect 2839 2005 2895 2007
rect 3287 2267 3343 2269
rect 3287 2007 3289 2267
rect 3289 2007 3341 2267
rect 3341 2007 3343 2267
rect 3287 2005 3343 2007
rect 3735 2267 3791 2269
rect 3735 2007 3737 2267
rect 3737 2007 3789 2267
rect 3789 2007 3791 2267
rect 3735 2005 3791 2007
rect 4183 2267 4239 2269
rect 4183 2007 4185 2267
rect 4185 2007 4237 2267
rect 4237 2007 4239 2267
rect 4183 2005 4239 2007
rect 4386 2267 4442 2269
rect 4386 2007 4388 2267
rect 4388 2007 4440 2267
rect 4440 2007 4442 2267
rect 4386 2005 4442 2007
rect 4589 2267 4645 2269
rect 4589 2007 4591 2267
rect 4591 2007 4643 2267
rect 4643 2007 4645 2267
rect 4589 2005 4645 2007
rect 5037 2267 5093 2269
rect 5037 2007 5039 2267
rect 5039 2007 5091 2267
rect 5091 2007 5093 2267
rect 5037 2005 5093 2007
rect 5485 2267 5541 2269
rect 5485 2007 5487 2267
rect 5487 2007 5539 2267
rect 5539 2007 5541 2267
rect 5485 2005 5541 2007
rect 5933 2267 5989 2269
rect 5933 2007 5935 2267
rect 5935 2007 5987 2267
rect 5987 2007 5989 2267
rect 5933 2005 5989 2007
rect 6381 2267 6437 2269
rect 6381 2007 6383 2267
rect 6383 2007 6435 2267
rect 6435 2007 6437 2267
rect 6381 2005 6437 2007
rect 6829 2267 6885 2269
rect 6829 2007 6831 2267
rect 6831 2007 6883 2267
rect 6883 2007 6885 2267
rect 6829 2005 6885 2007
rect 7042 2267 7202 2269
rect 7042 2007 7044 2267
rect 7044 2007 7200 2267
rect 7200 2007 7202 2267
rect 7042 2005 7202 2007
rect 1272 1476 1432 1478
rect 1272 1424 1274 1476
rect 1274 1424 1430 1476
rect 1430 1424 1432 1476
rect 1272 1422 1432 1424
rect 4600 1476 4760 1478
rect 4600 1424 4602 1476
rect 4602 1424 4758 1476
rect 4758 1424 4760 1476
rect 4600 1422 4760 1424
rect 128 1216 184 1218
rect 128 1164 130 1216
rect 130 1164 182 1216
rect 182 1164 184 1216
rect 128 1162 184 1164
rect 128 998 184 1000
rect 128 946 130 998
rect 130 946 182 998
rect 182 946 184 998
rect 128 944 184 946
rect 653 1205 709 1207
rect 653 1153 655 1205
rect 655 1153 707 1205
rect 707 1153 709 1205
rect 653 1151 709 1153
rect 653 987 709 989
rect 653 935 655 987
rect 655 935 707 987
rect 707 935 709 987
rect 653 933 709 935
rect 1101 1205 1157 1207
rect 1101 1153 1103 1205
rect 1103 1153 1155 1205
rect 1155 1153 1157 1205
rect 1101 1151 1157 1153
rect 1101 987 1157 989
rect 1101 935 1103 987
rect 1103 935 1155 987
rect 1155 935 1157 987
rect 1101 933 1157 935
rect 2517 1205 2573 1207
rect 2517 1153 2519 1205
rect 2519 1153 2571 1205
rect 2571 1153 2573 1205
rect 2517 1151 2573 1153
rect 2517 987 2573 989
rect 2517 935 2519 987
rect 2519 935 2571 987
rect 2571 935 2573 987
rect 2517 933 2573 935
rect 2965 1205 3021 1207
rect 2965 1153 2967 1205
rect 2967 1153 3019 1205
rect 3019 1153 3021 1205
rect 2965 1151 3021 1153
rect 2965 987 3021 989
rect 2965 935 2967 987
rect 2967 935 3019 987
rect 3019 935 3021 987
rect 2965 933 3021 935
rect 3213 1219 3269 1221
rect 3213 959 3215 1219
rect 3215 959 3267 1219
rect 3267 959 3269 1219
rect 3213 957 3269 959
rect 3661 1219 3717 1221
rect 3661 959 3663 1219
rect 3663 959 3715 1219
rect 3715 959 3717 1219
rect 3661 957 3717 959
rect 4986 1205 5042 1207
rect 4986 1153 4988 1205
rect 4988 1153 5040 1205
rect 5040 1153 5042 1205
rect 4986 1151 5042 1153
rect 4986 987 5042 989
rect 4986 935 4988 987
rect 4988 935 5040 987
rect 5040 935 5042 987
rect 4986 933 5042 935
rect 5227 1214 5283 1216
rect 5227 1162 5229 1214
rect 5229 1162 5281 1214
rect 5281 1162 5283 1214
rect 5227 1160 5283 1162
rect 5227 996 5283 998
rect 5227 944 5229 996
rect 5229 944 5281 996
rect 5281 944 5283 996
rect 5227 942 5283 944
rect 5675 1214 5731 1216
rect 5675 1162 5677 1214
rect 5677 1162 5729 1214
rect 5729 1162 5731 1214
rect 5675 1160 5731 1162
rect 5675 996 5731 998
rect 5675 944 5677 996
rect 5677 944 5729 996
rect 5729 944 5731 996
rect 5675 942 5731 944
rect 6123 1214 6179 1216
rect 6123 1162 6125 1214
rect 6125 1162 6177 1214
rect 6177 1162 6179 1214
rect 6123 1160 6179 1162
rect 6123 996 6179 998
rect 6123 944 6125 996
rect 6125 944 6177 996
rect 6177 944 6179 996
rect 6123 942 6179 944
rect 6571 1214 6627 1216
rect 6571 1162 6573 1214
rect 6573 1162 6625 1214
rect 6625 1162 6627 1214
rect 6571 1160 6627 1162
rect 6571 996 6627 998
rect 6571 944 6573 996
rect 6573 944 6625 996
rect 6625 944 6627 996
rect 6571 942 6627 944
rect 7096 1216 7152 1218
rect 7096 1164 7098 1216
rect 7098 1164 7150 1216
rect 7150 1164 7152 1216
rect 7096 1162 7152 1164
rect 7096 998 7152 1000
rect 7096 946 7098 998
rect 7098 946 7150 998
rect 7150 946 7152 998
rect 7096 944 7152 946
rect 128 514 184 516
rect 128 462 130 514
rect 130 462 182 514
rect 182 462 184 514
rect 128 460 184 462
rect 128 296 184 298
rect 128 244 130 296
rect 130 244 182 296
rect 182 244 184 296
rect 128 242 184 244
rect 653 514 709 516
rect 653 462 655 514
rect 655 462 707 514
rect 707 462 709 514
rect 653 460 709 462
rect 653 296 709 298
rect 653 244 655 296
rect 655 244 707 296
rect 707 244 709 296
rect 653 242 709 244
rect 1101 513 1157 515
rect 1101 461 1103 513
rect 1103 461 1155 513
rect 1155 461 1157 513
rect 1101 459 1157 461
rect 1101 327 1157 329
rect 1101 275 1103 327
rect 1103 275 1155 327
rect 1155 275 1157 327
rect 1101 273 1157 275
rect 2517 513 2573 515
rect 2517 461 2519 513
rect 2519 461 2571 513
rect 2571 461 2573 513
rect 2517 459 2573 461
rect 2517 327 2573 329
rect 2517 275 2519 327
rect 2519 275 2571 327
rect 2571 275 2573 327
rect 2517 273 2573 275
rect 2965 513 3021 515
rect 2965 461 2967 513
rect 2967 461 3019 513
rect 3019 461 3021 513
rect 2965 459 3021 461
rect 2965 327 3021 329
rect 2965 275 2967 327
rect 2967 275 3019 327
rect 3019 275 3021 327
rect 2965 273 3021 275
rect 3213 490 3269 492
rect 3213 230 3215 490
rect 3215 230 3267 490
rect 3267 230 3269 490
rect 3213 228 3269 230
rect 3661 490 3717 492
rect 3661 230 3663 490
rect 3663 230 3715 490
rect 3715 230 3717 490
rect 3661 228 3717 230
rect 668 55 724 56
rect 668 3 670 55
rect 670 3 722 55
rect 722 3 724 55
rect 668 0 724 3
rect 880 55 936 56
rect 880 3 882 55
rect 882 3 934 55
rect 934 3 936 55
rect 880 0 936 3
rect 4986 513 5042 515
rect 4986 461 4988 513
rect 4988 461 5040 513
rect 5040 461 5042 513
rect 4986 459 5042 461
rect 4986 327 5042 329
rect 4986 275 4988 327
rect 4988 275 5040 327
rect 5040 275 5042 327
rect 4986 273 5042 275
rect 5227 514 5283 516
rect 5227 462 5229 514
rect 5229 462 5281 514
rect 5281 462 5283 514
rect 5227 460 5283 462
rect 5227 296 5283 298
rect 5227 244 5229 296
rect 5229 244 5281 296
rect 5281 244 5283 296
rect 5227 242 5283 244
rect 5675 514 5731 516
rect 5675 462 5677 514
rect 5677 462 5729 514
rect 5729 462 5731 514
rect 5675 460 5731 462
rect 5675 296 5731 298
rect 5675 244 5677 296
rect 5677 244 5729 296
rect 5729 244 5731 296
rect 5675 242 5731 244
rect 6123 514 6179 516
rect 6123 462 6125 514
rect 6125 462 6177 514
rect 6177 462 6179 514
rect 6123 460 6179 462
rect 6123 296 6179 298
rect 6123 244 6125 296
rect 6125 244 6177 296
rect 6177 244 6179 296
rect 6123 242 6179 244
rect 6571 514 6627 516
rect 6571 462 6573 514
rect 6573 462 6625 514
rect 6625 462 6627 514
rect 6571 460 6627 462
rect 6571 296 6627 298
rect 6571 244 6573 296
rect 6573 244 6625 296
rect 6625 244 6627 296
rect 6571 242 6627 244
rect 7048 508 7208 510
rect 7048 248 7050 508
rect 7050 248 7206 508
rect 7206 248 7208 508
rect 7048 246 7208 248
<< metal3 >>
rect 91 3545 7407 3555
rect 91 3281 172 3545
rect 228 3281 620 3545
rect 676 3281 1943 3545
rect 1999 3281 2391 3545
rect 2447 3281 2839 3545
rect 2895 3281 3287 3545
rect 3343 3281 3735 3545
rect 3791 3281 4183 3545
rect 4239 3281 4386 3545
rect 4442 3281 4589 3545
rect 4645 3281 5037 3545
rect 5093 3281 5485 3545
rect 5541 3281 5933 3545
rect 5989 3281 6381 3545
rect 6437 3281 6829 3545
rect 6885 3281 7048 3545
rect 7208 3281 7407 3545
rect 91 3271 7407 3281
rect 2003 3042 2391 3057
rect 2003 2986 2013 3042
rect 2381 2986 2391 3042
rect 2003 2969 2391 2986
rect 91 2269 7407 2279
rect 91 2005 172 2269
rect 228 2005 620 2269
rect 676 2005 1068 2269
rect 1124 2005 1516 2269
rect 1572 2005 1720 2269
rect 1776 2005 1943 2269
rect 1999 2005 2391 2269
rect 2447 2005 2839 2269
rect 2895 2005 3287 2269
rect 3343 2005 3735 2269
rect 3791 2005 4183 2269
rect 4239 2005 4386 2269
rect 4442 2005 4589 2269
rect 4645 2005 5037 2269
rect 5093 2005 5485 2269
rect 5541 2005 5933 2269
rect 5989 2005 6381 2269
rect 6437 2005 6829 2269
rect 6885 2005 7042 2269
rect 7202 2005 7407 2269
rect 91 1995 7407 2005
rect 1262 1478 4770 1494
rect 1262 1422 1272 1478
rect 1432 1422 4600 1478
rect 4760 1422 4770 1478
rect 1262 1406 4770 1422
rect 91 1221 7407 1298
rect 91 1218 3213 1221
rect 91 1162 128 1218
rect 184 1207 3213 1218
rect 184 1162 653 1207
rect 91 1151 653 1162
rect 709 1151 1101 1207
rect 1157 1151 2517 1207
rect 2573 1151 2965 1207
rect 3021 1151 3213 1207
rect 91 1000 3213 1151
rect 91 944 128 1000
rect 184 989 3213 1000
rect 184 944 653 989
rect 91 933 653 944
rect 709 933 1101 989
rect 1157 933 2517 989
rect 2573 933 2965 989
rect 3021 957 3213 989
rect 3269 957 3661 1221
rect 3717 1218 7407 1221
rect 3717 1216 7096 1218
rect 3717 1207 5227 1216
rect 3717 1151 4986 1207
rect 5042 1160 5227 1207
rect 5283 1160 5675 1216
rect 5731 1160 6123 1216
rect 6179 1160 6571 1216
rect 6627 1162 7096 1216
rect 7152 1162 7407 1218
rect 6627 1160 7407 1162
rect 5042 1151 7407 1160
rect 3717 1000 7407 1151
rect 3717 998 7096 1000
rect 3717 989 5227 998
rect 3717 957 4986 989
rect 3021 933 4986 957
rect 5042 942 5227 989
rect 5283 942 5675 998
rect 5731 942 6123 998
rect 6179 942 6571 998
rect 6627 944 7096 998
rect 7152 944 7407 1000
rect 6627 942 7407 944
rect 5042 933 7407 942
rect 91 843 7407 933
rect 91 554 221 555
rect 616 554 746 555
rect 5190 554 5320 555
rect 5638 554 5768 555
rect 6086 554 6216 555
rect 6534 554 6664 555
rect 91 516 7407 554
rect 91 460 128 516
rect 184 460 653 516
rect 709 515 5227 516
rect 709 460 1101 515
rect 91 459 1101 460
rect 1157 459 2517 515
rect 2573 459 2965 515
rect 3021 492 4986 515
rect 3021 459 3213 492
rect 91 329 3213 459
rect 91 298 1101 329
rect 91 242 128 298
rect 184 242 653 298
rect 709 273 1101 298
rect 1157 273 2517 329
rect 2573 273 2965 329
rect 3021 273 3213 329
rect 709 242 3213 273
rect 91 228 3213 242
rect 3269 228 3661 492
rect 3717 459 4986 492
rect 5042 460 5227 515
rect 5283 460 5675 516
rect 5731 460 6123 516
rect 6179 460 6571 516
rect 6627 510 7407 516
rect 6627 460 7048 510
rect 5042 459 7048 460
rect 3717 329 7048 459
rect 3717 273 4986 329
rect 5042 298 7048 329
rect 5042 273 5227 298
rect 3717 242 5227 273
rect 5283 242 5675 298
rect 5731 242 6123 298
rect 6179 242 6571 298
rect 6627 246 7048 298
rect 7208 246 7407 510
rect 6627 242 7407 246
rect 3717 228 7407 242
rect 91 203 7407 228
rect 632 56 972 95
rect 632 0 668 56
rect 724 0 880 56
rect 936 0 972 56
rect 632 -38 972 0
use M1_NACTIVE$$202392620_256x8m81  M1_NACTIVE$$202392620_256x8m81_0
timestamp 1669390400
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M1_NACTIVE$$202392620_256x8m81  M1_NACTIVE$$202392620_256x8m81_1
timestamp 1669390400
transform 1 0 156 0 1 379
box 0 0 1 1
use M1_NACTIVE$$202392620_256x8m81  M1_NACTIVE$$202392620_256x8m81_2
timestamp 1669390400
transform 1 0 156 0 1 1081
box 0 0 1 1
use M1_NACTIVE4310590878124_256x8m81  M1_NACTIVE4310590878124_256x8m81_0
timestamp 1669390400
transform 1 0 1748 0 1 2132
box 0 0 1 1
use M1_NACTIVE4310590878124_256x8m81  M1_NACTIVE4310590878124_256x8m81_1
timestamp 1669390400
transform 1 0 4414 0 1 2132
box 0 0 1 1
use M1_NACTIVE4310590878164_256x8m81  M1_NACTIVE4310590878164_256x8m81_0
timestamp 1669390400
transform 1 0 7121 0 1 2132
box 0 0 1 1
use M1_PACTIVE4310590878136_256x8m81  M1_PACTIVE4310590878136_256x8m81_0
timestamp 1669390400
transform 1 0 4414 0 1 3408
box 0 0 1 1
use M1_PACTIVE4310590878163_256x8m81  M1_PACTIVE4310590878163_256x8m81_0
timestamp 1669390400
transform 1 0 7121 0 1 373
box 0 0 1 1
use M1_PACTIVE4310590878163_256x8m81  M1_PACTIVE4310590878163_256x8m81_1
timestamp 1669390400
transform 1 0 7121 0 1 3408
box 0 0 1 1
use M1_PACTIVE4310590878165_256x8m81  M1_PACTIVE4310590878165_256x8m81_0
timestamp 1669390400
transform 1 0 1427 0 1 3408
box -183 -136 183 136
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1669390400
transform 1 0 4678 0 1 1446
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_1
timestamp 1669390400
transform 1 0 5919 0 1 1656
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_2
timestamp 1669390400
transform 1 0 6373 0 1 1656
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_3
timestamp 1669390400
transform 1 0 6716 0 1 1656
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_4
timestamp 1669390400
transform 1 0 4039 0 1 -41
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_5
timestamp 1669390400
transform 1 0 4337 0 1 1407
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_6
timestamp 1669390400
transform 1 0 5243 0 1 709
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_7
timestamp 1669390400
transform 1 0 5477 0 1 1656
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_8
timestamp 1669390400
transform 1 0 4649 0 1 41
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_9
timestamp 1669390400
transform 1 0 1100 0 1 635
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_10
timestamp 1669390400
transform 1 0 2579 0 1 711
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_11
timestamp 1669390400
transform 1 0 2528 0 1 47
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_12
timestamp 1669390400
transform 1 0 3382 0 1 47
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_13
timestamp 1669390400
transform 1 0 1777 0 1 -224
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_14
timestamp 1669390400
transform 1 0 540 0 1 1663
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_15
timestamp 1669390400
transform 1 0 540 0 1 1406
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_16
timestamp 1669390400
transform 0 -1 1406 1 0 694
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_17
timestamp 1669390400
transform 1 0 822 0 1 61
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_18
timestamp 1669390400
transform 1 0 1696 0 1 2847
box 0 0 1 1
use M2_M1$$201262124_256x8m81  M2_M1$$201262124_256x8m81_0
timestamp 1669390400
transform 1 0 802 0 1 29
box 0 0 1 1
use M2_M1$$202395692_256x8m81  M2_M1$$202395692_256x8m81_0
timestamp 1669390400
transform 1 0 5014 0 1 394
box 0 0 1 1
use M2_M1$$202395692_256x8m81  M2_M1$$202395692_256x8m81_1
timestamp 1669390400
transform 1 0 2545 0 1 394
box 0 0 1 1
use M2_M1$$202395692_256x8m81  M2_M1$$202395692_256x8m81_2
timestamp 1669390400
transform 1 0 2993 0 1 394
box 0 0 1 1
use M2_M1$$202395692_256x8m81  M2_M1$$202395692_256x8m81_3
timestamp 1669390400
transform 1 0 1129 0 1 394
box 0 0 1 1
use M2_M1$$202396716_256x8m81  M2_M1$$202396716_256x8m81_0
timestamp 1669390400
transform 1 0 1636 0 1 703
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_0
timestamp 1669390400
transform 1 0 5703 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_1
timestamp 1669390400
transform 1 0 6151 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_2
timestamp 1669390400
transform 1 0 6599 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_3
timestamp 1669390400
transform 1 0 5255 0 -1 1079
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_4
timestamp 1669390400
transform 1 0 4121 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_5
timestamp 1669390400
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_6
timestamp 1669390400
transform 1 0 6599 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_7
timestamp 1669390400
transform 1 0 6151 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_8
timestamp 1669390400
transform 1 0 5703 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_9
timestamp 1669390400
transform 1 0 5255 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_10
timestamp 1669390400
transform 1 0 5014 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_11
timestamp 1669390400
transform 1 0 4790 0 1 336
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_12
timestamp 1669390400
transform 1 0 4790 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_13
timestamp 1669390400
transform 1 0 4121 0 1 336
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_14
timestamp 1669390400
transform 1 0 2545 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_15
timestamp 1669390400
transform 1 0 2993 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_16
timestamp 1669390400
transform 1 0 156 0 1 1081
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_17
timestamp 1669390400
transform 1 0 156 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_18
timestamp 1669390400
transform 1 0 681 0 1 1070
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_19
timestamp 1669390400
transform 1 0 681 0 1 379
box 0 0 1 1
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_20
timestamp 1669390400
transform 1 0 1129 0 1 1070
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_0
timestamp 1669390400
transform 1 0 3689 0 1 1089
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_1
timestamp 1669390400
transform 1 0 3689 0 1 360
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_2
timestamp 1669390400
transform 1 0 3241 0 1 360
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_3
timestamp 1669390400
transform 1 0 3241 0 1 1089
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_4
timestamp 1669390400
transform 1 0 2867 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_5
timestamp 1669390400
transform 1 0 2419 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_6
timestamp 1669390400
transform 1 0 1971 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_7
timestamp 1669390400
transform 1 0 3315 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_8
timestamp 1669390400
transform 1 0 1971 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_9
timestamp 1669390400
transform 1 0 2419 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_10
timestamp 1669390400
transform 1 0 2867 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_11
timestamp 1669390400
transform 1 0 3315 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_12
timestamp 1669390400
transform 1 0 1748 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_13
timestamp 1669390400
transform 1 0 200 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_14
timestamp 1669390400
transform 1 0 648 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_15
timestamp 1669390400
transform 1 0 648 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_16
timestamp 1669390400
transform 1 0 200 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_17
timestamp 1669390400
transform 1 0 1544 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_18
timestamp 1669390400
transform 1 0 1096 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_19
timestamp 1669390400
transform 1 0 6857 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_20
timestamp 1669390400
transform 1 0 6409 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_21
timestamp 1669390400
transform 1 0 4414 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_22
timestamp 1669390400
transform 1 0 4414 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_23
timestamp 1669390400
transform 1 0 4211 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_24
timestamp 1669390400
transform 1 0 3763 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_25
timestamp 1669390400
transform 1 0 4211 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_26
timestamp 1669390400
transform 1 0 3763 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_27
timestamp 1669390400
transform 1 0 5513 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_28
timestamp 1669390400
transform 1 0 5065 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_29
timestamp 1669390400
transform 1 0 4617 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_30
timestamp 1669390400
transform 1 0 5961 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_31
timestamp 1669390400
transform 1 0 6857 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_32
timestamp 1669390400
transform 1 0 6409 0 1 2137
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_33
timestamp 1669390400
transform 1 0 4617 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_34
timestamp 1669390400
transform 1 0 5065 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_35
timestamp 1669390400
transform 1 0 5513 0 1 3413
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_36
timestamp 1669390400
transform 1 0 5961 0 1 3413
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_0
timestamp 1669390400
transform 0 -1 4680 1 0 1450
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_1
timestamp 1669390400
transform 0 -1 456 1 0 -123
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_2
timestamp 1669390400
transform 0 -1 1352 1 0 1450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_0
timestamp 1669390400
transform 0 -1 2197 1 0 3014
box 0 0 1 1
use M2_M14310590878167_256x8m81  M2_M14310590878167_256x8m81_0
timestamp 1669390400
transform 1 0 7128 0 1 378
box 0 0 1 1
use M2_M14310590878167_256x8m81  M2_M14310590878167_256x8m81_1
timestamp 1669390400
transform 1 0 7128 0 1 3413
box 0 0 1 1
use M2_M14310590878167_256x8m81  M2_M14310590878167_256x8m81_2
timestamp 1669390400
transform 1 0 7122 0 1 2137
box 0 0 1 1
use M2_M14310590878168_256x8m81  M2_M14310590878168_256x8m81_0
timestamp 1669390400
transform 1 0 1433 0 1 3413
box -142 -142 142 142
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_0
timestamp 1669390400
transform 1 0 6599 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_1
timestamp 1669390400
transform 1 0 6151 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_2
timestamp 1669390400
transform 1 0 5255 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_3
timestamp 1669390400
transform 1 0 6599 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_4
timestamp 1669390400
transform 1 0 7124 0 1 1081
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_5
timestamp 1669390400
transform 1 0 5255 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_6
timestamp 1669390400
transform 1 0 5703 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_7
timestamp 1669390400
transform 1 0 6151 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_8
timestamp 1669390400
transform 1 0 5014 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_9
timestamp 1669390400
transform 1 0 5703 0 -1 1079
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_10
timestamp 1669390400
transform 1 0 2545 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_11
timestamp 1669390400
transform 1 0 2993 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_12
timestamp 1669390400
transform 1 0 156 0 1 1081
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_13
timestamp 1669390400
transform 1 0 156 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_14
timestamp 1669390400
transform 1 0 681 0 1 1070
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_15
timestamp 1669390400
transform 1 0 681 0 1 379
box 0 0 1 1
use M3_M2$$201252908_256x8m81  M3_M2$$201252908_256x8m81_16
timestamp 1669390400
transform 1 0 1129 0 1 1070
box 0 0 1 1
use M3_M2$$201255980_256x8m81  M3_M2$$201255980_256x8m81_0
timestamp 1669390400
transform 1 0 802 0 1 28
box 0 0 1 1
use M3_M2$$202397740_256x8m81  M3_M2$$202397740_256x8m81_0
timestamp 1669390400
transform 1 0 5014 0 1 394
box 0 0 1 1
use M3_M2$$202397740_256x8m81  M3_M2$$202397740_256x8m81_1
timestamp 1669390400
transform 1 0 2545 0 1 394
box 0 0 1 1
use M3_M2$$202397740_256x8m81  M3_M2$$202397740_256x8m81_2
timestamp 1669390400
transform 1 0 2993 0 1 394
box 0 0 1 1
use M3_M2$$202397740_256x8m81  M3_M2$$202397740_256x8m81_3
timestamp 1669390400
transform 1 0 1129 0 1 394
box 0 0 1 1
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_0
timestamp 1669390400
transform 1 0 4680 0 1 1450
box 0 0 1 1
use M3_M2431059087814_256x8m81  M3_M2431059087814_256x8m81_1
timestamp 1669390400
transform 1 0 1352 0 1 1450
box 0 0 1 1
use M3_M24310590878122_256x8m81  M3_M24310590878122_256x8m81_0
timestamp 1669390400
transform 0 -1 2197 1 0 3014
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_0
timestamp 1669390400
transform 1 0 3689 0 1 1089
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_1
timestamp 1669390400
transform 1 0 3689 0 1 360
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_2
timestamp 1669390400
transform 1 0 3241 0 1 1089
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_3
timestamp 1669390400
transform 1 0 3241 0 1 360
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_4
timestamp 1669390400
transform 1 0 1544 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_5
timestamp 1669390400
transform 1 0 1096 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_6
timestamp 1669390400
transform 1 0 1748 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_7
timestamp 1669390400
transform 1 0 648 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_8
timestamp 1669390400
transform 1 0 1971 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_9
timestamp 1669390400
transform 1 0 2419 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_10
timestamp 1669390400
transform 1 0 2867 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_11
timestamp 1669390400
transform 1 0 3315 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_12
timestamp 1669390400
transform 1 0 200 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_13
timestamp 1669390400
transform 1 0 200 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_14
timestamp 1669390400
transform 1 0 648 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_15
timestamp 1669390400
transform 1 0 1971 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_16
timestamp 1669390400
transform 1 0 2419 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_17
timestamp 1669390400
transform 1 0 2867 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_18
timestamp 1669390400
transform 1 0 3315 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_19
timestamp 1669390400
transform 1 0 4211 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_20
timestamp 1669390400
transform 1 0 3763 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_21
timestamp 1669390400
transform 1 0 4617 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_22
timestamp 1669390400
transform 1 0 5065 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_23
timestamp 1669390400
transform 1 0 5513 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_24
timestamp 1669390400
transform 1 0 5961 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_25
timestamp 1669390400
transform 1 0 6857 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_26
timestamp 1669390400
transform 1 0 6409 0 1 3413
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_27
timestamp 1669390400
transform 1 0 4211 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_28
timestamp 1669390400
transform 1 0 3763 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_29
timestamp 1669390400
transform 1 0 4617 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_30
timestamp 1669390400
transform 1 0 5065 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_31
timestamp 1669390400
transform 1 0 5513 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_32
timestamp 1669390400
transform 1 0 5961 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_33
timestamp 1669390400
transform 1 0 6857 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_34
timestamp 1669390400
transform 1 0 6409 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_35
timestamp 1669390400
transform 1 0 4414 0 1 2137
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_36
timestamp 1669390400
transform 1 0 4414 0 1 3413
box 0 0 1 1
use M3_M24310590878144_256x8m81  M3_M24310590878144_256x8m81_0
timestamp 1669390400
transform 1 0 1433 0 1 3413
box -142 -142 142 142
use M3_M24310590878166_256x8m81  M3_M24310590878166_256x8m81_0
timestamp 1669390400
transform 1 0 7128 0 1 378
box 0 0 1 1
use M3_M24310590878166_256x8m81  M3_M24310590878166_256x8m81_1
timestamp 1669390400
transform 1 0 7128 0 1 3413
box 0 0 1 1
use M3_M24310590878166_256x8m81  M3_M24310590878166_256x8m81_2
timestamp 1669390400
transform 1 0 7122 0 1 2137
box 0 0 1 1
use nmos_1p2$$202595372_256x8m81  nmos_1p2$$202595372_256x8m81_0
timestamp 1669390400
transform 1 0 2853 0 1 372
box -119 -73 177 264
use nmos_1p2$$202595372_256x8m81  nmos_1p2$$202595372_256x8m81_1
timestamp 1669390400
transform 1 0 2181 0 1 372
box -119 -73 177 264
use nmos_1p2$$202596396_256x8m81  nmos_1p2$$202596396_256x8m81_0
timestamp 1669390400
transform 1 0 2405 0 1 372
box -119 -73 177 264
use nmos_5p0431059087818_256x8m81  nmos_5p0431059087818_256x8m81_0
timestamp 1669390400
transform 1 0 4842 0 -1 440
box -88 -44 208 236
use nmos_5p0431059087818_256x8m81  nmos_5p0431059087818_256x8m81_1
timestamp 1669390400
transform 1 0 4618 0 -1 440
box -88 -44 208 236
use nmos_5p0431059087818_256x8m81  nmos_5p0431059087818_256x8m81_2
timestamp 1669390400
transform 1 0 509 0 1 213
box -88 -44 208 236
use nmos_5p0431059087818_256x8m81  nmos_5p0431059087818_256x8m81_3
timestamp 1669390400
transform 1 0 733 0 1 213
box -88 -44 208 236
use nmos_5p0431059087818_256x8m81  nmos_5p0431059087818_256x8m81_4
timestamp 1669390400
transform 1 0 1181 0 1 295
box -88 -44 208 236
use nmos_5p04310590878110_256x8m81  nmos_5p04310590878110_256x8m81_0
timestamp 1669390400
transform 1 0 1688 0 1 109
box -88 -44 208 498
use nmos_5p04310590878139_256x8m81  nmos_5p04310590878139_256x8m81_0
timestamp 1669390400
transform 1 0 3950 0 1 109
box -88 -44 432 498
use nmos_5p04310590878179_256x8m81  nmos_5p04310590878179_256x8m81_0
timestamp 1669390400
transform 1 0 4669 0 1 3214
box -88 -44 2224 428
use nmos_5p04310590878179_256x8m81  nmos_5p04310590878179_256x8m81_1
timestamp 1669390400
transform 1 0 2023 0 1 3214
box -88 -44 2224 428
use nmos_5p04310590878180_256x8m81  nmos_5p04310590878180_256x8m81_0
timestamp 1669390400
transform 1 0 3293 0 1 324
box -88 -44 432 284
use nmos_5p04310590878182_256x8m81  nmos_5p04310590878182_256x8m81_0
timestamp 1669390400
transform 1 0 252 0 1 3214
box -88 -44 656 444
use nmos_5p04310590878185_256x8m81  nmos_5p04310590878185_256x8m81_0
timestamp 1669390400
transform 1 0 5307 0 1 381
box -88 -44 1552 222
use pmos_1p2$$202586156_256x8m81  pmos_1p2$$202586156_256x8m81_0
timestamp 1669390400
transform 1 0 2405 0 1 843
box -286 -141 344 595
use pmos_1p2$$202587180_256x8m81  pmos_1p2$$202587180_256x8m81_0
timestamp 1669390400
transform 1 0 1719 0 1 843
box -286 -141 344 595
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_0
timestamp 1669390400
transform 1 0 4842 0 -1 1297
box -208 -120 328 574
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_1
timestamp 1669390400
transform 1 0 733 0 1 843
box -208 -120 328 574
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_2
timestamp 1669390400
transform 1 0 2822 0 1 843
box -208 -120 328 574
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_3
timestamp 1669390400
transform 1 0 509 0 1 843
box -208 -120 328 574
use pmos_5p04310590878114_256x8m81  pmos_5p04310590878114_256x8m81_4
timestamp 1669390400
transform 1 0 1181 0 1 843
box -208 -120 328 574
use pmos_5p04310590878120_256x8m81  pmos_5p04310590878120_256x8m81_0
timestamp 1669390400
transform 1 0 3950 0 1 843
box -208 -120 552 574
use pmos_5p04310590878141_256x8m81  pmos_5p04310590878141_256x8m81_0
timestamp 1669390400
transform 1 0 4510 0 -1 1297
box -208 -120 328 312
use pmos_5p04310590878141_256x8m81  pmos_5p04310590878141_256x8m81_1
timestamp 1669390400
transform 1 0 2036 0 1 843
box -208 -120 328 312
use pmos_5p04310590878181_256x8m81  pmos_5p04310590878181_256x8m81_0
timestamp 1669390400
transform 1 0 4669 0 1 1884
box -208 -120 2344 1064
use pmos_5p04310590878181_256x8m81  pmos_5p04310590878181_256x8m81_1
timestamp 1669390400
transform 1 0 2023 0 1 1884
box -208 -120 2344 1064
use pmos_5p04310590878183_256x8m81  pmos_5p04310590878183_256x8m81_0
timestamp 1669390400
transform 1 0 5307 0 1 843
box -208 -120 1672 560
use pmos_5p04310590878184_256x8m81  pmos_5p04310590878184_256x8m81_0
timestamp 1669390400
transform 1 0 3293 0 1 843
box -208 -120 552 688
use pmos_5p04310590878186_256x8m81  pmos_5p04310590878186_256x8m81_0
timestamp 1669390400
transform 1 0 252 0 1 1884
box -208 -120 1448 616
<< labels >>
rlabel metal1 s 481 1428 481 1428 4 wen
port 1 nsew
rlabel metal1 s 6626 3004 6626 3004 4 GWE
port 2 nsew
rlabel metal3 s 252 3479 252 3479 4 vss
port 3 nsew
flabel metal3 s 2212 3015 2212 3015 0 FreeSans 1000 0 0 0 IGWEN
port 4 nsew
rlabel metal3 s 252 2175 252 2175 4 vdd
port 5 nsew
rlabel metal3 s 252 379 252 379 4 vss
port 3 nsew
rlabel metal3 s 252 1070 252 1070 4 vdd
port 5 nsew
rlabel metal3 s 865 61 865 61 4 clk
port 6 nsew
<< properties >>
string GDS_END 1091078
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1068080
string path 23.850 7.250 6.310 7.250 
<< end >>
