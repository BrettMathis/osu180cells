magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -2355 -227 2354 228
<< nsubdiff >>
rect -2212 23 2212 80
rect -2212 -23 -2158 23
rect -2112 -23 -2000 23
rect -1954 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1954 23
rect 2000 -23 2112 23
rect 2158 -23 2212 23
rect -2212 -80 2212 -23
<< nsubdiffcont >>
rect -2158 -23 -2112 23
rect -2000 -23 -1954 23
rect -1841 -23 -1795 23
rect -1683 -23 -1637 23
rect -1525 -23 -1479 23
rect -1367 -23 -1321 23
rect -1209 -23 -1163 23
rect -1051 -23 -1005 23
rect -893 -23 -847 23
rect -735 -23 -689 23
rect -577 -23 -531 23
rect -418 -23 -372 23
rect -260 -23 -214 23
rect -102 -23 -56 23
rect 56 -23 102 23
rect 214 -23 260 23
rect 372 -23 418 23
rect 531 -23 577 23
rect 689 -23 735 23
rect 847 -23 893 23
rect 1005 -23 1051 23
rect 1163 -23 1209 23
rect 1321 -23 1367 23
rect 1479 -23 1525 23
rect 1637 -23 1683 23
rect 1795 -23 1841 23
rect 1954 -23 2000 23
rect 2112 -23 2158 23
<< metal1 >>
rect -2193 23 2192 60
rect -2193 -23 -2158 23
rect -2112 -23 -2000 23
rect -1954 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1954 23
rect 2000 -23 2112 23
rect 2158 -23 2192 23
rect -2193 -60 2192 -23
<< properties >>
string GDS_END 991240
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 989172
<< end >>
