magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 3670 870
<< pwell >>
rect -86 -86 3670 352
<< mvnmos >>
rect 124 68 324 232
rect 572 68 772 232
rect 1020 68 1220 232
rect 1468 68 1668 232
rect 1916 68 2116 232
rect 2364 68 2564 232
rect 2812 68 3012 232
rect 3260 68 3460 232
<< mvpmos >>
rect 124 472 324 716
rect 572 472 772 716
rect 1020 472 1220 716
rect 1468 472 1668 716
rect 1916 472 2116 716
rect 2364 472 2564 716
rect 2812 472 3012 716
rect 3260 472 3460 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 324 192 412 232
rect 324 146 353 192
rect 399 146 412 192
rect 324 68 412 146
rect 484 192 572 232
rect 484 146 497 192
rect 543 146 572 192
rect 484 68 572 146
rect 772 192 860 232
rect 772 146 801 192
rect 847 146 860 192
rect 772 68 860 146
rect 932 192 1020 232
rect 932 146 945 192
rect 991 146 1020 192
rect 932 68 1020 146
rect 1220 192 1308 232
rect 1220 146 1249 192
rect 1295 146 1308 192
rect 1220 68 1308 146
rect 1380 192 1468 232
rect 1380 146 1393 192
rect 1439 146 1468 192
rect 1380 68 1468 146
rect 1668 192 1756 232
rect 1668 146 1697 192
rect 1743 146 1756 192
rect 1668 68 1756 146
rect 1828 192 1916 232
rect 1828 146 1841 192
rect 1887 146 1916 192
rect 1828 68 1916 146
rect 2116 192 2204 232
rect 2116 146 2145 192
rect 2191 146 2204 192
rect 2116 68 2204 146
rect 2276 192 2364 232
rect 2276 146 2289 192
rect 2335 146 2364 192
rect 2276 68 2364 146
rect 2564 192 2652 232
rect 2564 146 2593 192
rect 2639 146 2652 192
rect 2564 68 2652 146
rect 2724 192 2812 232
rect 2724 146 2737 192
rect 2783 146 2812 192
rect 2724 68 2812 146
rect 3012 192 3100 232
rect 3012 146 3041 192
rect 3087 146 3100 192
rect 3012 68 3100 146
rect 3172 192 3260 232
rect 3172 146 3185 192
rect 3231 146 3260 192
rect 3172 68 3260 146
rect 3460 192 3548 232
rect 3460 146 3489 192
rect 3535 146 3548 192
rect 3460 68 3548 146
<< mvpdiff >>
rect 36 657 124 716
rect 36 517 49 657
rect 95 517 124 657
rect 36 472 124 517
rect 324 657 412 716
rect 324 517 353 657
rect 399 517 412 657
rect 324 472 412 517
rect 484 657 572 716
rect 484 517 497 657
rect 543 517 572 657
rect 484 472 572 517
rect 772 657 860 716
rect 772 517 801 657
rect 847 517 860 657
rect 772 472 860 517
rect 932 657 1020 716
rect 932 517 945 657
rect 991 517 1020 657
rect 932 472 1020 517
rect 1220 657 1308 716
rect 1220 517 1249 657
rect 1295 517 1308 657
rect 1220 472 1308 517
rect 1380 657 1468 716
rect 1380 517 1393 657
rect 1439 517 1468 657
rect 1380 472 1468 517
rect 1668 657 1756 716
rect 1668 517 1697 657
rect 1743 517 1756 657
rect 1668 472 1756 517
rect 1828 657 1916 716
rect 1828 517 1841 657
rect 1887 517 1916 657
rect 1828 472 1916 517
rect 2116 657 2204 716
rect 2116 517 2145 657
rect 2191 517 2204 657
rect 2116 472 2204 517
rect 2276 657 2364 716
rect 2276 517 2289 657
rect 2335 517 2364 657
rect 2276 472 2364 517
rect 2564 657 2652 716
rect 2564 517 2593 657
rect 2639 517 2652 657
rect 2564 472 2652 517
rect 2724 657 2812 716
rect 2724 517 2737 657
rect 2783 517 2812 657
rect 2724 472 2812 517
rect 3012 657 3100 716
rect 3012 517 3041 657
rect 3087 517 3100 657
rect 3012 472 3100 517
rect 3172 657 3260 716
rect 3172 517 3185 657
rect 3231 517 3260 657
rect 3172 472 3260 517
rect 3460 657 3548 716
rect 3460 517 3489 657
rect 3535 517 3548 657
rect 3460 472 3548 517
<< mvndiffc >>
rect 49 146 95 192
rect 353 146 399 192
rect 497 146 543 192
rect 801 146 847 192
rect 945 146 991 192
rect 1249 146 1295 192
rect 1393 146 1439 192
rect 1697 146 1743 192
rect 1841 146 1887 192
rect 2145 146 2191 192
rect 2289 146 2335 192
rect 2593 146 2639 192
rect 2737 146 2783 192
rect 3041 146 3087 192
rect 3185 146 3231 192
rect 3489 146 3535 192
<< mvpdiffc >>
rect 49 517 95 657
rect 353 517 399 657
rect 497 517 543 657
rect 801 517 847 657
rect 945 517 991 657
rect 1249 517 1295 657
rect 1393 517 1439 657
rect 1697 517 1743 657
rect 1841 517 1887 657
rect 2145 517 2191 657
rect 2289 517 2335 657
rect 2593 517 2639 657
rect 2737 517 2783 657
rect 3041 517 3087 657
rect 3185 517 3231 657
rect 3489 517 3535 657
<< polysilicon >>
rect 124 716 324 760
rect 572 716 772 760
rect 1020 716 1220 760
rect 1468 716 1668 760
rect 1916 716 2116 760
rect 2364 716 2564 760
rect 2812 716 3012 760
rect 3260 716 3460 760
rect 124 438 324 472
rect 124 392 160 438
rect 300 392 324 438
rect 124 375 324 392
rect 572 438 772 472
rect 572 392 608 438
rect 748 392 772 438
rect 572 375 772 392
rect 1020 438 1220 472
rect 1020 392 1056 438
rect 1196 392 1220 438
rect 1020 375 1220 392
rect 1468 438 1668 472
rect 1468 392 1504 438
rect 1644 392 1668 438
rect 1468 375 1668 392
rect 1916 438 2116 472
rect 1916 392 1952 438
rect 2092 392 2116 438
rect 1916 375 2116 392
rect 2364 438 2564 472
rect 2364 392 2400 438
rect 2540 392 2564 438
rect 2364 375 2564 392
rect 2812 438 3012 472
rect 2812 392 2848 438
rect 2988 392 3012 438
rect 2812 375 3012 392
rect 3260 438 3460 472
rect 3260 392 3296 438
rect 3436 392 3460 438
rect 3260 375 3460 392
rect 124 311 324 324
rect 124 265 152 311
rect 292 265 324 311
rect 124 232 324 265
rect 572 311 772 324
rect 572 265 600 311
rect 740 265 772 311
rect 572 232 772 265
rect 1020 311 1220 324
rect 1020 265 1048 311
rect 1188 265 1220 311
rect 1020 232 1220 265
rect 1468 311 1668 324
rect 1468 265 1496 311
rect 1636 265 1668 311
rect 1468 232 1668 265
rect 1916 311 2116 324
rect 1916 265 1944 311
rect 2084 265 2116 311
rect 1916 232 2116 265
rect 2364 311 2564 324
rect 2364 265 2392 311
rect 2532 265 2564 311
rect 2364 232 2564 265
rect 2812 311 3012 324
rect 2812 265 2840 311
rect 2980 265 3012 311
rect 2812 232 3012 265
rect 3260 311 3460 324
rect 3260 265 3288 311
rect 3428 265 3460 311
rect 3260 232 3460 265
rect 124 24 324 68
rect 572 24 772 68
rect 1020 24 1220 68
rect 1468 24 1668 68
rect 1916 24 2116 68
rect 2364 24 2564 68
rect 2812 24 3012 68
rect 3260 24 3460 68
<< polycontact >>
rect 160 392 300 438
rect 608 392 748 438
rect 1056 392 1196 438
rect 1504 392 1644 438
rect 1952 392 2092 438
rect 2400 392 2540 438
rect 2848 392 2988 438
rect 3296 392 3436 438
rect 152 265 292 311
rect 600 265 740 311
rect 1048 265 1188 311
rect 1496 265 1636 311
rect 1944 265 2084 311
rect 2392 265 2532 311
rect 2840 265 2980 311
rect 3288 265 3428 311
<< metal1 >>
rect 0 724 3584 844
rect 49 657 95 678
rect 49 311 95 517
rect 353 657 399 724
rect 353 498 399 517
rect 497 657 543 678
rect 146 392 160 438
rect 300 392 399 438
rect 49 265 152 311
rect 292 265 304 311
rect 49 192 95 209
rect 49 60 95 146
rect 353 192 399 392
rect 497 311 543 517
rect 801 657 847 724
rect 801 498 847 517
rect 945 657 991 678
rect 594 392 608 438
rect 748 392 847 438
rect 497 265 600 311
rect 740 265 752 311
rect 353 106 399 146
rect 497 192 543 209
rect 497 60 543 146
rect 801 192 847 392
rect 945 311 991 517
rect 1249 657 1295 724
rect 1249 498 1295 517
rect 1393 657 1439 678
rect 1042 392 1056 438
rect 1196 392 1295 438
rect 945 265 1048 311
rect 1188 265 1200 311
rect 801 106 847 146
rect 945 192 991 209
rect 945 60 991 146
rect 1249 192 1295 392
rect 1393 311 1439 517
rect 1697 657 1743 724
rect 1697 498 1743 517
rect 1841 657 1887 678
rect 1490 392 1504 438
rect 1644 392 1743 438
rect 1393 265 1496 311
rect 1636 265 1648 311
rect 1249 106 1295 146
rect 1393 192 1439 209
rect 1393 60 1439 146
rect 1697 192 1743 392
rect 1841 311 1887 517
rect 2145 657 2191 724
rect 2145 498 2191 517
rect 2289 657 2335 678
rect 1938 392 1952 438
rect 2092 392 2191 438
rect 1841 265 1944 311
rect 2084 265 2096 311
rect 1697 106 1743 146
rect 1841 192 1887 209
rect 1841 60 1887 146
rect 2145 192 2191 392
rect 2289 311 2335 517
rect 2593 657 2639 724
rect 2593 498 2639 517
rect 2737 657 2783 678
rect 2386 392 2400 438
rect 2540 392 2639 438
rect 2289 265 2392 311
rect 2532 265 2544 311
rect 2145 106 2191 146
rect 2289 192 2335 209
rect 2289 60 2335 146
rect 2593 192 2639 392
rect 2737 311 2783 517
rect 3041 657 3087 724
rect 3041 498 3087 517
rect 3185 657 3231 678
rect 2834 392 2848 438
rect 2988 392 3087 438
rect 2737 265 2840 311
rect 2980 265 2992 311
rect 2593 106 2639 146
rect 2737 192 2783 209
rect 2737 60 2783 146
rect 3041 192 3087 392
rect 3185 311 3231 517
rect 3489 657 3535 724
rect 3489 498 3535 517
rect 3282 392 3296 438
rect 3436 392 3535 438
rect 3185 265 3288 311
rect 3428 265 3440 311
rect 3041 106 3087 146
rect 3185 192 3231 209
rect 3185 60 3231 146
rect 3489 192 3535 392
rect 3489 106 3535 146
rect 0 -60 3584 60
<< labels >>
flabel metal1 s 0 724 3584 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 3185 60 3231 209 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3489 498 3535 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 3041 498 3087 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2593 498 2639 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2145 498 2191 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 498 1743 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 498 1295 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 498 847 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 2737 60 2783 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 209 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3584 60 1 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 784
string GDS_END 395038
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 385046
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
