* NGSPICE file created from ffra.ext - technology: gf180mcuC

.subckt ffra a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] ci[0] ci[1] ci[2] ci[3] ci[4]
+ ci[5] ci[6] ci[7] clk o[0] o[1] o[2] o[3] o[4] o[5] o[6] o[7] rst vdd vss
.ends

