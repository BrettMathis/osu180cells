magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 1630 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 700 190 760 360
rect 870 190 930 360
rect 1040 190 1100 360
rect 1210 190 1270 360
rect 1380 190 1440 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 700 1090 760 1430
rect 870 1090 930 1430
rect 1040 1090 1100 1430
rect 1210 1090 1270 1430
rect 1380 1090 1440 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 298 530 360
rect 420 252 452 298
rect 498 252 530 298
rect 420 190 530 252
rect 590 298 700 360
rect 590 252 622 298
rect 668 252 700 298
rect 590 190 700 252
rect 760 298 870 360
rect 760 252 792 298
rect 838 252 870 298
rect 760 190 870 252
rect 930 298 1040 360
rect 930 252 962 298
rect 1008 252 1040 298
rect 930 190 1040 252
rect 1100 298 1210 360
rect 1100 252 1132 298
rect 1178 252 1210 298
rect 1100 190 1210 252
rect 1270 298 1380 360
rect 1270 252 1302 298
rect 1348 252 1380 298
rect 1270 190 1380 252
rect 1440 298 1540 360
rect 1440 252 1472 298
rect 1518 252 1540 298
rect 1440 190 1540 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 700 1430
rect 590 1143 622 1377
rect 668 1143 700 1377
rect 590 1090 700 1143
rect 760 1377 870 1430
rect 760 1143 792 1377
rect 838 1143 870 1377
rect 760 1090 870 1143
rect 930 1377 1040 1430
rect 930 1143 962 1377
rect 1008 1143 1040 1377
rect 930 1090 1040 1143
rect 1100 1377 1210 1430
rect 1100 1143 1132 1377
rect 1178 1143 1210 1377
rect 1100 1090 1210 1143
rect 1270 1377 1380 1430
rect 1270 1143 1302 1377
rect 1348 1143 1380 1377
rect 1270 1090 1380 1143
rect 1440 1377 1540 1430
rect 1440 1143 1472 1377
rect 1518 1143 1540 1377
rect 1440 1090 1540 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 452 252 498 298
rect 622 252 668 298
rect 792 252 838 298
rect 962 252 1008 298
rect 1132 252 1178 298
rect 1302 252 1348 298
rect 1472 252 1518 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 792 1143 838 1377
rect 962 1143 1008 1377
rect 1132 1143 1178 1377
rect 1302 1143 1348 1377
rect 1472 1143 1518 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
rect 1290 1568 1380 1590
rect 1290 1522 1312 1568
rect 1358 1522 1380 1568
rect 1290 1500 1380 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 700 1430 760 1480
rect 870 1430 930 1480
rect 1040 1430 1100 1480
rect 1210 1430 1270 1480
rect 1380 1430 1440 1480
rect 190 1040 250 1090
rect 360 1040 420 1090
rect 530 1040 590 1090
rect 700 1040 760 1090
rect 870 1040 930 1090
rect 1040 1040 1100 1090
rect 1210 1040 1270 1090
rect 1380 1040 1440 1090
rect 190 990 1440 1040
rect 190 800 250 990
rect 160 780 250 800
rect 90 758 250 780
rect 90 712 112 758
rect 158 712 250 758
rect 90 690 250 712
rect 160 680 250 690
rect 190 450 250 680
rect 190 400 1440 450
rect 190 360 250 400
rect 360 360 420 400
rect 530 360 590 400
rect 700 360 760 400
rect 870 360 930 400
rect 1040 360 1100 400
rect 1210 360 1270 400
rect 1380 360 1440 400
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 700 140 760 190
rect 870 140 930 190
rect 1040 140 1100 190
rect 1210 140 1270 190
rect 1380 140 1440 190
<< polycontact >>
rect 112 712 158 758
<< metal1 >>
rect 0 1568 1630 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1630 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1630 1566
rect 0 1470 1630 1514
rect 110 1377 160 1470
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 1060 160 1143
rect 280 1377 330 1430
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 940 330 1143
rect 450 1377 500 1470
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1060 500 1143
rect 620 1377 670 1430
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 940 670 1143
rect 790 1377 840 1470
rect 790 1143 792 1377
rect 838 1143 840 1377
rect 790 1060 840 1143
rect 960 1377 1010 1430
rect 960 1143 962 1377
rect 1008 1143 1010 1377
rect 960 940 1010 1143
rect 1130 1377 1180 1470
rect 1130 1143 1132 1377
rect 1178 1143 1180 1377
rect 1130 1060 1180 1143
rect 1300 1377 1350 1430
rect 1300 1143 1302 1377
rect 1348 1143 1350 1377
rect 1300 940 1350 1143
rect 1470 1377 1520 1470
rect 1470 1143 1472 1377
rect 1518 1143 1520 1377
rect 1470 1060 1520 1143
rect 280 936 1350 940
rect 280 884 1294 936
rect 1346 884 1350 936
rect 280 860 1350 884
rect 80 758 180 760
rect 80 756 112 758
rect 80 704 104 756
rect 158 712 180 758
rect 156 704 180 712
rect 80 670 180 704
rect 280 460 330 860
rect 620 460 670 860
rect 960 460 1010 860
rect 1270 840 1350 860
rect 1300 460 1350 840
rect 280 380 1350 460
rect 110 298 160 360
rect 110 252 112 298
rect 158 252 160 298
rect 110 120 160 252
rect 280 298 330 380
rect 280 252 282 298
rect 328 252 330 298
rect 280 160 330 252
rect 450 298 500 360
rect 450 252 452 298
rect 498 252 500 298
rect 450 120 500 252
rect 620 298 670 380
rect 620 252 622 298
rect 668 252 670 298
rect 620 160 670 252
rect 790 298 840 360
rect 790 252 792 298
rect 838 252 840 298
rect 790 120 840 252
rect 960 298 1010 380
rect 960 252 962 298
rect 1008 252 1010 298
rect 960 160 1010 252
rect 1130 298 1180 360
rect 1130 252 1132 298
rect 1178 252 1180 298
rect 1130 120 1180 252
rect 1300 298 1350 380
rect 1300 252 1302 298
rect 1348 252 1350 298
rect 1300 160 1350 252
rect 1470 298 1520 360
rect 1470 252 1472 298
rect 1518 252 1520 298
rect 1470 120 1520 252
rect 0 106 1630 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1630 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1630 54
rect 0 -30 1630 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 1294 884 1346 936
rect 104 712 112 756
rect 112 712 156 756
rect 104 704 156 712
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1480 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1480 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1480 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1480 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1480 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1480 1390 1514
rect 100 1470 180 1480
rect 340 1470 420 1480
rect 580 1470 660 1480
rect 820 1470 900 1480
rect 1060 1470 1140 1480
rect 1300 1470 1380 1480
rect 1270 936 1370 950
rect 1270 884 1294 936
rect 1346 884 1370 936
rect 1270 840 1370 884
rect 80 756 180 770
rect 80 704 104 756
rect 156 704 180 756
rect 80 660 180 704
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 20 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 20 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 20 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 20 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 20 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 20 1390 54
rect 100 10 180 20
rect 340 10 420 20
rect 580 10 660 20
rect 820 10 900 20
rect 1060 10 1140 20
rect 1300 10 1380 20
<< labels >>
rlabel metal2 s 100 1470 180 1550 4 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 100 10 180 90 4 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 80 660 180 740 4 A
port 1 nsew signal input
rlabel metal2 s 1270 840 1370 920 4 Y
port 2 nsew signal output
rlabel metal1 s 80 670 180 730 1 A
port 1 nsew signal input
rlabel metal2 s 90 1480 190 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 340 1470 420 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 330 1480 430 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 580 1470 660 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 570 1480 670 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 820 1470 900 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 810 1480 910 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1060 1470 1140 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1050 1480 1150 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1300 1470 1380 1550 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 1290 1480 1390 1540 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 110 1060 160 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 450 1060 500 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 790 1060 840 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1130 1060 1180 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1470 1060 1520 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 1470 1630 1590 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 90 20 190 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 340 10 420 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 330 20 430 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 580 10 660 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 570 20 670 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 820 10 900 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 810 20 910 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1060 10 1140 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1050 20 1150 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1300 10 1380 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 1290 20 1390 80 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 110 -30 160 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 450 -30 500 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 790 -30 840 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1130 -30 1180 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 1470 -30 1520 330 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 -30 1630 90 1 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 280 160 330 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 620 160 670 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 960 160 1010 1400 1 Y
port 2 nsew signal output
rlabel metal1 s 280 380 1350 430 1 Y
port 2 nsew signal output
rlabel metal1 s 1270 840 1350 910 1 Y
port 2 nsew signal output
rlabel metal1 s 280 860 1350 910 1 Y
port 2 nsew signal output
rlabel metal1 s 1300 160 1350 1400 1 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 -30 1630 1590
string GDS_END 370242
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 357858
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
