magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 1044
<< mvndiff >>
rect -88 1031 0 1044
rect -88 985 -75 1031
rect -29 985 0 1031
rect -88 923 0 985
rect -88 877 -75 923
rect -29 877 0 923
rect -88 815 0 877
rect -88 769 -75 815
rect -29 769 0 815
rect -88 707 0 769
rect -88 661 -75 707
rect -29 661 0 707
rect -88 599 0 661
rect -88 553 -75 599
rect -29 553 0 599
rect -88 491 0 553
rect -88 445 -75 491
rect -29 445 0 491
rect -88 383 0 445
rect -88 337 -75 383
rect -29 337 0 383
rect -88 275 0 337
rect -88 229 -75 275
rect -29 229 0 275
rect -88 167 0 229
rect -88 121 -75 167
rect -29 121 0 167
rect -88 59 0 121
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1031 208 1044
rect 120 985 149 1031
rect 195 985 208 1031
rect 120 923 208 985
rect 120 877 149 923
rect 195 877 208 923
rect 120 815 208 877
rect 120 769 149 815
rect 195 769 208 815
rect 120 707 208 769
rect 120 661 149 707
rect 195 661 208 707
rect 120 599 208 661
rect 120 553 149 599
rect 195 553 208 599
rect 120 491 208 553
rect 120 445 149 491
rect 195 445 208 491
rect 120 383 208 445
rect 120 337 149 383
rect 195 337 208 383
rect 120 275 208 337
rect 120 229 149 275
rect 195 229 208 275
rect 120 167 208 229
rect 120 121 149 167
rect 195 121 208 167
rect 120 59 208 121
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 985 -29 1031
rect -75 877 -29 923
rect -75 769 -29 815
rect -75 661 -29 707
rect -75 553 -29 599
rect -75 445 -29 491
rect -75 337 -29 383
rect -75 229 -29 275
rect -75 121 -29 167
rect -75 13 -29 59
rect 149 985 195 1031
rect 149 877 195 923
rect 149 769 195 815
rect 149 661 195 707
rect 149 553 195 599
rect 149 445 195 491
rect 149 337 195 383
rect 149 229 195 275
rect 149 121 195 167
rect 149 13 195 59
<< polysilicon >>
rect 0 1044 120 1088
rect 0 -44 120 0
<< metal1 >>
rect -75 1031 -29 1044
rect -75 923 -29 985
rect -75 815 -29 877
rect -75 707 -29 769
rect -75 599 -29 661
rect -75 491 -29 553
rect -75 383 -29 445
rect -75 275 -29 337
rect -75 167 -29 229
rect -75 59 -29 121
rect -75 0 -29 13
rect 149 1031 195 1044
rect 149 923 195 985
rect 149 815 195 877
rect 149 707 195 769
rect 149 599 195 661
rect 149 491 195 553
rect 149 383 195 445
rect 149 275 195 337
rect 149 167 195 229
rect 149 59 195 121
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 522 -52 522 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 522 172 522 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 179060
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 176884
<< end >>
