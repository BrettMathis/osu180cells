magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
<< mvpmos >>
rect 124 610 224 939
rect 368 573 468 939
rect 582 573 682 939
rect 796 573 896 939
<< mvndiff >>
rect 36 297 124 333
rect 36 157 49 297
rect 95 157 124 297
rect 36 69 124 157
rect 244 297 348 333
rect 244 157 273 297
rect 319 157 348 297
rect 244 69 348 157
rect 468 274 572 333
rect 468 228 497 274
rect 543 228 572 274
rect 468 69 572 228
rect 692 203 796 333
rect 692 157 721 203
rect 767 157 796 203
rect 692 69 796 157
rect 916 297 1004 333
rect 916 157 945 297
rect 991 157 1004 297
rect 916 69 1004 157
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 610 124 721
rect 224 861 368 939
rect 224 721 293 861
rect 339 721 368 861
rect 224 610 368 721
rect 288 573 368 610
rect 468 573 582 939
rect 682 573 796 939
rect 896 861 984 939
rect 896 721 925 861
rect 971 721 984 861
rect 896 573 984 721
<< mvndiffc >>
rect 49 157 95 297
rect 273 157 319 297
rect 497 228 543 274
rect 721 157 767 203
rect 945 157 991 297
<< mvpdiffc >>
rect 49 721 95 861
rect 293 721 339 861
rect 925 721 971 861
<< polysilicon >>
rect 124 939 224 983
rect 368 939 468 983
rect 582 939 682 983
rect 796 939 896 983
rect 124 500 224 610
rect 124 454 137 500
rect 183 454 224 500
rect 124 377 224 454
rect 368 500 468 573
rect 368 454 381 500
rect 427 454 468 500
rect 368 377 468 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 377 682 454
rect 796 500 896 573
rect 796 454 809 500
rect 855 454 896 500
rect 796 377 896 454
rect 124 333 244 377
rect 348 333 468 377
rect 572 333 692 377
rect 796 333 916 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
<< polycontact >>
rect 137 454 183 500
rect 381 454 427 500
rect 595 454 641 500
rect 809 454 855 500
<< metal1 >>
rect 0 918 1120 1098
rect 49 861 95 918
rect 49 710 95 721
rect 293 861 339 872
rect 925 861 971 918
rect 339 721 530 766
rect 293 690 530 721
rect 925 710 971 721
rect 366 500 427 511
rect 126 454 137 500
rect 183 454 194 500
rect 126 354 194 454
rect 366 454 381 500
rect 366 354 427 454
rect 484 308 530 690
rect 584 454 595 500
rect 641 454 652 500
rect 584 354 652 454
rect 798 454 809 500
rect 855 454 866 500
rect 798 354 866 454
rect 49 297 95 308
rect 49 90 95 157
rect 273 297 319 308
rect 484 297 991 308
rect 484 274 945 297
rect 484 228 497 274
rect 543 262 945 274
rect 543 228 554 262
rect 721 203 767 214
rect 319 157 721 182
rect 273 136 767 157
rect 945 146 991 157
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 366 354 427 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 584 354 652 500 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 798 354 866 500 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 126 354 194 500 0 FreeSans 200 0 0 0 B
port 4 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 49 90 95 308 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 293 766 339 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
rlabel metal1 s 293 690 530 766 1 ZN
port 5 nsew default output
rlabel metal1 s 484 308 530 690 1 ZN
port 5 nsew default output
rlabel metal1 s 484 262 991 308 1 ZN
port 5 nsew default output
rlabel metal1 s 945 228 991 262 1 ZN
port 5 nsew default output
rlabel metal1 s 484 228 554 262 1 ZN
port 5 nsew default output
rlabel metal1 s 945 146 991 228 1 ZN
port 5 nsew default output
rlabel metal1 s 925 710 971 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 145026
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 141458
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
