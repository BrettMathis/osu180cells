magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 2550 870
<< pwell >>
rect -86 -86 2550 352
<< mvnmos >>
rect 124 79 244 172
rect 384 93 504 172
rect 552 93 672 172
rect 776 93 896 172
rect 944 93 1064 172
rect 1204 79 1324 172
rect 1388 79 1508 172
rect 1756 68 1876 232
rect 1980 68 2100 232
rect 2204 68 2324 232
<< mvpmos >>
rect 144 531 244 716
rect 384 590 484 716
rect 532 590 632 716
rect 736 590 836 716
rect 944 590 1044 716
rect 1204 531 1304 716
rect 1408 531 1508 716
rect 1776 472 1876 716
rect 2000 472 2100 716
rect 2204 472 2304 716
<< mvndiff >>
rect 36 152 124 172
rect 36 106 49 152
rect 95 106 124 152
rect 36 79 124 106
rect 244 152 384 172
rect 244 106 273 152
rect 319 106 384 152
rect 244 93 384 106
rect 504 93 552 172
rect 672 152 776 172
rect 672 106 701 152
rect 747 106 776 152
rect 672 93 776 106
rect 896 93 944 172
rect 1064 152 1204 172
rect 1064 106 1093 152
rect 1139 106 1204 152
rect 1064 93 1204 106
rect 244 79 324 93
rect 1124 79 1204 93
rect 1324 79 1388 172
rect 1508 152 1596 172
rect 1508 106 1537 152
rect 1583 106 1596 152
rect 1508 79 1596 106
rect 1668 168 1756 232
rect 1668 122 1681 168
rect 1727 122 1756 168
rect 1668 68 1756 122
rect 1876 168 1980 232
rect 1876 122 1905 168
rect 1951 122 1980 168
rect 1876 68 1980 122
rect 2100 168 2204 232
rect 2100 122 2129 168
rect 2175 122 2204 168
rect 2100 68 2204 122
rect 2324 168 2412 232
rect 2324 122 2353 168
rect 2399 122 2412 168
rect 2324 68 2412 122
<< mvpdiff >>
rect 56 665 144 716
rect 56 619 69 665
rect 115 619 144 665
rect 56 531 144 619
rect 244 665 384 716
rect 244 619 273 665
rect 319 619 384 665
rect 244 590 384 619
rect 484 590 532 716
rect 632 665 736 716
rect 632 619 661 665
rect 707 619 736 665
rect 632 590 736 619
rect 836 590 944 716
rect 1044 665 1204 716
rect 1044 619 1073 665
rect 1119 619 1204 665
rect 1044 590 1204 619
rect 244 531 324 590
rect 1124 531 1204 590
rect 1304 665 1408 716
rect 1304 619 1333 665
rect 1379 619 1408 665
rect 1304 531 1408 619
rect 1508 703 1596 716
rect 1508 563 1537 703
rect 1583 563 1596 703
rect 1508 531 1596 563
rect 1688 665 1776 716
rect 1688 525 1701 665
rect 1747 525 1776 665
rect 1688 472 1776 525
rect 1876 665 2000 716
rect 1876 525 1905 665
rect 1951 525 2000 665
rect 1876 472 2000 525
rect 2100 665 2204 716
rect 2100 525 2129 665
rect 2175 525 2204 665
rect 2100 472 2204 525
rect 2304 665 2392 716
rect 2304 525 2333 665
rect 2379 525 2392 665
rect 2304 472 2392 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 701 106 747 152
rect 1093 106 1139 152
rect 1537 106 1583 152
rect 1681 122 1727 168
rect 1905 122 1951 168
rect 2129 122 2175 168
rect 2353 122 2399 168
<< mvpdiffc >>
rect 69 619 115 665
rect 273 619 319 665
rect 661 619 707 665
rect 1073 619 1119 665
rect 1333 619 1379 665
rect 1537 563 1583 703
rect 1701 525 1747 665
rect 1905 525 1951 665
rect 2129 525 2175 665
rect 2333 525 2379 665
<< polysilicon >>
rect 144 716 244 760
rect 384 716 484 760
rect 532 716 632 760
rect 736 716 836 760
rect 944 716 1044 760
rect 1204 716 1304 760
rect 1408 716 1508 760
rect 1776 716 1876 760
rect 2000 716 2100 760
rect 2204 716 2304 760
rect 144 413 244 531
rect 124 302 244 413
rect 124 256 175 302
rect 221 256 244 302
rect 124 172 244 256
rect 384 414 484 590
rect 384 368 411 414
rect 457 368 484 414
rect 384 268 484 368
rect 532 516 632 590
rect 532 470 559 516
rect 605 470 632 516
rect 532 409 632 470
rect 736 516 836 590
rect 736 470 763 516
rect 809 470 836 516
rect 736 457 836 470
rect 944 516 1044 590
rect 944 470 981 516
rect 1027 470 1044 516
rect 944 467 1044 470
rect 532 363 896 409
rect 552 302 672 315
rect 384 172 504 268
rect 552 256 593 302
rect 639 256 672 302
rect 552 172 672 256
rect 776 172 896 363
rect 944 172 1064 467
rect 1204 444 1304 531
rect 1408 444 1508 531
rect 1204 291 1324 444
rect 1204 245 1241 291
rect 1287 245 1324 291
rect 1204 172 1324 245
rect 1388 415 1508 444
rect 1388 369 1411 415
rect 1457 369 1508 415
rect 1776 404 1876 472
rect 1388 172 1508 369
rect 1756 372 1876 404
rect 2000 385 2100 472
rect 2204 385 2304 472
rect 1756 326 1792 372
rect 1838 326 1876 372
rect 1756 232 1876 326
rect 1980 372 2324 385
rect 1980 326 2019 372
rect 2159 326 2324 372
rect 1980 313 2324 326
rect 1980 232 2100 313
rect 2204 232 2324 313
rect 124 35 244 79
rect 384 35 504 93
rect 552 35 672 93
rect 776 35 896 93
rect 944 35 1064 93
rect 1204 35 1324 79
rect 1388 35 1508 79
rect 1756 24 1876 68
rect 1980 24 2100 68
rect 2204 24 2324 68
<< polycontact >>
rect 175 256 221 302
rect 411 368 457 414
rect 559 470 605 516
rect 763 470 809 516
rect 981 470 1027 516
rect 593 256 639 302
rect 1241 245 1287 291
rect 1411 369 1457 415
rect 1792 326 1838 372
rect 2019 326 2159 372
<< metal1 >>
rect 0 724 2464 844
rect 38 665 115 676
rect 38 619 69 665
rect 38 516 115 619
rect 273 665 319 724
rect 1073 665 1119 724
rect 1526 703 1594 724
rect 632 619 661 665
rect 707 619 912 665
rect 273 600 319 619
rect 700 516 809 559
rect 38 470 559 516
rect 605 470 632 516
rect 700 470 763 516
rect 38 152 106 470
rect 193 414 654 424
rect 193 368 411 414
rect 457 368 654 414
rect 193 358 654 368
rect 700 312 809 470
rect 156 302 809 312
rect 156 256 175 302
rect 221 256 593 302
rect 639 256 809 302
rect 156 248 809 256
rect 864 291 912 619
rect 1073 600 1119 619
rect 1333 665 1379 676
rect 1333 516 1379 619
rect 1526 563 1537 703
rect 1583 563 1594 703
rect 1701 665 1747 676
rect 962 470 981 516
rect 1027 470 1594 516
rect 1008 415 1476 424
rect 1008 369 1411 415
rect 1457 369 1476 415
rect 1008 360 1476 369
rect 1526 372 1594 470
rect 1701 468 1747 525
rect 1905 665 1951 724
rect 1905 514 1951 525
rect 2128 665 2220 676
rect 2128 525 2129 665
rect 2175 525 2220 665
rect 2128 468 2220 525
rect 2333 665 2379 724
rect 2333 514 2379 525
rect 1701 422 1963 468
rect 2128 422 2332 468
rect 1917 372 1963 422
rect 1526 326 1792 372
rect 1838 326 1849 372
rect 1917 326 2019 372
rect 2159 326 2187 372
rect 864 245 1241 291
rect 1287 245 1306 291
rect 38 106 49 152
rect 95 106 106 152
rect 273 152 319 172
rect 864 152 912 245
rect 682 106 701 152
rect 747 106 912 152
rect 1093 152 1139 172
rect 1526 152 1594 326
rect 1917 276 1963 326
rect 2260 276 2332 422
rect 1526 106 1537 152
rect 1583 106 1594 152
rect 1681 230 1963 276
rect 1681 168 1727 230
rect 2128 226 2332 276
rect 1681 111 1727 122
rect 1905 168 1951 179
rect 273 60 319 106
rect 1093 60 1139 106
rect 1905 60 1951 122
rect 2128 168 2220 226
rect 2128 122 2129 168
rect 2175 122 2220 168
rect 2128 111 2220 122
rect 2353 168 2399 179
rect 2353 60 2399 122
rect 0 -60 2464 60
<< labels >>
flabel metal1 s 2128 468 2220 676 0 FreeSans 400 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2353 172 2399 179 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 1008 360 1476 424 0 FreeSans 400 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 724 2464 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 193 358 654 424 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel metal1 s 700 312 809 559 0 FreeSans 400 0 0 0 E
port 2 nsew clock input
rlabel metal1 s 156 248 809 312 1 E
port 2 nsew clock input
rlabel metal1 s 2128 422 2332 468 1 Q
port 4 nsew default output
rlabel metal1 s 2260 276 2332 422 1 Q
port 4 nsew default output
rlabel metal1 s 2128 226 2332 276 1 Q
port 4 nsew default output
rlabel metal1 s 2128 111 2220 226 1 Q
port 4 nsew default output
rlabel metal1 s 2333 600 2379 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1905 600 1951 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 600 1594 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1073 600 1119 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 600 319 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2333 563 2379 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1905 563 1951 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1526 563 1594 600 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2333 514 2379 563 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1905 514 1951 563 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1905 172 1951 179 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2353 60 2399 172 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1905 60 1951 172 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1093 60 1139 172 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 172 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string GDS_END 640520
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 634662
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
