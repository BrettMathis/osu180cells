magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -296 -137 586 284
<< polysilicon >>
rect -31 2526 89 2597
rect 193 2526 313 2597
rect -31 -71 89 -1
rect 193 -71 313 -1
use pmos_5p043105899832102_64x8m81  pmos_5p043105899832102_64x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 552 2646
<< properties >>
string GDS_END 1333714
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1333272
<< end >>
