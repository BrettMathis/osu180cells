magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -79 513 80 572
rect -79 467 -23 513
rect 23 467 80 513
rect -79 350 80 467
rect -79 304 -23 350
rect 23 304 80 350
rect -79 186 80 304
rect -79 140 -23 186
rect 23 140 80 186
rect -79 23 80 140
rect -79 -23 -23 23
rect 23 -23 80 23
rect -79 -140 80 -23
rect -79 -186 -23 -140
rect 23 -186 80 -140
rect -79 -304 80 -186
rect -79 -350 -23 -304
rect 23 -350 80 -304
rect -79 -467 80 -350
rect -79 -513 -23 -467
rect 23 -513 80 -467
rect -79 -572 80 -513
<< psubdiffcont >>
rect -23 467 23 513
rect -23 304 23 350
rect -23 140 23 186
rect -23 -23 23 23
rect -23 -186 23 -140
rect -23 -350 23 -304
rect -23 -513 23 -467
<< metal1 >>
rect -70 513 71 563
rect -70 467 -23 513
rect 23 467 71 513
rect -70 350 71 467
rect -70 304 -23 350
rect 23 304 71 350
rect -70 186 71 304
rect -70 140 -23 186
rect 23 140 71 186
rect -70 23 71 140
rect -70 -23 -23 23
rect 23 -23 71 23
rect -70 -140 71 -23
rect -70 -186 -23 -140
rect 23 -186 71 -140
rect -70 -304 71 -186
rect -70 -350 -23 -304
rect 23 -350 71 -304
rect -70 -467 71 -350
rect -70 -513 -23 -467
rect 23 -513 71 -467
rect -70 -563 71 -513
<< properties >>
string GDS_END 241202
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 240558
<< end >>
