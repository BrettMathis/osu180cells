magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 610 800 1230
<< nmos >>
rect 180 190 240 360
rect 350 190 410 360
rect 540 190 600 360
<< pmos >>
rect 210 700 270 1040
rect 330 700 390 1040
rect 520 700 580 1040
<< ndiff >>
rect 80 268 180 360
rect 80 222 102 268
rect 148 222 180 268
rect 80 190 180 222
rect 240 258 350 360
rect 240 212 272 258
rect 318 212 350 258
rect 240 190 350 212
rect 410 268 540 360
rect 410 222 452 268
rect 498 222 540 268
rect 410 190 540 222
rect 600 288 700 360
rect 600 242 632 288
rect 678 242 700 288
rect 600 190 700 242
<< pdiff >>
rect 110 987 210 1040
rect 110 753 132 987
rect 178 753 210 987
rect 110 700 210 753
rect 270 700 330 1040
rect 390 980 520 1040
rect 390 840 432 980
rect 478 840 520 980
rect 390 700 520 840
rect 580 988 680 1040
rect 580 942 612 988
rect 658 942 680 988
rect 580 770 680 942
rect 580 700 690 770
<< ndiffc >>
rect 102 222 148 268
rect 272 212 318 258
rect 452 222 498 268
rect 632 242 678 288
<< pdiffc >>
rect 132 753 178 987
rect 432 840 478 980
rect 612 942 658 988
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
<< nsubdiff >>
rect 90 1178 180 1200
rect 90 1132 112 1178
rect 158 1132 180 1178
rect 90 1110 180 1132
rect 330 1178 420 1200
rect 330 1132 352 1178
rect 398 1132 420 1178
rect 330 1110 420 1132
rect 570 1178 660 1200
rect 570 1132 592 1178
rect 638 1132 660 1178
rect 570 1110 660 1132
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
<< nsubdiffcont >>
rect 112 1132 158 1178
rect 352 1132 398 1178
rect 592 1132 638 1178
<< polysilicon >>
rect 210 1040 270 1090
rect 330 1040 390 1090
rect 520 1040 580 1090
rect 210 680 270 700
rect 160 640 270 680
rect 330 650 390 700
rect 160 520 220 640
rect 320 623 430 650
rect 320 577 357 623
rect 403 577 430 623
rect 320 550 430 577
rect 110 493 220 520
rect 110 447 147 493
rect 193 450 220 493
rect 330 450 390 550
rect 520 520 580 700
rect 470 493 600 520
rect 193 447 240 450
rect 110 420 240 447
rect 330 420 410 450
rect 470 447 497 493
rect 543 447 600 493
rect 470 420 600 447
rect 180 360 240 420
rect 350 360 410 420
rect 540 360 600 420
rect 180 140 240 190
rect 350 140 410 190
rect 540 140 600 190
<< polycontact >>
rect 357 577 403 623
rect 147 447 193 493
rect 497 447 543 493
<< metal1 >>
rect 0 1178 800 1230
rect 0 1132 112 1178
rect 158 1176 352 1178
rect 398 1176 592 1178
rect 638 1176 800 1178
rect 166 1132 352 1176
rect 406 1132 592 1176
rect 0 1124 114 1132
rect 166 1124 354 1132
rect 406 1124 594 1132
rect 646 1124 800 1176
rect 0 1110 800 1124
rect 130 987 180 1110
rect 130 753 132 987
rect 178 753 180 987
rect 130 700 180 753
rect 420 980 490 1040
rect 420 840 432 980
rect 478 840 490 980
rect 610 988 660 1110
rect 610 942 612 988
rect 658 942 660 988
rect 610 890 660 942
rect 420 760 490 840
rect 420 756 700 760
rect 420 704 624 756
rect 676 704 700 756
rect 420 700 700 704
rect 620 690 690 700
rect 330 626 430 630
rect 330 574 354 626
rect 406 574 430 626
rect 330 570 430 574
rect 120 496 220 500
rect 120 444 144 496
rect 196 444 220 496
rect 120 440 220 444
rect 470 496 570 500
rect 470 444 494 496
rect 546 444 570 496
rect 470 440 570 444
rect 100 330 510 380
rect 100 268 150 330
rect 100 222 102 268
rect 148 222 150 268
rect 100 190 150 222
rect 270 258 320 280
rect 270 212 272 258
rect 318 212 320 258
rect 270 120 320 212
rect 440 268 510 330
rect 440 222 452 268
rect 498 222 510 268
rect 440 190 510 222
rect 630 288 680 690
rect 630 242 632 288
rect 678 242 680 288
rect 630 190 680 242
rect 0 106 800 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 800 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 800 54
rect 0 0 800 52
<< via1 >>
rect 114 1132 158 1176
rect 158 1132 166 1176
rect 354 1132 398 1176
rect 398 1132 406 1176
rect 594 1132 638 1176
rect 638 1132 646 1176
rect 114 1124 166 1132
rect 354 1124 406 1132
rect 594 1124 646 1132
rect 624 704 676 756
rect 354 623 406 626
rect 354 577 357 623
rect 357 577 403 623
rect 403 577 406 623
rect 354 574 406 577
rect 144 493 196 496
rect 144 447 147 493
rect 147 447 193 493
rect 193 447 196 493
rect 144 444 196 447
rect 494 493 546 496
rect 494 447 497 493
rect 497 447 543 493
rect 543 447 546 493
rect 494 444 546 447
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
<< metal2 >>
rect 100 1180 180 1190
rect 340 1180 420 1190
rect 580 1180 660 1190
rect 90 1176 190 1180
rect 90 1124 114 1176
rect 166 1124 190 1176
rect 90 1120 190 1124
rect 330 1176 430 1180
rect 330 1124 354 1176
rect 406 1124 430 1176
rect 330 1120 430 1124
rect 570 1176 670 1180
rect 570 1124 594 1176
rect 646 1124 670 1176
rect 570 1120 670 1124
rect 100 1110 180 1120
rect 340 1110 420 1120
rect 580 1110 660 1120
rect 610 760 690 770
rect 600 756 700 760
rect 600 704 624 756
rect 676 704 700 756
rect 600 700 700 704
rect 610 690 690 700
rect 330 626 430 640
rect 330 574 354 626
rect 406 574 430 626
rect 330 560 430 574
rect 120 496 220 510
rect 120 444 144 496
rect 196 444 220 496
rect 120 430 220 444
rect 470 496 570 510
rect 470 444 494 496
rect 546 444 570 496
rect 470 430 570 444
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
<< labels >>
rlabel metal2 s 100 1110 180 1190 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 100 40 180 120 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 610 690 690 770 4 Y
port 1 nsew signal output
rlabel metal2 s 120 430 220 510 4 A0
port 2 nsew signal input
rlabel metal2 s 330 560 430 640 4 A1
port 3 nsew signal input
rlabel metal2 s 470 430 570 510 4 B
port 4 nsew signal input
rlabel metal1 s 120 440 220 500 1 A0
port 2 nsew signal input
rlabel metal1 s 330 570 430 630 1 A1
port 3 nsew signal input
rlabel metal1 s 470 440 570 500 1 B
port 4 nsew signal input
rlabel metal2 s 90 1120 190 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 340 1110 420 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 330 1120 430 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 1110 660 1190 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 570 1120 670 1180 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 130 700 180 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 610 890 660 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 1110 800 1230 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 270 0 320 280 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 0 0 800 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 600 700 700 760 1 Y
port 1 nsew signal output
rlabel metal1 s 420 700 490 1040 1 Y
port 1 nsew signal output
rlabel metal1 s 630 190 680 760 1 Y
port 1 nsew signal output
rlabel metal1 s 620 690 690 760 1 Y
port 1 nsew signal output
rlabel metal1 s 420 700 700 760 1 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 800 1230
string GDS_END 432138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 424990
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
