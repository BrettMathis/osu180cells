magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 302
<< mvpmos >>
rect 0 0 120 182
<< mvpdiff >>
rect -88 169 0 182
rect -88 123 -75 169
rect -29 123 0 169
rect -88 59 0 123
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 169 208 182
rect 120 123 149 169
rect 195 123 208 169
rect 120 59 208 123
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 123 -29 169
rect -75 13 -29 59
rect 149 123 195 169
rect 149 13 195 59
<< polysilicon >>
rect 0 182 120 226
rect 0 -44 120 0
<< metal1 >>
rect -75 169 -29 182
rect -75 59 -29 123
rect -75 0 -29 13
rect 149 169 195 182
rect 149 59 195 123
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 91 -52 91 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 91 172 91 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 147738
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 146522
<< end >>
