magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 0 1000 1620 1620
<< nmos >>
rect 190 190 250 360
rect 360 190 420 360
rect 530 190 590 360
rect 850 190 910 360
rect 1020 190 1080 360
rect 1190 190 1250 360
rect 1360 190 1420 360
<< pmos >>
rect 190 1090 250 1430
rect 360 1090 420 1430
rect 530 1090 590 1430
rect 850 1090 910 1430
rect 1020 1090 1080 1430
rect 1190 1090 1250 1430
rect 1360 1090 1420 1430
<< ndiff >>
rect 90 298 190 360
rect 90 252 112 298
rect 158 252 190 298
rect 90 190 190 252
rect 250 298 360 360
rect 250 252 282 298
rect 328 252 360 298
rect 250 190 360 252
rect 420 190 530 360
rect 590 298 690 360
rect 590 252 622 298
rect 668 252 690 298
rect 590 190 690 252
rect 750 298 850 360
rect 750 252 772 298
rect 818 252 850 298
rect 750 190 850 252
rect 910 338 1020 360
rect 910 292 942 338
rect 988 292 1020 338
rect 910 190 1020 292
rect 1080 298 1190 360
rect 1080 252 1112 298
rect 1158 252 1190 298
rect 1080 190 1190 252
rect 1250 298 1360 360
rect 1250 252 1282 298
rect 1328 252 1360 298
rect 1250 190 1360 252
rect 1420 298 1520 360
rect 1420 252 1452 298
rect 1498 252 1520 298
rect 1420 190 1520 252
<< pdiff >>
rect 90 1377 190 1430
rect 90 1143 112 1377
rect 158 1143 190 1377
rect 90 1090 190 1143
rect 250 1377 360 1430
rect 250 1143 282 1377
rect 328 1143 360 1377
rect 250 1090 360 1143
rect 420 1377 530 1430
rect 420 1143 452 1377
rect 498 1143 530 1377
rect 420 1090 530 1143
rect 590 1377 690 1430
rect 590 1143 622 1377
rect 668 1143 690 1377
rect 590 1090 690 1143
rect 750 1377 850 1430
rect 750 1143 772 1377
rect 818 1143 850 1377
rect 750 1090 850 1143
rect 910 1090 1020 1430
rect 1080 1377 1190 1430
rect 1080 1143 1112 1377
rect 1158 1143 1190 1377
rect 1080 1090 1190 1143
rect 1250 1377 1360 1430
rect 1250 1143 1282 1377
rect 1328 1143 1360 1377
rect 1250 1090 1360 1143
rect 1420 1377 1520 1430
rect 1420 1143 1452 1377
rect 1498 1143 1520 1377
rect 1420 1090 1520 1143
<< ndiffc >>
rect 112 252 158 298
rect 282 252 328 298
rect 622 252 668 298
rect 772 252 818 298
rect 942 292 988 338
rect 1112 252 1158 298
rect 1282 252 1328 298
rect 1452 252 1498 298
<< pdiffc >>
rect 112 1143 158 1377
rect 282 1143 328 1377
rect 452 1143 498 1377
rect 622 1143 668 1377
rect 772 1143 818 1377
rect 1112 1143 1158 1377
rect 1282 1143 1328 1377
rect 1452 1143 1498 1377
<< psubdiff >>
rect 90 98 180 120
rect 90 52 112 98
rect 158 52 180 98
rect 90 30 180 52
rect 330 98 420 120
rect 330 52 352 98
rect 398 52 420 98
rect 330 30 420 52
rect 570 98 660 120
rect 570 52 592 98
rect 638 52 660 98
rect 570 30 660 52
rect 810 98 900 120
rect 810 52 832 98
rect 878 52 900 98
rect 810 30 900 52
rect 1050 98 1140 120
rect 1050 52 1072 98
rect 1118 52 1140 98
rect 1050 30 1140 52
rect 1290 98 1380 120
rect 1290 52 1312 98
rect 1358 52 1380 98
rect 1290 30 1380 52
<< nsubdiff >>
rect 90 1568 180 1590
rect 90 1522 112 1568
rect 158 1522 180 1568
rect 90 1500 180 1522
rect 330 1568 420 1590
rect 330 1522 352 1568
rect 398 1522 420 1568
rect 330 1500 420 1522
rect 570 1568 660 1590
rect 570 1522 592 1568
rect 638 1522 660 1568
rect 570 1500 660 1522
rect 810 1568 900 1590
rect 810 1522 832 1568
rect 878 1522 900 1568
rect 810 1500 900 1522
rect 1050 1568 1140 1590
rect 1050 1522 1072 1568
rect 1118 1522 1140 1568
rect 1050 1500 1140 1522
rect 1290 1568 1380 1590
rect 1290 1522 1312 1568
rect 1358 1522 1380 1568
rect 1290 1500 1380 1522
<< psubdiffcont >>
rect 112 52 158 98
rect 352 52 398 98
rect 592 52 638 98
rect 832 52 878 98
rect 1072 52 1118 98
rect 1312 52 1358 98
<< nsubdiffcont >>
rect 112 1522 158 1568
rect 352 1522 398 1568
rect 592 1522 638 1568
rect 832 1522 878 1568
rect 1072 1522 1118 1568
rect 1312 1522 1358 1568
<< polysilicon >>
rect 190 1430 250 1480
rect 360 1430 420 1480
rect 530 1430 590 1480
rect 850 1430 910 1480
rect 1020 1430 1080 1480
rect 1190 1430 1250 1480
rect 1360 1430 1420 1480
rect 190 1040 250 1090
rect 190 1013 310 1040
rect 190 967 237 1013
rect 283 967 310 1013
rect 190 940 310 967
rect 190 360 250 940
rect 360 780 420 1090
rect 300 753 420 780
rect 300 707 327 753
rect 373 707 420 753
rect 300 680 420 707
rect 360 360 420 680
rect 530 650 590 1090
rect 850 780 910 1090
rect 780 753 910 780
rect 780 707 807 753
rect 853 707 910 753
rect 780 680 910 707
rect 470 623 590 650
rect 470 577 497 623
rect 543 577 590 623
rect 470 550 590 577
rect 530 360 590 550
rect 850 360 910 680
rect 1020 650 1080 1090
rect 1190 1040 1250 1090
rect 1190 1013 1310 1040
rect 1190 967 1237 1013
rect 1283 967 1310 1013
rect 1190 940 1310 967
rect 1020 623 1140 650
rect 1020 577 1067 623
rect 1113 577 1140 623
rect 1020 550 1140 577
rect 1020 360 1080 550
rect 1190 360 1250 940
rect 1360 780 1420 1090
rect 1300 753 1420 780
rect 1300 707 1327 753
rect 1373 707 1420 753
rect 1300 680 1420 707
rect 1360 360 1420 680
rect 190 140 250 190
rect 360 140 420 190
rect 530 140 590 190
rect 850 140 910 190
rect 1020 140 1080 190
rect 1190 140 1250 190
rect 1360 140 1420 190
<< polycontact >>
rect 237 967 283 1013
rect 327 707 373 753
rect 807 707 853 753
rect 497 577 543 623
rect 1237 967 1283 1013
rect 1067 577 1113 623
rect 1327 707 1373 753
<< metal1 >>
rect 0 1568 1620 1620
rect 0 1522 112 1568
rect 158 1566 352 1568
rect 398 1566 592 1568
rect 638 1566 832 1568
rect 878 1566 1072 1568
rect 1118 1566 1312 1568
rect 1358 1566 1620 1568
rect 166 1522 352 1566
rect 406 1522 592 1566
rect 646 1522 832 1566
rect 886 1522 1072 1566
rect 1126 1522 1312 1566
rect 0 1514 114 1522
rect 166 1514 354 1522
rect 406 1514 594 1522
rect 646 1514 834 1522
rect 886 1514 1074 1522
rect 1126 1514 1314 1522
rect 1366 1514 1620 1566
rect 0 1500 1620 1514
rect 110 1377 160 1430
rect 110 1143 112 1377
rect 158 1143 160 1377
rect 110 500 160 1143
rect 280 1377 330 1500
rect 280 1143 282 1377
rect 328 1143 330 1377
rect 280 1090 330 1143
rect 450 1377 500 1430
rect 450 1143 452 1377
rect 498 1143 500 1377
rect 450 1020 500 1143
rect 620 1377 670 1500
rect 620 1143 622 1377
rect 668 1143 670 1377
rect 620 1090 670 1143
rect 770 1377 820 1500
rect 770 1143 772 1377
rect 818 1143 820 1377
rect 770 1090 820 1143
rect 1110 1377 1160 1430
rect 1110 1143 1112 1377
rect 1158 1143 1160 1377
rect 210 1016 700 1020
rect 210 1013 624 1016
rect 210 967 237 1013
rect 283 967 624 1013
rect 210 964 624 967
rect 676 964 700 1016
rect 210 960 700 964
rect 300 756 400 760
rect 300 704 324 756
rect 376 704 400 756
rect 300 700 400 704
rect 470 626 570 630
rect 470 574 494 626
rect 546 574 570 626
rect 470 570 570 574
rect 80 496 180 500
rect 80 444 104 496
rect 156 444 180 496
rect 80 440 180 444
rect 110 298 160 440
rect 110 252 112 298
rect 158 252 160 298
rect 110 190 160 252
rect 280 298 330 360
rect 280 252 282 298
rect 328 252 330 298
rect 280 120 330 252
rect 620 298 670 960
rect 1110 760 1160 1143
rect 1280 1377 1330 1500
rect 1280 1143 1282 1377
rect 1328 1143 1330 1377
rect 1280 1090 1330 1143
rect 1450 1377 1500 1430
rect 1450 1143 1452 1377
rect 1498 1143 1500 1377
rect 1450 1030 1500 1143
rect 1450 1020 1520 1030
rect 1210 1016 1310 1020
rect 1210 964 1234 1016
rect 1286 964 1310 1016
rect 1210 960 1310 964
rect 1440 1016 1540 1020
rect 1440 964 1464 1016
rect 1516 964 1540 1016
rect 1440 960 1540 964
rect 1450 950 1520 960
rect 780 756 880 760
rect 780 704 804 756
rect 856 704 880 756
rect 1110 753 1400 760
rect 1110 750 1327 753
rect 780 700 880 704
rect 940 707 1327 750
rect 1373 707 1400 753
rect 940 700 1400 707
rect 620 252 622 298
rect 668 252 670 298
rect 620 190 670 252
rect 770 298 820 380
rect 770 252 772 298
rect 818 252 820 298
rect 940 338 990 700
rect 1040 626 1140 630
rect 1040 574 1064 626
rect 1116 574 1140 626
rect 1040 570 1140 574
rect 940 292 942 338
rect 988 292 990 338
rect 940 270 990 292
rect 1110 298 1160 380
rect 770 220 820 252
rect 1110 252 1112 298
rect 1158 252 1160 298
rect 1110 220 1160 252
rect 770 170 1160 220
rect 1280 298 1330 360
rect 1280 252 1282 298
rect 1328 252 1330 298
rect 1280 120 1330 252
rect 1450 298 1500 950
rect 1450 252 1452 298
rect 1498 252 1500 298
rect 1450 190 1500 252
rect 0 106 1620 120
rect 0 98 114 106
rect 166 98 354 106
rect 406 98 594 106
rect 646 98 834 106
rect 886 98 1074 106
rect 1126 98 1314 106
rect 0 52 112 98
rect 166 54 352 98
rect 406 54 592 98
rect 646 54 832 98
rect 886 54 1072 98
rect 1126 54 1312 98
rect 1366 54 1620 106
rect 158 52 352 54
rect 398 52 592 54
rect 638 52 832 54
rect 878 52 1072 54
rect 1118 52 1312 54
rect 1358 52 1620 54
rect 0 0 1620 52
<< via1 >>
rect 114 1522 158 1566
rect 158 1522 166 1566
rect 354 1522 398 1566
rect 398 1522 406 1566
rect 594 1522 638 1566
rect 638 1522 646 1566
rect 834 1522 878 1566
rect 878 1522 886 1566
rect 1074 1522 1118 1566
rect 1118 1522 1126 1566
rect 1314 1522 1358 1566
rect 1358 1522 1366 1566
rect 114 1514 166 1522
rect 354 1514 406 1522
rect 594 1514 646 1522
rect 834 1514 886 1522
rect 1074 1514 1126 1522
rect 1314 1514 1366 1522
rect 624 964 676 1016
rect 324 753 376 756
rect 324 707 327 753
rect 327 707 373 753
rect 373 707 376 753
rect 324 704 376 707
rect 494 623 546 626
rect 494 577 497 623
rect 497 577 543 623
rect 543 577 546 623
rect 494 574 546 577
rect 104 444 156 496
rect 1234 1013 1286 1016
rect 1234 967 1237 1013
rect 1237 967 1283 1013
rect 1283 967 1286 1013
rect 1234 964 1286 967
rect 1464 964 1516 1016
rect 804 753 856 756
rect 804 707 807 753
rect 807 707 853 753
rect 853 707 856 753
rect 804 704 856 707
rect 1064 623 1116 626
rect 1064 577 1067 623
rect 1067 577 1113 623
rect 1113 577 1116 623
rect 1064 574 1116 577
rect 114 98 166 106
rect 354 98 406 106
rect 594 98 646 106
rect 834 98 886 106
rect 1074 98 1126 106
rect 1314 98 1366 106
rect 114 54 158 98
rect 158 54 166 98
rect 354 54 398 98
rect 398 54 406 98
rect 594 54 638 98
rect 638 54 646 98
rect 834 54 878 98
rect 878 54 886 98
rect 1074 54 1118 98
rect 1118 54 1126 98
rect 1314 54 1358 98
rect 1358 54 1366 98
<< metal2 >>
rect 100 1570 180 1580
rect 340 1570 420 1580
rect 580 1570 660 1580
rect 820 1570 900 1580
rect 1060 1570 1140 1580
rect 1300 1570 1380 1580
rect 90 1566 190 1570
rect 90 1514 114 1566
rect 166 1514 190 1566
rect 90 1510 190 1514
rect 330 1566 430 1570
rect 330 1514 354 1566
rect 406 1514 430 1566
rect 330 1510 430 1514
rect 570 1566 670 1570
rect 570 1514 594 1566
rect 646 1514 670 1566
rect 570 1510 670 1514
rect 810 1566 910 1570
rect 810 1514 834 1566
rect 886 1514 910 1566
rect 810 1510 910 1514
rect 1050 1566 1150 1570
rect 1050 1514 1074 1566
rect 1126 1514 1150 1566
rect 1050 1510 1150 1514
rect 1290 1566 1390 1570
rect 1290 1514 1314 1566
rect 1366 1514 1390 1566
rect 1290 1510 1390 1514
rect 100 1500 180 1510
rect 340 1500 420 1510
rect 580 1500 660 1510
rect 820 1500 900 1510
rect 1060 1500 1140 1510
rect 1300 1500 1380 1510
rect 600 1020 700 1030
rect 1210 1020 1310 1030
rect 600 1016 1310 1020
rect 600 964 624 1016
rect 676 964 1234 1016
rect 1286 964 1310 1016
rect 600 960 1310 964
rect 600 950 700 960
rect 1210 950 1310 960
rect 1440 1016 1540 1030
rect 1440 964 1464 1016
rect 1516 964 1540 1016
rect 1440 950 1540 964
rect 300 760 400 770
rect 780 760 880 770
rect 300 756 880 760
rect 300 704 324 756
rect 376 704 804 756
rect 856 704 880 756
rect 300 700 880 704
rect 300 690 400 700
rect 780 690 880 700
rect 470 630 570 640
rect 1040 630 1140 640
rect 470 626 1140 630
rect 470 574 494 626
rect 546 574 1064 626
rect 1116 574 1140 626
rect 470 570 1140 574
rect 470 560 570 570
rect 1040 560 1140 570
rect 80 496 180 510
rect 80 444 104 496
rect 156 444 180 496
rect 80 430 180 444
rect 100 110 180 120
rect 340 110 420 120
rect 580 110 660 120
rect 820 110 900 120
rect 1060 110 1140 120
rect 1300 110 1380 120
rect 90 106 190 110
rect 90 54 114 106
rect 166 54 190 106
rect 90 50 190 54
rect 330 106 430 110
rect 330 54 354 106
rect 406 54 430 106
rect 330 50 430 54
rect 570 106 670 110
rect 570 54 594 106
rect 646 54 670 106
rect 570 50 670 54
rect 810 106 910 110
rect 810 54 834 106
rect 886 54 910 106
rect 810 50 910 54
rect 1050 106 1150 110
rect 1050 54 1074 106
rect 1126 54 1150 106
rect 1050 50 1150 54
rect 1290 106 1390 110
rect 1290 54 1314 106
rect 1366 54 1390 106
rect 1290 50 1390 54
rect 100 40 180 50
rect 340 40 420 50
rect 580 40 660 50
rect 820 40 900 50
rect 1060 40 1140 50
rect 1300 40 1380 50
<< labels >>
rlabel metal2 s 100 40 180 120 4 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 100 1500 180 1580 4 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 300 690 400 770 4 A
port 1 nsew signal input
rlabel metal2 s 470 560 570 640 4 B
port 2 nsew signal input
rlabel metal2 s 1440 950 1540 1030 4 S
port 3 nsew signal output
rlabel metal2 s 80 430 180 510 4 CO
port 4 nsew signal output
rlabel metal2 s 300 700 880 760 1 A
port 1 nsew signal input
rlabel metal2 s 780 690 880 770 1 A
port 1 nsew signal input
rlabel metal1 s 300 700 400 760 1 A
port 1 nsew signal input
rlabel metal1 s 780 700 880 760 1 A
port 1 nsew signal input
rlabel metal2 s 470 570 1140 630 1 B
port 2 nsew signal input
rlabel metal2 s 1040 560 1140 640 1 B
port 2 nsew signal input
rlabel metal1 s 470 570 570 630 1 B
port 2 nsew signal input
rlabel metal1 s 1040 570 1140 630 1 B
port 2 nsew signal input
rlabel metal1 s 110 190 160 1430 1 CO
port 4 nsew signal output
rlabel metal1 s 80 440 180 500 1 CO
port 4 nsew signal output
rlabel metal1 s 1450 190 1500 1430 1 S
port 3 nsew signal output
rlabel metal1 s 1450 950 1520 1030 1 S
port 3 nsew signal output
rlabel metal1 s 1440 960 1540 1020 1 S
port 3 nsew signal output
rlabel metal2 s 90 1510 190 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 340 1500 420 1580 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 330 1510 430 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 580 1500 660 1580 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 570 1510 670 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 820 1500 900 1580 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 810 1510 910 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1060 1500 1140 1580 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1050 1510 1150 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1300 1500 1380 1580 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 1290 1510 1390 1570 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 280 1090 330 1620 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 620 1090 670 1620 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 770 1090 820 1620 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 1280 1090 1330 1620 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal1 s 0 1500 1620 1620 1 VDD
port 10 nsew power bidirectional abutment
rlabel metal2 s 90 50 190 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 340 40 420 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 330 50 430 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 580 40 660 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 570 50 670 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 820 40 900 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 810 50 910 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1060 40 1140 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1050 50 1150 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1300 40 1380 120 1 VSS
port 11 nsew ground bidirectional
rlabel metal2 s 1290 50 1390 110 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 280 0 330 360 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 1280 0 1330 360 1 VSS
port 11 nsew ground bidirectional
rlabel metal1 s 0 0 1620 120 1 VSS
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1620 1620
string GDS_END 39936
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_12T/gds/gf180mcu_osu_sc_12T.gds
string GDS_START 25556
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
