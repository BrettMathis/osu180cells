magic
tech gf180mcuB
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -81 820 81 825
rect -81 792 -76 820
rect -48 792 -14 820
rect 14 792 48 820
rect 76 792 81 820
rect -81 758 81 792
rect -81 730 -76 758
rect -48 730 -14 758
rect 14 730 48 758
rect 76 730 81 758
rect -81 696 81 730
rect -81 668 -76 696
rect -48 668 -14 696
rect 14 668 48 696
rect 76 668 81 696
rect -81 634 81 668
rect -81 606 -76 634
rect -48 606 -14 634
rect 14 606 48 634
rect 76 606 81 634
rect -81 572 81 606
rect -81 544 -76 572
rect -48 544 -14 572
rect 14 544 48 572
rect 76 544 81 572
rect -81 510 81 544
rect -81 482 -76 510
rect -48 482 -14 510
rect 14 482 48 510
rect 76 482 81 510
rect -81 448 81 482
rect -81 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 81 448
rect -81 386 81 420
rect -81 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 81 386
rect -81 324 81 358
rect -81 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 81 324
rect -81 262 81 296
rect -81 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 81 262
rect -81 200 81 234
rect -81 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 81 200
rect -81 138 81 172
rect -81 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 81 138
rect -81 76 81 110
rect -81 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 81 76
rect -81 14 81 48
rect -81 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 81 14
rect -81 -48 81 -14
rect -81 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 81 -48
rect -81 -110 81 -76
rect -81 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 81 -110
rect -81 -172 81 -138
rect -81 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 81 -172
rect -81 -234 81 -200
rect -81 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 81 -234
rect -81 -296 81 -262
rect -81 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 81 -296
rect -81 -358 81 -324
rect -81 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 81 -358
rect -81 -420 81 -386
rect -81 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 81 -420
rect -81 -482 81 -448
rect -81 -510 -76 -482
rect -48 -510 -14 -482
rect 14 -510 48 -482
rect 76 -510 81 -482
rect -81 -544 81 -510
rect -81 -572 -76 -544
rect -48 -572 -14 -544
rect 14 -572 48 -544
rect 76 -572 81 -544
rect -81 -606 81 -572
rect -81 -634 -76 -606
rect -48 -634 -14 -606
rect 14 -634 48 -606
rect 76 -634 81 -606
rect -81 -668 81 -634
rect -81 -696 -76 -668
rect -48 -696 -14 -668
rect 14 -696 48 -668
rect 76 -696 81 -668
rect -81 -730 81 -696
rect -81 -758 -76 -730
rect -48 -758 -14 -730
rect 14 -758 48 -730
rect 76 -758 81 -730
rect -81 -792 81 -758
rect -81 -820 -76 -792
rect -48 -820 -14 -792
rect 14 -820 48 -792
rect 76 -820 81 -792
rect -81 -825 81 -820
<< via2 >>
rect -76 792 -48 820
rect -14 792 14 820
rect 48 792 76 820
rect -76 730 -48 758
rect -14 730 14 758
rect 48 730 76 758
rect -76 668 -48 696
rect -14 668 14 696
rect 48 668 76 696
rect -76 606 -48 634
rect -14 606 14 634
rect 48 606 76 634
rect -76 544 -48 572
rect -14 544 14 572
rect 48 544 76 572
rect -76 482 -48 510
rect -14 482 14 510
rect 48 482 76 510
rect -76 420 -48 448
rect -14 420 14 448
rect 48 420 76 448
rect -76 358 -48 386
rect -14 358 14 386
rect 48 358 76 386
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect -76 -386 -48 -358
rect -14 -386 14 -358
rect 48 -386 76 -358
rect -76 -448 -48 -420
rect -14 -448 14 -420
rect 48 -448 76 -420
rect -76 -510 -48 -482
rect -14 -510 14 -482
rect 48 -510 76 -482
rect -76 -572 -48 -544
rect -14 -572 14 -544
rect 48 -572 76 -544
rect -76 -634 -48 -606
rect -14 -634 14 -606
rect 48 -634 76 -606
rect -76 -696 -48 -668
rect -14 -696 14 -668
rect 48 -696 76 -668
rect -76 -758 -48 -730
rect -14 -758 14 -730
rect 48 -758 76 -730
rect -76 -820 -48 -792
rect -14 -820 14 -792
rect 48 -820 76 -792
<< metal3 >>
rect -81 820 81 825
rect -81 792 -76 820
rect -48 792 -14 820
rect 14 792 48 820
rect 76 792 81 820
rect -81 758 81 792
rect -81 730 -76 758
rect -48 730 -14 758
rect 14 730 48 758
rect 76 730 81 758
rect -81 696 81 730
rect -81 668 -76 696
rect -48 668 -14 696
rect 14 668 48 696
rect 76 668 81 696
rect -81 634 81 668
rect -81 606 -76 634
rect -48 606 -14 634
rect 14 606 48 634
rect 76 606 81 634
rect -81 572 81 606
rect -81 544 -76 572
rect -48 544 -14 572
rect 14 544 48 572
rect 76 544 81 572
rect -81 510 81 544
rect -81 482 -76 510
rect -48 482 -14 510
rect 14 482 48 510
rect 76 482 81 510
rect -81 448 81 482
rect -81 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 81 448
rect -81 386 81 420
rect -81 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 81 386
rect -81 324 81 358
rect -81 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 81 324
rect -81 262 81 296
rect -81 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 81 262
rect -81 200 81 234
rect -81 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 81 200
rect -81 138 81 172
rect -81 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 81 138
rect -81 76 81 110
rect -81 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 81 76
rect -81 14 81 48
rect -81 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 81 14
rect -81 -48 81 -14
rect -81 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 81 -48
rect -81 -110 81 -76
rect -81 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 81 -110
rect -81 -172 81 -138
rect -81 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 81 -172
rect -81 -234 81 -200
rect -81 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 81 -234
rect -81 -296 81 -262
rect -81 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 81 -296
rect -81 -358 81 -324
rect -81 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 81 -358
rect -81 -420 81 -386
rect -81 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 81 -420
rect -81 -482 81 -448
rect -81 -510 -76 -482
rect -48 -510 -14 -482
rect 14 -510 48 -482
rect 76 -510 81 -482
rect -81 -544 81 -510
rect -81 -572 -76 -544
rect -48 -572 -14 -544
rect 14 -572 48 -544
rect 76 -572 81 -544
rect -81 -606 81 -572
rect -81 -634 -76 -606
rect -48 -634 -14 -606
rect 14 -634 48 -606
rect 76 -634 81 -606
rect -81 -668 81 -634
rect -81 -696 -76 -668
rect -48 -696 -14 -668
rect 14 -696 48 -668
rect 76 -696 81 -668
rect -81 -730 81 -696
rect -81 -758 -76 -730
rect -48 -758 -14 -730
rect 14 -758 48 -730
rect 76 -758 81 -730
rect -81 -792 81 -758
rect -81 -820 -76 -792
rect -48 -820 -14 -792
rect 14 -820 48 -792
rect 76 -820 81 -792
rect -81 -825 81 -820
<< properties >>
string GDS_END 755712
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 750396
<< end >>
