magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 278 92 308
rect 0 226 20 278
rect 72 226 92 278
rect 0 92 92 226
rect 0 40 20 92
rect 72 40 92 92
rect 0 0 92 40
<< via1 >>
rect 20 226 72 278
rect 20 40 72 92
<< metal2 >>
rect 0 280 92 308
rect 0 224 18 280
rect 74 224 92 280
rect 0 94 92 224
rect 0 38 18 94
rect 74 38 92 94
rect 0 0 92 38
<< via2 >>
rect 18 278 74 280
rect 18 226 20 278
rect 20 226 72 278
rect 72 226 74 278
rect 18 224 74 226
rect 18 92 74 94
rect 18 40 20 92
rect 20 40 72 92
rect 72 40 74 92
rect 18 38 74 40
<< metal3 >>
rect 0 280 93 308
rect 0 224 18 280
rect 74 224 93 280
rect 0 94 93 224
rect 0 38 18 94
rect 74 38 93 94
rect 0 -1 93 38
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 0
box 0 0 1 1
use via2_x2_R90_128x8m81  via2_x2_R90_128x8m81_0
timestamp 1669390400
transform 1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 308872
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 308780
<< end >>
