magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 224 844
rect 28 162 95 542
rect 0 -60 224 60
<< labels >>
rlabel metal1 s 28 162 95 542 6 I
port 1 nsew default input
rlabel metal1 s 0 724 224 844 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -60 224 60 8 VSS
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 784
string LEFclass core ANTENNACELL
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1223506
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1222028
<< end >>
