magic
tech gf180mcuC
timestamp 1669390400
<< metal1 >>
rect 0 111 80 123
rect 13 70 18 111
rect 42 76 49 104
rect 61 89 66 111
rect 42 70 70 76
rect 62 69 69 70
rect 33 57 43 63
rect 12 44 22 50
rect 47 44 57 50
rect 27 12 32 28
rect 63 19 68 69
rect 0 0 80 12
<< obsm1 >>
rect 10 33 51 38
rect 10 19 15 33
rect 44 19 51 33
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 61 76 69 77
rect 60 70 70 76
rect 61 69 69 70
rect 33 56 43 64
rect 12 43 22 51
rect 47 43 57 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 s 12 43 22 51 6 A0
port 2 nsew signal input
rlabel metal1 s 12 44 22 50 6 A0
port 2 nsew signal input
rlabel metal2 s 33 56 43 64 6 A1
port 3 nsew signal input
rlabel metal1 s 33 57 43 63 6 A1
port 3 nsew signal input
rlabel metal2 s 47 43 57 51 6 B
port 4 nsew signal input
rlabel metal1 s 47 44 57 50 6 B
port 4 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal1 s 13 70 18 123 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal1 s 61 89 66 123 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal1 s 0 111 80 123 6 VDD
port 9 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 10 nsew ground bidirectional
rlabel metal1 s 27 0 32 28 6 VSS
port 10 nsew ground bidirectional
rlabel metal1 s 0 0 80 12 6 VSS
port 10 nsew ground bidirectional
rlabel metal2 s 61 69 69 77 6 Y
port 1 nsew signal output
rlabel metal2 s 60 70 70 76 6 Y
port 1 nsew signal output
rlabel metal1 s 42 70 49 104 6 Y
port 1 nsew signal output
rlabel metal1 s 63 19 68 76 6 Y
port 1 nsew signal output
rlabel metal1 s 62 69 69 76 6 Y
port 1 nsew signal output
rlabel metal1 s 42 70 70 76 6 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 432138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_osu_sc_9T/gds/gf180mcu_osu_sc_9T.gds
string GDS_START 424990
<< end >>
