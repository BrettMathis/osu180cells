magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -530 4793 759 5011
rect -530 3964 4955 4793
rect -530 3963 4956 3964
rect -530 2692 5175 3963
rect -530 2672 4573 2692
rect 2599 2671 4573 2672
rect 2600 2602 4573 2671
rect -530 624 -82 713
rect 3535 624 4165 625
rect 4848 624 5175 679
rect -530 55 5175 624
rect -530 -24 -82 55
<< psubdiff >>
rect -352 5539 -268 5558
rect -352 5211 -333 5539
rect -287 5211 -268 5539
rect -352 5192 -268 5211
rect -389 2191 86 2250
rect -389 2145 -333 2191
rect -287 2145 -175 2191
rect -129 2145 -17 2191
rect 29 2145 86 2191
rect -389 2027 86 2145
rect -389 1981 -333 2027
rect -287 1981 -175 2027
rect -129 1981 -17 2027
rect 29 1981 86 2027
rect -389 1922 86 1981
rect 4560 2191 5035 2250
rect 4560 2145 4616 2191
rect 4662 2145 4774 2191
rect 4820 2145 4932 2191
rect 4978 2145 5035 2191
rect 4560 2027 5035 2145
rect 4560 1981 4616 2027
rect 4662 1981 4774 2027
rect 4820 1981 4932 2027
rect 4978 1981 5035 2027
rect 4560 1922 5035 1981
rect -468 1088 -151 1148
rect -468 1042 -412 1088
rect -366 1042 -254 1088
rect -208 1042 -151 1088
rect -468 983 -151 1042
rect 4718 1088 5035 1148
rect 4718 1042 4774 1088
rect 4820 1042 4932 1088
rect 4978 1042 5035 1088
rect 4718 983 5035 1042
<< nsubdiff >>
rect -387 388 -232 445
rect -387 342 -333 388
rect -287 342 -232 388
rect -387 285 -232 342
<< psubdiffcont >>
rect -333 5211 -287 5539
rect -333 2145 -287 2191
rect -175 2145 -129 2191
rect -17 2145 29 2191
rect -333 1981 -287 2027
rect -175 1981 -129 2027
rect -17 1981 29 2027
rect 4616 2145 4662 2191
rect 4774 2145 4820 2191
rect 4932 2145 4978 2191
rect 4616 1981 4662 2027
rect 4774 1981 4820 2027
rect 4932 1981 4978 2027
rect -412 1042 -366 1088
rect -254 1042 -208 1088
rect 4774 1042 4820 1088
rect 4932 1042 4978 1088
<< nsubdiffcont >>
rect -333 342 -287 388
<< polysilicon >>
rect 159 4903 279 5523
rect 383 4903 503 5523
rect 1074 5460 1194 5532
rect 1298 5460 1418 5532
rect 1522 5460 1642 5532
rect 1746 5460 1866 5532
rect 1970 5460 2090 5532
rect 2270 5520 3499 5580
rect 1074 4934 1194 5005
rect 1298 4934 1418 5005
rect 1522 4934 1642 5005
rect 1746 4934 1866 5005
rect 1970 4934 2090 5005
rect 661 4888 2090 4934
rect 661 4842 735 4888
rect 781 4873 2090 4888
rect 781 4842 854 4873
rect 661 4796 854 4842
rect 1074 4708 1194 4873
rect 1298 4708 1418 4873
rect 1522 4708 1642 4873
rect 2270 4772 2328 5520
rect 2483 5460 2603 5520
rect 2707 5460 2827 5520
rect 2931 5460 3051 5520
rect 3155 5460 3275 5520
rect 3379 5460 3499 5520
rect 3892 5460 4012 5532
rect 4116 5460 4236 5532
rect 4340 5460 4460 5532
rect 4564 5460 4684 5532
rect 2483 4932 2603 5005
rect 2707 4932 2827 5005
rect 2931 4932 3051 5005
rect 3155 4932 3275 5005
rect 3379 4932 3499 5005
rect 3892 4834 4012 5005
rect 1746 4712 2328 4772
rect 2014 4683 2328 4712
rect 2548 4788 4012 4834
rect 2548 4742 2623 4788
rect 2669 4742 2781 4788
rect 2827 4742 2939 4788
rect 2985 4742 3097 4788
rect 3143 4742 3255 4788
rect 3301 4759 4012 4788
rect 4116 4759 4236 5005
rect 4340 4759 4460 5005
rect 4564 4759 4684 5005
rect 3301 4742 4684 4759
rect 2548 4698 4684 4742
rect 2549 4696 3376 4698
rect 2014 4607 2206 4683
rect 2014 4561 2087 4607
rect 2133 4561 2206 4607
rect 2014 4443 2206 4561
rect 2014 4397 2087 4443
rect 2133 4397 2206 4443
rect 2014 4351 2206 4397
rect 159 4072 503 4118
rect 159 4026 298 4072
rect 344 4026 503 4072
rect 159 3980 503 4026
rect 2796 3788 2974 3807
rect 2796 3742 2815 3788
rect 2955 3742 2974 3788
rect 2796 3723 2974 3742
rect 391 2749 510 2790
rect 615 2749 734 2790
rect 839 2749 958 2790
rect 1063 2749 1182 2790
rect 1287 2749 1406 2790
rect 1511 2749 1630 2790
rect 1735 2749 1854 2790
rect 166 2709 2302 2749
rect 166 2690 2477 2709
rect 166 2688 2318 2690
rect 390 2323 510 2688
rect 614 2323 734 2688
rect 838 2323 958 2688
rect 1062 2323 1182 2688
rect 1286 2323 1406 2688
rect 1510 2323 1630 2688
rect 1734 2644 2318 2688
rect 2458 2644 2477 2690
rect 1734 2625 2477 2644
rect 1734 2323 1854 2625
rect 2182 2433 2302 2452
rect 2182 2387 2217 2433
rect 2263 2387 2302 2433
rect 2854 2422 2974 2712
rect 2182 2335 2302 2387
rect 2630 2361 2974 2422
rect 2854 2332 2974 2361
rect 3078 2332 3198 2712
rect 3302 2449 3422 2712
rect 3750 2671 3870 2712
rect 3975 2671 4094 2712
rect 4199 2671 4318 2672
rect 3750 2651 4318 2671
rect 3568 2632 4318 2651
rect 3568 2586 3587 2632
rect 3633 2611 4318 2632
rect 3633 2586 3870 2611
rect 3568 2568 3870 2586
rect 3568 2567 3652 2568
rect 3302 2403 3332 2449
rect 3378 2403 3422 2449
rect 3302 2365 3422 2403
rect 3303 2332 3422 2365
rect 3750 2332 3870 2568
rect 3974 2332 4094 2611
rect 2406 1577 2526 1665
rect 2406 1576 2527 1577
rect 3078 1576 3198 1688
rect 2406 1531 3198 1576
rect 2406 1516 2786 1531
rect 2713 1485 2786 1516
rect 2832 1516 3198 1531
rect 2832 1485 2905 1516
rect 2713 1440 2905 1485
rect 246 1336 439 1381
rect 246 1290 320 1336
rect 366 1290 439 1336
rect 246 1259 439 1290
rect 887 1336 1080 1381
rect 887 1290 961 1336
rect 1007 1290 1080 1336
rect 887 1259 1080 1290
rect 171 1198 1186 1259
rect 171 602 291 1198
rect 395 602 515 1198
rect 619 602 739 1198
rect 843 602 963 1198
rect 1067 602 1186 1198
rect 4251 1105 4370 1177
rect 1616 756 1736 883
rect 1305 737 1736 756
rect 1305 691 1324 737
rect 1370 691 1736 737
rect 1305 672 1736 691
rect 1616 514 1736 672
rect 1840 796 1960 861
rect 2341 815 2460 874
rect 1840 750 1859 796
rect 1905 750 1960 796
rect 1840 514 1960 750
rect 2029 796 2460 815
rect 2029 750 2048 796
rect 2094 750 2460 796
rect 2029 731 2460 750
rect 2340 683 2460 731
rect 2341 514 2460 683
rect 2565 735 2685 876
rect 3065 874 3184 883
rect 3065 754 3185 874
rect 2565 689 2584 735
rect 2630 689 2685 735
rect 2565 514 2685 689
rect 2796 735 3185 754
rect 2796 689 2815 735
rect 2861 689 3185 735
rect 2796 670 3185 689
rect 3065 514 3185 670
rect 3289 735 3409 871
rect 3790 754 3910 874
rect 3289 689 3308 735
rect 3354 689 3409 735
rect 3289 514 3409 689
rect 3495 735 3910 754
rect 3495 689 3514 735
rect 3560 689 3910 735
rect 4251 713 4371 874
rect 3495 670 3910 689
rect 3790 514 3910 670
rect 4188 694 4595 713
rect 4188 648 4207 694
rect 4253 648 4595 694
rect 4188 629 4595 648
rect 4251 514 4371 629
rect 4475 514 4595 629
rect 3790 273 3910 346
<< polycontact >>
rect 735 4842 781 4888
rect 2623 4742 2669 4788
rect 2781 4742 2827 4788
rect 2939 4742 2985 4788
rect 3097 4742 3143 4788
rect 3255 4742 3301 4788
rect 2087 4561 2133 4607
rect 2087 4397 2133 4443
rect 298 4026 344 4072
rect 2815 3742 2955 3788
rect 2318 2644 2458 2690
rect 2217 2387 2263 2433
rect 3587 2586 3633 2632
rect 3332 2403 3378 2449
rect 2786 1485 2832 1531
rect 320 1290 366 1336
rect 961 1290 1007 1336
rect 1324 691 1370 737
rect 1859 750 1905 796
rect 2048 750 2094 796
rect 2584 689 2630 735
rect 2815 689 2861 735
rect 3308 689 3354 735
rect 3514 689 3560 735
rect 4207 648 4253 694
<< metal1 >>
rect -344 5539 -276 5550
rect -344 5211 -333 5539
rect -287 5211 -276 5539
rect 1190 5530 3574 5597
rect 1190 5451 1305 5530
rect -344 5200 -276 5211
rect 308 5120 354 5451
rect 1189 5268 1305 5451
rect 1635 5145 1751 5530
rect 2083 5145 2199 5530
rect 2632 5145 2678 5530
rect 3080 5145 3126 5530
rect 3528 5315 3574 5530
rect 4007 5530 4569 5580
rect 308 5045 763 5120
rect 308 4689 354 5045
rect 691 4924 763 5045
rect 691 4888 815 4924
rect 691 4842 735 4888
rect 781 4842 815 4888
rect 2408 4843 2454 5104
rect 2856 4843 2902 5104
rect 3304 4843 3350 5104
rect 691 4805 815 4842
rect 1187 4811 3350 4843
rect 1187 4759 2313 4811
rect 2365 4759 2493 4811
rect 2545 4788 3350 4811
rect 2545 4759 2623 4788
rect 1187 4742 2623 4759
rect 2669 4742 2781 4788
rect 2827 4742 2939 4788
rect 2985 4742 3097 4788
rect 3143 4742 3255 4788
rect 3301 4742 3350 4788
rect 1187 4723 3350 4742
rect 1187 4481 1303 4723
rect 1635 4585 1751 4723
rect 2589 4705 3350 4723
rect 2054 4617 2166 4643
rect 2053 4607 2166 4617
rect 2053 4576 2087 4607
rect 2053 4524 2073 4576
rect 2133 4561 2166 4607
rect 2125 4524 2166 4561
rect 2053 4443 2166 4524
rect 2053 4397 2087 4443
rect 2133 4397 2166 4443
rect 2053 4390 2166 4397
rect 2053 4338 2073 4390
rect 2125 4360 2166 4390
rect 2125 4338 2145 4360
rect 2053 4298 2145 4338
rect 263 4072 378 4108
rect 263 4026 298 4072
rect 344 4026 378 4072
rect 263 4000 378 4026
rect 843 4000 1152 4022
rect 263 3948 881 4000
rect 933 3948 1061 4000
rect 1113 3948 1152 4000
rect 263 3925 1152 3948
rect 2665 4018 2781 4358
rect 3111 4018 3227 4379
rect 3559 4018 3675 4379
rect 4007 4018 4123 5530
rect 4453 4018 4569 5530
rect 2665 3898 4569 4018
rect 54 3721 2412 3841
rect 2778 3796 3086 3818
rect 2778 3788 2816 3796
rect 2868 3788 2996 3796
rect 2778 3742 2815 3788
rect 2955 3744 2996 3788
rect 3048 3744 3086 3796
rect 2955 3742 3086 3744
rect 2778 3722 3086 3742
rect 54 3325 170 3721
rect 505 3365 620 3721
rect 953 3365 1068 3721
rect 1400 3365 1516 3721
rect 1848 3365 1964 3721
rect 2296 3472 2412 3721
rect 281 2633 396 2866
rect 729 2633 844 2866
rect 1177 2633 1292 2866
rect 1624 2719 1740 2866
rect 2072 2719 2188 3336
rect 1624 2633 2188 2719
rect 281 2599 2188 2633
rect 2294 2718 2592 2741
rect 2294 2690 2330 2718
rect 2382 2690 2592 2718
rect 2294 2644 2318 2690
rect 2458 2644 2592 2690
rect 2968 2672 3084 2803
rect 3451 2672 3497 2803
rect 2968 2671 3085 2672
rect 3451 2671 3533 2672
rect 281 2513 1740 2599
rect 2294 2583 2592 2644
rect 2744 2632 3655 2671
rect 2744 2586 3587 2632
rect 3633 2586 3655 2632
rect -380 2191 77 2240
rect -380 2145 -333 2191
rect -287 2145 -175 2191
rect -129 2145 -17 2191
rect 29 2145 77 2191
rect 281 2187 396 2513
rect 729 2187 844 2513
rect 1177 2187 1292 2513
rect 1624 2187 1740 2513
rect 2744 2552 3655 2586
rect 2181 2449 2489 2471
rect 2181 2433 2219 2449
rect 2181 2387 2217 2433
rect 2271 2397 2399 2449
rect 2451 2397 2489 2449
rect 2263 2387 2489 2397
rect 2181 2375 2489 2387
rect -380 2027 77 2145
rect -380 1981 -333 2027
rect -287 1981 -175 2027
rect -129 1981 -17 2027
rect 29 1981 77 2027
rect -380 1931 77 1981
rect 505 1762 620 2186
rect 953 1762 1068 2186
rect 1400 1762 1516 2186
rect 1870 1762 1942 2035
rect 2744 1765 2860 2552
rect 3083 2449 3391 2471
rect 3083 2397 3121 2449
rect 3173 2397 3301 2449
rect 3378 2403 3391 2449
rect 3353 2397 3391 2403
rect 3083 2375 3391 2397
rect 3864 2162 3980 2842
rect 4569 2191 5026 2240
rect 4569 2145 4616 2191
rect 4662 2145 4774 2191
rect 4820 2145 4932 2191
rect 4978 2145 5026 2191
rect 4569 2027 5026 2145
rect 4569 1981 4616 2027
rect 4662 1981 4774 2027
rect 4820 1981 4932 2027
rect 4978 1981 5026 2027
rect 4569 1931 5026 1981
rect 4574 1786 4955 1826
rect 505 1688 1942 1762
rect 4574 1734 4611 1786
rect 4663 1734 4823 1786
rect 4875 1734 4955 1786
rect 74 1568 414 1608
rect 864 1604 4470 1608
rect 74 1516 112 1568
rect 164 1516 324 1568
rect 376 1516 414 1568
rect 74 1390 414 1516
rect 860 1584 4470 1604
rect 860 1532 890 1584
rect 942 1532 1076 1584
rect 1128 1532 4191 1584
rect 4243 1532 4377 1584
rect 4429 1532 4470 1584
rect 860 1531 4470 1532
rect 860 1512 2786 1531
rect 864 1511 2786 1512
rect 2752 1485 2786 1511
rect 2832 1511 4470 1531
rect 4574 1568 4955 1734
rect 4574 1516 4611 1568
rect 4663 1516 4823 1568
rect 4875 1516 4955 1568
rect 2832 1485 2867 1511
rect 2752 1471 2867 1485
rect 4574 1391 4955 1516
rect 4574 1390 4956 1391
rect -374 1350 5025 1390
rect -374 1298 112 1350
rect 164 1336 324 1350
rect 376 1336 4611 1350
rect 164 1298 320 1336
rect 376 1298 961 1336
rect -374 1290 320 1298
rect 366 1290 961 1298
rect 1007 1298 4611 1336
rect 4663 1298 4823 1350
rect 4875 1298 5025 1350
rect 1007 1290 5025 1298
rect -374 1253 5025 1290
rect -460 1088 -160 1139
rect -460 1042 -412 1088
rect -366 1042 -254 1088
rect -208 1042 -160 1088
rect -460 992 -160 1042
rect 72 1121 164 1161
rect 72 1069 92 1121
rect 144 1069 164 1121
rect -277 991 -262 992
rect 72 935 164 1069
rect 492 1121 584 1161
rect 492 1069 512 1121
rect 564 1069 584 1121
rect 72 883 92 935
rect 144 883 164 935
rect 72 842 164 883
rect 320 762 366 1017
rect 492 935 584 1069
rect 964 1121 1056 1161
rect 964 1069 984 1121
rect 1036 1069 1056 1121
rect 492 883 512 935
rect 564 883 584 935
rect 492 842 584 883
rect 768 762 814 1017
rect 964 935 1056 1069
rect 1216 1154 1604 1155
rect 1216 1132 1729 1154
rect 1216 1080 1459 1132
rect 1511 1080 1639 1132
rect 1691 1080 1729 1132
rect 1216 1058 1729 1080
rect 1820 1121 1916 1161
rect 1820 1069 1840 1121
rect 1892 1069 1916 1121
rect 964 883 984 935
rect 1036 883 1056 935
rect 964 842 1056 883
rect 1216 762 1262 1017
rect 1541 826 1587 1004
rect 1820 935 1916 1069
rect 2481 1121 2573 1161
rect 2481 1069 2501 1121
rect 2553 1069 2573 1121
rect 1820 883 1840 935
rect 1892 883 1916 935
rect 1989 884 2109 1004
rect 1820 842 1916 883
rect 1504 786 1596 826
rect 320 737 1413 762
rect 320 691 1324 737
rect 1370 691 1413 737
rect 320 643 1413 691
rect 1504 734 1524 786
rect 1576 734 1596 786
rect 1848 796 1916 842
rect 1848 750 1859 796
rect 1905 750 1916 796
rect 1848 739 1916 750
rect 2037 796 2109 884
rect 2037 750 2048 796
rect 2094 750 2109 796
rect 320 461 366 643
rect 732 642 814 643
rect 1180 642 1262 643
rect 768 461 814 642
rect 1216 461 1262 642
rect 1504 600 1596 734
rect 1504 548 1524 600
rect 1576 548 1596 600
rect 1504 507 1596 548
rect -367 388 -252 425
rect -367 342 -333 388
rect -287 342 -252 388
rect 1541 355 1587 507
rect 2037 355 2109 750
rect 2228 746 2300 978
rect 2481 935 2573 1069
rect 3204 1121 3296 1161
rect 3204 1069 3224 1121
rect 3276 1069 3296 1121
rect 2481 883 2501 935
rect 2553 883 2573 935
rect 2481 842 2573 883
rect 2762 746 2834 978
rect 2950 858 3023 978
rect 2951 746 3023 858
rect 3204 935 3296 1069
rect 3929 1121 4021 1161
rect 3929 1069 3949 1121
rect 4001 1069 4021 1121
rect 3204 883 3224 935
rect 3276 883 3296 935
rect 3204 842 3296 883
rect 3438 858 3571 978
rect 2228 735 2641 746
rect 2228 689 2584 735
rect 2630 689 2641 735
rect 2228 678 2641 689
rect 2762 735 2872 746
rect 2762 689 2815 735
rect 2861 689 2872 735
rect 2762 678 2872 689
rect 2951 735 3365 746
rect 2951 689 3308 735
rect 3354 689 3365 735
rect 2951 678 3365 689
rect 3503 735 3571 858
rect 3503 689 3514 735
rect 3560 689 3571 735
rect 2228 355 2300 678
rect 2762 355 2834 678
rect 2951 347 3023 678
rect 3503 536 3571 689
rect 3459 347 3571 536
rect -367 305 -252 342
rect 3715 334 3761 1004
rect 3929 935 4021 1069
rect 3929 883 3949 935
rect 4001 883 4021 935
rect 3929 842 4021 883
rect 4153 1121 4245 1161
rect 4153 1069 4173 1121
rect 4225 1069 4245 1121
rect 4153 935 4245 1069
rect 4153 883 4173 935
rect 4225 883 4245 935
rect 4153 842 4245 883
rect 4377 1053 4469 1093
rect 4377 1001 4397 1053
rect 4449 1001 4469 1053
rect 4377 867 4469 1001
rect 4726 1088 5026 1139
rect 4726 1042 4774 1088
rect 4820 1042 4932 1088
rect 4978 1042 5026 1088
rect 4726 992 5026 1042
rect 4909 991 4924 992
rect 4377 815 4397 867
rect 4449 815 4469 867
rect 4377 774 4469 815
rect 3979 694 4287 713
rect 3979 693 4207 694
rect 3979 641 4009 693
rect 4061 641 4195 693
rect 4253 648 4287 694
rect 4247 641 4287 648
rect 3979 621 4287 641
rect 4400 205 4446 774
<< via1 >>
rect 2313 4759 2365 4811
rect 2493 4759 2545 4811
rect 2073 4561 2087 4576
rect 2087 4561 2125 4576
rect 2073 4524 2125 4561
rect 2073 4338 2125 4390
rect 881 3948 933 4000
rect 1061 3948 1113 4000
rect 2816 3788 2868 3796
rect 2816 3744 2868 3788
rect 2996 3744 3048 3796
rect 2330 2690 2382 2718
rect 2330 2666 2382 2690
rect 2219 2433 2271 2449
rect 2219 2397 2263 2433
rect 2263 2397 2271 2433
rect 2399 2397 2451 2449
rect 3121 2397 3173 2449
rect 3301 2403 3332 2449
rect 3332 2403 3353 2449
rect 3301 2397 3353 2403
rect 4611 1734 4663 1786
rect 4823 1734 4875 1786
rect 112 1516 164 1568
rect 324 1516 376 1568
rect 890 1532 942 1584
rect 1076 1532 1128 1584
rect 4191 1532 4243 1584
rect 4377 1532 4429 1584
rect 4611 1516 4663 1568
rect 4823 1516 4875 1568
rect 112 1298 164 1350
rect 324 1336 376 1350
rect 324 1298 366 1336
rect 366 1298 376 1336
rect 4611 1298 4663 1350
rect 4823 1298 4875 1350
rect 92 1069 144 1121
rect 512 1069 564 1121
rect 92 883 144 935
rect 984 1069 1036 1121
rect 512 883 564 935
rect 1459 1080 1511 1132
rect 1639 1080 1691 1132
rect 1840 1069 1892 1121
rect 984 883 1036 935
rect 2501 1069 2553 1121
rect 1840 883 1892 935
rect 1524 734 1576 786
rect 1524 548 1576 600
rect 3224 1069 3276 1121
rect 2501 883 2553 935
rect 3949 1069 4001 1121
rect 3224 883 3276 935
rect 3949 883 4001 935
rect 4173 1069 4225 1121
rect 4173 883 4225 935
rect 4397 1001 4449 1053
rect 4397 815 4449 867
rect 4009 641 4061 693
rect 4195 648 4207 693
rect 4207 648 4247 693
rect 4195 641 4247 648
<< metal2 >>
rect 2275 4833 2364 4834
rect 2275 4811 2583 4833
rect 2275 4759 2313 4811
rect 2365 4759 2493 4811
rect 2545 4759 2583 4811
rect 2275 4737 2583 4759
rect 2053 4576 2146 4616
rect 2053 4524 2073 4576
rect 2125 4524 2146 4576
rect 2053 4390 2146 4524
rect 2053 4338 2073 4390
rect 2125 4338 2146 4390
rect 860 4000 1134 4040
rect 860 3948 881 4000
rect 933 3948 1061 4000
rect 1113 3948 1134 4000
rect 860 3907 1134 3948
rect 199 1608 294 1609
rect 74 1570 414 1608
rect 74 1514 110 1570
rect 166 1514 322 1570
rect 378 1514 414 1570
rect 74 1352 414 1514
rect 860 1604 954 3907
rect 2053 3805 2146 4338
rect 2275 3997 2364 4737
rect 2275 3905 2867 3997
rect 2777 3818 2867 3905
rect 2053 3708 2685 3805
rect 2777 3796 3086 3818
rect 2777 3744 2816 3796
rect 2868 3744 2996 3796
rect 3048 3744 3086 3796
rect 2777 3722 3086 3744
rect 2777 3721 2867 3722
rect 2590 3707 2685 3708
rect 2295 2738 2422 2739
rect 2189 2720 2497 2738
rect 2189 2664 2217 2720
rect 2273 2718 2403 2720
rect 2273 2666 2330 2718
rect 2382 2666 2403 2718
rect 2273 2664 2403 2666
rect 2459 2664 2497 2720
rect 2189 2646 2497 2664
rect 2591 2472 2685 3707
rect 1635 2471 3280 2472
rect 1635 2449 3391 2471
rect 1635 2397 2219 2449
rect 2271 2397 2399 2449
rect 2451 2397 3121 2449
rect 3173 2397 3301 2449
rect 3353 2397 3391 2449
rect 1635 2375 3391 2397
rect 860 1584 1168 1604
rect 860 1532 890 1584
rect 942 1532 1076 1584
rect 1128 1532 1168 1584
rect 860 1512 1168 1532
rect 860 1511 954 1512
rect 74 1296 110 1352
rect 166 1296 322 1352
rect 378 1296 414 1352
rect 74 1257 414 1296
rect 72 1150 164 1161
rect 492 1150 584 1161
rect 964 1150 1056 1161
rect 1421 1154 1510 1155
rect 1635 1154 1729 2375
rect 4574 1788 4955 1826
rect 4574 1732 4609 1788
rect 4665 1732 4821 1788
rect 4877 1732 4955 1788
rect 4376 1604 4470 1608
rect 4161 1584 4470 1604
rect 4161 1532 4191 1584
rect 4243 1532 4377 1584
rect 4429 1532 4470 1584
rect 4161 1512 4470 1532
rect 72 1121 165 1150
rect 72 1112 92 1121
rect 144 1112 165 1121
rect 72 1056 90 1112
rect 146 1056 165 1112
rect 72 935 165 1056
rect 72 926 92 935
rect 144 926 165 935
rect 72 870 90 926
rect 146 870 165 926
rect 72 831 165 870
rect 492 1121 585 1150
rect 492 1112 512 1121
rect 564 1112 585 1121
rect 492 1056 510 1112
rect 566 1056 585 1112
rect 492 935 585 1056
rect 492 926 512 935
rect 564 926 585 935
rect 492 870 510 926
rect 566 870 585 926
rect 492 831 585 870
rect 964 1121 1057 1150
rect 964 1112 984 1121
rect 1036 1112 1057 1121
rect 964 1056 982 1112
rect 1038 1056 1057 1112
rect 1421 1132 1729 1154
rect 1421 1080 1459 1132
rect 1511 1080 1639 1132
rect 1691 1080 1729 1132
rect 1421 1058 1729 1080
rect 1820 1150 1912 1161
rect 2481 1150 2573 1161
rect 3204 1150 3296 1161
rect 3929 1150 4021 1161
rect 4153 1150 4245 1161
rect 1820 1121 1913 1150
rect 1820 1112 1840 1121
rect 1892 1112 1913 1121
rect 964 935 1057 1056
rect 964 926 984 935
rect 1036 926 1057 935
rect 964 870 982 926
rect 1038 870 1057 926
rect 964 831 1057 870
rect 1820 1056 1838 1112
rect 1894 1056 1913 1112
rect 1820 935 1913 1056
rect 1820 926 1840 935
rect 1892 926 1913 935
rect 1820 870 1838 926
rect 1894 870 1913 926
rect 1820 831 1913 870
rect 2481 1121 2574 1150
rect 2481 1112 2501 1121
rect 2553 1112 2574 1121
rect 2481 1056 2499 1112
rect 2555 1056 2574 1112
rect 2481 935 2574 1056
rect 2481 926 2501 935
rect 2553 926 2574 935
rect 2481 870 2499 926
rect 2555 870 2574 926
rect 2481 831 2574 870
rect 3204 1121 3297 1150
rect 3204 1112 3224 1121
rect 3276 1112 3297 1121
rect 3204 1056 3222 1112
rect 3278 1056 3297 1112
rect 3204 935 3297 1056
rect 3204 926 3224 935
rect 3276 926 3297 935
rect 3204 870 3222 926
rect 3278 870 3297 926
rect 3204 831 3297 870
rect 3929 1121 4022 1150
rect 3929 1112 3949 1121
rect 4001 1112 4022 1121
rect 3929 1056 3947 1112
rect 4003 1056 4022 1112
rect 3929 935 4022 1056
rect 3929 926 3949 935
rect 4001 926 4022 935
rect 3929 870 3947 926
rect 4003 870 4022 926
rect 3929 831 4022 870
rect 4153 1121 4246 1150
rect 4153 1112 4173 1121
rect 4225 1112 4246 1121
rect 4153 1056 4171 1112
rect 4227 1056 4246 1112
rect 4153 935 4246 1056
rect 4153 926 4173 935
rect 4225 926 4246 935
rect 4153 870 4171 926
rect 4227 870 4246 926
rect 4153 831 4246 870
rect 4376 1053 4470 1512
rect 4574 1570 4955 1732
rect 4574 1514 4609 1570
rect 4665 1514 4821 1570
rect 4877 1514 4955 1570
rect 4574 1352 4955 1514
rect 4574 1296 4609 1352
rect 4665 1296 4821 1352
rect 4877 1296 4955 1352
rect 4574 1257 4955 1296
rect 4376 1001 4397 1053
rect 4449 1001 4470 1053
rect 4376 867 4470 1001
rect 1504 786 1596 826
rect 1504 734 1524 786
rect 1576 734 1596 786
rect 4376 815 4397 867
rect 4449 815 4470 867
rect 4376 777 4470 815
rect 4377 775 4469 777
rect 1504 717 1596 734
rect 1504 713 3989 717
rect 1504 693 4287 713
rect 1504 641 4009 693
rect 4061 641 4195 693
rect 4247 641 4287 693
rect 1504 621 4287 641
rect 1504 620 3989 621
rect 1504 600 1596 620
rect 1504 548 1524 600
rect 1576 548 1596 600
rect 1504 508 1596 548
<< via2 >>
rect 110 1568 166 1570
rect 110 1516 112 1568
rect 112 1516 164 1568
rect 164 1516 166 1568
rect 110 1514 166 1516
rect 322 1568 378 1570
rect 322 1516 324 1568
rect 324 1516 376 1568
rect 376 1516 378 1568
rect 322 1514 378 1516
rect 2217 2664 2273 2720
rect 2403 2664 2459 2720
rect 110 1350 166 1352
rect 110 1298 112 1350
rect 112 1298 164 1350
rect 164 1298 166 1350
rect 110 1296 166 1298
rect 322 1350 378 1352
rect 322 1298 324 1350
rect 324 1298 376 1350
rect 376 1298 378 1350
rect 322 1296 378 1298
rect 4609 1786 4665 1788
rect 4609 1734 4611 1786
rect 4611 1734 4663 1786
rect 4663 1734 4665 1786
rect 4609 1732 4665 1734
rect 4821 1786 4877 1788
rect 4821 1734 4823 1786
rect 4823 1734 4875 1786
rect 4875 1734 4877 1786
rect 4821 1732 4877 1734
rect 90 1069 92 1112
rect 92 1069 144 1112
rect 144 1069 146 1112
rect 90 1056 146 1069
rect 90 883 92 926
rect 92 883 144 926
rect 144 883 146 926
rect 90 870 146 883
rect 510 1069 512 1112
rect 512 1069 564 1112
rect 564 1069 566 1112
rect 510 1056 566 1069
rect 510 883 512 926
rect 512 883 564 926
rect 564 883 566 926
rect 510 870 566 883
rect 982 1069 984 1112
rect 984 1069 1036 1112
rect 1036 1069 1038 1112
rect 982 1056 1038 1069
rect 982 883 984 926
rect 984 883 1036 926
rect 1036 883 1038 926
rect 982 870 1038 883
rect 1838 1069 1840 1112
rect 1840 1069 1892 1112
rect 1892 1069 1894 1112
rect 1838 1056 1894 1069
rect 1838 883 1840 926
rect 1840 883 1892 926
rect 1892 883 1894 926
rect 1838 870 1894 883
rect 2499 1069 2501 1112
rect 2501 1069 2553 1112
rect 2553 1069 2555 1112
rect 2499 1056 2555 1069
rect 2499 883 2501 926
rect 2501 883 2553 926
rect 2553 883 2555 926
rect 2499 870 2555 883
rect 3222 1069 3224 1112
rect 3224 1069 3276 1112
rect 3276 1069 3278 1112
rect 3222 1056 3278 1069
rect 3222 883 3224 926
rect 3224 883 3276 926
rect 3276 883 3278 926
rect 3222 870 3278 883
rect 3947 1069 3949 1112
rect 3949 1069 4001 1112
rect 4001 1069 4003 1112
rect 3947 1056 4003 1069
rect 3947 883 3949 926
rect 3949 883 4001 926
rect 4001 883 4003 926
rect 3947 870 4003 883
rect 4171 1069 4173 1112
rect 4173 1069 4225 1112
rect 4225 1069 4227 1112
rect 4171 1056 4227 1069
rect 4171 883 4173 926
rect 4173 883 4225 926
rect 4225 883 4227 926
rect 4171 870 4227 883
rect 4609 1568 4665 1570
rect 4609 1516 4611 1568
rect 4611 1516 4663 1568
rect 4663 1516 4665 1568
rect 4609 1514 4665 1516
rect 4821 1568 4877 1570
rect 4821 1516 4823 1568
rect 4823 1516 4875 1568
rect 4875 1516 4877 1568
rect 4821 1514 4877 1516
rect 4609 1350 4665 1352
rect 4609 1298 4611 1350
rect 4611 1298 4663 1350
rect 4663 1298 4665 1350
rect 4609 1296 4665 1298
rect 4821 1350 4877 1352
rect 4821 1298 4823 1350
rect 4823 1298 4875 1350
rect 4875 1298 4877 1350
rect 4821 1296 4877 1298
<< metal3 >>
rect -358 5127 5125 5655
rect -361 3105 5001 4467
rect 3875 2741 3970 2742
rect 4326 2741 4419 2742
rect 2189 2720 4419 2741
rect 2189 2664 2217 2720
rect 2273 2664 2403 2720
rect 2459 2664 4419 2720
rect 2189 2645 4419 2664
rect -361 1933 5001 2547
rect -374 1788 5025 1826
rect -374 1732 4609 1788
rect 4665 1732 4821 1788
rect 4877 1732 5025 1788
rect -374 1570 5025 1732
rect -374 1514 110 1570
rect 166 1514 322 1570
rect 378 1514 4609 1570
rect 4665 1514 4821 1570
rect 4877 1514 5025 1570
rect -374 1352 5025 1514
rect -374 1296 110 1352
rect 166 1296 322 1352
rect 378 1296 4609 1352
rect 4665 1296 4821 1352
rect 4877 1296 5025 1352
rect -374 1257 5025 1296
rect -361 1112 5001 1150
rect -361 1056 90 1112
rect 146 1056 510 1112
rect 566 1056 982 1112
rect 1038 1056 1838 1112
rect 1894 1056 2499 1112
rect 2555 1056 3222 1112
rect 3278 1056 3947 1112
rect 4003 1056 4171 1112
rect 4227 1056 5001 1112
rect -361 926 5001 1056
rect -361 870 90 926
rect 146 870 510 926
rect 566 870 982 926
rect 1038 870 1838 926
rect 1894 870 2499 926
rect 2555 870 3222 926
rect 3278 870 3947 926
rect 4003 870 4171 926
rect 4227 870 5001 926
rect -361 718 5001 870
rect -361 126 5021 581
use M1_NWELL$$44998700_256x8m81  M1_NWELL$$44998700_256x8m81_0
timestamp 1669390400
transform 1 0 -310 0 -1 365
box 0 0 1 1
use M1_NWELL$$44999724_256x8m81  M1_NWELL$$44999724_256x8m81_0
timestamp 1669390400
transform 1 0 4876 0 1 3328
box -300 -636 300 636
use M1_NWELL$$45000748_256x8m81  M1_NWELL$$45000748_256x8m81_0
timestamp 1669390400
transform 1 0 -310 0 1 3328
box -220 -636 221 636
use M1_PACTIVE4310590878130_256x8m81  M1_PACTIVE4310590878130_256x8m81_0
timestamp 1669390400
transform 1 0 -310 0 1 5375
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1669390400
transform 1 0 984 0 1 1313
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1669390400
transform 1 0 343 0 1 1313
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1669390400
transform 1 0 321 0 1 4049
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1669390400
transform 1 0 758 0 1 4865
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_0
timestamp 1669390400
transform 1 0 2110 0 1 4502
box 0 0 1 1
use M1_POLY2$$45109292_256x8m81  M1_POLY2$$45109292_256x8m81_0
timestamp 1669390400
transform 1 0 2962 0 1 4765
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1669390400
transform 1 0 3610 0 1 2609
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_1
timestamp 1669390400
transform 1 0 2607 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_2
timestamp 1669390400
transform 1 0 2838 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_3
timestamp 1669390400
transform 1 0 3331 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_4
timestamp 1669390400
transform 1 0 3537 0 1 712
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_5
timestamp 1669390400
transform 1 0 4230 0 1 671
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_6
timestamp 1669390400
transform 1 0 3355 0 1 2426
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_7
timestamp 1669390400
transform 1 0 1882 0 1 773
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_8
timestamp 1669390400
transform 1 0 2071 0 1 773
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_9
timestamp 1669390400
transform 1 0 1347 0 1 714
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_10
timestamp 1669390400
transform 1 0 2240 0 1 2410
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1669390400
transform 1 0 2885 0 1 3765
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_1
timestamp 1669390400
transform 1 0 2388 0 1 2667
box 0 0 1 1
use M1_PSUB$$44997676_256x8m81  M1_PSUB$$44997676_256x8m81_0
timestamp 1669390400
transform 1 0 4797 0 -1 2086
box 0 0 1 1
use M1_PSUB$$44997676_256x8m81  M1_PSUB$$44997676_256x8m81_1
timestamp 1669390400
transform 1 0 -152 0 -1 2086
box 0 0 1 1
use M1_PSUB$$45110316_285_256x8m81  M1_PSUB$$45110316_285_256x8m81_0
timestamp 1669390400
transform 1 0 4876 0 -1 1065
box 0 0 1 1
use M1_PSUB$$45110316_285_256x8m81  M1_PSUB$$45110316_285_256x8m81_1
timestamp 1669390400
transform 1 0 -310 0 -1 1065
box 0 0 1 1
use M2_M1$$43374636_256x8m81  M2_M1$$43374636_256x8m81_0
timestamp 1669390400
transform 1 0 244 0 1 1433
box 0 0 1 1
use M2_M1$$45002796_256x8m81  M2_M1$$45002796_256x8m81_0
timestamp 1669390400
transform 1 0 3063 0 1 1324
box -1119 -67 1119 66
use M2_M1$$45003820_256x8m81  M2_M1$$45003820_256x8m81_0
timestamp 1669390400
transform 1 0 4743 0 1 1542
box 0 0 1 1
use M2_M1c$$203396140_256x8m81  M2_M1c$$203396140_256x8m81_0
timestamp 1669390400
transform 1 0 997 0 1 3974
box 0 0 1 1
use M3_M2$$45005868_256x8m81  M3_M2$$45005868_256x8m81_0
timestamp 1669390400
transform 1 0 3063 0 1 1324
box -1119 -67 1119 67
use M3_M2$$45006892_256x8m81  M3_M2$$45006892_256x8m81_0
timestamp 1669390400
transform 1 0 4743 0 1 1542
box 0 0 1 1
use M3_M2$$45008940_256x8m81  M3_M2$$45008940_256x8m81_0
timestamp 1669390400
transform 1 0 244 0 1 1433
box 0 0 1 1
use nmos_1p2$$45100076_256x8m81  nmos_1p2$$45100076_256x8m81_0
timestamp 1669390400
transform -1 0 4063 0 -1 2301
box -119 -74 401 595
use nmos_1p2$$45101100_256x8m81  nmos_1p2$$45101100_256x8m81_0
timestamp 1669390400
transform 1 0 202 0 1 855
box -119 -74 1073 300
use nmos_1p2$$45102124_256x8m81  nmos_1p2$$45102124_256x8m81_0
timestamp 1669390400
transform -1 0 1823 0 -1 2301
box -119 -74 1521 527
use nmos_1p2$$45103148_256x8m81  nmos_1p2$$45103148_256x8m81_0
timestamp 1669390400
transform -1 0 3391 0 -1 2301
box -119 -74 1297 645
use nmos_5p04310590878112_256x8m81  nmos_5p04310590878112_256x8m81_0
timestamp 1669390400
transform -1 0 4684 0 1 5006
box -88 -44 880 498
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_0
timestamp 1669390400
transform 1 0 3065 0 1 884
box -88 -44 432 164
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_1
timestamp 1669390400
transform 1 0 1616 0 1 884
box -88 -44 432 164
use nmos_5p04310590878123_256x8m81  nmos_5p04310590878123_256x8m81_2
timestamp 1669390400
transform 1 0 2341 0 1 884
box -88 -44 432 164
use nmos_5p04310590878126_256x8m81  nmos_5p04310590878126_256x8m81_0
timestamp 1669390400
transform 1 0 1074 0 1 5006
box -88 -44 1104 498
use nmos_5p04310590878126_256x8m81  nmos_5p04310590878126_256x8m81_1
timestamp 1669390400
transform 1 0 2483 0 1 5006
box -88 -44 1104 498
use nmos_5p04310590878131_256x8m81  nmos_5p04310590878131_256x8m81_0
timestamp 1669390400
transform -1 0 503 0 1 5223
box -88 -44 432 272
use nmos_5p04310590878132_256x8m81  nmos_5p04310590878132_256x8m81_0
timestamp 1669390400
transform 1 0 3790 0 1 884
box -88 -44 208 164
use nmos_5p04310590878133_256x8m81  nmos_5p04310590878133_256x8m81_0
timestamp 1669390400
transform 1 0 4251 0 1 818
box -88 -44 208 332
use pmos_1p2$$45095980_256x8m81  pmos_1p2$$45095980_256x8m81_0
timestamp 1669390400
transform -1 0 4653 0 1 4090
box -286 -142 2360 686
use pmos_1p2$$46281772_256x8m81  pmos_1p2$$46281772_256x8m81_0
timestamp 1669390400
transform -1 0 4287 0 -1 3650
box -286 -142 792 1028
use pmos_1p2$$46281772_256x8m81  pmos_1p2$$46281772_256x8m81_1
timestamp 1669390400
transform -1 0 3391 0 -1 3650
box -286 -142 792 1028
use pmos_1p2$$46282796_256x8m81  pmos_1p2$$46282796_256x8m81_0
timestamp 1669390400
transform 1 0 202 0 1 118
box -286 -142 1240 595
use pmos_1p2$$46283820_256x8m81  pmos_1p2$$46283820_256x8m81_0
timestamp 1669390400
transform -1 0 2271 0 -1 3629
box -286 -142 2360 958
use pmos_1p2$$46284844_256x8m81  pmos_1p2$$46284844_256x8m81_0
timestamp 1669390400
transform 1 0 4282 0 1 197
box -286 -142 568 482
use pmos_1p2$$46285868_256x8m81  pmos_1p2$$46285868_256x8m81_0
timestamp 1669390400
transform 1 0 1777 0 1 4198
box -286 -142 344 595
use pmos_1p2$$46286892_256x8m81  pmos_1p2$$46286892_256x8m81_0
timestamp 1669390400
transform 1 0 1105 0 1 4198
box -286 -142 792 595
use pmos_1p2$$46287916_256x8m81  pmos_1p2$$46287916_256x8m81_0
timestamp 1669390400
transform -1 0 472 0 1 4189
box -286 -142 568 822
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_0
timestamp 1669390400
transform 1 0 3065 0 1 296
box -208 -120 552 360
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_1
timestamp 1669390400
transform 1 0 1616 0 1 296
box -208 -120 552 360
use pmos_5p04310590878125_256x8m81  pmos_5p04310590878125_256x8m81_2
timestamp 1669390400
transform 1 0 2341 0 1 296
box -208 -120 552 360
use pmos_5p04310590878138_256x8m81  pmos_5p04310590878138_256x8m81_0
timestamp 1669390400
transform 1 0 3790 0 1 334
box -208 -120 328 360
use po_m1_256x8m81  po_m1_256x8m81_0
timestamp 1669390400
transform 1 0 2743 0 1 1440
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1669390400
transform -1 0 3744 0 -1 2251
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1669390400
transform 1 0 3189 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1669390400
transform 1 0 2466 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1669390400
transform -1 0 3522 0 -1 2251
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1669390400
transform 1 0 4909 0 1 830
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1669390400
transform 1 0 4909 0 1 1934
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1669390400
transform 1 0 4601 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1669390400
transform 1 0 4148 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1669390400
transform 1 0 3942 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1669390400
transform -1 0 4190 0 -1 2251
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1669390400
transform 1 0 72 0 1 194
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1669390400
transform -1 0 -264 0 -1 555
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1669390400
transform -1 0 1506 0 -1 2251
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1669390400
transform 1 0 -356 0 1 830
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1669390400
transform 1 0 -356 0 1 1934
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1669390400
transform 1 0 1741 0 1 127
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1669390400
transform 1 0 968 0 1 190
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1669390400
transform 1 0 521 0 1 192
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1669390400
transform -1 0 2174 0 -1 2251
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_19
timestamp 1669390400
transform -1 0 1950 0 -1 4409
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_20
timestamp 1669390400
transform 1 0 -356 0 1 3106
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_21
timestamp 1669390400
transform -1 0 -264 0 -1 5550
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_22
timestamp 1669390400
transform -1 0 105 0 -1 5531
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_23
timestamp 1669390400
transform -1 0 153 0 -1 4409
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_24
timestamp 1669390400
transform -1 0 1065 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_25
timestamp 1669390400
transform -1 0 1504 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_26
timestamp 1669390400
transform -1 0 1970 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_27
timestamp 1669390400
transform -1 0 601 0 -1 5531
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_28
timestamp 1669390400
transform -1 0 601 0 -1 4409
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_29
timestamp 1669390400
transform -1 0 1067 0 -1 4452
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_30
timestamp 1669390400
transform -1 0 1504 0 -1 4409
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_31
timestamp 1669390400
transform -1 0 105 0 -1 3636
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_32
timestamp 1669390400
transform -1 0 1504 0 -1 3636
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_33
timestamp 1669390400
transform 1 0 -356 0 1 3684
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_34
timestamp 1669390400
transform 1 0 4909 0 1 3106
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_35
timestamp 1669390400
transform 1 0 4909 0 1 3573
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_36
timestamp 1669390400
transform -1 0 3742 0 -1 3575
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_37
timestamp 1669390400
transform -1 0 4192 0 -1 3575
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_38
timestamp 1669390400
transform -1 0 3298 0 -1 3575
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_39
timestamp 1669390400
transform -1 0 2868 0 -1 3575
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_40
timestamp 1669390400
transform -1 0 2556 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_41
timestamp 1669390400
transform -1 0 2993 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_42
timestamp 1669390400
transform -1 0 3435 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_43
timestamp 1669390400
transform -1 0 3889 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_44
timestamp 1669390400
transform -1 0 4335 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_45
timestamp 1669390400
transform -1 0 4783 0 -1 4434
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_46
timestamp 1669390400
transform -1 0 3887 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_47
timestamp 1669390400
transform -1 0 4333 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_48
timestamp 1669390400
transform -1 0 4785 0 -1 5445
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_49
timestamp 1669390400
transform -1 0 4418 0 -1 2963
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_50
timestamp 1669390400
transform -1 0 3968 0 -1 2963
box 0 -1 93 308
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_51
timestamp 1669390400
transform -1 0 2389 0 -1 3593
box 0 -1 93 308
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1669390400
transform 0 -1 2422 1 0 2646
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1669390400
transform 1 0 4377 0 1 775
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1669390400
transform 1 0 2481 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1669390400
transform 1 0 3204 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1669390400
transform 1 0 3929 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1669390400
transform 1 0 4153 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_5
timestamp 1669390400
transform 1 0 1504 0 1 508
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_6
timestamp 1669390400
transform 1 0 1820 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_7
timestamp 1669390400
transform 1 0 72 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_8
timestamp 1669390400
transform 1 0 492 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_9
timestamp 1669390400
transform 1 0 964 0 1 843
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_10
timestamp 1669390400
transform -1 0 2145 0 -1 4616
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1669390400
transform 0 -1 4469 1 0 1512
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1669390400
transform 0 -1 4287 1 0 621
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1669390400
transform 0 -1 1168 1 0 1512
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_0
timestamp 1669390400
transform 0 1 3083 -1 0 2471
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_1
timestamp 1669390400
transform 0 1 1421 -1 0 1154
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_2
timestamp 1669390400
transform 0 1 2778 -1 0 3818
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_3
timestamp 1669390400
transform 0 1 2181 -1 0 2471
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_4
timestamp 1669390400
transform 0 1 2275 -1 0 4833
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_0
timestamp 1669390400
transform 1 0 3204 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_1
timestamp 1669390400
transform 1 0 2481 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_2
timestamp 1669390400
transform 1 0 3929 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_3
timestamp 1669390400
transform 1 0 4153 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_4
timestamp 1669390400
transform 1 0 964 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_5
timestamp 1669390400
transform 1 0 492 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_6
timestamp 1669390400
transform 1 0 72 0 1 832
box 0 0 1 1
use via2_x2_256x8m81  via2_x2_256x8m81_7
timestamp 1669390400
transform 1 0 1820 0 1 832
box 0 0 1 1
use via2_x2_R90_256x8m81  via2_x2_R90_256x8m81_0
timestamp 1669390400
transform 0 -1 2497 1 0 2646
box 0 0 1 1
<< labels >>
rlabel metal1 s 1456 2584 1456 2584 4 pcb
port 1 nsew
rlabel metal1 s 4066 5565 4066 5565 4 se
port 2 nsew
rlabel metal3 s 2398 3802 2398 3802 4 vdd
port 3 nsew
rlabel metal3 s 2163 5443 2163 5443 4 vss
port 4 nsew
rlabel metal3 s 2288 1061 2288 1061 4 vss
port 4 nsew
rlabel metal3 s 248 1437 248 1437 4 men
port 5 nsew
rlabel metal3 s 2288 2151 2288 2151 4 vss
port 4 nsew
rlabel metal3 s 1489 379 1489 379 4 vdd
port 3 nsew
<< properties >>
string GDS_END 495216
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 476246
string path 20.320 27.120 20.320 27.785 22.565 27.785 22.565 26.905 
<< end >>
