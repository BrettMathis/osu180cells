magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 377 5014 870
rect -86 352 1249 377
rect 2000 352 5014 377
<< pwell >>
rect 1249 352 2000 377
rect -86 -86 5014 352
<< mvnmos >>
rect 124 156 244 228
rect 348 156 468 228
rect 516 156 636 228
rect 740 156 860 228
rect 908 156 1028 228
rect 1168 135 1288 228
rect 1631 139 1751 232
rect 2043 158 2163 230
rect 2267 158 2387 230
rect 2435 158 2555 230
rect 2698 158 2818 230
rect 2936 158 3056 230
rect 3160 158 3280 230
rect 3420 69 3540 232
rect 3644 69 3764 232
rect 4012 69 4132 232
rect 4236 69 4356 232
rect 4460 69 4580 232
rect 4684 69 4804 232
<< mvpmos >>
rect 124 502 224 628
rect 348 502 448 628
rect 496 502 596 628
rect 700 502 800 628
rect 888 502 988 628
rect 1188 502 1288 686
rect 1651 497 1751 660
rect 2032 502 2132 628
rect 2246 502 2346 628
rect 2424 502 2524 628
rect 2716 502 2818 628
rect 2950 502 3050 628
rect 3164 502 3264 628
rect 3404 472 3504 715
rect 3644 472 3744 715
rect 4032 472 4132 715
rect 4246 472 4346 715
rect 4480 472 4580 715
rect 4694 472 4794 715
<< mvndiff >>
rect 1348 244 1424 257
rect 1348 228 1361 244
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 228
rect 636 215 740 228
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 228
rect 1028 215 1168 228
rect 1028 169 1070 215
rect 1116 169 1168 215
rect 1028 156 1168 169
rect 1088 135 1168 156
rect 1288 198 1361 228
rect 1407 198 1424 244
rect 1811 244 1883 257
rect 1811 232 1824 244
rect 1288 135 1424 198
rect 1543 198 1631 232
rect 1543 152 1556 198
rect 1602 152 1631 198
rect 1543 139 1631 152
rect 1751 198 1824 232
rect 1870 198 1883 244
rect 3340 230 3420 232
rect 1751 139 1883 198
rect 1955 217 2043 230
rect 1955 171 1968 217
rect 2014 171 2043 217
rect 1955 158 2043 171
rect 2163 217 2267 230
rect 2163 171 2192 217
rect 2238 171 2267 217
rect 2163 158 2267 171
rect 2387 158 2435 230
rect 2555 217 2698 230
rect 2555 171 2607 217
rect 2653 171 2698 217
rect 2555 158 2698 171
rect 2818 217 2936 230
rect 2818 171 2857 217
rect 2903 171 2936 217
rect 2818 158 2936 171
rect 3056 217 3160 230
rect 3056 171 3085 217
rect 3131 171 3160 217
rect 3056 158 3160 171
rect 3280 158 3420 230
rect 3340 69 3420 158
rect 3540 128 3644 232
rect 3540 82 3569 128
rect 3615 82 3644 128
rect 3540 69 3644 82
rect 3764 172 3852 232
rect 3764 126 3793 172
rect 3839 126 3852 172
rect 3764 69 3852 126
rect 3924 171 4012 232
rect 3924 125 3937 171
rect 3983 125 4012 171
rect 3924 69 4012 125
rect 4132 188 4236 232
rect 4132 142 4161 188
rect 4207 142 4236 188
rect 4132 69 4236 142
rect 4356 171 4460 232
rect 4356 125 4385 171
rect 4431 125 4460 171
rect 4356 69 4460 125
rect 4580 188 4684 232
rect 4580 142 4609 188
rect 4655 142 4684 188
rect 4580 69 4684 142
rect 4804 171 4892 232
rect 4804 125 4833 171
rect 4879 125 4892 171
rect 4804 69 4892 125
<< mvpdiff >>
rect 1048 686 1120 701
rect 1512 716 1586 729
rect 1048 682 1188 686
rect 1048 636 1061 682
rect 1107 636 1188 682
rect 1048 628 1188 636
rect 36 590 124 628
rect 36 544 49 590
rect 95 544 124 590
rect 36 502 124 544
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 502 348 569
rect 448 502 496 628
rect 596 587 700 628
rect 596 541 625 587
rect 671 541 700 587
rect 596 502 700 541
rect 800 502 888 628
rect 988 502 1188 628
rect 1288 561 1376 686
rect 1288 515 1317 561
rect 1363 515 1376 561
rect 1288 502 1376 515
rect 1512 670 1525 716
rect 1571 670 1586 716
rect 1512 660 1586 670
rect 1512 497 1651 660
rect 1751 561 1839 660
rect 2584 645 2656 658
rect 2584 628 2597 645
rect 1751 515 1780 561
rect 1826 515 1839 561
rect 1751 497 1839 515
rect 1944 595 2032 628
rect 1944 549 1957 595
rect 2003 549 2032 595
rect 1944 502 2032 549
rect 2132 563 2246 628
rect 2132 517 2171 563
rect 2217 517 2246 563
rect 2132 502 2246 517
rect 2346 502 2424 628
rect 2524 599 2597 628
rect 2643 628 2656 645
rect 3324 628 3404 715
rect 2643 599 2716 628
rect 2524 502 2716 599
rect 2818 563 2950 628
rect 2818 517 2865 563
rect 2911 517 2950 563
rect 2818 502 2950 517
rect 3050 563 3164 628
rect 3050 517 3089 563
rect 3135 517 3164 563
rect 3050 502 3164 517
rect 3264 502 3404 628
rect 3324 472 3404 502
rect 3504 702 3644 715
rect 3504 562 3553 702
rect 3599 562 3644 702
rect 3504 472 3644 562
rect 3744 658 3852 715
rect 3744 612 3793 658
rect 3839 612 3852 658
rect 3744 547 3852 612
rect 3744 501 3793 547
rect 3839 501 3852 547
rect 3744 472 3852 501
rect 3944 679 4032 715
rect 3944 633 3957 679
rect 4003 633 4032 679
rect 3944 560 4032 633
rect 3944 514 3957 560
rect 4003 514 4032 560
rect 3944 472 4032 514
rect 4132 662 4246 715
rect 4132 616 4171 662
rect 4217 616 4246 662
rect 4132 557 4246 616
rect 4132 511 4171 557
rect 4217 511 4246 557
rect 4132 472 4246 511
rect 4346 679 4480 715
rect 4346 633 4389 679
rect 4435 633 4480 679
rect 4346 560 4480 633
rect 4346 514 4389 560
rect 4435 514 4480 560
rect 4346 472 4480 514
rect 4580 662 4694 715
rect 4580 616 4614 662
rect 4660 616 4694 662
rect 4580 557 4694 616
rect 4580 511 4614 557
rect 4660 511 4694 557
rect 4580 472 4694 511
rect 4794 679 4882 715
rect 4794 633 4823 679
rect 4869 633 4882 679
rect 4794 560 4882 633
rect 4794 514 4823 560
rect 4869 514 4882 560
rect 4794 472 4882 514
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1070 169 1116 215
rect 1361 198 1407 244
rect 1556 152 1602 198
rect 1824 198 1870 244
rect 1968 171 2014 217
rect 2192 171 2238 217
rect 2607 171 2653 217
rect 2857 171 2903 217
rect 3085 171 3131 217
rect 3569 82 3615 128
rect 3793 126 3839 172
rect 3937 125 3983 171
rect 4161 142 4207 188
rect 4385 125 4431 171
rect 4609 142 4655 188
rect 4833 125 4879 171
<< mvpdiffc >>
rect 1061 636 1107 682
rect 49 544 95 590
rect 263 569 309 615
rect 625 541 671 587
rect 1317 515 1363 561
rect 1525 670 1571 716
rect 1780 515 1826 561
rect 1957 549 2003 595
rect 2171 517 2217 563
rect 2597 599 2643 645
rect 2865 517 2911 563
rect 3089 517 3135 563
rect 3553 562 3599 702
rect 3793 612 3839 658
rect 3793 501 3839 547
rect 3957 633 4003 679
rect 3957 514 4003 560
rect 4171 616 4217 662
rect 4171 511 4217 557
rect 4389 633 4435 679
rect 4389 514 4435 560
rect 4614 616 4660 662
rect 4614 511 4660 557
rect 4823 633 4869 679
rect 4823 514 4869 560
<< polysilicon >>
rect 124 720 800 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 700 628 800 720
rect 888 628 988 692
rect 1188 686 1288 730
rect 1651 720 3050 760
rect 1651 660 1751 720
rect 124 432 224 502
rect 124 351 244 432
rect 124 305 150 351
rect 196 305 244 351
rect 124 228 244 305
rect 348 351 448 502
rect 348 305 374 351
rect 420 305 448 351
rect 496 403 596 502
rect 700 458 800 502
rect 888 458 988 502
rect 496 357 509 403
rect 555 371 596 403
rect 908 434 988 458
rect 1188 442 1288 502
rect 2032 628 2132 672
rect 2246 628 2346 720
rect 2424 628 2524 672
rect 2716 628 2818 672
rect 2950 628 3050 720
rect 3404 715 3504 759
rect 3644 715 3744 759
rect 4032 715 4132 759
rect 4246 715 4346 759
rect 4480 715 4580 759
rect 4694 715 4794 759
rect 3164 628 3264 672
rect 908 388 926 434
rect 972 388 988 434
rect 555 357 860 371
rect 496 325 860 357
rect 348 272 448 305
rect 348 228 468 272
rect 516 228 636 272
rect 740 228 860 325
rect 908 272 988 388
rect 1168 424 1288 442
rect 1651 432 1751 497
rect 1651 427 1674 432
rect 1168 378 1209 424
rect 1255 378 1288 424
rect 908 228 1028 272
rect 1168 228 1288 378
rect 1631 386 1674 427
rect 1720 386 1751 432
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1631 232 1751 386
rect 2032 451 2132 502
rect 2246 458 2346 502
rect 2424 460 2524 502
rect 2032 405 2065 451
rect 2111 405 2132 451
rect 2032 389 2132 405
rect 2424 414 2455 460
rect 2501 442 2524 460
rect 2501 414 2555 442
rect 2032 343 2352 389
rect 2424 386 2555 414
rect 2267 292 2352 343
rect 2043 230 2163 274
rect 2267 230 2387 292
rect 2435 230 2555 386
rect 2716 340 2818 502
rect 2950 442 3050 502
rect 3164 469 3264 502
rect 2950 402 3109 442
rect 3164 423 3192 469
rect 3238 423 3264 469
rect 3404 428 3504 472
rect 3164 410 3264 423
rect 2716 294 2736 340
rect 2782 294 2818 340
rect 3068 362 3109 402
rect 3420 405 3504 428
rect 3068 322 3220 362
rect 2716 276 2818 294
rect 2698 230 2818 276
rect 2936 309 3016 322
rect 2936 263 2957 309
rect 3003 274 3016 309
rect 3160 274 3220 322
rect 3003 263 3056 274
rect 2936 230 3056 263
rect 3160 230 3280 274
rect 3420 265 3442 405
rect 3488 276 3504 405
rect 3644 439 3744 472
rect 3644 299 3669 439
rect 3715 299 3744 439
rect 3644 276 3744 299
rect 4032 406 4132 472
rect 4032 276 4053 406
rect 3488 265 3540 276
rect 3420 232 3540 265
rect 3644 232 3764 276
rect 4012 266 4053 276
rect 4099 396 4132 406
rect 4246 396 4346 472
rect 4480 396 4580 472
rect 4694 396 4794 472
rect 4099 343 4794 396
rect 4099 266 4132 343
rect 4012 232 4132 266
rect 4236 276 4346 343
rect 4480 276 4580 343
rect 4236 232 4356 276
rect 4460 232 4580 276
rect 4684 276 4794 343
rect 4684 232 4804 276
rect 1168 91 1288 135
rect 124 24 636 64
rect 1631 70 1751 139
rect 2043 70 2163 158
rect 2267 114 2387 158
rect 2435 114 2555 158
rect 2698 114 2818 158
rect 2936 107 3056 158
rect 3160 114 3280 158
rect 1631 24 2163 70
rect 3420 25 3540 69
rect 3644 25 3764 69
rect 4012 25 4132 69
rect 4236 25 4356 69
rect 4460 25 4580 69
rect 4684 25 4804 69
<< polycontact >>
rect 150 305 196 351
rect 374 305 420 351
rect 509 357 555 403
rect 926 388 972 434
rect 1209 378 1255 424
rect 1674 386 1720 432
rect 2065 405 2111 451
rect 2455 414 2501 460
rect 3192 423 3238 469
rect 2736 294 2782 340
rect 2957 263 3003 309
rect 3442 265 3488 405
rect 3669 299 3715 439
rect 4053 266 4099 406
<< metal1 >>
rect 0 724 4928 844
rect 252 615 320 724
rect 1050 682 1118 724
rect 1050 636 1061 682
rect 1107 636 1118 682
rect 1514 716 1582 724
rect 1514 670 1525 716
rect 1571 670 1582 716
rect 49 590 95 603
rect 252 569 263 615
rect 309 569 320 615
rect 1175 624 1464 664
rect 1674 624 2003 670
rect 1175 618 1720 624
rect 1175 587 1221 618
rect 49 523 95 544
rect 606 541 625 587
rect 671 541 1221 587
rect 1418 578 1720 618
rect 1957 595 2003 624
rect 1317 561 1363 572
rect 49 477 555 523
rect 1780 561 1826 572
rect 1363 515 1720 532
rect 1317 486 1720 515
rect 49 215 95 477
rect 49 158 95 169
rect 141 351 206 431
rect 141 305 150 351
rect 196 305 206 351
rect 141 120 206 305
rect 365 351 430 431
rect 365 305 374 351
rect 420 305 430 351
rect 509 403 555 477
rect 682 434 1036 443
rect 682 388 926 434
rect 972 388 1036 434
rect 682 359 1036 388
rect 1093 424 1326 438
rect 1093 378 1209 424
rect 1255 378 1326 424
rect 1093 359 1326 378
rect 509 325 555 357
rect 273 215 319 228
rect 273 60 319 169
rect 365 120 430 305
rect 885 261 1252 307
rect 885 215 931 261
rect 654 169 665 215
rect 711 169 931 215
rect 1059 169 1070 215
rect 1116 169 1127 215
rect 1059 60 1127 169
rect 1206 152 1252 261
rect 1372 255 1418 486
rect 1674 432 1720 486
rect 1674 375 1720 386
rect 1957 538 2003 549
rect 2065 630 2498 678
rect 1780 410 1826 515
rect 2065 451 2111 630
rect 1780 405 2065 410
rect 1780 364 2111 405
rect 2171 563 2217 574
rect 1350 244 1418 255
rect 1350 198 1361 244
rect 1407 198 1418 244
rect 1464 261 1721 307
rect 1464 152 1510 261
rect 1206 106 1510 152
rect 1556 198 1602 209
rect 1556 60 1602 152
rect 1675 152 1721 261
rect 1813 255 1859 364
rect 2171 340 2217 517
rect 2452 553 2498 630
rect 2586 645 2654 724
rect 3542 702 3610 724
rect 2586 599 2597 645
rect 2643 599 2654 645
rect 2734 632 3249 678
rect 2734 553 2780 632
rect 2452 506 2780 553
rect 2865 563 2911 574
rect 2865 460 2911 517
rect 2440 414 2455 460
rect 2501 414 2911 460
rect 2171 294 2736 340
rect 2782 294 2793 340
rect 1813 244 1881 255
rect 1813 198 1824 244
rect 1870 198 1881 244
rect 1968 217 2014 228
rect 1968 152 2014 171
rect 2192 217 2238 294
rect 2857 217 2903 414
rect 2957 309 3003 632
rect 2957 252 3003 263
rect 3085 563 3135 574
rect 3085 517 3089 563
rect 3085 355 3135 517
rect 3181 469 3249 632
rect 3542 562 3553 702
rect 3599 562 3610 702
rect 3957 679 4003 724
rect 3542 560 3610 562
rect 3793 658 3839 669
rect 3793 547 3839 612
rect 3181 423 3192 469
rect 3238 423 3249 469
rect 3181 414 3249 423
rect 3331 463 3726 510
rect 3331 355 3377 463
rect 3658 439 3726 463
rect 3085 308 3377 355
rect 3439 405 3491 416
rect 2192 160 2238 171
rect 2596 171 2607 217
rect 2653 171 2664 217
rect 1675 106 2014 152
rect 2596 60 2664 171
rect 2857 160 2903 171
rect 3085 217 3135 308
rect 3131 171 3135 217
rect 3439 265 3442 405
rect 3488 265 3491 405
rect 3658 299 3669 439
rect 3715 299 3726 439
rect 3658 292 3726 299
rect 3793 359 3839 501
rect 4389 679 4435 724
rect 3957 560 4003 633
rect 3957 492 4003 514
rect 4152 662 4236 678
rect 4152 616 4171 662
rect 4217 616 4236 662
rect 4152 557 4236 616
rect 4152 511 4171 557
rect 4217 511 4236 557
rect 4152 432 4236 511
rect 4823 679 4869 724
rect 4389 560 4435 633
rect 4389 492 4435 514
rect 4596 662 4680 678
rect 4596 616 4614 662
rect 4660 616 4680 662
rect 4596 557 4680 616
rect 4596 511 4614 557
rect 4660 511 4680 557
rect 4596 432 4680 511
rect 4823 560 4869 633
rect 4823 492 4869 514
rect 4049 406 4103 417
rect 4049 359 4053 406
rect 3793 313 4053 359
rect 3439 246 3491 265
rect 3793 246 3839 313
rect 4049 266 4053 313
rect 4099 266 4103 406
rect 4049 255 4103 266
rect 4152 348 4680 432
rect 3439 199 3839 246
rect 3085 160 3135 171
rect 3793 172 3839 199
rect 3569 128 3615 145
rect 3793 115 3839 126
rect 3937 171 3983 190
rect 3569 60 3615 82
rect 3937 60 3983 125
rect 4152 188 4236 348
rect 4152 142 4161 188
rect 4207 142 4236 188
rect 4152 123 4236 142
rect 4385 171 4431 190
rect 4385 60 4431 125
rect 4596 188 4680 348
rect 4596 142 4609 188
rect 4655 142 4680 188
rect 4596 123 4680 142
rect 4833 171 4879 190
rect 4833 60 4879 125
rect 0 -60 4928 60
<< labels >>
flabel metal1 s 4596 432 4680 678 0 FreeSans 400 0 0 0 Q
port 5 nsew default output
flabel metal1 s 141 120 206 431 0 FreeSans 400 0 0 0 SE
port 2 nsew default input
flabel metal1 s 365 120 430 431 0 FreeSans 400 0 0 0 SI
port 3 nsew default input
flabel metal1 s 0 724 4928 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1093 359 1326 438 0 FreeSans 400 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 682 359 1036 443 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel metal1 s 273 217 319 228 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4152 432 4236 678 1 Q
port 5 nsew default output
rlabel metal1 s 4152 348 4680 432 1 Q
port 5 nsew default output
rlabel metal1 s 4596 123 4680 348 1 Q
port 5 nsew default output
rlabel metal1 s 4152 123 4236 348 1 Q
port 5 nsew default output
rlabel metal1 s 4823 670 4869 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 670 4435 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 670 4003 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3542 670 3610 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 670 2654 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1514 670 1582 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 670 1118 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4823 636 4869 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 636 4435 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 636 4003 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3542 636 3610 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 636 2654 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 636 1118 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 636 320 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4823 599 4869 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 599 4435 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 599 4003 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3542 599 3610 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 599 2654 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 599 320 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4823 569 4869 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 569 4435 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 569 4003 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3542 569 3610 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4823 560 4869 569 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 560 4435 569 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 560 4003 569 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3542 560 3610 569 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4823 492 4869 560 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4389 492 4435 560 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3957 492 4003 560 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2596 215 2664 217 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 215 319 217 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 209 2664 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 209 1127 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 209 319 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 190 2664 209 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 190 1602 209 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 190 1127 209 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 190 319 209 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4833 145 4879 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4385 145 4431 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3937 145 3983 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 145 2664 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 145 1602 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 145 1127 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 145 319 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4833 60 4879 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4385 60 4431 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3937 60 3983 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3569 60 3615 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 60 2664 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 60 1602 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 60 1127 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 145 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4928 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4928 784
string GDS_END 206642
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 196466
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
