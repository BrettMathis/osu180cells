magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -65 2202 65 2243
rect -65 2150 -26 2202
rect 26 2150 65 2202
rect -65 1985 65 2150
rect -65 1933 -26 1985
rect 26 1933 65 1985
rect -65 1767 65 1933
rect -65 1715 -26 1767
rect 26 1715 65 1767
rect -65 1549 65 1715
rect -65 1497 -26 1549
rect 26 1497 65 1549
rect -65 1332 65 1497
rect -65 1280 -26 1332
rect 26 1280 65 1332
rect -65 1114 65 1280
rect -65 1062 -26 1114
rect 26 1062 65 1114
rect -65 897 65 1062
rect -65 845 -26 897
rect 26 845 65 897
rect -65 679 65 845
rect -65 627 -26 679
rect 26 627 65 679
rect -65 461 65 627
rect -65 409 -26 461
rect 26 409 65 461
rect -65 244 65 409
rect -65 192 -26 244
rect 26 192 65 244
rect -65 26 65 192
rect -65 -26 -26 26
rect 26 -26 65 26
rect -65 -192 65 -26
rect -65 -244 -26 -192
rect 26 -244 65 -192
rect -65 -409 65 -244
rect -65 -461 -26 -409
rect 26 -461 65 -409
rect -65 -627 65 -461
rect -65 -679 -26 -627
rect 26 -679 65 -627
rect -65 -845 65 -679
rect -65 -897 -26 -845
rect 26 -897 65 -845
rect -65 -1062 65 -897
rect -65 -1114 -26 -1062
rect 26 -1114 65 -1062
rect -65 -1280 65 -1114
rect -65 -1332 -26 -1280
rect 26 -1332 65 -1280
rect -65 -1497 65 -1332
rect -65 -1549 -26 -1497
rect 26 -1549 65 -1497
rect -65 -1715 65 -1549
rect -65 -1767 -26 -1715
rect 26 -1767 65 -1715
rect -65 -1933 65 -1767
rect -65 -1985 -26 -1933
rect 26 -1985 65 -1933
rect -65 -2150 65 -1985
rect -65 -2202 -26 -2150
rect 26 -2202 65 -2150
rect -65 -2243 65 -2202
<< via1 >>
rect -26 2150 26 2202
rect -26 1933 26 1985
rect -26 1715 26 1767
rect -26 1497 26 1549
rect -26 1280 26 1332
rect -26 1062 26 1114
rect -26 845 26 897
rect -26 627 26 679
rect -26 409 26 461
rect -26 192 26 244
rect -26 -26 26 26
rect -26 -244 26 -192
rect -26 -461 26 -409
rect -26 -679 26 -627
rect -26 -897 26 -845
rect -26 -1114 26 -1062
rect -26 -1332 26 -1280
rect -26 -1549 26 -1497
rect -26 -1767 26 -1715
rect -26 -1985 26 -1933
rect -26 -2202 26 -2150
<< metal2 >>
rect -64 2202 65 2243
rect -64 2150 -26 2202
rect 26 2150 65 2202
rect -64 1985 65 2150
rect -64 1933 -26 1985
rect 26 1933 65 1985
rect -64 1767 65 1933
rect -64 1715 -26 1767
rect 26 1715 65 1767
rect -64 1549 65 1715
rect -64 1497 -26 1549
rect 26 1497 65 1549
rect -64 1332 65 1497
rect -64 1280 -26 1332
rect 26 1280 65 1332
rect -64 1114 65 1280
rect -64 1062 -26 1114
rect 26 1062 65 1114
rect -64 897 65 1062
rect -64 845 -26 897
rect 26 845 65 897
rect -64 679 65 845
rect -64 627 -26 679
rect 26 627 65 679
rect -64 461 65 627
rect -64 409 -26 461
rect 26 409 65 461
rect -64 244 65 409
rect -64 192 -26 244
rect 26 192 65 244
rect -64 26 65 192
rect -64 -26 -26 26
rect 26 -26 65 26
rect -64 -192 65 -26
rect -64 -244 -26 -192
rect 26 -244 65 -192
rect -64 -409 65 -244
rect -64 -461 -26 -409
rect 26 -461 65 -409
rect -64 -627 65 -461
rect -64 -679 -26 -627
rect 26 -679 65 -627
rect -64 -845 65 -679
rect -64 -897 -26 -845
rect 26 -897 65 -845
rect -64 -1062 65 -897
rect -64 -1114 -26 -1062
rect 26 -1114 65 -1062
rect -64 -1280 65 -1114
rect -64 -1332 -26 -1280
rect 26 -1332 65 -1280
rect -64 -1497 65 -1332
rect -64 -1549 -26 -1497
rect 26 -1549 65 -1497
rect -64 -1715 65 -1549
rect -64 -1767 -26 -1715
rect 26 -1767 65 -1715
rect -64 -1933 65 -1767
rect -64 -1985 -26 -1933
rect 26 -1985 65 -1933
rect -64 -2150 65 -1985
rect -64 -2202 -26 -2150
rect 26 -2202 65 -2150
rect -64 -2243 65 -2202
<< properties >>
string GDS_END 673640
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 672164
<< end >>
