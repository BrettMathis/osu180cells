magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect 85432 578 85816 46102
<< metal1 >>
rect 0 403 1000 46294
<< metal2 >>
rect 424 403 1424 45776
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB43105899832108_64x8m81  M1_PSUB43105899832108_64x8m81_0
timestamp 1669390400
transform -1 0 85672 0 1 45688
box -42 -42 85602 414
use M1_PSUB43105899832108_64x8m81  M1_PSUB43105899832108_64x8m81_1
timestamp 1669390400
transform -1 0 85672 0 1 620
box -42 -42 85602 414
use M1_PSUB43105899832109_64x8m81  M1_PSUB43105899832109_64x8m81_0
timestamp 1669390400
transform 1 0 85474 0 1 1140
box -42 -42 342 44442
use M1_PSUB43105899832109_64x8m81  M1_PSUB43105899832109_64x8m81_1
timestamp 1669390400
transform 1 0 112 0 1 1140
box -42 -42 342 44442
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2255308
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2254652
string path 4.620 11.160 4.620 0.000 
<< end >>
