magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4006 1094
<< pwell >>
rect -86 -86 4006 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 217 836 333
rect 884 217 1004 333
rect 1108 217 1228 333
rect 1276 217 1396 333
rect 1576 217 1696 333
rect 1800 217 1920 333
rect 2024 217 2144 333
rect 2192 217 2312 333
rect 2460 69 2580 333
rect 2684 69 2804 333
rect 2908 69 3028 333
rect 3132 69 3252 333
rect 3356 69 3476 333
rect 3580 69 3700 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 756 573 856 773
rect 904 573 1004 773
rect 1148 573 1248 773
rect 1296 573 1396 773
rect 1576 573 1676 773
rect 1799 573 1899 773
rect 2084 573 2184 773
rect 2240 573 2340 773
rect 2488 573 2588 939
rect 2692 573 2792 939
rect 2896 573 2996 939
rect 3100 573 3200 939
rect 3304 573 3404 939
rect 3508 573 3608 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 276 716 333
rect 628 230 641 276
rect 687 230 716 276
rect 628 217 716 230
rect 836 217 884 333
rect 1004 320 1108 333
rect 1004 274 1033 320
rect 1079 274 1108 320
rect 1004 217 1108 274
rect 1228 217 1276 333
rect 1396 217 1576 333
rect 1696 320 1800 333
rect 1696 274 1725 320
rect 1771 274 1800 320
rect 1696 217 1800 274
rect 1920 320 2024 333
rect 1920 274 1949 320
rect 1995 274 2024 320
rect 1920 217 2024 274
rect 2144 217 2192 333
rect 2312 222 2460 333
rect 2312 217 2385 222
rect 1456 127 1516 217
rect 1445 119 1516 127
rect 1445 114 1517 119
rect 1445 68 1458 114
rect 1504 68 1517 114
rect 2372 82 2385 217
rect 2431 82 2460 222
rect 2372 69 2460 82
rect 2580 320 2684 333
rect 2580 180 2609 320
rect 2655 180 2684 320
rect 2580 69 2684 180
rect 2804 222 2908 333
rect 2804 82 2833 222
rect 2879 82 2908 222
rect 2804 69 2908 82
rect 3028 320 3132 333
rect 3028 180 3057 320
rect 3103 180 3132 320
rect 3028 69 3132 180
rect 3252 222 3356 333
rect 3252 82 3281 222
rect 3327 82 3356 222
rect 3252 69 3356 82
rect 3476 314 3580 333
rect 3476 174 3505 314
rect 3551 174 3580 314
rect 3476 69 3580 174
rect 3700 222 3788 333
rect 3700 82 3729 222
rect 3775 82 3788 222
rect 3700 69 3788 82
rect 1445 55 1517 68
<< mvpdiff >>
rect 624 932 696 945
rect 56 836 144 849
rect 56 696 69 836
rect 115 696 144 836
rect 56 573 144 696
rect 244 836 348 849
rect 244 790 273 836
rect 319 790 348 836
rect 244 573 348 790
rect 448 632 536 849
rect 448 586 477 632
rect 523 586 536 632
rect 448 573 536 586
rect 624 792 637 932
rect 683 792 696 932
rect 2400 926 2488 939
rect 624 773 696 792
rect 2400 786 2413 926
rect 2459 786 2488 926
rect 2400 773 2488 786
rect 624 573 756 773
rect 856 573 904 773
rect 1004 632 1148 773
rect 1004 586 1033 632
rect 1079 586 1148 632
rect 1004 573 1148 586
rect 1248 573 1296 773
rect 1396 760 1576 773
rect 1396 620 1425 760
rect 1471 620 1576 760
rect 1396 573 1576 620
rect 1676 726 1799 773
rect 1676 586 1724 726
rect 1770 586 1799 726
rect 1676 573 1799 586
rect 1899 726 2084 773
rect 1899 586 1949 726
rect 1995 586 2084 726
rect 1899 573 2084 586
rect 2184 573 2240 773
rect 2340 573 2488 773
rect 2588 726 2692 939
rect 2588 586 2617 726
rect 2663 586 2692 726
rect 2588 573 2692 586
rect 2792 926 2896 939
rect 2792 786 2821 926
rect 2867 786 2896 926
rect 2792 573 2896 786
rect 2996 726 3100 939
rect 2996 586 3025 726
rect 3071 586 3100 726
rect 2996 573 3100 586
rect 3200 926 3304 939
rect 3200 786 3229 926
rect 3275 786 3304 926
rect 3200 573 3304 786
rect 3404 726 3508 939
rect 3404 586 3433 726
rect 3479 586 3508 726
rect 3404 573 3508 586
rect 3608 926 3696 939
rect 3608 786 3637 926
rect 3683 786 3696 926
rect 3608 573 3696 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 230 687 276
rect 1033 274 1079 320
rect 1725 274 1771 320
rect 1949 274 1995 320
rect 1458 68 1504 114
rect 2385 82 2431 222
rect 2609 180 2655 320
rect 2833 82 2879 222
rect 3057 180 3103 320
rect 3281 82 3327 222
rect 3505 174 3551 314
rect 3729 82 3775 222
<< mvpdiffc >>
rect 69 696 115 836
rect 273 790 319 836
rect 477 586 523 632
rect 637 792 683 932
rect 2413 786 2459 926
rect 1033 586 1079 632
rect 1425 620 1471 760
rect 1724 586 1770 726
rect 1949 586 1995 726
rect 2617 586 2663 726
rect 2821 786 2867 926
rect 3025 586 3071 726
rect 3229 786 3275 926
rect 3433 586 3479 726
rect 3637 786 3683 926
<< polysilicon >>
rect 2488 939 2588 983
rect 2692 939 2792 983
rect 2896 939 2996 983
rect 3100 939 3200 983
rect 3304 939 3404 983
rect 3508 939 3608 983
rect 144 849 244 893
rect 348 849 448 893
rect 1148 865 1899 905
rect 1148 852 1248 865
rect 756 773 856 817
rect 904 773 1004 817
rect 1148 806 1161 852
rect 1207 806 1248 852
rect 1148 773 1248 806
rect 1296 773 1396 817
rect 1576 773 1676 817
rect 1799 773 1899 865
rect 2084 773 2184 817
rect 2240 773 2340 817
rect 144 504 244 573
rect 144 458 157 504
rect 203 458 244 504
rect 144 377 244 458
rect 124 333 244 377
rect 348 433 448 573
rect 756 540 856 573
rect 756 494 769 540
rect 815 494 856 540
rect 756 481 856 494
rect 348 412 836 433
rect 348 366 361 412
rect 407 393 836 412
rect 407 366 468 393
rect 348 333 468 366
rect 716 333 836 393
rect 904 412 1004 573
rect 1148 529 1248 573
rect 904 377 926 412
rect 884 366 926 377
rect 972 366 1004 412
rect 1296 412 1396 573
rect 1296 377 1337 412
rect 884 333 1004 366
rect 1108 333 1228 377
rect 1276 366 1337 377
rect 1383 366 1396 412
rect 1276 333 1396 366
rect 1576 540 1676 573
rect 1576 494 1589 540
rect 1635 494 1676 540
rect 1576 377 1676 494
rect 1799 485 1899 573
rect 2084 540 2184 573
rect 2084 529 2125 540
rect 2112 494 2125 529
rect 2171 494 2184 540
rect 1799 445 2064 485
rect 2112 481 2184 494
rect 2240 529 2340 573
rect 2488 540 2588 573
rect 2024 377 2064 445
rect 2240 412 2312 529
rect 2240 377 2253 412
rect 1576 333 1696 377
rect 1800 333 1920 377
rect 2024 333 2144 377
rect 2192 366 2253 377
rect 2299 366 2312 412
rect 2488 494 2501 540
rect 2547 494 2588 540
rect 2488 456 2588 494
rect 2692 456 2792 573
rect 2896 529 2996 573
rect 2488 393 2792 456
rect 2488 377 2580 393
rect 2192 333 2312 366
rect 2460 333 2580 377
rect 2684 377 2792 393
rect 2908 465 2996 529
rect 3100 465 3200 573
rect 3304 465 3404 573
rect 3508 465 3608 573
rect 2908 452 3700 465
rect 2908 406 2921 452
rect 2967 406 3125 452
rect 3171 406 3331 452
rect 3377 406 3700 452
rect 2908 393 3700 406
rect 2684 333 2804 377
rect 2908 333 3028 393
rect 3132 333 3252 393
rect 3356 333 3476 393
rect 3580 333 3700 393
rect 124 131 244 175
rect 348 131 468 175
rect 716 173 836 217
rect 884 173 1004 217
rect 1108 184 1228 217
rect 1108 138 1121 184
rect 1167 138 1228 184
rect 1276 173 1396 217
rect 1108 125 1228 138
rect 1576 173 1696 217
rect 1800 184 1920 217
rect 1800 138 1813 184
rect 1859 138 1920 184
rect 2024 173 2144 217
rect 2192 173 2312 217
rect 1800 125 1920 138
rect 2460 25 2580 69
rect 2684 25 2804 69
rect 2908 25 3028 69
rect 3132 25 3252 69
rect 3356 25 3476 69
rect 3580 25 3700 69
<< polycontact >>
rect 1161 806 1207 852
rect 157 458 203 504
rect 769 494 815 540
rect 361 366 407 412
rect 926 366 972 412
rect 1337 366 1383 412
rect 1589 494 1635 540
rect 2125 494 2171 540
rect 2253 366 2299 412
rect 2501 494 2547 540
rect 2921 406 2967 452
rect 3125 406 3171 452
rect 3331 406 3377 452
rect 1121 138 1167 184
rect 1813 138 1859 184
<< metal1 >>
rect 0 932 3920 1098
rect 0 918 637 932
rect 69 836 115 847
rect 262 836 330 918
rect 262 790 273 836
rect 319 790 330 836
rect 683 926 3920 932
rect 683 918 2413 926
rect 637 781 683 792
rect 1161 852 1207 863
rect 1161 735 1207 806
rect 115 696 1207 735
rect 69 689 1207 696
rect 1425 760 1471 918
rect 2459 918 2821 926
rect 2413 775 2459 786
rect 2867 918 3229 926
rect 2821 775 2867 786
rect 3275 918 3637 926
rect 3229 775 3275 786
rect 3683 918 3920 926
rect 3637 775 3683 786
rect 69 685 407 689
rect 142 504 301 542
rect 142 458 157 504
rect 203 458 301 504
rect 142 447 301 458
rect 361 412 407 685
rect 477 632 523 643
rect 477 551 523 586
rect 1033 632 1079 643
rect 1425 609 1471 620
rect 1724 726 1771 737
rect 1033 551 1079 586
rect 1770 586 1771 726
rect 477 540 815 551
rect 477 505 769 540
rect 49 366 361 401
rect 769 379 815 494
rect 1033 540 1635 551
rect 1033 494 1589 540
rect 1033 483 1635 494
rect 49 355 407 366
rect 49 320 95 355
rect 49 263 95 274
rect 497 333 815 379
rect 497 320 543 333
rect 497 263 543 274
rect 641 276 687 287
rect 273 234 319 245
rect 273 90 319 188
rect 641 90 687 230
rect 769 184 815 333
rect 926 412 978 423
rect 972 366 978 412
rect 926 242 978 366
rect 1033 320 1079 483
rect 1724 423 1771 586
rect 1337 412 1771 423
rect 1383 366 1771 412
rect 1337 355 1771 366
rect 1033 263 1079 274
rect 1725 320 1771 355
rect 1725 263 1771 274
rect 1949 726 2387 737
rect 1995 691 2387 726
rect 1949 320 1995 586
rect 1949 263 1995 274
rect 2125 540 2171 551
rect 2341 540 2387 691
rect 2617 726 2663 737
rect 2341 494 2501 540
rect 2547 494 2558 540
rect 2125 217 2171 494
rect 2617 463 2663 586
rect 3025 726 3071 737
rect 3433 726 3554 737
rect 3071 586 3433 621
rect 3479 586 3554 726
rect 3025 575 3554 586
rect 2617 452 3377 463
rect 2617 423 2921 452
rect 2253 412 2921 423
rect 2299 406 2921 412
rect 2967 406 3125 452
rect 3171 406 3331 452
rect 2299 395 3377 406
rect 2299 366 2662 395
rect 2253 355 2662 366
rect 2609 320 2662 355
rect 3423 331 3554 575
rect 1133 184 2171 217
rect 769 138 1121 184
rect 1167 171 1813 184
rect 1167 138 1178 171
rect 1802 138 1813 171
rect 1859 138 2171 184
rect 2385 222 2431 233
rect 1458 114 1504 125
rect 0 68 1458 90
rect 1504 82 2385 90
rect 2655 180 2662 320
rect 3057 320 3554 331
rect 2609 169 2662 180
rect 2833 222 2879 233
rect 2431 82 2833 90
rect 3103 314 3554 320
rect 3103 279 3505 314
rect 3057 169 3103 180
rect 3281 222 3327 233
rect 2879 82 3281 90
rect 3502 174 3505 279
rect 3551 174 3554 314
rect 3502 163 3554 174
rect 3729 222 3775 233
rect 3327 82 3729 90
rect 3775 82 3920 90
rect 1504 68 3920 82
rect 0 -90 3920 68
<< labels >>
flabel metal1 s 142 447 301 542 0 FreeSans 200 0 0 0 CLK
port 2 nsew clock input
flabel metal1 s 926 242 978 423 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3433 621 3554 737 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3920 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 641 245 687 287 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3025 621 3071 737 1 Q
port 3 nsew default output
rlabel metal1 s 3025 575 3554 621 1 Q
port 3 nsew default output
rlabel metal1 s 3423 331 3554 575 1 Q
port 3 nsew default output
rlabel metal1 s 3057 279 3554 331 1 Q
port 3 nsew default output
rlabel metal1 s 3502 169 3554 279 1 Q
port 3 nsew default output
rlabel metal1 s 3057 169 3103 279 1 Q
port 3 nsew default output
rlabel metal1 s 3502 163 3554 169 1 Q
port 3 nsew default output
rlabel metal1 s 3637 790 3683 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3229 790 3275 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2821 790 2867 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2413 790 2459 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1425 790 1471 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 637 790 683 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 262 790 330 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3637 781 3683 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3229 781 3275 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2821 781 2867 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2413 781 2459 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1425 781 1471 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 637 781 683 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3637 775 3683 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3229 775 3275 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2821 775 2867 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2413 775 2459 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1425 775 1471 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1425 609 1471 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3729 125 3775 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3281 125 3327 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2833 125 2879 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2385 125 2431 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 641 125 687 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3729 90 3775 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3281 90 3327 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2833 90 2879 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2385 90 2431 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1458 90 1504 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3920 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 1008
string GDS_END 593174
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 584544
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
