magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -1119 26 1119 66
rect -1119 -26 -1080 26
rect -1028 -26 -870 26
rect -818 -26 -659 26
rect -607 -26 -448 26
rect -396 -26 -237 26
rect -185 -26 -26 26
rect 26 -26 185 26
rect 237 -26 396 26
rect 448 -26 607 26
rect 659 -26 818 26
rect 870 -26 1028 26
rect 1080 -26 1119 26
rect -1119 -67 1119 -26
<< via1 >>
rect -1080 -26 -1028 26
rect -870 -26 -818 26
rect -659 -26 -607 26
rect -448 -26 -396 26
rect -237 -26 -185 26
rect -26 -26 26 26
rect 185 -26 237 26
rect 396 -26 448 26
rect 607 -26 659 26
rect 818 -26 870 26
rect 1028 -26 1080 26
<< metal2 >>
rect -1118 26 1119 66
rect -1118 -26 -1080 26
rect -1028 -26 -870 26
rect -818 -26 -659 26
rect -607 -26 -448 26
rect -396 -26 -237 26
rect -185 -26 -26 26
rect 26 -26 185 26
rect 237 -26 396 26
rect 448 -26 607 26
rect 659 -26 818 26
rect 870 -26 1028 26
rect 1080 -26 1119 26
rect -1118 -67 1119 -26
<< properties >>
string GDS_END 205056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 204220
<< end >>
