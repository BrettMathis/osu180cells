magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 568
rect 224 0 344 568
rect 448 0 568 568
rect 672 0 792 568
rect 896 0 1016 568
rect 1120 0 1240 568
rect 1344 0 1464 568
rect 1568 0 1688 568
<< mvndiff >>
rect -88 555 0 568
rect -88 509 -75 555
rect -29 509 0 555
rect -88 431 0 509
rect -88 385 -75 431
rect -29 385 0 431
rect -88 307 0 385
rect -88 261 -75 307
rect -29 261 0 307
rect -88 183 0 261
rect -88 137 -75 183
rect -29 137 0 183
rect -88 59 0 137
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 555 224 568
rect 120 509 149 555
rect 195 509 224 555
rect 120 431 224 509
rect 120 385 149 431
rect 195 385 224 431
rect 120 307 224 385
rect 120 261 149 307
rect 195 261 224 307
rect 120 183 224 261
rect 120 137 149 183
rect 195 137 224 183
rect 120 59 224 137
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 555 448 568
rect 344 509 373 555
rect 419 509 448 555
rect 344 431 448 509
rect 344 385 373 431
rect 419 385 448 431
rect 344 307 448 385
rect 344 261 373 307
rect 419 261 448 307
rect 344 183 448 261
rect 344 137 373 183
rect 419 137 448 183
rect 344 59 448 137
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 555 672 568
rect 568 509 597 555
rect 643 509 672 555
rect 568 431 672 509
rect 568 385 597 431
rect 643 385 672 431
rect 568 307 672 385
rect 568 261 597 307
rect 643 261 672 307
rect 568 183 672 261
rect 568 137 597 183
rect 643 137 672 183
rect 568 59 672 137
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 555 896 568
rect 792 509 821 555
rect 867 509 896 555
rect 792 431 896 509
rect 792 385 821 431
rect 867 385 896 431
rect 792 307 896 385
rect 792 261 821 307
rect 867 261 896 307
rect 792 183 896 261
rect 792 137 821 183
rect 867 137 896 183
rect 792 59 896 137
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 555 1120 568
rect 1016 509 1045 555
rect 1091 509 1120 555
rect 1016 431 1120 509
rect 1016 385 1045 431
rect 1091 385 1120 431
rect 1016 307 1120 385
rect 1016 261 1045 307
rect 1091 261 1120 307
rect 1016 183 1120 261
rect 1016 137 1045 183
rect 1091 137 1120 183
rect 1016 59 1120 137
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 555 1344 568
rect 1240 509 1269 555
rect 1315 509 1344 555
rect 1240 431 1344 509
rect 1240 385 1269 431
rect 1315 385 1344 431
rect 1240 307 1344 385
rect 1240 261 1269 307
rect 1315 261 1344 307
rect 1240 183 1344 261
rect 1240 137 1269 183
rect 1315 137 1344 183
rect 1240 59 1344 137
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 555 1568 568
rect 1464 509 1493 555
rect 1539 509 1568 555
rect 1464 431 1568 509
rect 1464 385 1493 431
rect 1539 385 1568 431
rect 1464 307 1568 385
rect 1464 261 1493 307
rect 1539 261 1568 307
rect 1464 183 1568 261
rect 1464 137 1493 183
rect 1539 137 1568 183
rect 1464 59 1568 137
rect 1464 13 1493 59
rect 1539 13 1568 59
rect 1464 0 1568 13
rect 1688 555 1776 568
rect 1688 509 1717 555
rect 1763 509 1776 555
rect 1688 431 1776 509
rect 1688 385 1717 431
rect 1763 385 1776 431
rect 1688 307 1776 385
rect 1688 261 1717 307
rect 1763 261 1776 307
rect 1688 183 1776 261
rect 1688 137 1717 183
rect 1763 137 1776 183
rect 1688 59 1776 137
rect 1688 13 1717 59
rect 1763 13 1776 59
rect 1688 0 1776 13
<< mvndiffc >>
rect -75 509 -29 555
rect -75 385 -29 431
rect -75 261 -29 307
rect -75 137 -29 183
rect -75 13 -29 59
rect 149 509 195 555
rect 149 385 195 431
rect 149 261 195 307
rect 149 137 195 183
rect 149 13 195 59
rect 373 509 419 555
rect 373 385 419 431
rect 373 261 419 307
rect 373 137 419 183
rect 373 13 419 59
rect 597 509 643 555
rect 597 385 643 431
rect 597 261 643 307
rect 597 137 643 183
rect 597 13 643 59
rect 821 509 867 555
rect 821 385 867 431
rect 821 261 867 307
rect 821 137 867 183
rect 821 13 867 59
rect 1045 509 1091 555
rect 1045 385 1091 431
rect 1045 261 1091 307
rect 1045 137 1091 183
rect 1045 13 1091 59
rect 1269 509 1315 555
rect 1269 385 1315 431
rect 1269 261 1315 307
rect 1269 137 1315 183
rect 1269 13 1315 59
rect 1493 509 1539 555
rect 1493 385 1539 431
rect 1493 261 1539 307
rect 1493 137 1539 183
rect 1493 13 1539 59
rect 1717 509 1763 555
rect 1717 385 1763 431
rect 1717 261 1763 307
rect 1717 137 1763 183
rect 1717 13 1763 59
<< polysilicon >>
rect 0 568 120 612
rect 224 568 344 612
rect 448 568 568 612
rect 672 568 792 612
rect 896 568 1016 612
rect 1120 568 1240 612
rect 1344 568 1464 612
rect 1568 568 1688 612
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
<< metal1 >>
rect -75 555 -29 568
rect -75 431 -29 509
rect -75 307 -29 385
rect -75 183 -29 261
rect -75 59 -29 137
rect -75 0 -29 13
rect 149 555 195 568
rect 149 431 195 509
rect 149 307 195 385
rect 149 183 195 261
rect 149 59 195 137
rect 149 0 195 13
rect 373 555 419 568
rect 373 431 419 509
rect 373 307 419 385
rect 373 183 419 261
rect 373 59 419 137
rect 373 0 419 13
rect 597 555 643 568
rect 597 431 643 509
rect 597 307 643 385
rect 597 183 643 261
rect 597 59 643 137
rect 597 0 643 13
rect 821 555 867 568
rect 821 431 867 509
rect 821 307 867 385
rect 821 183 867 261
rect 821 59 867 137
rect 821 0 867 13
rect 1045 555 1091 568
rect 1045 431 1091 509
rect 1045 307 1091 385
rect 1045 183 1091 261
rect 1045 59 1091 137
rect 1045 0 1091 13
rect 1269 555 1315 568
rect 1269 431 1315 509
rect 1269 307 1315 385
rect 1269 183 1315 261
rect 1269 59 1315 137
rect 1269 0 1315 13
rect 1493 555 1539 568
rect 1493 431 1539 509
rect 1493 307 1539 385
rect 1493 183 1539 261
rect 1493 59 1539 137
rect 1493 0 1539 13
rect 1717 555 1763 568
rect 1717 431 1763 509
rect 1717 307 1763 385
rect 1717 183 1763 261
rect 1717 59 1763 137
rect 1717 0 1763 13
<< labels >>
flabel metal1 s -52 284 -52 284 0 FreeSans 200 0 0 0 S
flabel metal1 s 1740 284 1740 284 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 284 172 284 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 284 396 284 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 284 620 284 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 284 844 284 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 284 1068 284 0 FreeSans 200 0 0 0 D
flabel metal1 s 1292 284 1292 284 0 FreeSans 200 0 0 0 S
flabel metal1 s 1516 284 1516 284 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 70938
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 64488
<< end >>
