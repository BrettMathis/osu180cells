magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 6583 29008 9560 29932
rect 13849 29658 15116 29948
rect 13849 29581 15441 29658
rect 10186 29017 10786 29089
rect 13850 29008 15441 29581
rect 6583 28958 8962 29008
rect 16520 28976 21087 29903
<< mvndiff >>
rect 2123 28860 2278 29248
rect 25490 28860 25646 29248
<< mvpsubdiff >>
rect 15782 29782 16254 29839
rect 15782 29736 15837 29782
rect 15883 29736 15995 29782
rect 16041 29736 16153 29782
rect 16199 29736 16254 29782
rect 15782 29679 16254 29736
<< mvnsubdiff >>
rect 13985 29782 14931 29839
rect 13985 29736 14040 29782
rect 14086 29736 14198 29782
rect 14244 29736 14356 29782
rect 14402 29736 14514 29782
rect 14560 29736 14673 29782
rect 14719 29736 14831 29782
rect 14877 29736 14931 29782
rect 13985 29679 14931 29736
<< mvpsubdiffcont >>
rect 15837 29736 15883 29782
rect 15995 29736 16041 29782
rect 16153 29736 16199 29782
<< mvnsubdiffcont >>
rect 14040 29736 14086 29782
rect 14198 29736 14244 29782
rect 14356 29736 14402 29782
rect 14514 29736 14560 29782
rect 14673 29736 14719 29782
rect 14831 29736 14877 29782
<< polysilicon >>
rect 13623 29716 13801 29735
rect 13623 29670 13642 29716
rect 13782 29670 13801 29716
rect 15364 29764 15467 29783
rect 15364 29718 15390 29764
rect 15436 29718 15467 29764
rect 13623 29651 13801 29670
rect 6556 29496 6690 29616
rect 9314 29518 9448 29623
rect 6556 29392 6659 29496
rect 6374 29272 6690 29392
rect 9314 29378 9358 29518
rect 9404 29378 9448 29518
rect 11998 29431 12082 29450
rect 11998 29392 12017 29431
rect 9314 29273 9448 29378
rect 11043 29272 11385 29392
rect 11914 29291 12017 29392
rect 12063 29291 12082 29431
rect 11914 29272 12082 29291
rect 13664 29273 13768 29651
rect 15364 29392 15467 29718
rect 18271 29506 18355 29616
rect 13915 29272 13986 29392
rect 15305 29272 15467 29392
rect 15583 29471 15667 29490
rect 15583 29331 15602 29471
rect 15648 29392 15667 29471
rect 15648 29331 15755 29392
rect 15583 29272 15755 29331
rect 16255 29272 16656 29392
rect 17975 29272 18045 29392
rect 18271 29366 18290 29506
rect 18336 29366 18355 29506
rect 18271 29272 18355 29366
rect 21010 29392 21113 29616
rect 21010 29272 21325 29392
rect 23347 29272 23417 29392
<< polycontact >>
rect 13642 29670 13782 29716
rect 15390 29718 15436 29764
rect 9358 29378 9404 29518
rect 12017 29291 12063 29431
rect 15602 29331 15648 29471
rect 18290 29366 18336 29506
<< metal1 >>
rect 2123 29116 4017 29767
rect 4324 29452 6336 29839
rect 6728 29706 7700 29746
rect 6728 29654 6766 29706
rect 6818 29654 6977 29706
rect 7029 29654 7188 29706
rect 7240 29654 7399 29706
rect 7451 29654 7610 29706
rect 7662 29654 7700 29706
rect 6728 29614 7700 29654
rect 11385 29731 11913 29819
rect 11385 29679 11575 29731
rect 11627 29679 11755 29731
rect 11807 29679 11913 29731
rect 9323 29518 9439 29585
rect 6482 29388 6767 29508
rect 4335 29245 5307 29285
rect 6482 29277 6598 29388
rect 9323 29378 9358 29518
rect 9404 29378 9439 29518
rect 10338 29508 10888 29515
rect 10337 29474 10888 29508
rect 10337 29422 10376 29474
rect 10428 29422 10587 29474
rect 10639 29422 10798 29474
rect 10850 29422 10888 29474
rect 10337 29388 10888 29422
rect 11385 29513 11913 29679
rect 13531 29782 14912 29819
rect 15755 29818 16283 29819
rect 13531 29778 14040 29782
rect 13531 29726 14033 29778
rect 14086 29736 14198 29782
rect 14244 29778 14356 29782
rect 14085 29726 14244 29736
rect 14296 29736 14356 29778
rect 14402 29778 14514 29782
rect 14402 29736 14455 29778
rect 14296 29726 14455 29736
rect 14507 29736 14514 29778
rect 14560 29736 14673 29782
rect 14719 29736 14831 29782
rect 14877 29736 14912 29782
rect 14507 29726 14912 29736
rect 13531 29717 14912 29726
rect 13531 29665 13569 29717
rect 13621 29716 13781 29717
rect 13621 29670 13642 29716
rect 13833 29699 14912 29717
rect 15061 29782 16283 29818
rect 15061 29778 15837 29782
rect 15061 29726 15100 29778
rect 15152 29726 15311 29778
rect 15363 29764 15522 29778
rect 15363 29726 15390 29764
rect 15061 29718 15390 29726
rect 15436 29726 15522 29764
rect 15574 29726 15733 29778
rect 15785 29736 15837 29778
rect 15883 29736 15995 29782
rect 16041 29736 16153 29782
rect 16199 29736 16283 29782
rect 20112 29740 20874 29746
rect 15785 29726 16283 29736
rect 15436 29718 16283 29726
rect 13833 29686 14545 29699
rect 13833 29685 14040 29686
rect 15061 29685 16283 29718
rect 13621 29665 13781 29670
rect 13833 29665 13871 29685
rect 13531 29624 13871 29665
rect 11385 29461 11575 29513
rect 11627 29461 11755 29513
rect 11807 29461 11913 29513
rect 15591 29471 15659 29482
rect 11385 29421 11913 29461
rect 12006 29431 12334 29468
rect 10338 29382 10888 29388
rect 4335 29193 4373 29245
rect 4425 29193 4584 29245
rect 4636 29193 4795 29245
rect 4847 29193 5006 29245
rect 5058 29193 5217 29245
rect 5269 29193 5307 29245
rect 4335 29153 5307 29193
rect 6240 29157 6598 29277
rect 6728 29243 7700 29283
rect 6728 29191 6766 29243
rect 6818 29191 6977 29243
rect 7029 29191 7188 29243
rect 7240 29191 7399 29243
rect 7451 29191 7610 29243
rect 7662 29191 7700 29243
rect 6728 29151 7700 29191
rect 9323 29277 9439 29378
rect 12006 29291 12017 29431
rect 12063 29422 12334 29431
rect 13509 29422 14174 29468
rect 15591 29467 15602 29471
rect 12063 29291 12074 29422
rect 15268 29421 15602 29467
rect 15591 29331 15602 29421
rect 15648 29331 15659 29471
rect 15755 29388 16283 29685
rect 16656 29706 20942 29740
rect 16656 29654 20151 29706
rect 20203 29654 20362 29706
rect 20414 29654 20573 29706
rect 20625 29654 20784 29706
rect 20836 29654 20942 29706
rect 16656 29620 20942 29654
rect 16656 29436 17974 29620
rect 20112 29613 20874 29620
rect 18279 29506 18347 29517
rect 15591 29320 15659 29331
rect 18279 29366 18290 29506
rect 18336 29366 18347 29506
rect 20898 29421 21184 29467
rect 18279 29355 18347 29366
rect 12006 29280 12074 29291
rect 9323 29157 11913 29277
rect 12294 29243 13478 29284
rect 18279 29277 18346 29355
rect 12294 29191 12333 29243
rect 12385 29191 12544 29243
rect 12596 29191 12755 29243
rect 12807 29191 12966 29243
rect 13018 29191 13177 29243
rect 13229 29191 13387 29243
rect 13439 29191 13478 29243
rect 13570 29198 14174 29244
rect 12294 29150 13478 29191
rect 15755 29157 18346 29277
rect 20112 29243 20874 29283
rect 20112 29191 20151 29243
rect 20203 29191 20362 29243
rect 20414 29191 20573 29243
rect 20625 29191 20784 29243
rect 20836 29191 20874 29243
rect 21067 29243 21184 29421
rect 21324 29402 23346 29819
rect 22366 29243 23338 29283
rect 21067 29197 21425 29243
rect 20112 29150 20874 29191
rect 22366 29191 22404 29243
rect 22456 29191 22615 29243
rect 22667 29191 22826 29243
rect 22878 29191 23037 29243
rect 23089 29191 23248 29243
rect 23300 29191 23338 29243
rect 22366 29151 23338 29191
rect 23751 29116 25646 29767
rect 2123 28865 2278 29116
rect 25490 28865 25646 29116
<< via1 >>
rect 6766 29654 6818 29706
rect 6977 29654 7029 29706
rect 7188 29654 7240 29706
rect 7399 29654 7451 29706
rect 7610 29654 7662 29706
rect 11575 29679 11627 29731
rect 11755 29679 11807 29731
rect 10376 29422 10428 29474
rect 10587 29422 10639 29474
rect 10798 29422 10850 29474
rect 14033 29736 14040 29778
rect 14040 29736 14085 29778
rect 14033 29726 14085 29736
rect 14244 29726 14296 29778
rect 14455 29726 14507 29778
rect 13569 29665 13621 29717
rect 13781 29716 13833 29717
rect 13781 29670 13782 29716
rect 13782 29670 13833 29716
rect 15100 29726 15152 29778
rect 15311 29726 15363 29778
rect 15522 29726 15574 29778
rect 15733 29726 15785 29778
rect 13781 29665 13833 29670
rect 11575 29461 11627 29513
rect 11755 29461 11807 29513
rect 4373 29193 4425 29245
rect 4584 29193 4636 29245
rect 4795 29193 4847 29245
rect 5006 29193 5058 29245
rect 5217 29193 5269 29245
rect 6766 29191 6818 29243
rect 6977 29191 7029 29243
rect 7188 29191 7240 29243
rect 7399 29191 7451 29243
rect 7610 29191 7662 29243
rect 20151 29654 20203 29706
rect 20362 29654 20414 29706
rect 20573 29654 20625 29706
rect 20784 29654 20836 29706
rect 12333 29191 12385 29243
rect 12544 29191 12596 29243
rect 12755 29191 12807 29243
rect 12966 29191 13018 29243
rect 13177 29191 13229 29243
rect 13387 29191 13439 29243
rect 20151 29191 20203 29243
rect 20362 29191 20414 29243
rect 20573 29191 20625 29243
rect 20784 29191 20836 29243
rect 22404 29191 22456 29243
rect 22615 29191 22667 29243
rect 22826 29191 22878 29243
rect 23037 29191 23089 29243
rect 23248 29191 23300 29243
<< metal2 >>
rect 2092 28813 4211 29876
rect 5550 29728 6347 29801
rect 5550 29672 5611 29728
rect 5667 29672 5822 29728
rect 5878 29672 6033 29728
rect 6089 29672 6244 29728
rect 6300 29672 6347 29728
rect 4334 29247 5307 29286
rect 4334 29191 4371 29247
rect 4427 29191 4582 29247
rect 4638 29191 4793 29247
rect 4849 29191 5004 29247
rect 5060 29191 5215 29247
rect 5271 29191 5307 29247
rect 4334 29153 5307 29191
rect 5550 28813 6347 29672
rect 6451 29706 7738 29801
rect 6451 29654 6766 29706
rect 6818 29654 6977 29706
rect 7029 29654 7188 29706
rect 7240 29654 7399 29706
rect 7451 29654 7610 29706
rect 7662 29654 7738 29706
rect 6451 29243 7738 29654
rect 6451 29191 6766 29243
rect 6818 29191 6977 29243
rect 7029 29191 7188 29243
rect 7240 29191 7399 29243
rect 7451 29191 7610 29243
rect 7662 29191 7738 29243
rect 6451 28813 7738 29191
rect 8186 29245 9066 29284
rect 8186 29189 8222 29245
rect 8278 29189 8433 29245
rect 8489 29189 8644 29245
rect 8700 29189 8855 29245
rect 8911 29189 9066 29245
rect 8186 28813 9066 29189
rect 9591 28813 10186 29801
rect 10276 29474 10941 29801
rect 10276 29422 10376 29474
rect 10428 29422 10587 29474
rect 10639 29422 10798 29474
rect 10850 29422 10941 29474
rect 10276 28813 10941 29422
rect 11537 29731 11846 29801
rect 13994 29778 14545 29819
rect 11537 29728 11575 29731
rect 11627 29728 11755 29731
rect 11807 29728 11846 29731
rect 11537 29672 11573 29728
rect 11629 29672 11753 29728
rect 11809 29672 11846 29728
rect 11537 29513 11846 29672
rect 13531 29717 13871 29758
rect 13531 29665 13569 29717
rect 13621 29665 13781 29717
rect 13833 29665 13871 29717
rect 13531 29624 13871 29665
rect 13994 29726 14033 29778
rect 14085 29726 14244 29778
rect 14296 29726 14455 29778
rect 14507 29726 14545 29778
rect 11537 29461 11575 29513
rect 11627 29461 11755 29513
rect 11807 29461 11846 29513
rect 11537 28813 11846 29461
rect 12294 29245 13478 29284
rect 12294 29189 12331 29245
rect 12387 29189 12542 29245
rect 12598 29189 12753 29245
rect 12809 29189 12964 29245
rect 13020 29189 13175 29245
rect 13231 29189 13385 29245
rect 13441 29189 13478 29245
rect 12294 29150 13478 29189
rect 13994 29238 14545 29726
rect 13994 29182 14031 29238
rect 14087 29182 14242 29238
rect 14298 29182 14453 29238
rect 14509 29182 14545 29238
rect 13994 29144 14545 29182
rect 15026 29778 15887 29819
rect 15026 29726 15100 29778
rect 15152 29726 15311 29778
rect 15363 29726 15522 29778
rect 15574 29726 15733 29778
rect 15785 29726 15887 29778
rect 12040 28828 12639 28964
rect 12040 28772 12100 28828
rect 12156 28772 12311 28828
rect 12367 28772 12522 28828
rect 12578 28772 12639 28828
rect 15026 28813 15887 29726
rect 20112 29706 21313 29801
rect 20112 29654 20151 29706
rect 20203 29654 20362 29706
rect 20414 29654 20573 29706
rect 20625 29654 20784 29706
rect 20836 29654 21313 29706
rect 20112 29243 21313 29654
rect 20112 29191 20151 29243
rect 20203 29191 20362 29243
rect 20414 29191 20573 29243
rect 20625 29191 20784 29243
rect 20836 29191 21313 29243
rect 20112 28813 21313 29191
rect 21421 29728 22236 29819
rect 21421 29672 21458 29728
rect 21514 29672 21669 29728
rect 21725 29672 21880 29728
rect 21936 29672 22091 29728
rect 22147 29672 22236 29728
rect 21421 28813 22236 29672
rect 22365 29245 23338 29284
rect 22365 29189 22402 29245
rect 22458 29189 22613 29245
rect 22669 29189 22824 29245
rect 22880 29189 23035 29245
rect 23091 29189 23246 29245
rect 23302 29189 23338 29245
rect 22365 29151 23338 29189
rect 23549 28813 25677 29876
rect 12040 28699 12639 28772
rect 8561 -21 8691 112
rect 12841 -164 12971 -31
rect 13219 -164 13348 -31
rect 13597 -164 13726 -31
rect 13974 -164 14104 -31
rect 14352 -164 14481 -31
rect 14730 -164 14859 -31
rect 16882 -164 17011 -31
rect 17260 -164 17389 -31
rect 17637 -164 17767 -31
rect 18015 -164 18144 -31
rect 18393 -164 18522 -31
rect 18770 -164 18900 -31
rect 19148 -164 19277 -31
rect 19526 -164 19655 -31
<< via2 >>
rect 5611 29672 5667 29728
rect 5822 29672 5878 29728
rect 6033 29672 6089 29728
rect 6244 29672 6300 29728
rect 4371 29245 4427 29247
rect 4371 29193 4373 29245
rect 4373 29193 4425 29245
rect 4425 29193 4427 29245
rect 4371 29191 4427 29193
rect 4582 29245 4638 29247
rect 4582 29193 4584 29245
rect 4584 29193 4636 29245
rect 4636 29193 4638 29245
rect 4582 29191 4638 29193
rect 4793 29245 4849 29247
rect 4793 29193 4795 29245
rect 4795 29193 4847 29245
rect 4847 29193 4849 29245
rect 4793 29191 4849 29193
rect 5004 29245 5060 29247
rect 5004 29193 5006 29245
rect 5006 29193 5058 29245
rect 5058 29193 5060 29245
rect 5004 29191 5060 29193
rect 5215 29245 5271 29247
rect 5215 29193 5217 29245
rect 5217 29193 5269 29245
rect 5269 29193 5271 29245
rect 5215 29191 5271 29193
rect 8222 29189 8278 29245
rect 8433 29189 8489 29245
rect 8644 29189 8700 29245
rect 8855 29189 8911 29245
rect 11573 29679 11575 29728
rect 11575 29679 11627 29728
rect 11627 29679 11629 29728
rect 11573 29672 11629 29679
rect 11753 29679 11755 29728
rect 11755 29679 11807 29728
rect 11807 29679 11809 29728
rect 11753 29672 11809 29679
rect 12331 29243 12387 29245
rect 12331 29191 12333 29243
rect 12333 29191 12385 29243
rect 12385 29191 12387 29243
rect 12331 29189 12387 29191
rect 12542 29243 12598 29245
rect 12542 29191 12544 29243
rect 12544 29191 12596 29243
rect 12596 29191 12598 29243
rect 12542 29189 12598 29191
rect 12753 29243 12809 29245
rect 12753 29191 12755 29243
rect 12755 29191 12807 29243
rect 12807 29191 12809 29243
rect 12753 29189 12809 29191
rect 12964 29243 13020 29245
rect 12964 29191 12966 29243
rect 12966 29191 13018 29243
rect 13018 29191 13020 29243
rect 12964 29189 13020 29191
rect 13175 29243 13231 29245
rect 13175 29191 13177 29243
rect 13177 29191 13229 29243
rect 13229 29191 13231 29243
rect 13175 29189 13231 29191
rect 13385 29243 13441 29245
rect 13385 29191 13387 29243
rect 13387 29191 13439 29243
rect 13439 29191 13441 29243
rect 13385 29189 13441 29191
rect 14031 29182 14087 29238
rect 14242 29182 14298 29238
rect 14453 29182 14509 29238
rect 12100 28772 12156 28828
rect 12311 28772 12367 28828
rect 12522 28772 12578 28828
rect 21458 29672 21514 29728
rect 21669 29672 21725 29728
rect 21880 29672 21936 29728
rect 22091 29672 22147 29728
rect 22402 29243 22458 29245
rect 22402 29191 22404 29243
rect 22404 29191 22456 29243
rect 22456 29191 22458 29243
rect 22402 29189 22458 29191
rect 22613 29243 22669 29245
rect 22613 29191 22615 29243
rect 22615 29191 22667 29243
rect 22667 29191 22669 29243
rect 22613 29189 22669 29191
rect 22824 29243 22880 29245
rect 22824 29191 22826 29243
rect 22826 29191 22878 29243
rect 22878 29191 22880 29243
rect 22824 29189 22880 29191
rect 23035 29243 23091 29245
rect 23035 29191 23037 29243
rect 23037 29191 23089 29243
rect 23089 29191 23091 29243
rect 23035 29189 23091 29191
rect 23246 29243 23302 29245
rect 23246 29191 23248 29243
rect 23248 29191 23300 29243
rect 23300 29191 23302 29243
rect 23246 29189 23302 29191
<< metal3 >>
rect 69 29633 199 29767
rect 1725 29728 25945 29801
rect 1725 29672 5611 29728
rect 5667 29672 5822 29728
rect 5878 29672 6033 29728
rect 6089 29672 6244 29728
rect 6300 29672 11573 29728
rect 11629 29672 11753 29728
rect 11809 29672 21458 29728
rect 21514 29672 21669 29728
rect 21725 29672 21880 29728
rect 21936 29672 22091 29728
rect 22147 29672 25945 29728
rect 1725 29599 25945 29672
rect -1 29173 128 29307
rect 1725 29247 5307 29341
rect 1725 29191 4371 29247
rect 4427 29191 4582 29247
rect 4638 29191 4793 29247
rect 4849 29191 5004 29247
rect 5060 29191 5215 29247
rect 5271 29191 5307 29247
rect 1725 29139 5307 29191
rect 8186 29245 13478 29284
rect 8186 29189 8222 29245
rect 8278 29189 8433 29245
rect 8489 29189 8644 29245
rect 8700 29189 8855 29245
rect 8911 29189 12331 29245
rect 12387 29189 12542 29245
rect 12598 29189 12753 29245
rect 12809 29189 12964 29245
rect 13020 29189 13175 29245
rect 13231 29189 13385 29245
rect 13441 29189 13478 29245
rect 13994 29238 14545 29277
rect 13994 29203 14031 29238
rect 8186 29150 13478 29189
rect 13993 29182 14031 29203
rect 14087 29182 14242 29238
rect 14298 29182 14453 29238
rect 14509 29182 14545 29238
rect 13993 29144 14545 29182
rect 22365 29245 25945 29341
rect 22365 29189 22402 29245
rect 22458 29189 22613 29245
rect 22669 29189 22824 29245
rect 22880 29189 23035 29245
rect 23091 29189 23246 29245
rect 23302 29189 25945 29245
rect 69 28733 199 28867
rect 12063 28828 12615 28867
rect 13993 28832 14092 29144
rect 22365 29139 25945 29189
rect 27640 29173 27769 29307
rect 12063 28772 12100 28828
rect 12156 28772 12311 28828
rect 12367 28772 12522 28828
rect 12578 28772 12615 28828
rect 12063 28733 12615 28772
rect -1 28273 128 28407
rect 27640 28273 27769 28407
rect -1 27393 128 27527
rect 27640 27393 27769 27527
rect -1 26473 128 26607
rect 27640 26473 27769 26607
rect -1 25593 128 25727
rect 27640 25593 27769 25727
rect -1 24673 128 24807
rect 27640 24673 27769 24807
rect -1 23793 128 23927
rect 27640 23793 27769 23927
rect -1 22873 128 23007
rect 27640 22873 27769 23007
rect -1 21993 128 22127
rect 27640 21993 27769 22127
rect -1 21073 128 21207
rect 27640 21073 27769 21207
rect -1 20193 128 20327
rect 27640 20193 27769 20327
rect -1 19273 128 19407
rect 27640 19273 27769 19407
rect -1 18393 128 18527
rect 27640 18393 27769 18527
rect -1 17473 128 17607
rect 27640 17473 27769 17607
rect -1 16593 128 16727
rect 27640 16593 27769 16727
rect -1 15673 128 15807
rect 27640 15673 27769 15807
rect -1 14793 128 14927
rect 27640 14793 27769 14927
rect -1 13873 128 14007
rect 27640 13873 27769 14007
rect -1 12993 128 13127
rect 27640 12993 27769 13127
rect -1 12073 128 12207
rect 27640 12073 27769 12207
rect -1 11193 128 11327
rect 27640 11193 27769 11327
rect -1 10273 128 10407
rect 27640 10273 27769 10407
rect -1 9393 128 9527
rect 27640 9393 27769 9527
rect -1 8473 128 8607
rect 27640 8473 27769 8607
rect -1 7593 128 7727
rect 27640 7593 27769 7727
rect -1 6673 128 6807
rect 27640 6673 27769 6807
rect -1 5793 128 5927
rect 27640 5793 27769 5927
rect -1 4873 128 5007
rect 27640 4873 27769 5007
rect -1 3993 128 4127
rect 27640 3993 27769 4127
rect -1 3073 128 3207
rect 27640 3073 27769 3207
rect -1 2193 128 2327
rect 27640 2193 27769 2327
rect -1 1273 128 1407
rect 27640 1273 27769 1407
rect -1 393 128 527
rect 27640 393 27769 527
use M1_NACTIVE$$203393068_256x8m81  M1_NACTIVE$$203393068_256x8m81_0
timestamp 1669390400
transform 1 0 14063 0 1 29759
box 0 0 1 1
use M1_NWELL$$204218412_256x8m81  M1_NWELL$$204218412_256x8m81_0
timestamp 1669390400
transform -1 0 25568 0 1 29686
box -221 -717 1960 228
use M1_NWELL$$204218412_256x8m81  M1_NWELL$$204218412_256x8m81_1
timestamp 1669390400
transform 1 0 2200 0 1 29686
box -221 -717 1960 228
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_0
timestamp 1669390400
transform 1 0 11463 0 1 29759
box -78 -80 1817 80
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_1
timestamp 1669390400
transform 1 0 21475 0 1 29759
box -78 -80 1817 80
use M1_PACTIVE$$204148780_256x8m81  M1_PACTIVE$$204148780_256x8m81_2
timestamp 1669390400
transform 1 0 4390 0 1 29759
box -78 -80 1817 80
use M1_PACTIVE$$204149804_256x8m81  M1_PACTIVE$$204149804_256x8m81_0
timestamp 1669390400
transform 1 0 15860 0 1 29759
box 0 0 1 1
use M1_POLY2$$204150828_256x8m81  M1_POLY2$$204150828_256x8m81_0
timestamp 1669390400
transform 1 0 9381 0 1 29448
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1669390400
transform 1 0 15413 0 1 29741
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1669390400
transform 0 -1 13712 1 0 29693
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_1
timestamp 1669390400
transform 1 0 15625 0 1 29401
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_2
timestamp 1669390400
transform 1 0 18313 0 1 29436
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_3
timestamp 1669390400
transform 1 0 12040 0 1 29361
box 0 0 1 1
use M2_M1$$201262124_256x8m81  M2_M1$$201262124_256x8m81_0
timestamp 1669390400
transform 1 0 13701 0 1 29691
box 0 0 1 1
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_0
timestamp 1669390400
transform 1 0 10402 0 1 29448
box 0 0 1 1
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_1
timestamp 1669390400
transform 1 0 14059 0 1 29752
box 0 0 1 1
use M2_M1$$204139564_256x8m81  M2_M1$$204139564_256x8m81_0
timestamp 1669390400
transform 1 0 11601 0 1 29705
box 0 0 1 1
use M2_M1$$204140588_256x8m81  M2_M1$$204140588_256x8m81_0
timestamp 1669390400
transform 1 0 12359 0 1 29217
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_0
timestamp 1669390400
transform 1 0 15126 0 1 29752
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_1
timestamp 1669390400
transform 1 0 20177 0 1 29680
box 0 0 1 1
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_2
timestamp 1669390400
transform 1 0 20177 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_0
timestamp 1669390400
transform 1 0 6792 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_1
timestamp 1669390400
transform 1 0 22430 0 1 29217
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_2
timestamp 1669390400
transform 1 0 4399 0 1 29219
box 0 0 1 1
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_3
timestamp 1669390400
transform 1 0 6792 0 1 29680
box 0 0 1 1
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_0
timestamp 1669390400
transform -1 0 25612 0 1 29700
box -65 -502 1751 67
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_1
timestamp 1669390400
transform 1 0 2156 0 1 29700
box -65 -502 1751 67
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_0
timestamp 1669390400
transform 1 0 21486 0 1 29700
box -65 -284 697 67
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_1
timestamp 1669390400
transform 1 0 5639 0 1 29700
box -65 -284 697 67
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_0
timestamp 1669390400
transform 1 0 5639 0 1 29700
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_1
timestamp 1669390400
transform 1 0 8250 0 1 29217
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_2
timestamp 1669390400
transform 1 0 21486 0 1 29700
box 0 0 1 1
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_3
timestamp 1669390400
transform 1 0 21486 0 1 29700
box 0 0 1 1
use M3_M2$$204143660_256x8m81  M3_M2$$204143660_256x8m81_0
timestamp 1669390400
transform 1 0 11601 0 1 29700
box 0 0 1 1
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_0
timestamp 1669390400
transform 1 0 22430 0 1 29217
box 0 0 1 1
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_1
timestamp 1669390400
transform 1 0 4399 0 1 29219
box 0 0 1 1
use M3_M2$$204145708_256x8m81  M3_M2$$204145708_256x8m81_0
timestamp 1669390400
transform 1 0 12359 0 1 29217
box 0 0 1 1
use M3_M2$$204146732_256x8m81  M3_M2$$204146732_256x8m81_0
timestamp 1669390400
transform 1 0 14059 0 1 29210
box 0 0 1 1
use M3_M2$$204147756_256x8m81  M3_M2$$204147756_256x8m81_0
timestamp 1669390400
transform 1 0 12339 0 1 28800
box 0 0 1 1
use nmos_1p2$$204213292_R90_256x8m81  nmos_1p2$$204213292_R90_256x8m81_0
timestamp 1669390400
transform 0 -1 6346 1 0 29303
box -119 -71 177 2091
use nmos_1p2$$204215340_256x8m81  nmos_1p2$$204215340_256x8m81_0
timestamp 1669390400
transform 0 -1 13604 -1 0 29362
box -119 -71 177 1389
use nmos_5p04310590878199_256x8m81  nmos_5p04310590878199_256x8m81_0
timestamp 1669390400
transform 0 -1 23346 1 0 29272
box -88 -44 208 2066
use nmos_5p043105908781111_256x8m81  nmos_5p043105908781111_256x8m81_0
timestamp 1669390400
transform 0 -1 16283 1 0 29272
box -88 -44 208 572
use nmos_5p043105908781111_256x8m81  nmos_5p043105908781111_256x8m81_1
timestamp 1669390400
transform 0 -1 11913 1 0 29272
box -88 -44 208 572
use pmos_1p2$$204216364_256x8m81  pmos_1p2$$204216364_256x8m81_0
timestamp 1669390400
transform 0 -1 20950 1 0 29303
box -296 -137 586 2646
use pmos_1p2$$204216364_256x8m81  pmos_1p2$$204216364_256x8m81_1
timestamp 1669390400
transform 0 -1 9245 1 0 29303
box -296 -137 586 2646
use pmos_1p2$$204217388_256x8m81  pmos_1p2$$204217388_256x8m81_0
timestamp 1669390400
transform 0 -1 11004 1 0 29303
box -295 -137 355 1454
use pmos_5p043105908781101_256x8m81  pmos_5p043105908781101_256x8m81_0
timestamp 1669390400
transform 0 -1 15304 1 0 29272
box -208 -120 328 1438
use pmos_5p043105908781101_256x8m81  pmos_5p043105908781101_256x8m81_1
timestamp 1669390400
transform 0 -1 17974 1 0 29272
box -208 -120 328 1438
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_0
timestamp 1669390400
transform 0 -1 2203 -1 0 28950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_1
timestamp 1669390400
transform 0 -1 2203 -1 0 27150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_2
timestamp 1669390400
transform 0 -1 2203 -1 0 25350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_3
timestamp 1669390400
transform 0 -1 2203 -1 0 23550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_4
timestamp 1669390400
transform 0 -1 2203 -1 0 21750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_5
timestamp 1669390400
transform 0 -1 2203 -1 0 19950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_6
timestamp 1669390400
transform 0 -1 2203 -1 0 18150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_7
timestamp 1669390400
transform 0 -1 2203 -1 0 16350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_8
timestamp 1669390400
transform 0 -1 2203 -1 0 14550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_9
timestamp 1669390400
transform 0 -1 2203 -1 0 12750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_10
timestamp 1669390400
transform 0 -1 2203 -1 0 10950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_11
timestamp 1669390400
transform 0 -1 2203 -1 0 9150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_12
timestamp 1669390400
transform 0 -1 2203 -1 0 7350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_13
timestamp 1669390400
transform 0 -1 2203 -1 0 5550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_14
timestamp 1669390400
transform 0 -1 2203 -1 0 3750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_15
timestamp 1669390400
transform 0 -1 2203 -1 0 1950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_16
timestamp 1669390400
transform 0 1 25566 -1 0 28950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_17
timestamp 1669390400
transform 0 1 25566 -1 0 27150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_18
timestamp 1669390400
transform 0 1 25566 -1 0 25350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_19
timestamp 1669390400
transform 0 1 25566 -1 0 23550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_20
timestamp 1669390400
transform 0 1 25566 -1 0 21750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_21
timestamp 1669390400
transform 0 1 25566 -1 0 19950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_22
timestamp 1669390400
transform 0 1 25566 -1 0 18150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_23
timestamp 1669390400
transform 0 1 25566 -1 0 16350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_24
timestamp 1669390400
transform 0 1 25566 -1 0 14550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_25
timestamp 1669390400
transform 0 1 25566 -1 0 12750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_26
timestamp 1669390400
transform 0 1 25566 -1 0 10950
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_27
timestamp 1669390400
transform 0 1 25566 -1 0 9150
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_28
timestamp 1669390400
transform 0 1 25566 -1 0 7350
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_29
timestamp 1669390400
transform 0 1 25566 -1 0 5550
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_30
timestamp 1669390400
transform 0 1 25566 -1 0 3750
box -60 -407 2159 6582
use pmoscap_W2_5_477_R270_256x8m81  pmoscap_W2_5_477_R270_256x8m81_31
timestamp 1669390400
transform 0 1 25566 -1 0 1950
box -60 -407 2159 6582
use pmoscap_W2_5_R270_256x8m81  pmoscap_W2_5_R270_256x8m81_0
timestamp 1669390400
transform 0 -1 2203 -1 0 29850
box -60 -407 1259 3251
use pmoscap_W2_5_R270_256x8m81  pmoscap_W2_5_R270_256x8m81_1
timestamp 1669390400
transform 0 1 25566 -1 0 29850
box -60 -407 1259 3251
use xdec32_256x8m81  xdec32_256x8m81_0
timestamp 1669390400
transform 1 0 1726 0 1 0
box 0 -228 24219 29028
<< labels >>
rlabel metal3 s 27705 29240 27705 29240 4 DRWL
port 1 nsew
rlabel metal3 s 27705 28340 27705 28340 4 RWL[31]
port 2 nsew
rlabel metal3 s 27705 27460 27705 27460 4 RWL[30]
port 3 nsew
rlabel metal3 s 27705 26540 27705 26540 4 RWL[29]
port 4 nsew
rlabel metal3 s 27705 25660 27705 25660 4 RWL[28]
port 5 nsew
rlabel metal3 s 27705 24740 27705 24740 4 RWL[27]
port 6 nsew
rlabel metal3 s 27705 23860 27705 23860 4 RWL[26]
port 7 nsew
rlabel metal3 s 27705 22940 27705 22940 4 RWL[25]
port 8 nsew
rlabel metal3 s 27705 22060 27705 22060 4 RWL[24]
port 9 nsew
rlabel metal3 s 27705 21140 27705 21140 4 RWL[23]
port 10 nsew
rlabel metal3 s 27705 20260 27705 20260 4 RWL[22]
port 11 nsew
rlabel metal3 s 27705 19340 27705 19340 4 RWL[21]
port 12 nsew
rlabel metal3 s 27705 5860 27705 5860 4 RWL[6]
port 13 nsew
rlabel metal3 s 27705 4060 27705 4060 4 RWL[4]
port 14 nsew
rlabel metal3 s 27705 2260 27705 2260 4 RWL[2]
port 15 nsew
rlabel metal3 s 27705 460 27705 460 4 RWL[0]
port 16 nsew
rlabel metal3 s 27705 1340 27705 1340 4 RWL[1]
port 17 nsew
rlabel metal3 s 27705 3140 27705 3140 4 RWL[3]
port 18 nsew
rlabel metal3 s 27705 4940 27705 4940 4 RWL[5]
port 19 nsew
rlabel metal3 s 27705 6740 27705 6740 4 RWL[7]
port 20 nsew
rlabel metal3 s 27705 7660 27705 7660 4 RWL[8]
port 21 nsew
rlabel metal3 s 27705 8540 27705 8540 4 RWL[9]
port 22 nsew
rlabel metal3 s 27705 9460 27705 9460 4 RWL[10]
port 23 nsew
rlabel metal3 s 27705 10340 27705 10340 4 RWL[11]
port 24 nsew
rlabel metal3 s 27705 11260 27705 11260 4 RWL[12]
port 25 nsew
rlabel metal3 s 27705 12140 27705 12140 4 RWL[13]
port 26 nsew
rlabel metal3 s 27705 13060 27705 13060 4 RWL[14]
port 27 nsew
rlabel metal3 s 27705 13940 27705 13940 4 RWL[15]
port 28 nsew
rlabel metal3 s 27705 14860 27705 14860 4 RWL[16]
port 29 nsew
rlabel metal3 s 27705 15740 27705 15740 4 RWL[17]
port 30 nsew
rlabel metal3 s 27705 16660 27705 16660 4 RWL[18]
port 31 nsew
rlabel metal3 s 27705 17540 27705 17540 4 RWL[19]
port 32 nsew
rlabel metal3 s 27705 18460 27705 18460 4 RWL[20]
port 33 nsew
rlabel metal3 s 64 26540 64 26540 4 LWL[29]
port 34 nsew
rlabel metal3 s 64 27460 64 27460 4 LWL[30]
port 35 nsew
rlabel metal3 s 64 28340 64 28340 4 LWL[31]
port 36 nsew
rlabel metal3 s 64 17540 64 17540 4 LWL[19]
port 37 nsew
rlabel metal3 s 64 18460 64 18460 4 LWL[20]
port 38 nsew
rlabel metal3 s 64 19340 64 19340 4 LWL[21]
port 39 nsew
rlabel metal3 s 64 20260 64 20260 4 LWL[22]
port 40 nsew
rlabel metal3 s 64 21140 64 21140 4 LWL[23]
port 41 nsew
rlabel metal3 s 64 22060 64 22060 4 LWL[24]
port 42 nsew
rlabel metal3 s 64 22940 64 22940 4 LWL[25]
port 43 nsew
rlabel metal3 s 64 23860 64 23860 4 LWL[26]
port 44 nsew
rlabel metal3 s 64 24740 64 24740 4 LWL[27]
port 45 nsew
rlabel metal3 s 64 25660 64 25660 4 LWL[28]
port 46 nsew
rlabel metal3 s 64 9460 64 9460 4 LWL[10]
port 47 nsew
rlabel metal3 s 64 10340 64 10340 4 LWL[11]
port 48 nsew
rlabel metal3 s 64 11260 64 11260 4 LWL[12]
port 49 nsew
rlabel metal3 s 64 12140 64 12140 4 LWL[13]
port 50 nsew
rlabel metal3 s 64 13060 64 13060 4 LWL[14]
port 51 nsew
rlabel metal3 s 64 13940 64 13940 4 LWL[15]
port 52 nsew
rlabel metal3 s 64 14860 64 14860 4 LWL[16]
port 53 nsew
rlabel metal3 s 64 15740 64 15740 4 LWL[17]
port 54 nsew
rlabel metal3 s 64 16660 64 16660 4 LWL[18]
port 55 nsew
rlabel metal3 s 64 4940 64 4940 4 LWL[5]
port 56 nsew
rlabel metal3 s 64 4060 64 4060 4 LWL[4]
port 57 nsew
rlabel metal3 s 64 3140 64 3140 4 LWL[3]
port 58 nsew
rlabel metal3 s 64 2260 64 2260 4 LWL[2]
port 59 nsew
rlabel metal3 s 64 1340 64 1340 4 LWL[1]
port 60 nsew
rlabel metal3 s 64 460 64 460 4 LWL[0]
port 61 nsew
rlabel metal3 s 64 7660 64 7660 4 LWL[8]
port 62 nsew
rlabel metal3 s 64 8540 64 8540 4 LWL[9]
port 63 nsew
rlabel metal3 s 64 5860 64 5860 4 LWL[6]
port 64 nsew
rlabel metal3 s 64 6740 64 6740 4 LWL[7]
port 65 nsew
rlabel metal3 s 134 29700 134 29700 4 vss
port 66 nsew
rlabel metal3 s 134 28800 134 28800 4 vdd
port 67 nsew
rlabel metal3 s 64 29240 64 29240 4 DLWL
port 68 nsew
rlabel metal2 s 14794 -97 14794 -97 4 xb[0]
port 69 nsew
rlabel metal2 s 14417 -97 14417 -97 4 xb[1]
port 70 nsew
rlabel metal2 s 14039 -97 14039 -97 4 xb[2]
port 71 nsew
rlabel metal2 s 13661 -97 13661 -97 4 xb[3]
port 72 nsew
rlabel metal2 s 16947 -97 16947 -97 4 xa[7]
port 73 nsew
rlabel metal2 s 17324 -97 17324 -97 4 xa[6]
port 74 nsew
rlabel metal2 s 17702 -97 17702 -97 4 xa[5]
port 75 nsew
rlabel metal2 s 18080 -97 18080 -97 4 xa[4]
port 76 nsew
rlabel metal2 s 19591 -97 19591 -97 4 xa[0]
port 77 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 78 nsew
rlabel metal2 s 18457 -97 18457 -97 4 xa[3]
port 79 nsew
rlabel metal2 s 18835 -97 18835 -97 4 xa[2]
port 80 nsew
rlabel metal2 s 19213 -97 19213 -97 4 xa[1]
port 81 nsew
rlabel metal2 s 13284 -97 13284 -97 4 xc[0]
port 82 nsew
rlabel metal2 s 12906 -97 12906 -97 4 xc[1]
port 83 nsew
<< properties >>
string GDS_END 2364906
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2346134
<< end >>
