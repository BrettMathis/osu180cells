magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 918 6384 1098
rect 301 769 347 918
rect 972 874 1040 918
rect 1380 874 1448 918
rect 1788 874 1856 918
rect 2256 874 2324 918
rect 2700 881 2768 918
rect 3108 881 3176 918
rect 3516 881 3584 918
rect 3924 881 3992 918
rect 4332 881 4400 918
rect 4740 881 4808 918
rect 5148 881 5216 918
rect 5556 881 5624 918
rect 2904 673 5818 835
rect 5975 776 6021 918
rect 109 466 315 542
rect 1060 430 2425 542
rect 5706 330 5818 673
rect 5706 327 6101 330
rect 2919 173 6101 327
rect 273 90 319 139
rect 854 90 922 125
rect 1340 90 1408 127
rect 1788 90 1856 127
rect 2236 90 2304 127
rect 2681 90 2756 127
rect 3132 90 3200 127
rect 3580 90 3648 127
rect 4028 90 4096 127
rect 4476 90 4544 127
rect 4924 90 4992 127
rect 5372 90 5440 127
rect 5820 90 5888 127
rect 6279 90 6325 232
rect 0 -90 6384 90
<< obsm1 >>
rect 97 634 143 750
rect 585 689 2540 828
rect 881 666 2540 689
rect 97 588 719 634
rect 361 320 407 588
rect 673 483 719 588
rect 789 437 835 643
rect 38 274 407 320
rect 629 391 835 437
rect 629 298 675 391
rect 881 331 927 666
rect 2471 551 2540 666
rect 2471 494 5524 551
rect 497 217 675 298
rect 721 263 927 331
rect 2771 373 5555 432
rect 2771 330 2829 373
rect 1127 217 2829 330
rect 497 173 2829 217
rect 497 171 1173 173
rect 497 136 543 171
<< labels >>
rlabel metal1 s 109 466 315 542 6 EN
port 1 nsew default input
rlabel metal1 s 1060 430 2425 542 6 I
port 2 nsew default input
rlabel metal1 s 2904 673 5818 835 6 Z
port 3 nsew default output
rlabel metal1 s 5706 330 5818 673 6 Z
port 3 nsew default output
rlabel metal1 s 5706 327 6101 330 6 Z
port 3 nsew default output
rlabel metal1 s 2919 173 6101 327 6 Z
port 3 nsew default output
rlabel metal1 s 0 918 6384 1098 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5975 881 6021 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5556 881 5624 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5148 881 5216 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4740 881 4808 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4332 881 4400 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3924 881 3992 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3516 881 3584 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3108 881 3176 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2700 881 2768 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2256 881 2324 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1788 881 1856 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1380 881 1448 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 972 881 1040 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 881 347 918 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5975 874 6021 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2256 874 2324 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1788 874 1856 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1380 874 1448 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 972 874 1040 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 874 347 881 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5975 776 6021 874 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 776 347 874 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 301 769 347 776 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6279 139 6325 232 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6279 127 6325 139 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 139 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6279 125 6325 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5820 125 5888 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5372 125 5440 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4924 125 4992 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4476 125 4544 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4028 125 4096 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3580 125 3648 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3132 125 3200 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2681 125 2756 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2236 125 2304 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1788 125 1856 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1340 125 1408 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6279 90 6325 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5820 90 5888 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5372 90 5440 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4924 90 4992 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4476 90 4544 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4028 90 4096 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3580 90 3648 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3132 90 3200 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2681 90 2756 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2236 90 2304 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1788 90 1856 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1340 90 1408 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 854 90 922 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 6384 90 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6384 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1354310
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1341602
<< end >>
