magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 6048 844
rect 252 569 320 724
rect 1075 577 1121 724
rect 1518 670 1586 724
rect 2602 689 2670 724
rect 3240 689 3312 724
rect 141 119 206 430
rect 273 60 319 228
rect 365 119 430 430
rect 682 353 878 431
rect 1026 353 1326 431
rect 1110 60 1156 205
rect 1573 60 1619 209
rect 4093 583 4139 724
rect 2756 60 2828 183
rect 4121 242 4228 438
rect 4526 594 4594 724
rect 4498 353 4686 431
rect 4953 506 4999 724
rect 5157 531 5236 676
rect 5361 600 5407 724
rect 5517 531 5617 676
rect 5769 600 5815 724
rect 5157 477 5908 531
rect 5851 307 5908 477
rect 4372 60 4440 215
rect 5170 241 5908 307
rect 5011 60 5057 185
rect 5170 122 5287 241
rect 5459 60 5505 185
rect 5627 122 5739 241
rect 5907 60 5953 185
rect 0 -60 6048 60
<< obsm1 >>
rect 49 523 95 608
rect 654 549 824 595
rect 1217 632 1472 678
rect 778 531 824 549
rect 1217 531 1263 632
rect 1426 624 1472 632
rect 1641 632 1967 678
rect 2253 643 2556 678
rect 2716 643 3194 678
rect 3358 643 3655 678
rect 2253 632 3655 643
rect 1641 624 1687 632
rect 1426 578 1687 624
rect 49 477 571 523
rect 778 484 1263 531
rect 1322 524 1368 578
rect 1322 477 1707 524
rect 49 156 95 477
rect 525 307 571 477
rect 926 307 972 350
rect 525 261 972 307
rect 1018 252 1248 298
rect 1389 257 1435 477
rect 1661 382 1707 477
rect 1777 407 1823 578
rect 1921 477 1967 632
rect 2510 597 2762 632
rect 3148 597 3404 632
rect 2160 459 2206 574
rect 2336 551 2440 555
rect 2832 551 2920 556
rect 2336 505 2920 551
rect 2992 551 3080 556
rect 3472 551 3558 556
rect 2992 505 3558 551
rect 2160 413 3181 459
rect 1777 360 2079 407
rect 1018 215 1064 252
rect 650 169 1064 215
rect 1202 152 1248 252
rect 1367 198 1435 257
rect 1481 259 1736 306
rect 1481 152 1527 259
rect 1202 106 1527 152
rect 1690 152 1736 259
rect 1830 198 1898 360
rect 1985 152 2031 196
rect 1690 106 2031 152
rect 2209 124 2255 413
rect 3265 367 3333 505
rect 3609 407 3655 632
rect 3705 632 4047 678
rect 2325 275 2371 340
rect 2459 321 3333 367
rect 3705 361 3751 632
rect 3909 445 3955 567
rect 4001 537 4047 632
rect 4185 632 4463 678
rect 4185 537 4231 632
rect 4001 491 4231 537
rect 2325 229 2920 275
rect 2874 152 2920 229
rect 3265 198 3333 321
rect 3388 152 3434 349
rect 3489 315 3751 361
rect 3797 399 4037 445
rect 3489 198 3557 315
rect 3797 244 3843 399
rect 3714 198 3843 244
rect 3889 152 3935 353
rect 2874 106 3935 152
rect 3991 192 4037 399
rect 4286 431 4354 586
rect 4416 548 4463 632
rect 4640 632 4898 678
rect 4640 548 4686 632
rect 4416 502 4686 548
rect 4280 385 4354 431
rect 4280 192 4326 385
rect 4402 307 4448 440
rect 4738 307 4806 586
rect 4852 382 4898 632
rect 4989 365 5745 419
rect 4989 307 5035 365
rect 4402 261 5035 307
rect 3991 143 4326 192
rect 4867 131 4913 261
<< labels >>
rlabel metal1 s 682 353 878 431 6 D
port 1 nsew default input
rlabel metal1 s 4498 353 4686 431 6 RN
port 2 nsew default input
rlabel metal1 s 141 119 206 430 6 SE
port 3 nsew default input
rlabel metal1 s 4121 242 4228 438 6 SETN
port 4 nsew default input
rlabel metal1 s 365 119 430 430 6 SI
port 5 nsew default input
rlabel metal1 s 1026 353 1326 431 6 CLK
port 6 nsew clock input
rlabel metal1 s 5517 531 5617 676 6 Q
port 7 nsew default output
rlabel metal1 s 5157 531 5236 676 6 Q
port 7 nsew default output
rlabel metal1 s 5157 477 5908 531 6 Q
port 7 nsew default output
rlabel metal1 s 5851 307 5908 477 6 Q
port 7 nsew default output
rlabel metal1 s 5170 241 5908 307 6 Q
port 7 nsew default output
rlabel metal1 s 5627 122 5739 241 6 Q
port 7 nsew default output
rlabel metal1 s 5170 122 5287 241 6 Q
port 7 nsew default output
rlabel metal1 s 0 724 6048 844 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5769 689 5815 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5361 689 5407 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 689 4999 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 689 4594 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 689 4139 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3240 689 3312 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2602 689 2670 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1518 689 1586 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 689 1121 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 689 320 724 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5769 670 5815 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5361 670 5407 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 670 4999 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 670 4594 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 670 4139 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1518 670 1586 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 670 1121 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 689 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5769 600 5815 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5361 600 5407 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 600 4999 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 600 4594 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 600 4139 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 600 1121 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 600 320 670 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 594 4999 600 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 594 4594 600 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 594 4139 600 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 594 1121 600 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 594 320 600 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 583 4999 594 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 583 4139 594 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 583 1121 594 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 583 320 594 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 577 4999 583 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 577 1121 583 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 577 320 583 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 569 4999 577 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 577 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4953 506 4999 569 6 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 273 215 319 228 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 209 4440 215 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 209 319 215 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 205 4440 209 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 205 1619 209 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 205 319 209 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 185 4440 205 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 185 1619 205 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 185 1156 205 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 185 319 205 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5907 183 5953 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5459 183 5505 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5011 183 5057 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 183 4440 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 183 1619 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 183 1156 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 185 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5907 60 5953 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5459 60 5505 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5011 60 5057 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 60 4440 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2756 60 2828 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 60 1619 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 60 1156 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6048 60 8 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6048 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 275880
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 263098
<< end >>
