* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_addf_1 A B CI CO S
X0 a_110_109 A VDD VDD pmos_3p3 w=34 l=6
X1 S a_161_19 VDD VDD pmos_3p3 w=34 l=6
X2 S a_161_19 VSS VSS nmos_3p3 w=17 l=6
X3 VDD CI a_195_109 VDD pmos_3p3 w=34 l=6
X4 a_195_19 B a_178_19 VSS nmos_3p3 w=17 l=6
X5 a_76_109 B a_59_19 VDD pmos_3p3 w=34 l=6
X6 VDD A a_76_109 VDD pmos_3p3 w=34 l=6
X7 a_59_19 CI a_9_109 VDD pmos_3p3 w=34 l=6
X8 a_178_19 A a_161_19 VSS nmos_3p3 w=17 l=6
X9 a_9_109 B VDD VDD pmos_3p3 w=34 l=6
X10 a_110_19 CI VSS VSS nmos_3p3 w=17 l=6
X11 VDD A a_9_109 VDD pmos_3p3 w=34 l=6
X12 a_59_19 CI a_9_19 VSS nmos_3p3 w=17 l=6
X13 VSS B a_110_19 VSS nmos_3p3 w=17 l=6
X14 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X15 CO a_59_19 VSS VSS nmos_3p3 w=17 l=6
X16 VSS CI a_195_19 VSS nmos_3p3 w=17 l=6
X17 CO a_59_19 VDD VDD pmos_3p3 w=34 l=6
X18 VSS A a_76_19 VSS nmos_3p3 w=17 l=6
X19 a_161_19 a_59_19 a_110_19 VSS nmos_3p3 w=17 l=6
X20 a_76_19 B a_59_19 VSS nmos_3p3 w=17 l=6
X21 a_178_109 A a_161_19 VDD pmos_3p3 w=34 l=6
X22 a_195_109 B a_178_109 VDD pmos_3p3 w=34 l=6
X23 a_9_19 B VSS VSS nmos_3p3 w=17 l=6
X24 a_110_19 A VSS VSS nmos_3p3 w=17 l=6
X25 a_161_19 a_59_19 a_110_109 VDD pmos_3p3 w=34 l=6
X26 VDD B a_110_109 VDD pmos_3p3 w=34 l=6
X27 a_110_109 CI VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_addh_1 A B S CO
X0 VDD B a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 A VDD VDD pmos_3p3 w=34 l=6
X2 VDD a_19_14 CO VDD pmos_3p3 w=34 l=6
X3 a_19_14 B a_42_19 VSS nmos_3p3 w=17 l=6
X4 S a_91_19 VSS VSS nmos_3p3 w=17 l=6
X5 VSS a_19_14 CO VSS nmos_3p3 w=17 l=6
X6 S a_91_19 VDD VDD pmos_3p3 w=34 l=6
X7 a_91_19 B a_91_109 VDD pmos_3p3 w=34 l=6
X8 VDD a_19_14 a_91_19 VDD pmos_3p3 w=34 l=6
X9 a_91_109 A VDD VDD pmos_3p3 w=34 l=6
X10 a_91_19 A a_75_19 VSS nmos_3p3 w=17 l=6
X11 a_42_19 A VSS VSS nmos_3p3 w=17 l=6
X12 VSS a_19_14 a_75_19 VSS nmos_3p3 w=17 l=6
X13 a_75_19 B a_91_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_and2_1 A B Y
X0 Y a_12_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD B a_12_19 VDD pmos_3p3 w=34 l=6
X2 a_12_19 A VDD VDD pmos_3p3 w=34 l=6
X3 Y a_12_19 VSS VSS nmos_3p3 w=17 l=6
X4 a_28_19 A a_12_19 VSS nmos_3p3 w=17 l=6
X5 VSS B a_28_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_aoi21_1 Y A0 A1 B
X0 Y B a_9_109 VDD pmos_3p3 w=34 l=6
X1 a_9_109 A1 VDD VDD pmos_3p3 w=34 l=6
X2 VDD A0 a_9_109 VDD pmos_3p3 w=34 l=6
X3 VSS B Y VSS nmos_3p3 w=17 l=6
X4 a_28_19 A0 VSS VSS nmos_3p3 w=17 l=6
X5 Y A1 a_28_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_1 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X2 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X3 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_2 A Y
X0 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X1 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X2 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X3 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X4 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X5 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_4 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X2 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X3 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X4 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X5 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X6 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X7 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X8 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X9 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_8 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X2 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X3 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X4 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X5 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X6 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X7 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X8 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X9 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X10 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X11 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X12 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X13 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X14 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X15 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X16 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X17 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_16 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X2 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X3 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X4 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X5 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X6 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X7 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X8 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X9 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X10 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X11 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X12 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X13 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X14 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X15 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X16 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X17 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X18 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X19 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X20 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X21 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X22 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X23 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X24 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X25 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X26 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X27 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X28 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X29 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X30 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X31 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X32 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X33 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
C0 VDD Y 2.051450fF
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_1 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X2 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X3 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_2 A Y
X0 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X1 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X2 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X3 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X4 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X5 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_4 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X2 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X3 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X4 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X5 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X6 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X7 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X8 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X9 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_8 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X2 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X3 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X4 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X5 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X6 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X7 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X8 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X9 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X10 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X11 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X12 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X13 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X14 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X15 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X16 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X17 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkbuf_16 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X2 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X3 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X4 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X5 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X6 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X7 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X8 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X9 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X10 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X11 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X12 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X13 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X14 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X15 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X16 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X17 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X18 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X19 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X20 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X21 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X22 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X23 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X24 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X25 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X26 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X27 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X28 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X29 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X30 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X31 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X32 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X33 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
C0 VDD Y 2.051450fF
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkinv_1 A Y
X0 Y A VDD VDD pmos_3p3 w=34 l=6
X1 Y A VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkinv_2 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 Y A VSS VSS nmos_3p3 w=17 l=6
X3 VSS A Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkinv_4 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 VDD A Y VDD pmos_3p3 w=34 l=6
X3 Y A VDD VDD pmos_3p3 w=34 l=6
X4 Y A VSS VSS nmos_3p3 w=17 l=6
X5 Y A VSS VSS nmos_3p3 w=17 l=6
X6 VSS A Y VSS nmos_3p3 w=17 l=6
X7 VSS A Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkinv_8 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 VDD A Y VDD pmos_3p3 w=34 l=6
X2 Y A VDD VDD pmos_3p3 w=34 l=6
X3 Y A VDD VDD pmos_3p3 w=34 l=6
X4 VDD A Y VDD pmos_3p3 w=34 l=6
X5 VSS A Y VSS nmos_3p3 w=17 l=6
X6 Y A VDD VDD pmos_3p3 w=34 l=6
X7 Y A VSS VSS nmos_3p3 w=17 l=6
X8 Y A VSS VSS nmos_3p3 w=17 l=6
X9 Y A VSS VSS nmos_3p3 w=17 l=6
X10 Y A VSS VSS nmos_3p3 w=17 l=6
X11 VSS A Y VSS nmos_3p3 w=17 l=6
X12 VSS A Y VSS nmos_3p3 w=17 l=6
X13 VSS A Y VSS nmos_3p3 w=17 l=6
X14 Y A VDD VDD pmos_3p3 w=34 l=6
X15 VDD A Y VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_clkinv_16 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 Y A VSS VSS nmos_3p3 w=17 l=6
X3 VDD A Y VDD pmos_3p3 w=34 l=6
X4 Y A VSS VSS nmos_3p3 w=17 l=6
X5 VDD A Y VDD pmos_3p3 w=34 l=6
X6 Y A VDD VDD pmos_3p3 w=34 l=6
X7 Y A VDD VDD pmos_3p3 w=34 l=6
X8 VSS A Y VSS nmos_3p3 w=17 l=6
X9 VDD A Y VDD pmos_3p3 w=34 l=6
X10 VSS A Y VSS nmos_3p3 w=17 l=6
X11 Y A VDD VDD pmos_3p3 w=34 l=6
X12 Y A VSS VSS nmos_3p3 w=17 l=6
X13 Y A VSS VSS nmos_3p3 w=17 l=6
X14 Y A VSS VSS nmos_3p3 w=17 l=6
X15 Y A VSS VSS nmos_3p3 w=17 l=6
X16 VSS A Y VSS nmos_3p3 w=17 l=6
X17 VSS A Y VSS nmos_3p3 w=17 l=6
X18 Y A VSS VSS nmos_3p3 w=17 l=6
X19 Y A VSS VSS nmos_3p3 w=17 l=6
X20 VSS A Y VSS nmos_3p3 w=17 l=6
X21 VDD A Y VDD pmos_3p3 w=34 l=6
X22 Y A VDD VDD pmos_3p3 w=34 l=6
X23 VSS A Y VSS nmos_3p3 w=17 l=6
X24 VSS A Y VSS nmos_3p3 w=17 l=6
X25 VSS A Y VSS nmos_3p3 w=17 l=6
X26 Y A VDD VDD pmos_3p3 w=34 l=6
X27 VDD A Y VDD pmos_3p3 w=34 l=6
X28 Y A VDD VDD pmos_3p3 w=34 l=6
X29 VDD A Y VDD pmos_3p3 w=34 l=6
X30 VDD A Y VDD pmos_3p3 w=34 l=6
X31 Y A VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dff_1 D Q QN CLK
X0 a_75_109 a_52_14 a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 CLK a_42_109 VDD pmos_3p3 w=34 l=6
X2 a_135_68 a_114_19 VDD VDD pmos_3p3 w=34 l=6
X3 Q QN VSS VSS nmos_3p3 w=17 l=6
X4 a_131_19 a_52_14 a_114_19 VSS nmos_3p3 w=17 l=6
X5 a_42_109 D VDD VDD pmos_3p3 w=34 l=6
X6 a_135_68 a_114_19 VSS VSS nmos_3p3 w=17 l=6
X7 VDD a_19_14 a_9_19 VDD pmos_3p3 w=34 l=6
X8 a_75_19 CLK a_19_14 VSS nmos_3p3 w=17 l=6
X9 VSS a_135_68 a_131_19 VSS nmos_3p3 w=17 l=6
X10 a_19_14 a_52_14 a_42_19 VSS nmos_3p3 w=17 l=6
X11 VSS a_19_14 a_9_19 VSS nmos_3p3 w=17 l=6
X12 a_52_14 CLK VDD VDD pmos_3p3 w=34 l=6
X13 VDD a_135_68 a_131_109 VDD pmos_3p3 w=34 l=6
X14 a_131_109 CLK a_114_19 VDD pmos_3p3 w=34 l=6
X15 VSS a_135_68 QN VSS nmos_3p3 w=17 l=6
X16 a_114_19 a_52_14 a_103_109 VDD pmos_3p3 w=34 l=6
X17 a_114_19 CLK a_103_19 VSS nmos_3p3 w=17 l=6
X18 a_52_14 CLK VSS VSS nmos_3p3 w=17 l=6
X19 a_103_109 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X20 a_42_19 D VSS VSS nmos_3p3 w=17 l=6
X21 VDD a_9_19 a_75_109 VDD pmos_3p3 w=34 l=6
X22 a_103_19 a_9_19 VSS VSS nmos_3p3 w=17 l=6
X23 Q QN VDD VDD pmos_3p3 w=34 l=6
X24 VDD a_135_68 QN VDD pmos_3p3 w=34 l=6
X25 VSS a_9_19 a_75_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dffn_1 D Q QN CLKN
X0 a_75_109 a_52_14 a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 CLKN a_42_109 VDD pmos_3p3 w=34 l=6
X2 a_135_68 a_114_19 VDD VDD pmos_3p3 w=34 l=6
X3 Q QN VSS VSS nmos_3p3 w=17 l=6
X4 a_131_19 a_52_14 a_114_19 VSS nmos_3p3 w=17 l=6
X5 a_42_109 D VDD VDD pmos_3p3 w=34 l=6
X6 a_135_68 a_114_19 VSS VSS nmos_3p3 w=17 l=6
X7 VDD a_19_14 a_9_19 VDD pmos_3p3 w=34 l=6
X8 a_75_19 CLKN a_19_14 VSS nmos_3p3 w=17 l=6
X9 VSS a_135_68 a_131_19 VSS nmos_3p3 w=17 l=6
X10 a_19_14 a_52_14 a_42_19 VSS nmos_3p3 w=17 l=6
X11 VSS a_19_14 a_9_19 VSS nmos_3p3 w=17 l=6
X12 a_52_14 CLKN VDD VDD pmos_3p3 w=34 l=6
X13 VDD a_135_68 a_131_109 VDD pmos_3p3 w=34 l=6
X14 a_131_109 CLKN a_114_19 VDD pmos_3p3 w=34 l=6
X15 VSS a_135_68 QN VSS nmos_3p3 w=17 l=6
X16 a_114_19 a_52_14 a_103_109 VDD pmos_3p3 w=34 l=6
X17 a_114_19 CLKN a_103_19 VSS nmos_3p3 w=17 l=6
X18 a_52_14 CLKN VSS VSS nmos_3p3 w=17 l=6
X19 a_103_109 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X20 a_42_19 D VSS VSS nmos_3p3 w=17 l=6
X21 VDD a_9_19 a_75_109 VDD pmos_3p3 w=34 l=6
X22 a_103_19 a_9_19 VSS VSS nmos_3p3 w=17 l=6
X23 Q QN VDD VDD pmos_3p3 w=34 l=6
X24 VDD a_135_68 QN VDD pmos_3p3 w=34 l=6
X25 VSS a_9_19 a_75_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dffsr_1 D SN RN Q QN CLK
X0 a_156_109 a_133_14 a_82_14 VDD pmos_3p3 w=34 l=6
X1 VSS a_41_109 a_156_19 VSS nmos_3p3 w=17 l=6
X2 a_82_14 CLK a_123_109 VDD pmos_3p3 w=34 l=6
X3 a_212_109 CLK a_195_19 VDD pmos_3p3 w=34 l=6
X4 VSS a_25_19 a_216_68 VSS nmos_3p3 w=17 l=6
X5 a_195_19 CLK a_184_19 VSS nmos_3p3 w=17 l=6
X6 a_133_14 CLK VSS VSS nmos_3p3 w=17 l=6
X7 a_216_68 SN a_275_19 VSS nmos_3p3 w=17 l=6
X8 a_25_19 RN VDD VDD pmos_3p3 w=34 l=6
X9 a_123_109 D VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_216_68 QN VDD pmos_3p3 w=34 l=6
X11 Q QN VDD VDD pmos_3p3 w=34 l=6
X12 a_41_109 a_25_19 VSS VSS nmos_3p3 w=17 l=6
X13 a_25_19 RN VSS VSS nmos_3p3 w=17 l=6
X14 a_82_14 a_133_14 a_123_19 VSS nmos_3p3 w=17 l=6
X15 a_256_109 SN VDD VDD pmos_3p3 w=34 l=6
X16 a_275_19 a_195_19 VSS VSS nmos_3p3 w=17 l=6
X17 VDD a_195_19 a_256_109 VDD pmos_3p3 w=34 l=6
X18 a_212_19 a_133_14 a_195_19 VSS nmos_3p3 w=17 l=6
X19 a_216_68 a_25_19 a_256_109 VDD pmos_3p3 w=34 l=6
X20 VSS a_216_68 a_212_19 VSS nmos_3p3 w=17 l=6
X21 a_77_19 SN a_41_109 VSS nmos_3p3 w=17 l=6
X22 a_57_109 a_82_14 VDD VDD pmos_3p3 w=34 l=6
X23 a_57_109 a_25_19 a_41_109 VDD pmos_3p3 w=34 l=6
X24 VDD SN a_57_109 VDD pmos_3p3 w=34 l=6
X25 a_195_19 a_133_14 a_184_109 VDD pmos_3p3 w=34 l=6
X26 Q QN VSS VSS nmos_3p3 w=17 l=6
X27 a_184_109 a_41_109 VDD VDD pmos_3p3 w=34 l=6
X28 VSS a_82_14 a_77_19 VSS nmos_3p3 w=17 l=6
X29 a_156_19 CLK a_82_14 VSS nmos_3p3 w=17 l=6
X30 VDD a_41_109 a_156_109 VDD pmos_3p3 w=34 l=6
X31 a_133_14 CLK VDD VDD pmos_3p3 w=34 l=6
X32 a_123_19 D VSS VSS nmos_3p3 w=17 l=6
X33 VDD a_216_68 a_212_109 VDD pmos_3p3 w=34 l=6
X34 a_184_19 a_41_109 VSS VSS nmos_3p3 w=17 l=6
X35 VSS a_216_68 QN VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dlat_1 D CLK Q
X0 a_52_92 CLK VDD VDD pmos_3p3 w=34 l=6
X1 a_46_19 D VSS VSS nmos_3p3 w=17 l=6
X2 a_20_14 CLK a_46_19 VSS nmos_3p3 w=17 l=6
X3 VSS a_10_19 a_127_19 VSS nmos_3p3 w=17 l=6
X4 VDD a_10_19 a_77_109 VDD pmos_3p3 w=34 l=6
X5 a_77_109 CLK a_20_14 VDD pmos_3p3 w=34 l=6
X6 a_20_14 a_52_92 a_43_109 VDD pmos_3p3 w=34 l=6
X7 VDD a_20_14 a_10_19 VDD pmos_3p3 w=34 l=6
X8 a_43_109 D VDD VDD pmos_3p3 w=34 l=6
X9 Q a_127_19 VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_10_19 a_127_19 VDD pmos_3p3 w=34 l=6
X11 a_77_19 a_52_92 a_20_14 VSS nmos_3p3 w=17 l=6
X12 Q a_127_19 VSS VSS nmos_3p3 w=17 l=6
X13 VSS a_10_19 a_77_19 VSS nmos_3p3 w=17 l=6
X14 a_52_92 CLK VSS VSS nmos_3p3 w=17 l=6
X15 VSS a_20_14 a_10_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dlatn_1 D Q CLKN
X0 a_52_92 CLKN VDD VDD pmos_3p3 w=34 l=6
X1 a_46_19 D VSS VSS nmos_3p3 w=17 l=6
X2 a_20_14 CLKN a_46_19 VSS nmos_3p3 w=17 l=6
X3 VSS a_10_19 a_127_19 VSS nmos_3p3 w=17 l=6
X4 VDD a_10_19 a_77_109 VDD pmos_3p3 w=34 l=6
X5 a_77_109 CLKN a_20_14 VDD pmos_3p3 w=34 l=6
X6 a_20_14 a_52_92 a_43_109 VDD pmos_3p3 w=34 l=6
X7 VDD a_20_14 a_10_19 VDD pmos_3p3 w=34 l=6
X8 a_43_109 D VDD VDD pmos_3p3 w=34 l=6
X9 Q a_127_19 VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_10_19 a_127_19 VDD pmos_3p3 w=34 l=6
X11 a_77_19 a_52_92 a_20_14 VSS nmos_3p3 w=17 l=6
X12 Q a_127_19 VSS VSS nmos_3p3 w=17 l=6
X13 VSS a_10_19 a_77_19 VSS nmos_3p3 w=17 l=6
X14 a_52_92 CLKN VSS VSS nmos_3p3 w=17 l=6
X15 VSS a_20_14 a_10_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_1
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_2
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_4
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_8
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_16
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_inv_1 A Y
X0 Y A VDD VDD pmos_3p3 w=34 l=6
X1 Y A VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_inv_2 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 Y A VSS VSS nmos_3p3 w=17 l=6
X3 VSS A Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_inv_4 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 VDD A Y VDD pmos_3p3 w=34 l=6
X3 Y A VDD VDD pmos_3p3 w=34 l=6
X4 Y A VSS VSS nmos_3p3 w=17 l=6
X5 Y A VSS VSS nmos_3p3 w=17 l=6
X6 VSS A Y VSS nmos_3p3 w=17 l=6
X7 VSS A Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_inv_8 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 VDD A Y VDD pmos_3p3 w=34 l=6
X2 Y A VDD VDD pmos_3p3 w=34 l=6
X3 Y A VDD VDD pmos_3p3 w=34 l=6
X4 VDD A Y VDD pmos_3p3 w=34 l=6
X5 VSS A Y VSS nmos_3p3 w=17 l=6
X6 Y A VDD VDD pmos_3p3 w=34 l=6
X7 Y A VSS VSS nmos_3p3 w=17 l=6
X8 Y A VSS VSS nmos_3p3 w=17 l=6
X9 Y A VSS VSS nmos_3p3 w=17 l=6
X10 Y A VSS VSS nmos_3p3 w=17 l=6
X11 VSS A Y VSS nmos_3p3 w=17 l=6
X12 VSS A Y VSS nmos_3p3 w=17 l=6
X13 VSS A Y VSS nmos_3p3 w=17 l=6
X14 Y A VDD VDD pmos_3p3 w=34 l=6
X15 VDD A Y VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_inv_16 A Y
X0 VDD A Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 Y A VSS VSS nmos_3p3 w=17 l=6
X3 VDD A Y VDD pmos_3p3 w=34 l=6
X4 Y A VSS VSS nmos_3p3 w=17 l=6
X5 VDD A Y VDD pmos_3p3 w=34 l=6
X6 Y A VDD VDD pmos_3p3 w=34 l=6
X7 Y A VDD VDD pmos_3p3 w=34 l=6
X8 VSS A Y VSS nmos_3p3 w=17 l=6
X9 VDD A Y VDD pmos_3p3 w=34 l=6
X10 VSS A Y VSS nmos_3p3 w=17 l=6
X11 Y A VDD VDD pmos_3p3 w=34 l=6
X12 Y A VSS VSS nmos_3p3 w=17 l=6
X13 Y A VSS VSS nmos_3p3 w=17 l=6
X14 Y A VSS VSS nmos_3p3 w=17 l=6
X15 Y A VSS VSS nmos_3p3 w=17 l=6
X16 VSS A Y VSS nmos_3p3 w=17 l=6
X17 VSS A Y VSS nmos_3p3 w=17 l=6
X18 Y A VSS VSS nmos_3p3 w=17 l=6
X19 Y A VSS VSS nmos_3p3 w=17 l=6
X20 VSS A Y VSS nmos_3p3 w=17 l=6
X21 VDD A Y VDD pmos_3p3 w=34 l=6
X22 Y A VDD VDD pmos_3p3 w=34 l=6
X23 VSS A Y VSS nmos_3p3 w=17 l=6
X24 VSS A Y VSS nmos_3p3 w=17 l=6
X25 VSS A Y VSS nmos_3p3 w=17 l=6
X26 Y A VDD VDD pmos_3p3 w=34 l=6
X27 VDD A Y VDD pmos_3p3 w=34 l=6
X28 Y A VDD VDD pmos_3p3 w=34 l=6
X29 VDD A Y VDD pmos_3p3 w=34 l=6
X30 VDD A Y VDD pmos_3p3 w=34 l=6
X31 Y A VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_mux2_1 Y Sel A B
X0 B a_25_19 Y VDD pmos_3p3 w=34 l=6
X1 Y Sel A VDD pmos_3p3 w=34 l=6
X2 a_25_19 Sel VDD VDD pmos_3p3 w=34 l=6
X3 Y a_25_19 A VSS nmos_3p3 w=17 l=6
X4 a_25_19 Sel VSS VSS nmos_3p3 w=17 l=6
X5 B Sel Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_nand2_1 A B Y
X0 VDD B Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 a_28_19 A Y VSS nmos_3p3 w=17 l=6
X3 VSS B a_28_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_nor2_1 A Y B
X0 Y B a_25_109 VDD pmos_3p3 w=34 l=6
X1 a_25_109 A VDD VDD pmos_3p3 w=34 l=6
X2 Y A VSS VSS nmos_3p3 w=17 l=6
X3 VSS B Y VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_oai21_1 Y A0 A1 B
X0 Y B a_8_19 VSS nmos_3p3 w=17 l=6
X1 VSS A0 a_8_19 VSS nmos_3p3 w=17 l=6
X2 a_27_109 A0 VDD VDD pmos_3p3 w=34 l=6
X3 VDD B Y VDD pmos_3p3 w=34 l=6
X4 Y A1 a_27_109 VDD pmos_3p3 w=34 l=6
X5 a_8_19 A1 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_or2_1 B A Y
X0 VDD B a_25_109 VDD pmos_3p3 w=34 l=6
X1 a_25_109 A a_9_109 VDD pmos_3p3 w=34 l=6
X2 Y a_9_109 VSS VSS nmos_3p3 w=17 l=6
X3 a_9_109 A VSS VSS nmos_3p3 w=17 l=6
X4 Y a_9_109 VDD VDD pmos_3p3 w=34 l=6
X5 VSS B a_9_109 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_tiehi Y
X0 Y a_19_14 VDD VDD pmos_3p3 w=34 l=6
X1 a_19_14 a_19_14 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_tielo Y
X0 a_19_14 a_19_14 VDD VDD pmos_3p3 w=34 l=6
X1 Y a_19_14 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_xnor2_1 A Y B
X0 Y a_47_14 a_42_19 VSS nmos_3p3 w=17 l=6
X1 VDD B a_76_109 VDD pmos_3p3 w=34 l=6
X2 a_47_14 B VDD VDD pmos_3p3 w=34 l=6
X3 Y a_47_14 a_42_109 VDD pmos_3p3 w=34 l=6
X4 a_76_109 A Y VDD pmos_3p3 w=34 l=6
X5 a_42_109 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X6 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X7 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X8 a_76_19 a_9_19 Y VSS nmos_3p3 w=17 l=6
X9 a_42_19 A VSS VSS nmos_3p3 w=17 l=6
X10 a_47_14 B VSS VSS nmos_3p3 w=17 l=6
X11 VSS B a_76_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_xor2_1 A Y B
X0 Y B a_42_19 VSS nmos_3p3 w=17 l=6
X1 VDD B a_76_109 VDD pmos_3p3 w=34 l=6
X2 a_47_94 B VDD VDD pmos_3p3 w=34 l=6
X3 Y a_47_94 a_42_109 VDD pmos_3p3 w=34 l=6
X4 a_76_109 a_9_19 Y VDD pmos_3p3 w=34 l=6
X5 a_42_109 A VDD VDD pmos_3p3 w=34 l=6
X6 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X7 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X8 a_76_19 a_9_19 Y VSS nmos_3p3 w=17 l=6
X9 a_42_19 A VSS VSS nmos_3p3 w=17 l=6
X10 a_47_94 B VSS VSS nmos_3p3 w=17 l=6
X11 VSS a_47_94 a_76_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary


******* EOF

