magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 2203 2345 3203 47857
rect 87011 2345 88011 47857
<< metal2 >>
rect 2627 2345 3627 47857
rect 86587 2345 87587 47839
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_0
timestamp 1669390400
transform 1 0 59432 0 1 2876
box -162 -224 162 224
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_1
timestamp 1669390400
transform 1 0 60052 0 1 4068
box -162 -224 162 224
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_2
timestamp 1669390400
transform 1 0 29524 0 1 2876
box -162 -224 162 224
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_3
timestamp 1669390400
transform 1 0 28915 0 1 4068
box -162 -224 162 224
use M3_M2431058998327_64x8m81  M3_M2431058998327_64x8m81_0
timestamp 1669390400
transform 1 0 60052 0 1 4068
box -162 -224 162 224
use M3_M2431058998327_64x8m81  M3_M2431058998327_64x8m81_1
timestamp 1669390400
transform 1 0 28915 0 1 4068
box -162 -224 162 224
use power_route_01_64x8m81  power_route_01_64x8m81_0
timestamp 1669390400
transform -1 0 85469 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_1
timestamp 1669390400
transform -1 0 25893 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_2
timestamp 1669390400
transform 1 0 9233 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_3
timestamp 1669390400
transform 1 0 20033 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_4
timestamp 1669390400
transform 1 0 14633 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_5
timestamp 1669390400
transform 1 0 63409 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_6
timestamp 1669390400
transform 1 0 79609 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_7
timestamp 1669390400
transform 1 0 74209 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_8
timestamp 1669390400
transform 1 0 68809 0 1 46214
box -511 0 1714 2425
use power_route_01_64x8m81  power_route_01_64x8m81_9
timestamp 1669390400
transform 1 0 3833 0 1 46214
box -511 0 1714 2425
use power_route_02_a_64x8m81  power_route_02_a_64x8m81_0
timestamp 1669390400
transform 1 0 -1418 0 1 41689
box 3339 -250 30611 1350
use power_route_02_a_64x8m81  power_route_02_a_64x8m81_1
timestamp 1669390400
transform 1 0 -1418 0 1 45289
box 3339 -250 30611 1350
use power_route_02_a_64x8m81  power_route_02_a_64x8m81_2
timestamp 1669390400
transform 1 0 -1418 0 1 43489
box 3339 -250 30611 1350
use power_route_02_a_64x8m81  power_route_02_a_64x8m81_3
timestamp 1669390400
transform 1 0 -1418 0 1 38089
box 3339 -250 30611 1350
use power_route_02_a_64x8m81  power_route_02_a_64x8m81_4
timestamp 1669390400
transform 1 0 -1418 0 1 39889
box 3339 -250 30611 1350
use power_route_02_b_64x8m81  power_route_02_b_64x8m81_0
timestamp 1669390400
transform -1 0 91632 0 1 39889
box 3339 -250 30290 1350
use power_route_02_b_64x8m81  power_route_02_b_64x8m81_1
timestamp 1669390400
transform -1 0 91632 0 1 41689
box 3339 -250 30290 1350
use power_route_02_b_64x8m81  power_route_02_b_64x8m81_2
timestamp 1669390400
transform -1 0 91632 0 1 43489
box 3339 -250 30290 1350
use power_route_02_b_64x8m81  power_route_02_b_64x8m81_3
timestamp 1669390400
transform -1 0 91632 0 1 45289
box 3339 -250 30290 1350
use power_route_02_b_64x8m81  power_route_02_b_64x8m81_4
timestamp 1669390400
transform -1 0 91632 0 1 38089
box 3339 -250 30290 1350
use power_route_04_64x8m81  power_route_04_64x8m81_0
timestamp 1669390400
transform -1 0 91632 0 1 244
box 3339 2101 6632 47613
use power_route_04_64x8m81  power_route_04_64x8m81_1
timestamp 1669390400
transform 1 0 -1418 0 1 244
box 3339 2101 6632 47613
use power_route_05_64x8m81  power_route_05_64x8m81_0
timestamp 1669390400
transform 1 0 19656 0 1 230
box -8 2115 1235 7462
use power_route_05_64x8m81  power_route_05_64x8m81_1
timestamp 1669390400
transform 1 0 68432 0 1 230
box -8 2115 1235 7462
use power_route_05_64x8m81  power_route_05_64x8m81_2
timestamp 1669390400
transform 1 0 79232 0 1 230
box -8 2115 1235 7462
use power_route_05_64x8m81  power_route_05_64x8m81_3
timestamp 1669390400
transform 1 0 8856 0 1 230
box -8 2115 1235 7462
use power_route_06_64x8m81  power_route_06_64x8m81_0
timestamp 1669390400
transform 1 0 61241 0 1 230
box -7 2115 1234 18431
use power_route_06_64x8m81  power_route_06_64x8m81_1
timestamp 1669390400
transform 1 0 26784 0 1 230
box -7 2115 1234 18431
use power_route_07_64x8m81  power_route_07_64x8m81_0
timestamp 1669390400
transform 1 0 40746 0 1 230
box -8 3065 1235 7462
use power_route_07_64x8m81  power_route_07_64x8m81_1
timestamp 1669390400
transform 1 0 38926 0 1 230
box -8 3065 1235 7462
<< properties >>
string GDS_END 2272018
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2269944
string path 15.635 239.285 15.635 11.725 
<< end >>
