magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect -31 1318 89 1389
rect -31 -71 89 -1
use nmos_5p043105908781100_256x8m81  nmos_5p043105908781100_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -88 -44 208 1362
<< properties >>
string GDS_END 1886448
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1886196
<< end >>
