magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal2 >>
rect -7 7964 217 18431
rect -7 7908 16 7964
rect 72 7908 140 7964
rect 196 7908 217 7964
rect -7 7840 217 7908
rect -7 7784 16 7840
rect 72 7784 140 7840
rect 196 7784 217 7840
rect -7 7716 217 7784
rect -7 7660 16 7716
rect 72 7660 140 7716
rect 196 7660 217 7716
rect -7 5680 217 7660
rect -7 5624 16 5680
rect 72 5624 140 5680
rect 196 5624 217 5680
rect -7 5556 217 5624
rect -7 5500 16 5556
rect 72 5500 140 5556
rect 196 5500 217 5556
rect -7 5432 217 5500
rect -7 5376 16 5432
rect 72 5376 140 5432
rect 196 5376 217 5432
rect -7 4667 217 5376
rect -7 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 217 4667
rect -7 4543 217 4611
rect -7 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 217 4543
rect -7 4419 217 4487
rect -7 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 217 4419
rect -7 2115 217 4363
rect 495 7366 719 16012
rect 495 7310 516 7366
rect 572 7310 640 7366
rect 696 7310 719 7366
rect 495 7242 719 7310
rect 495 7186 516 7242
rect 572 7186 640 7242
rect 696 7186 719 7242
rect 495 7118 719 7186
rect 495 7062 516 7118
rect 572 7062 640 7118
rect 696 7062 719 7118
rect 495 6403 719 7062
rect 495 6347 516 6403
rect 572 6347 640 6403
rect 696 6347 719 6403
rect 495 6279 719 6347
rect 495 6223 516 6279
rect 572 6223 640 6279
rect 696 6223 719 6279
rect 495 6155 719 6223
rect 495 6099 516 6155
rect 572 6099 640 6155
rect 696 6099 719 6155
rect 495 3065 719 6099
rect 1010 7964 1234 18431
rect 1010 7908 1033 7964
rect 1089 7908 1157 7964
rect 1213 7908 1234 7964
rect 1010 7840 1234 7908
rect 1010 7784 1033 7840
rect 1089 7784 1157 7840
rect 1213 7784 1234 7840
rect 1010 7716 1234 7784
rect 1010 7660 1033 7716
rect 1089 7660 1157 7716
rect 1213 7660 1234 7716
rect 1010 5680 1234 7660
rect 1010 5624 1033 5680
rect 1089 5624 1157 5680
rect 1213 5624 1234 5680
rect 1010 5556 1234 5624
rect 1010 5500 1033 5556
rect 1089 5500 1157 5556
rect 1213 5500 1234 5556
rect 1010 5432 1234 5500
rect 1010 5376 1033 5432
rect 1089 5376 1157 5432
rect 1213 5376 1234 5432
rect 1010 4667 1234 5376
rect 1010 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1234 4667
rect 1010 4543 1234 4611
rect 1010 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1234 4543
rect 1010 4419 1234 4487
rect 1010 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1234 4419
rect 1010 2115 1234 4363
<< via2 >>
rect 16 7908 72 7964
rect 140 7908 196 7964
rect 16 7784 72 7840
rect 140 7784 196 7840
rect 16 7660 72 7716
rect 140 7660 196 7716
rect 16 5624 72 5680
rect 140 5624 196 5680
rect 16 5500 72 5556
rect 140 5500 196 5556
rect 16 5376 72 5432
rect 140 5376 196 5432
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 516 7310 572 7366
rect 640 7310 696 7366
rect 516 7186 572 7242
rect 640 7186 696 7242
rect 516 7062 572 7118
rect 640 7062 696 7118
rect 516 6347 572 6403
rect 640 6347 696 6403
rect 516 6223 572 6279
rect 640 6223 696 6279
rect 516 6099 572 6155
rect 640 6099 696 6155
rect 1033 7908 1089 7964
rect 1157 7908 1213 7964
rect 1033 7784 1089 7840
rect 1157 7784 1213 7840
rect 1033 7660 1089 7716
rect 1157 7660 1213 7716
rect 1033 5624 1089 5680
rect 1157 5624 1213 5680
rect 1033 5500 1089 5556
rect 1157 5500 1213 5556
rect 1033 5376 1089 5432
rect 1157 5376 1213 5432
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 6 7964 206 7974
rect 6 7908 16 7964
rect 72 7908 140 7964
rect 196 7908 206 7964
rect 6 7840 206 7908
rect 6 7784 16 7840
rect 72 7784 140 7840
rect 196 7784 206 7840
rect 6 7716 206 7784
rect 6 7660 16 7716
rect 72 7660 140 7716
rect 196 7660 206 7716
rect 6 7650 206 7660
rect 1023 7964 1223 7974
rect 1023 7908 1033 7964
rect 1089 7908 1157 7964
rect 1213 7908 1223 7964
rect 1023 7840 1223 7908
rect 1023 7784 1033 7840
rect 1089 7784 1157 7840
rect 1213 7784 1223 7840
rect 1023 7716 1223 7784
rect 1023 7660 1033 7716
rect 1089 7660 1157 7716
rect 1213 7660 1223 7716
rect 1023 7650 1223 7660
rect 506 7366 706 7376
rect 506 7310 516 7366
rect 572 7310 640 7366
rect 696 7310 706 7366
rect 506 7242 706 7310
rect 506 7186 516 7242
rect 572 7186 640 7242
rect 696 7186 706 7242
rect 506 7118 706 7186
rect 506 7062 516 7118
rect 572 7062 640 7118
rect 696 7062 706 7118
rect 506 7052 706 7062
rect 506 6403 706 6413
rect 506 6347 516 6403
rect 572 6347 640 6403
rect 696 6347 706 6403
rect 506 6279 706 6347
rect 506 6223 516 6279
rect 572 6223 640 6279
rect 696 6223 706 6279
rect 506 6155 706 6223
rect 506 6099 516 6155
rect 572 6099 640 6155
rect 696 6099 706 6155
rect 506 6089 706 6099
rect 6 5680 206 5690
rect 6 5624 16 5680
rect 72 5624 140 5680
rect 196 5624 206 5680
rect 6 5556 206 5624
rect 6 5500 16 5556
rect 72 5500 140 5556
rect 196 5500 206 5556
rect 6 5432 206 5500
rect 6 5376 16 5432
rect 72 5376 140 5432
rect 196 5376 206 5432
rect 6 5366 206 5376
rect 1023 5680 1223 5690
rect 1023 5624 1033 5680
rect 1089 5624 1157 5680
rect 1213 5624 1223 5680
rect 1023 5556 1223 5624
rect 1023 5500 1033 5556
rect 1089 5500 1157 5556
rect 1213 5500 1223 5556
rect 1023 5432 1223 5500
rect 1023 5376 1033 5432
rect 1089 5376 1157 5432
rect 1213 5376 1223 5432
rect 1023 5366 1223 5376
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_0
timestamp 1669390400
transform 1 0 1120 0 1 2599
box -100 -472 100 472
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_1
timestamp 1669390400
transform 1 0 103 0 1 2599
box -100 -472 100 472
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 6251
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_1
timestamp 1669390400
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_2
timestamp 1669390400
transform 1 0 106 0 1 5528
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_3
timestamp 1669390400
transform 1 0 1123 0 1 5528
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_4
timestamp 1669390400
transform 1 0 606 0 1 7214
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_5
timestamp 1669390400
transform 1 0 1123 0 1 7812
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_6
timestamp 1669390400
transform 1 0 106 0 1 7812
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_7
timestamp 1669390400
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_0
timestamp 1669390400
transform 1 0 106 0 1 9127
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_1
timestamp 1669390400
transform 1 0 106 0 1 13016
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_2
timestamp 1669390400
transform 1 0 1123 0 1 13016
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_3
timestamp 1669390400
transform 1 0 106 0 1 12329
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_4
timestamp 1669390400
transform 1 0 1123 0 1 12329
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_5
timestamp 1669390400
transform 1 0 106 0 1 17993
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_6
timestamp 1669390400
transform 1 0 1123 0 1 17993
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_7
timestamp 1669390400
transform 1 0 106 0 1 17306
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_8
timestamp 1669390400
transform 1 0 1123 0 1 17306
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_9
timestamp 1669390400
transform 1 0 106 0 1 16622
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_10
timestamp 1669390400
transform 1 0 1123 0 1 16622
box -100 -286 100 286
use M3_M24310590878172_256x8m81  M3_M24310590878172_256x8m81_11
timestamp 1669390400
transform 1 0 1123 0 1 9127
box -100 -286 100 286
use M3_M24310590878173_256x8m81  M3_M24310590878173_256x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 14944
box -100 -906 100 906
use M3_M24310590878174_256x8m81  M3_M24310590878174_256x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 10647
box -100 -596 100 596
use M3_M24310590878175_256x8m81  M3_M24310590878175_256x8m81_0
timestamp 1669390400
transform 1 0 606 0 1 3575
box -100 -472 100 472
<< properties >>
string GDS_END 1923520
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1922024
<< end >>
