magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 2550 870
<< pwell >>
rect -86 -86 2550 352
<< mvnmos >>
rect 124 87 244 179
rect 384 87 504 165
rect 752 86 872 165
rect 920 86 1040 165
rect 1144 86 1264 165
rect 1404 86 1524 179
rect 1628 86 1748 179
rect 1996 68 2116 232
rect 2220 68 2340 232
<< mvpmos >>
rect 124 532 224 716
rect 384 591 484 716
rect 772 590 872 716
rect 920 590 1020 716
rect 1124 590 1224 716
rect 1364 531 1464 716
rect 1568 531 1668 716
rect 2016 472 2116 716
rect 2220 472 2320 716
<< mvndiff >>
rect 36 152 124 179
rect 36 106 49 152
rect 95 106 124 152
rect 36 87 124 106
rect 244 165 324 179
rect 1908 192 1996 232
rect 1324 165 1404 179
rect 244 152 384 165
rect 244 106 273 152
rect 319 106 384 152
rect 244 87 384 106
rect 504 152 592 165
rect 504 106 533 152
rect 579 106 592 152
rect 504 87 592 106
rect 664 152 752 165
rect 664 106 677 152
rect 723 106 752 152
rect 664 86 752 106
rect 872 86 920 165
rect 1040 152 1144 165
rect 1040 106 1069 152
rect 1115 106 1144 152
rect 1040 86 1144 106
rect 1264 86 1404 165
rect 1524 152 1628 179
rect 1524 106 1553 152
rect 1599 106 1628 152
rect 1524 86 1628 106
rect 1748 152 1836 179
rect 1748 106 1777 152
rect 1823 106 1836 152
rect 1748 86 1836 106
rect 1908 146 1921 192
rect 1967 146 1996 192
rect 1908 68 1996 146
rect 2116 192 2220 232
rect 2116 146 2145 192
rect 2191 146 2220 192
rect 2116 68 2220 146
rect 2340 192 2428 232
rect 2340 146 2369 192
rect 2415 146 2428 192
rect 2340 68 2428 146
<< mvpdiff >>
rect 36 667 124 716
rect 36 621 49 667
rect 95 621 124 667
rect 36 532 124 621
rect 224 667 384 716
rect 224 621 273 667
rect 319 621 384 667
rect 224 591 384 621
rect 484 667 592 716
rect 484 621 533 667
rect 579 621 592 667
rect 484 591 592 621
rect 684 674 772 716
rect 684 628 697 674
rect 743 628 772 674
rect 224 532 324 591
rect 684 590 772 628
rect 872 590 920 716
rect 1020 674 1124 716
rect 1020 628 1049 674
rect 1095 628 1124 674
rect 1020 590 1124 628
rect 1224 590 1364 716
rect 1284 531 1364 590
rect 1464 703 1568 716
rect 1464 563 1493 703
rect 1539 563 1568 703
rect 1464 531 1568 563
rect 1668 626 1756 716
rect 1668 580 1697 626
rect 1743 580 1756 626
rect 1668 531 1756 580
rect 1928 665 2016 716
rect 1928 525 1941 665
rect 1987 525 2016 665
rect 1928 472 2016 525
rect 2116 665 2220 716
rect 2116 525 2145 665
rect 2191 525 2220 665
rect 2116 472 2220 525
rect 2320 665 2408 716
rect 2320 525 2349 665
rect 2395 525 2408 665
rect 2320 472 2408 525
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 533 106 579 152
rect 677 106 723 152
rect 1069 106 1115 152
rect 1553 106 1599 152
rect 1777 106 1823 152
rect 1921 146 1967 192
rect 2145 146 2191 192
rect 2369 146 2415 192
<< mvpdiffc >>
rect 49 621 95 667
rect 273 621 319 667
rect 533 621 579 667
rect 697 628 743 674
rect 1049 628 1095 674
rect 1493 563 1539 703
rect 1697 580 1743 626
rect 1941 525 1987 665
rect 2145 525 2191 665
rect 2349 525 2395 665
<< polysilicon >>
rect 124 716 224 760
rect 384 716 484 760
rect 772 716 872 760
rect 920 716 1020 760
rect 1124 716 1224 760
rect 1364 716 1464 760
rect 1568 716 1668 760
rect 2016 716 2116 760
rect 2220 716 2320 760
rect 124 433 224 532
rect 384 526 484 591
rect 384 513 695 526
rect 384 467 636 513
rect 682 467 695 513
rect 384 454 695 467
rect 124 415 244 433
rect 124 369 179 415
rect 225 369 244 415
rect 124 179 244 369
rect 384 278 504 454
rect 772 352 872 590
rect 920 513 1020 590
rect 920 467 947 513
rect 993 467 1020 513
rect 1124 551 1224 590
rect 1124 505 1151 551
rect 1197 505 1224 551
rect 1124 492 1224 505
rect 920 444 1020 467
rect 1364 461 1464 531
rect 920 404 1264 444
rect 384 232 415 278
rect 461 232 504 278
rect 384 165 504 232
rect 752 295 872 352
rect 752 249 789 295
rect 835 249 872 295
rect 752 165 872 249
rect 920 259 1040 272
rect 920 213 957 259
rect 1003 213 1040 259
rect 920 165 1040 213
rect 1144 165 1264 404
rect 1364 415 1391 461
rect 1437 415 1464 461
rect 1568 419 1668 531
rect 1364 316 1464 415
rect 1404 294 1464 316
rect 1628 357 1668 419
rect 2016 357 2116 472
rect 2220 357 2320 472
rect 1628 311 2340 357
rect 1628 295 1748 311
rect 1404 179 1524 294
rect 1628 249 1651 295
rect 1697 249 1748 295
rect 1628 179 1748 249
rect 1996 232 2116 311
rect 2220 232 2340 311
rect 124 42 244 87
rect 384 42 504 87
rect 752 42 872 86
rect 920 42 1040 86
rect 1144 42 1264 86
rect 1404 42 1524 86
rect 1628 42 1748 86
rect 1996 24 2116 68
rect 2220 24 2340 68
<< polycontact >>
rect 636 467 682 513
rect 179 369 225 415
rect 947 467 993 513
rect 1151 505 1197 551
rect 415 232 461 278
rect 789 249 835 295
rect 957 213 1003 259
rect 1391 415 1437 461
rect 1651 249 1697 295
<< metal1 >>
rect 0 724 2464 844
rect 38 667 115 678
rect 38 621 49 667
rect 95 621 115 667
rect 38 278 115 621
rect 273 667 319 724
rect 273 610 319 621
rect 522 667 579 678
rect 522 621 533 667
rect 354 424 430 550
rect 165 415 430 424
rect 165 369 179 415
rect 225 369 430 415
rect 165 360 430 369
rect 522 417 579 621
rect 697 674 743 724
rect 1482 703 1550 724
rect 1020 628 1049 674
rect 1095 628 1301 674
rect 697 617 743 628
rect 1151 551 1197 562
rect 625 467 636 513
rect 682 467 947 513
rect 993 467 1020 513
rect 1151 417 1197 505
rect 522 371 1197 417
rect 38 232 415 278
rect 461 232 472 278
rect 38 152 115 232
rect 38 106 49 152
rect 95 106 115 152
rect 273 152 319 163
rect 522 152 590 371
rect 670 295 886 312
rect 670 249 789 295
rect 835 249 886 295
rect 670 248 886 249
rect 522 106 533 152
rect 579 106 590 152
rect 677 152 723 165
rect 800 110 886 248
rect 957 259 1003 371
rect 957 202 1003 213
rect 1255 295 1301 628
rect 1482 563 1493 703
rect 1539 563 1550 703
rect 1941 665 1987 724
rect 1482 561 1550 563
rect 1697 626 1743 645
rect 1697 461 1743 580
rect 1941 506 1987 525
rect 2132 665 2216 676
rect 2132 525 2145 665
rect 2191 525 2216 665
rect 1364 415 1391 461
rect 1437 415 1834 461
rect 1255 249 1651 295
rect 1697 249 1716 295
rect 1255 152 1301 249
rect 1040 106 1069 152
rect 1115 106 1301 152
rect 1553 152 1599 179
rect 1766 152 1834 415
rect 1766 106 1777 152
rect 1823 106 1834 152
rect 1921 192 1967 211
rect 273 60 319 106
rect 677 60 723 106
rect 1553 60 1599 106
rect 1921 60 1967 146
rect 2132 192 2216 525
rect 2349 665 2395 724
rect 2349 506 2395 525
rect 2132 146 2145 192
rect 2191 146 2216 192
rect 2132 106 2216 146
rect 2369 192 2415 211
rect 2369 60 2415 146
rect 0 -60 2464 60
<< labels >>
flabel metal1 s 2132 106 2216 676 0 FreeSans 400 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 724 2464 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2369 179 2415 211 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 670 248 886 312 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel metal1 s 354 424 430 550 0 FreeSans 400 0 0 0 E
port 2 nsew clock input
rlabel metal1 s 800 110 886 248 1 D
port 1 nsew default input
rlabel metal1 s 165 360 430 424 1 E
port 2 nsew clock input
rlabel metal1 s 2349 617 2395 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 617 1987 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 617 1550 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 697 617 743 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 617 319 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 610 2395 617 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 610 1987 617 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 610 1550 617 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 610 319 617 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 561 2395 610 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 561 1987 610 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 561 1550 610 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 506 2395 561 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 506 1987 561 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1921 179 1967 211 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 165 2415 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 165 1967 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 165 1599 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 163 2415 165 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 163 1967 165 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 163 1599 165 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 163 723 165 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 60 2415 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 60 1967 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 60 1599 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 60 723 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 163 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string GDS_END 580594
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 574928
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
