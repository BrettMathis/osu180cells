magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -286 -142 344 3179
<< polysilicon >>
rect -31 3039 88 3111
rect -31 -74 88 -1
use pmos_5p04310590878167_256x8m81  pmos_5p04310590878167_256x8m81_0
timestamp 1669390400
transform 1 0 -31 0 1 0
box -208 -120 328 3160
<< properties >>
string GDS_END 367676
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 367362
<< end >>
