magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 1232 844
rect 264 632 310 724
rect 672 632 718 724
rect 132 232 204 458
rect 356 232 428 458
rect 573 232 652 458
rect 672 60 718 153
rect 896 130 990 676
rect 1116 506 1162 724
rect 1120 60 1166 153
rect 0 -60 1232 60
<< obsm1 >>
rect 49 582 117 671
rect 49 531 850 582
rect 257 173 303 531
rect 804 289 850 531
rect 47 127 303 173
<< labels >>
rlabel metal1 s 132 232 204 458 6 A1
port 1 nsew default input
rlabel metal1 s 356 232 428 458 6 A2
port 2 nsew default input
rlabel metal1 s 573 232 652 458 6 A3
port 3 nsew default input
rlabel metal1 s 896 130 990 676 6 Z
port 4 nsew default output
rlabel metal1 s 0 724 1232 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1116 632 1162 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 672 632 718 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 264 632 310 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1116 506 1162 632 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1120 60 1166 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 672 60 718 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1232 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1232 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1203138
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1199666
<< end >>
