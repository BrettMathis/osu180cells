magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -1977 186 1977 246
rect -1977 140 -1920 186
rect -1874 140 -1762 186
rect -1716 140 -1604 186
rect -1558 140 -1446 186
rect -1400 140 -1288 186
rect -1242 140 -1130 186
rect -1084 140 -972 186
rect -926 140 -814 186
rect -768 140 -656 186
rect -610 140 -497 186
rect -451 140 -339 186
rect -293 140 -181 186
rect -135 140 -23 186
rect 23 140 135 186
rect 181 140 293 186
rect 339 140 451 186
rect 497 140 610 186
rect 656 140 768 186
rect 814 140 926 186
rect 972 140 1084 186
rect 1130 140 1242 186
rect 1288 140 1400 186
rect 1446 140 1558 186
rect 1604 140 1716 186
rect 1762 140 1874 186
rect 1920 140 1977 186
rect -1977 23 1977 140
rect -1977 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 1977 23
rect -1977 -140 1977 -23
rect -1977 -186 -1920 -140
rect -1874 -186 -1762 -140
rect -1716 -186 -1604 -140
rect -1558 -186 -1446 -140
rect -1400 -186 -1288 -140
rect -1242 -186 -1130 -140
rect -1084 -186 -972 -140
rect -926 -186 -814 -140
rect -768 -186 -656 -140
rect -610 -186 -497 -140
rect -451 -186 -339 -140
rect -293 -186 -181 -140
rect -135 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1242 -140
rect 1288 -186 1400 -140
rect 1446 -186 1558 -140
rect 1604 -186 1716 -140
rect 1762 -186 1874 -140
rect 1920 -186 1977 -140
rect -1977 -245 1977 -186
<< psubdiffcont >>
rect -1920 140 -1874 186
rect -1762 140 -1716 186
rect -1604 140 -1558 186
rect -1446 140 -1400 186
rect -1288 140 -1242 186
rect -1130 140 -1084 186
rect -972 140 -926 186
rect -814 140 -768 186
rect -656 140 -610 186
rect -497 140 -451 186
rect -339 140 -293 186
rect -181 140 -135 186
rect -23 140 23 186
rect 135 140 181 186
rect 293 140 339 186
rect 451 140 497 186
rect 610 140 656 186
rect 768 140 814 186
rect 926 140 972 186
rect 1084 140 1130 186
rect 1242 140 1288 186
rect 1400 140 1446 186
rect 1558 140 1604 186
rect 1716 140 1762 186
rect 1874 140 1920 186
rect -1920 -23 -1874 23
rect -1762 -23 -1716 23
rect -1604 -23 -1558 23
rect -1446 -23 -1400 23
rect -1288 -23 -1242 23
rect -1130 -23 -1084 23
rect -972 -23 -926 23
rect -814 -23 -768 23
rect -656 -23 -610 23
rect -497 -23 -451 23
rect -339 -23 -293 23
rect -181 -23 -135 23
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect 1242 -23 1288 23
rect 1400 -23 1446 23
rect 1558 -23 1604 23
rect 1716 -23 1762 23
rect 1874 -23 1920 23
rect -1920 -186 -1874 -140
rect -1762 -186 -1716 -140
rect -1604 -186 -1558 -140
rect -1446 -186 -1400 -140
rect -1288 -186 -1242 -140
rect -1130 -186 -1084 -140
rect -972 -186 -926 -140
rect -814 -186 -768 -140
rect -656 -186 -610 -140
rect -497 -186 -451 -140
rect -339 -186 -293 -140
rect -181 -186 -135 -140
rect -23 -186 23 -140
rect 135 -186 181 -140
rect 293 -186 339 -140
rect 451 -186 497 -140
rect 610 -186 656 -140
rect 768 -186 814 -140
rect 926 -186 972 -140
rect 1084 -186 1130 -140
rect 1242 -186 1288 -140
rect 1400 -186 1446 -140
rect 1558 -186 1604 -140
rect 1716 -186 1762 -140
rect 1874 -186 1920 -140
<< metal1 >>
rect -1969 186 1968 237
rect -1969 140 -1920 186
rect -1874 140 -1762 186
rect -1716 140 -1604 186
rect -1558 140 -1446 186
rect -1400 140 -1288 186
rect -1242 140 -1130 186
rect -1084 140 -972 186
rect -926 140 -814 186
rect -768 140 -656 186
rect -610 140 -497 186
rect -451 140 -339 186
rect -293 140 -181 186
rect -135 140 -23 186
rect 23 140 135 186
rect 181 140 293 186
rect 339 140 451 186
rect 497 140 610 186
rect 656 140 768 186
rect 814 140 926 186
rect 972 140 1084 186
rect 1130 140 1242 186
rect 1288 140 1400 186
rect 1446 140 1558 186
rect 1604 140 1716 186
rect 1762 140 1874 186
rect 1920 140 1968 186
rect -1969 23 1968 140
rect -1969 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 1968 23
rect -1969 -140 1968 -23
rect -1969 -186 -1920 -140
rect -1874 -186 -1762 -140
rect -1716 -186 -1604 -140
rect -1558 -186 -1446 -140
rect -1400 -186 -1288 -140
rect -1242 -186 -1130 -140
rect -1084 -186 -972 -140
rect -926 -186 -814 -140
rect -768 -186 -656 -140
rect -610 -186 -497 -140
rect -451 -186 -339 -140
rect -293 -186 -181 -140
rect -135 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1242 -140
rect 1288 -186 1400 -140
rect 1446 -186 1558 -140
rect 1604 -186 1716 -140
rect 1762 -186 1874 -140
rect 1920 -186 1968 -140
rect -1969 -237 1968 -186
<< properties >>
string GDS_END 1076718
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1071722
<< end >>
