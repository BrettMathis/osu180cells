magic
tech gf180mcuC
magscale 1 5
timestamp 1669390400
<< metal2 >>
rect -81 448 81 453
rect -81 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 81 448
rect -81 386 81 420
rect -81 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 81 386
rect -81 324 81 358
rect -81 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 81 324
rect -81 262 81 296
rect -81 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 81 262
rect -81 200 81 234
rect -81 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 81 200
rect -81 138 81 172
rect -81 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 81 138
rect -81 76 81 110
rect -81 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 81 76
rect -81 14 81 48
rect -81 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 81 14
rect -81 -48 81 -14
rect -81 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 81 -48
rect -81 -110 81 -76
rect -81 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 81 -110
rect -81 -172 81 -138
rect -81 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 81 -172
rect -81 -234 81 -200
rect -81 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 81 -234
rect -81 -296 81 -262
rect -81 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 81 -296
rect -81 -358 81 -324
rect -81 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 81 -358
rect -81 -420 81 -386
rect -81 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 81 -420
rect -81 -453 81 -448
<< via2 >>
rect -76 420 -48 448
rect -14 420 14 448
rect 48 420 76 448
rect -76 358 -48 386
rect -14 358 14 386
rect 48 358 76 386
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect -76 -386 -48 -358
rect -14 -386 14 -358
rect 48 -386 76 -358
rect -76 -448 -48 -420
rect -14 -448 14 -420
rect 48 -448 76 -420
<< metal3 >>
rect -81 448 81 453
rect -81 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 81 448
rect -81 386 81 420
rect -81 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 81 386
rect -81 324 81 358
rect -81 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 81 324
rect -81 262 81 296
rect -81 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 81 262
rect -81 200 81 234
rect -81 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 81 200
rect -81 138 81 172
rect -81 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 81 138
rect -81 76 81 110
rect -81 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 81 76
rect -81 14 81 48
rect -81 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 81 14
rect -81 -48 81 -14
rect -81 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 81 -48
rect -81 -110 81 -76
rect -81 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 81 -110
rect -81 -172 81 -138
rect -81 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 81 -172
rect -81 -234 81 -200
rect -81 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 81 -234
rect -81 -296 81 -262
rect -81 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 81 -296
rect -81 -358 81 -324
rect -81 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 81 -358
rect -81 -420 81 -386
rect -81 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 81 -420
rect -81 -453 81 -448
<< properties >>
string GDS_END 717312
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 714300
<< end >>
