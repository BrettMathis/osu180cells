magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -221 -1860 221 1860
<< nsubdiff >>
rect -78 1656 77 1713
rect -78 1610 -23 1656
rect 23 1610 77 1656
rect -78 1492 77 1610
rect -78 1446 -23 1492
rect 23 1446 77 1492
rect -78 1329 77 1446
rect -78 1283 -23 1329
rect 23 1283 77 1329
rect -78 1166 77 1283
rect -78 1120 -23 1166
rect 23 1120 77 1166
rect -78 1003 77 1120
rect -78 957 -23 1003
rect 23 957 77 1003
rect -78 839 77 957
rect -78 793 -23 839
rect 23 793 77 839
rect -78 676 77 793
rect -78 630 -23 676
rect 23 630 77 676
rect -78 513 77 630
rect -78 467 -23 513
rect 23 467 77 513
rect -78 350 77 467
rect -78 304 -23 350
rect 23 304 77 350
rect -78 186 77 304
rect -78 140 -23 186
rect 23 140 77 186
rect -78 23 77 140
rect -78 -23 -23 23
rect 23 -23 77 23
rect -78 -140 77 -23
rect -78 -186 -23 -140
rect 23 -186 77 -140
rect -78 -304 77 -186
rect -78 -350 -23 -304
rect 23 -350 77 -304
rect -78 -467 77 -350
rect -78 -513 -23 -467
rect 23 -513 77 -467
rect -78 -630 77 -513
rect -78 -676 -23 -630
rect 23 -676 77 -630
rect -78 -793 77 -676
rect -78 -839 -23 -793
rect 23 -839 77 -793
rect -78 -957 77 -839
rect -78 -1003 -23 -957
rect 23 -1003 77 -957
rect -78 -1120 77 -1003
rect -78 -1166 -23 -1120
rect 23 -1166 77 -1120
rect -78 -1283 77 -1166
rect -78 -1329 -23 -1283
rect 23 -1329 77 -1283
rect -78 -1446 77 -1329
rect -78 -1492 -23 -1446
rect 23 -1492 77 -1446
rect -78 -1610 77 -1492
rect -78 -1656 -23 -1610
rect 23 -1656 77 -1610
rect -78 -1712 77 -1656
<< nsubdiffcont >>
rect -23 1610 23 1656
rect -23 1446 23 1492
rect -23 1283 23 1329
rect -23 1120 23 1166
rect -23 957 23 1003
rect -23 793 23 839
rect -23 630 23 676
rect -23 467 23 513
rect -23 304 23 350
rect -23 140 23 186
rect -23 -23 23 23
rect -23 -186 23 -140
rect -23 -350 23 -304
rect -23 -513 23 -467
rect -23 -676 23 -630
rect -23 -839 23 -793
rect -23 -1003 23 -957
rect -23 -1166 23 -1120
rect -23 -1329 23 -1283
rect -23 -1492 23 -1446
rect -23 -1656 23 -1610
<< metal1 >>
rect -58 1656 58 1692
rect -58 1610 -23 1656
rect 23 1610 58 1656
rect -58 1492 58 1610
rect -58 1446 -23 1492
rect 23 1446 58 1492
rect -58 1329 58 1446
rect -58 1283 -23 1329
rect 23 1283 58 1329
rect -58 1166 58 1283
rect -58 1120 -23 1166
rect 23 1120 58 1166
rect -58 1003 58 1120
rect -58 957 -23 1003
rect 23 957 58 1003
rect -58 839 58 957
rect -58 793 -23 839
rect 23 793 58 839
rect -58 676 58 793
rect -58 630 -23 676
rect 23 630 58 676
rect -58 513 58 630
rect -58 467 -23 513
rect 23 467 58 513
rect -58 350 58 467
rect -58 304 -23 350
rect 23 304 58 350
rect -58 186 58 304
rect -58 140 -23 186
rect 23 140 58 186
rect -58 23 58 140
rect -58 -23 -23 23
rect 23 -23 58 23
rect -58 -140 58 -23
rect -58 -186 -23 -140
rect 23 -186 58 -140
rect -58 -304 58 -186
rect -58 -350 -23 -304
rect 23 -350 58 -304
rect -58 -467 58 -350
rect -58 -513 -23 -467
rect 23 -513 58 -467
rect -58 -630 58 -513
rect -58 -676 -23 -630
rect 23 -676 58 -630
rect -58 -793 58 -676
rect -58 -839 -23 -793
rect 23 -839 58 -793
rect -58 -957 58 -839
rect -58 -1003 -23 -957
rect 23 -1003 58 -957
rect -58 -1120 58 -1003
rect -58 -1166 -23 -1120
rect 23 -1166 58 -1120
rect -58 -1283 58 -1166
rect -58 -1329 -23 -1283
rect 23 -1329 58 -1283
rect -58 -1446 58 -1329
rect -58 -1492 -23 -1446
rect 23 -1492 58 -1446
rect -58 -1610 58 -1492
rect -58 -1656 -23 -1610
rect 23 -1656 58 -1610
rect -58 -1692 58 -1656
<< properties >>
string GDS_END 166542
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 164922
<< end >>
