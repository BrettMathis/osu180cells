magic
tech gf180mcuC
magscale 1 10
timestamp 1669650257
<< checkpaint >>
rect 44000 44000 73000 73000
<< metal3 >>
rect 46000 59461 49000 71000
tri 49000 59461 50249 60710 sw
tri 46000 58747 46714 59461 ne
rect 46714 58747 50249 59461
tri 50249 58747 50963 59461 sw
tri 46714 54498 50963 58747 ne
tri 50963 54498 55212 58747 sw
tri 50963 50249 55212 54498 ne
tri 55212 50249 59461 54498 sw
tri 55212 46000 59461 50249 ne
tri 59461 49000 60710 50249 sw
rect 59461 46000 71000 49000
<< end >>
